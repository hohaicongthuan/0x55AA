module layer_10_featuremap_259(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3978b012),
	.w1(32'hbbd4a3af),
	.w2(32'h3ae4058c),
	.w3(32'h38763971),
	.w4(32'h3a4ffea4),
	.w5(32'h396e5717),
	.w6(32'hbb2c6cd3),
	.w7(32'h38da2dfc),
	.w8(32'hbb5e4459),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c7f08),
	.w1(32'hbbb83186),
	.w2(32'hbc017fba),
	.w3(32'hbb9dba9a),
	.w4(32'hbb50522d),
	.w5(32'hbc06f2c4),
	.w6(32'hbbfd2bb3),
	.w7(32'hbb41240a),
	.w8(32'hbc4f3ae0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0cf3c),
	.w1(32'h3c50822c),
	.w2(32'h3afaa0aa),
	.w3(32'hba278d31),
	.w4(32'h3b127f4a),
	.w5(32'h3b02632d),
	.w6(32'h3c835571),
	.w7(32'h3c23a30d),
	.w8(32'h3b27dacb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89f1d0),
	.w1(32'h3b3886c7),
	.w2(32'hbb136868),
	.w3(32'h3b163671),
	.w4(32'h3b97bda9),
	.w5(32'h3b45cff4),
	.w6(32'h3ba3d4bc),
	.w7(32'hbb183719),
	.w8(32'hbc199f9c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a670039),
	.w1(32'h3b7c7bee),
	.w2(32'h3c9ed8ce),
	.w3(32'h3a9588f7),
	.w4(32'h3b0fb9d7),
	.w5(32'hbb746602),
	.w6(32'h3c65b2fe),
	.w7(32'hbb8a61ac),
	.w8(32'hbb451b75),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e8b2f),
	.w1(32'hbbf7021e),
	.w2(32'h3b666b62),
	.w3(32'hbb93ec5f),
	.w4(32'h3b2f1d27),
	.w5(32'h3a20f747),
	.w6(32'hba21df55),
	.w7(32'h3bc52ccb),
	.w8(32'hbb27c321),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3fc04),
	.w1(32'hbbc0a25a),
	.w2(32'hbbf759f5),
	.w3(32'hba4922ae),
	.w4(32'hbb3dda4b),
	.w5(32'hbc27548a),
	.w6(32'hbb57b8a2),
	.w7(32'hbbb0b40b),
	.w8(32'hbbe36e2c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb903ebe0),
	.w1(32'hbbec8c04),
	.w2(32'hbbab0974),
	.w3(32'hbc3866e9),
	.w4(32'hbbbe3af1),
	.w5(32'hbb60b0cb),
	.w6(32'hbc4afa1e),
	.w7(32'hbc3f7e8b),
	.w8(32'hbbbbc93b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b2d1d),
	.w1(32'hbb08da7e),
	.w2(32'h3a55025f),
	.w3(32'h39dac550),
	.w4(32'hba01fcb9),
	.w5(32'hbab51e6a),
	.w6(32'hbb0ee7c9),
	.w7(32'hbade95f3),
	.w8(32'hbb297516),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0af83),
	.w1(32'hbc1f6a0d),
	.w2(32'hbb876e2f),
	.w3(32'hbc1e240b),
	.w4(32'h3b34a4ca),
	.w5(32'hbc175814),
	.w6(32'hbbe5cf66),
	.w7(32'h3991524e),
	.w8(32'hbc6183fb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae12fbf),
	.w1(32'hbbb2b3be),
	.w2(32'h3b7bd30c),
	.w3(32'hbc1547da),
	.w4(32'h3b77761e),
	.w5(32'hbbc9f779),
	.w6(32'h3aa6bd55),
	.w7(32'h3c00a9a1),
	.w8(32'hbb679de1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24f248),
	.w1(32'h3ac84b07),
	.w2(32'hbc308aa7),
	.w3(32'hbbd03d4e),
	.w4(32'hbbd55111),
	.w5(32'hbbf8256a),
	.w6(32'hbbd09ff5),
	.w7(32'h3a8368dd),
	.w8(32'hbbba4615),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90a4b2),
	.w1(32'h3babec1c),
	.w2(32'hbbfc752d),
	.w3(32'h3a2c7643),
	.w4(32'hbbe1262c),
	.w5(32'hbc00306f),
	.w6(32'h3af557ce),
	.w7(32'hbbb9ef48),
	.w8(32'hbc3133d9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1afc65),
	.w1(32'h3b66c32f),
	.w2(32'hbb939726),
	.w3(32'h3ab14f09),
	.w4(32'h3a94b65c),
	.w5(32'hba64c17a),
	.w6(32'h3bde8ce2),
	.w7(32'hbb87e81e),
	.w8(32'hbb00e129),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85dc36),
	.w1(32'h39572c31),
	.w2(32'hbb87f979),
	.w3(32'h3a9c9ff0),
	.w4(32'h3baa8bf0),
	.w5(32'h3b456f76),
	.w6(32'hbb6f2ebc),
	.w7(32'h3b677229),
	.w8(32'h3ac95750),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f10891),
	.w1(32'hbc89991d),
	.w2(32'hbc92f4f4),
	.w3(32'hbc782c79),
	.w4(32'h3afdd481),
	.w5(32'hbb8fe545),
	.w6(32'hbc971383),
	.w7(32'hbc39434b),
	.w8(32'hbbd49876),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a21fd),
	.w1(32'hb9361b2b),
	.w2(32'h3b0363f0),
	.w3(32'hbadbb0a9),
	.w4(32'hba9c88e5),
	.w5(32'h3b6251fa),
	.w6(32'hbb77590b),
	.w7(32'hbade9df6),
	.w8(32'h3b5732bc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e52ea),
	.w1(32'h3ba5287d),
	.w2(32'h3aa05101),
	.w3(32'h3a2cbd0f),
	.w4(32'hb7bbdd46),
	.w5(32'hbca1804d),
	.w6(32'h3b6c4c9d),
	.w7(32'h3bf0ba66),
	.w8(32'hbc167465),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b1052),
	.w1(32'hbc0e7aef),
	.w2(32'hbb690a79),
	.w3(32'hbc0c8ae8),
	.w4(32'hbb601975),
	.w5(32'h3b73cb71),
	.w6(32'hbba9a578),
	.w7(32'hb899fcbf),
	.w8(32'hbbcd8d91),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea942b),
	.w1(32'h3bc83873),
	.w2(32'h3b81de6d),
	.w3(32'h3af743f4),
	.w4(32'hb873b494),
	.w5(32'h3bb36ac1),
	.w6(32'h3c961f14),
	.w7(32'h3b640eab),
	.w8(32'h3c427c7c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9963b6),
	.w1(32'hbc72f447),
	.w2(32'hbc2673ba),
	.w3(32'hbc98b2cf),
	.w4(32'h3b3e2b9a),
	.w5(32'h3b35de3e),
	.w6(32'hbca0e61c),
	.w7(32'hbc088a78),
	.w8(32'hbb86f301),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2bafc),
	.w1(32'h39222814),
	.w2(32'h38c63bdf),
	.w3(32'h3a6858a3),
	.w4(32'h3bfffac8),
	.w5(32'hbb8a1270),
	.w6(32'hbbcaa1d3),
	.w7(32'h3b338c98),
	.w8(32'hbc025e95),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaadcd5),
	.w1(32'hbbd08f8a),
	.w2(32'hbc8366ca),
	.w3(32'hbc8056ee),
	.w4(32'h3ba0c0af),
	.w5(32'hbcba9f81),
	.w6(32'hbc66d09e),
	.w7(32'hb9c80410),
	.w8(32'hbcf8ffd0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28a9b6),
	.w1(32'hbc85084d),
	.w2(32'h3b1a9784),
	.w3(32'hbcd2f4e6),
	.w4(32'h3bec694b),
	.w5(32'hbc39b6ab),
	.w6(32'hbceeae1c),
	.w7(32'hba1c07af),
	.w8(32'hbcd55cc9),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc2b5f),
	.w1(32'hbb50a7fc),
	.w2(32'hbb737389),
	.w3(32'hbc7a0e32),
	.w4(32'h3b854730),
	.w5(32'h3c221cce),
	.w6(32'hbca80fd0),
	.w7(32'hba9af1b7),
	.w8(32'h3bc35b76),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c196cfd),
	.w1(32'h3b8ea3f8),
	.w2(32'hbbd59ed3),
	.w3(32'h3b71614b),
	.w4(32'hbb85ceb7),
	.w5(32'h3b27210b),
	.w6(32'h3981528f),
	.w7(32'hbc1a4182),
	.w8(32'h3adaaf5c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3986ba),
	.w1(32'hb9e45e99),
	.w2(32'hbbd3f407),
	.w3(32'h3ba2f8f7),
	.w4(32'h39d7981b),
	.w5(32'hbb01a486),
	.w6(32'h3b7fe4fd),
	.w7(32'hbb98ed33),
	.w8(32'hbb83a8ad),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbababf4e),
	.w1(32'hbb2315c8),
	.w2(32'hba6eb09e),
	.w3(32'hbb3cc5c9),
	.w4(32'h3a8edfc4),
	.w5(32'h3c51a3c2),
	.w6(32'hbb3b8205),
	.w7(32'hbb1c931d),
	.w8(32'h3bd8f90a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8944a9),
	.w1(32'h3b9db5a9),
	.w2(32'h3bd21854),
	.w3(32'h3b606368),
	.w4(32'h3ba4fedd),
	.w5(32'h3c7b71c8),
	.w6(32'h3c7be041),
	.w7(32'h3c13d346),
	.w8(32'h3c8ec5f4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bdc65),
	.w1(32'h3d07eedb),
	.w2(32'h3c813fd1),
	.w3(32'h3cd5853c),
	.w4(32'h3ca7a3e9),
	.w5(32'hbb6ac430),
	.w6(32'h3cd9da21),
	.w7(32'h3c4f99c3),
	.w8(32'hbc13f88a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe19862),
	.w1(32'hbbfd4566),
	.w2(32'hbc1d9295),
	.w3(32'h3b8db296),
	.w4(32'hbaa1a547),
	.w5(32'hbc17e7c7),
	.w6(32'h3bfd2261),
	.w7(32'hbb4d8bbd),
	.w8(32'h3aadf95a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0721c5),
	.w1(32'h3bc984b7),
	.w2(32'h3bab685a),
	.w3(32'hbc2df619),
	.w4(32'hbc01dca9),
	.w5(32'hbbbae9e5),
	.w6(32'h3a21f7b0),
	.w7(32'h3a866a2b),
	.w8(32'h3c3d49da),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2cc3f),
	.w1(32'hbc32d541),
	.w2(32'hbc5b90d6),
	.w3(32'h3bdb9096),
	.w4(32'h3af62396),
	.w5(32'h39d91ce0),
	.w6(32'h3b18c2de),
	.w7(32'hbb2d408a),
	.w8(32'hbb7476b9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05ec65),
	.w1(32'h3aeb7903),
	.w2(32'hbacd86ae),
	.w3(32'hbab16427),
	.w4(32'h3ba4ff6e),
	.w5(32'hbb91d465),
	.w6(32'hbba66d34),
	.w7(32'h3c4a4581),
	.w8(32'hbc219c11),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a6768),
	.w1(32'h3ada9da9),
	.w2(32'h3c3e44ea),
	.w3(32'hbb83a1dd),
	.w4(32'hba204bce),
	.w5(32'hb87d7d15),
	.w6(32'h3bd643c2),
	.w7(32'h3c094388),
	.w8(32'hbab86185),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a1894),
	.w1(32'hbbf7c90c),
	.w2(32'hb9da0d1b),
	.w3(32'hbc42ccb2),
	.w4(32'hbabb4def),
	.w5(32'h384139cc),
	.w6(32'hbc86d671),
	.w7(32'hbafb51ad),
	.w8(32'hbb8da0b3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fdfd7),
	.w1(32'h3bb393ea),
	.w2(32'hbc976c04),
	.w3(32'hbb044b20),
	.w4(32'h3b85947f),
	.w5(32'hb9f2ae47),
	.w6(32'h3c01a8ae),
	.w7(32'h3ca00e22),
	.w8(32'hba789d35),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a1c86),
	.w1(32'h3b8d221a),
	.w2(32'hbbe826ff),
	.w3(32'hbc10d028),
	.w4(32'h3c53afd3),
	.w5(32'h3c68fbb3),
	.w6(32'hbc3bb84e),
	.w7(32'h3bc84efd),
	.w8(32'hbb5dd4e4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d4c36),
	.w1(32'h3b75d1cd),
	.w2(32'h3b93b243),
	.w3(32'hbb9fcb8b),
	.w4(32'hbb3e37f6),
	.w5(32'h3bd180d2),
	.w6(32'h39af6776),
	.w7(32'h3c7e352d),
	.w8(32'hbb463df1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a913cf9),
	.w1(32'hba243b21),
	.w2(32'h3bd82784),
	.w3(32'h3b1fbc90),
	.w4(32'h3c80f5c1),
	.w5(32'h3acde233),
	.w6(32'hbc04c134),
	.w7(32'h3bcdfd5b),
	.w8(32'hbb85761a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e79b3),
	.w1(32'h3ba6b521),
	.w2(32'h3b4261b4),
	.w3(32'h3b7d4b78),
	.w4(32'h3b0bc5ae),
	.w5(32'h3c0857d1),
	.w6(32'h3bd2c18d),
	.w7(32'h3bd81904),
	.w8(32'h3bc0b7fa),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c021b50),
	.w1(32'h3a89be1d),
	.w2(32'hbb197996),
	.w3(32'h394de8d6),
	.w4(32'hbb1e9404),
	.w5(32'h3adf9eb4),
	.w6(32'hbb610595),
	.w7(32'hbbd9280f),
	.w8(32'h3b910704),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ad3c4),
	.w1(32'h39904335),
	.w2(32'hbb037e57),
	.w3(32'hba3b1211),
	.w4(32'h3c0847af),
	.w5(32'hbba06356),
	.w6(32'h3c0d4485),
	.w7(32'h3c177fa0),
	.w8(32'hbb4e4a02),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18ffe2),
	.w1(32'h3ad8bb96),
	.w2(32'hbc71c5a3),
	.w3(32'hbb8fa836),
	.w4(32'hbb9cb615),
	.w5(32'hbc3cbd80),
	.w6(32'h3c45d24a),
	.w7(32'hbc1839ad),
	.w8(32'hbc85b0d3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2621ce),
	.w1(32'h39085aae),
	.w2(32'hbc32b380),
	.w3(32'hbc2c742b),
	.w4(32'h3ba92097),
	.w5(32'hba1c40cf),
	.w6(32'hbc025355),
	.w7(32'hbaa9dede),
	.w8(32'hbc178f2c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed401e),
	.w1(32'h3b3cdb7d),
	.w2(32'hbbc2d782),
	.w3(32'hbbda2e55),
	.w4(32'h3b8244f0),
	.w5(32'hbbd28455),
	.w6(32'hbc5b9ae9),
	.w7(32'hbb8863fd),
	.w8(32'hbc32a265),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f1958),
	.w1(32'hb99ae574),
	.w2(32'hbc27ace2),
	.w3(32'hbc3167e0),
	.w4(32'hbb6e2649),
	.w5(32'h3a64bfe4),
	.w6(32'hbc224320),
	.w7(32'hbc09643a),
	.w8(32'hbc2f1b68),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83d730),
	.w1(32'hbbecd99b),
	.w2(32'hbb9cdc46),
	.w3(32'hbc0967bd),
	.w4(32'hbc84bb18),
	.w5(32'hbc898b6b),
	.w6(32'hbc895b4f),
	.w7(32'hbc84601e),
	.w8(32'hbc7dd03c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba63c6b),
	.w1(32'hbb071d07),
	.w2(32'hbc388ae9),
	.w3(32'h3adb30a4),
	.w4(32'hbbec493f),
	.w5(32'h3b815beb),
	.w6(32'h3aafc11c),
	.w7(32'hbb87e980),
	.w8(32'hbb69023d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9864b1),
	.w1(32'hbba8c004),
	.w2(32'hbb178107),
	.w3(32'h3aba6671),
	.w4(32'h3b5d2947),
	.w5(32'hbaf1cc79),
	.w6(32'hbc08fc95),
	.w7(32'hba95c87c),
	.w8(32'hbc105e3c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb460b6),
	.w1(32'hbc2c7d8f),
	.w2(32'h3a169e4f),
	.w3(32'hbb6cd653),
	.w4(32'h3b7772c6),
	.w5(32'hba5f1bce),
	.w6(32'hbb913243),
	.w7(32'hba215e3d),
	.w8(32'hbac97eee),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc507b4c),
	.w1(32'h39fb575e),
	.w2(32'hbafbe8ff),
	.w3(32'hbc0bae8e),
	.w4(32'hbb502bc5),
	.w5(32'hbc20dd7d),
	.w6(32'h3a9f8590),
	.w7(32'hbb2eb7bd),
	.w8(32'hbc24edfb),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977b144),
	.w1(32'hbbbb8852),
	.w2(32'h3b51294b),
	.w3(32'hbc1afeee),
	.w4(32'h3b5b34bc),
	.w5(32'hbb8613a9),
	.w6(32'hbb4b6f52),
	.w7(32'h3b752e14),
	.w8(32'hbc03bc57),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab73185),
	.w1(32'hbb401c40),
	.w2(32'hbbc8cf72),
	.w3(32'h3a7299e5),
	.w4(32'h3ad400b4),
	.w5(32'hbc1b5582),
	.w6(32'hbc45a87c),
	.w7(32'hbaffe7fa),
	.w8(32'hbca91eac),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c48c6),
	.w1(32'hbaedb054),
	.w2(32'hbba788ae),
	.w3(32'hbb9fa512),
	.w4(32'hbc1c72b5),
	.w5(32'hbb5fa4a2),
	.w6(32'hb873d830),
	.w7(32'hbc219aaf),
	.w8(32'hbbb05334),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba571479),
	.w1(32'h385d77c8),
	.w2(32'h3bc5f419),
	.w3(32'hbbd67c82),
	.w4(32'hbb04f4a9),
	.w5(32'h3afc8700),
	.w6(32'h3c0ae362),
	.w7(32'hbacef2a0),
	.w8(32'hbae68bd3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4de713),
	.w1(32'h3c05660d),
	.w2(32'h3ada6b8c),
	.w3(32'h3b70dabe),
	.w4(32'hbb79cea7),
	.w5(32'hbb96200a),
	.w6(32'h3c10426e),
	.w7(32'hba7c787f),
	.w8(32'hbc0654d6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a009543),
	.w1(32'h3c375377),
	.w2(32'hba2a788d),
	.w3(32'h3c39384d),
	.w4(32'hbab751bc),
	.w5(32'h3c05d90b),
	.w6(32'h3ca47406),
	.w7(32'h3929ec75),
	.w8(32'h3b2ba134),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27fdce),
	.w1(32'h3b0b1a5e),
	.w2(32'h3aee3698),
	.w3(32'h3b88142c),
	.w4(32'h3b97c0c9),
	.w5(32'hbbb14d9d),
	.w6(32'hbbcc8ca8),
	.w7(32'hbb2ced69),
	.w8(32'hbc6091c2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc443964),
	.w1(32'h3b62e16f),
	.w2(32'hbae48399),
	.w3(32'h3b5795a6),
	.w4(32'hba980f76),
	.w5(32'h3c323b48),
	.w6(32'h3b624cf0),
	.w7(32'h3b2e74d2),
	.w8(32'h39f94da1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e406d),
	.w1(32'hbb9e7ebf),
	.w2(32'hbaab3d6e),
	.w3(32'h3c0b1c4c),
	.w4(32'hbb88f926),
	.w5(32'hba7861ae),
	.w6(32'h3c16484b),
	.w7(32'h3c4070d7),
	.w8(32'h3bb4183d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd37c),
	.w1(32'h3b2075b0),
	.w2(32'hb9eaae5f),
	.w3(32'hbb3ee5d2),
	.w4(32'h3a1e4c63),
	.w5(32'hbc59e523),
	.w6(32'h3a047b35),
	.w7(32'hbc0762d6),
	.w8(32'hbc66ce4a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8e78b),
	.w1(32'h3b451d3c),
	.w2(32'h3bca6015),
	.w3(32'hbbf58129),
	.w4(32'hbbb9460f),
	.w5(32'h3b8c2582),
	.w6(32'hba8051b0),
	.w7(32'hbb145ac4),
	.w8(32'hba0a71b9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a835808),
	.w1(32'h3c661aaf),
	.w2(32'h3c0e9474),
	.w3(32'h3c40c5b3),
	.w4(32'h3b7fa133),
	.w5(32'h3c046020),
	.w6(32'h3c97fd2c),
	.w7(32'h3bb23cdb),
	.w8(32'h3b97f867),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c30c3),
	.w1(32'h3c2f31b0),
	.w2(32'h3c83a1aa),
	.w3(32'h3becf0df),
	.w4(32'h3b0ebb13),
	.w5(32'hbc476770),
	.w6(32'h3cad0280),
	.w7(32'h3b652fed),
	.w8(32'hbc0c986a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1f8e7),
	.w1(32'hba880150),
	.w2(32'h3b0f2e6f),
	.w3(32'hbc0b6d00),
	.w4(32'hbbd705fe),
	.w5(32'hbc3b08bc),
	.w6(32'h3a411a6c),
	.w7(32'hbb1fc83f),
	.w8(32'hbc0fcc43),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840f47),
	.w1(32'h3a39b34e),
	.w2(32'hbbcc59c9),
	.w3(32'hbbb76f23),
	.w4(32'hbb679a41),
	.w5(32'hbba7dbe5),
	.w6(32'h383d256d),
	.w7(32'hbb04a40a),
	.w8(32'hbb7f491f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba552fd7),
	.w1(32'h3b7690b3),
	.w2(32'hbc59f3fa),
	.w3(32'h3bb61e6d),
	.w4(32'hbb85d9df),
	.w5(32'hbbcbcf01),
	.w6(32'h3b3dd240),
	.w7(32'hbc08a1d2),
	.w8(32'hbc604b12),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1497b),
	.w1(32'hbb37839a),
	.w2(32'hbc50e557),
	.w3(32'hbb05bfc4),
	.w4(32'h3b655ec6),
	.w5(32'hbbeaf513),
	.w6(32'h38ac2ccc),
	.w7(32'hbba0fd4f),
	.w8(32'hbbc902ff),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5717ce),
	.w1(32'h3bbc0ab1),
	.w2(32'hbbd97510),
	.w3(32'hbbff9c61),
	.w4(32'h3cab1014),
	.w5(32'h3b193b86),
	.w6(32'hbcd0506d),
	.w7(32'h3c445bae),
	.w8(32'hbc108850),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e760b4),
	.w1(32'hbaf76837),
	.w2(32'hbbd51334),
	.w3(32'h3b28b9b7),
	.w4(32'h3aa9a120),
	.w5(32'h3c3d2f23),
	.w6(32'h3b416a3a),
	.w7(32'hbb319890),
	.w8(32'h3b82c46c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c4f5a),
	.w1(32'hbc5dce4f),
	.w2(32'hbbd11622),
	.w3(32'hbc4bb498),
	.w4(32'hbc3a7179),
	.w5(32'hbb92dfaa),
	.w6(32'hbc843475),
	.w7(32'hbc473ccc),
	.w8(32'h3b129e3d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc008142),
	.w1(32'h3b97b0ee),
	.w2(32'h3c3af008),
	.w3(32'hbbebdfac),
	.w4(32'hbb80e68f),
	.w5(32'h3be7f4ea),
	.w6(32'hbb595e92),
	.w7(32'hbc3a7a14),
	.w8(32'h3aaf14c6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826d9e),
	.w1(32'h3b55d845),
	.w2(32'h39c98317),
	.w3(32'h3b890a90),
	.w4(32'hbb69d6b5),
	.w5(32'hbc5f7761),
	.w6(32'h3b5607bb),
	.w7(32'h3bff0e7c),
	.w8(32'hbc4dd458),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c517b),
	.w1(32'hbc05deca),
	.w2(32'h3b27bf9e),
	.w3(32'hbba3c4ae),
	.w4(32'h3bad7f8d),
	.w5(32'hbb95d2cc),
	.w6(32'h3a5135a1),
	.w7(32'h3c3cd848),
	.w8(32'hbba88112),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb19655),
	.w1(32'h3b53d8b3),
	.w2(32'h3ab99d0d),
	.w3(32'hbb70bf9c),
	.w4(32'hbb80ddc0),
	.w5(32'hbbb52136),
	.w6(32'h3b313b69),
	.w7(32'h3b55cb9f),
	.w8(32'hbc3f4fad),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc023f52),
	.w1(32'hbb344969),
	.w2(32'hbc28c4cc),
	.w3(32'hba264da2),
	.w4(32'h3b30703a),
	.w5(32'hbc3eb15f),
	.w6(32'h3ba3a4dc),
	.w7(32'h3a719192),
	.w8(32'hbbde2fb8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc529964),
	.w1(32'h3a7bc880),
	.w2(32'hbaddcc8e),
	.w3(32'hbc80134f),
	.w4(32'h39f6b89b),
	.w5(32'hbbcf65d4),
	.w6(32'hbc2777ea),
	.w7(32'hbb8a709e),
	.w8(32'hbbd29cf8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4338b7),
	.w1(32'hbbb5d402),
	.w2(32'hbbed8b30),
	.w3(32'hbbaf0211),
	.w4(32'hb985a2c1),
	.w5(32'hbb913cf2),
	.w6(32'hbbf0aa66),
	.w7(32'hbba9d28a),
	.w8(32'hbc0bdff6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b082fcf),
	.w1(32'hbb1b40d9),
	.w2(32'hbada9ed0),
	.w3(32'h3a03af21),
	.w4(32'hbb0949c0),
	.w5(32'h3bec201e),
	.w6(32'h3aa6c6dc),
	.w7(32'h3b2eca10),
	.w8(32'h3ac1f46a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacfb12),
	.w1(32'h3af65508),
	.w2(32'hb9f509b2),
	.w3(32'h3bec4ca3),
	.w4(32'h3c0d4c17),
	.w5(32'hbad10473),
	.w6(32'hbb29d54b),
	.w7(32'hba748d88),
	.w8(32'h3aba19f2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf053f8),
	.w1(32'hbb3fb9cf),
	.w2(32'hbb9237b2),
	.w3(32'hbc09dd6a),
	.w4(32'hbb4b99d4),
	.w5(32'hbbba37d2),
	.w6(32'hbb999b4e),
	.w7(32'h3b28b4e0),
	.w8(32'hbbb3a2a6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fa358),
	.w1(32'hb9d41d75),
	.w2(32'hbbe3ae3f),
	.w3(32'h3bc09e07),
	.w4(32'h3bd3aa8b),
	.w5(32'hbba3f8e2),
	.w6(32'h3c64a140),
	.w7(32'hbb3ed173),
	.w8(32'hbb788245),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfd7b4),
	.w1(32'h38ad0b62),
	.w2(32'h3c20dcb1),
	.w3(32'h3ba58692),
	.w4(32'h3c06e793),
	.w5(32'hbaa8dbf2),
	.w6(32'h3bd15499),
	.w7(32'h3b99b375),
	.w8(32'hbba17615),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50f697),
	.w1(32'hbb09f256),
	.w2(32'hbc0e21f5),
	.w3(32'h3a6aa48e),
	.w4(32'h3b2fc556),
	.w5(32'hbb849185),
	.w6(32'h3b58a896),
	.w7(32'hbb109c72),
	.w8(32'hbb54d705),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d4b4d),
	.w1(32'h3b5614a6),
	.w2(32'hbac2ab38),
	.w3(32'hb937857c),
	.w4(32'hbba18c57),
	.w5(32'hb9e92c1d),
	.w6(32'h3c6bb99c),
	.w7(32'hbbdad86e),
	.w8(32'hba7345ce),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf54971),
	.w1(32'h3b8539f4),
	.w2(32'hba94824f),
	.w3(32'hbbfbe272),
	.w4(32'hbaa5aeca),
	.w5(32'h3abd8674),
	.w6(32'hbc07a73c),
	.w7(32'hbc11a072),
	.w8(32'hbbb8874a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66af27),
	.w1(32'hb9db4718),
	.w2(32'h3b3f4615),
	.w3(32'hba5cefbe),
	.w4(32'h392d32ba),
	.w5(32'hbaf11299),
	.w6(32'h3c04f3d5),
	.w7(32'h3bc802d7),
	.w8(32'hbba56f92),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb690e0),
	.w1(32'hbbd1d334),
	.w2(32'hbb4a6146),
	.w3(32'hbb1f3e71),
	.w4(32'h3b97a283),
	.w5(32'h3c400b6c),
	.w6(32'hbc4481b0),
	.w7(32'h3a96ad34),
	.w8(32'h3c9e30b4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f945d),
	.w1(32'h3c050ce2),
	.w2(32'hbae5d729),
	.w3(32'h3c678e08),
	.w4(32'h3a550057),
	.w5(32'hbc74128b),
	.w6(32'h3b829bc9),
	.w7(32'hbbd0bf08),
	.w8(32'hbca37f10),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11c61d),
	.w1(32'h3b2f3307),
	.w2(32'h3c4b8d87),
	.w3(32'h3bc4eaf5),
	.w4(32'h3cb4245c),
	.w5(32'h3cf788f5),
	.w6(32'hbc50da0b),
	.w7(32'h3c823c8f),
	.w8(32'h3d395f5c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc723b),
	.w1(32'h3ca4685a),
	.w2(32'h3b3ee06f),
	.w3(32'h3cce702b),
	.w4(32'h3c58b703),
	.w5(32'hbbf5900f),
	.w6(32'h3ccbf4b4),
	.w7(32'hbad602b6),
	.w8(32'hbc3e6e03),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf787a6),
	.w1(32'h3c419d23),
	.w2(32'h3bce8577),
	.w3(32'hbba6bb9c),
	.w4(32'h3c0c6064),
	.w5(32'hbb8e280d),
	.w6(32'hba908771),
	.w7(32'h3b4aa236),
	.w8(32'hbbb3ce9a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec2e9d),
	.w1(32'h3c958625),
	.w2(32'hbc33165a),
	.w3(32'h3c8842a7),
	.w4(32'hbbb9ae79),
	.w5(32'h3b602b94),
	.w6(32'h3c87aa90),
	.w7(32'hbb8b19c1),
	.w8(32'h3b24718c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e42cf5),
	.w1(32'hbbd864eb),
	.w2(32'hbc0e3190),
	.w3(32'hbb214c5e),
	.w4(32'hbaf37a5b),
	.w5(32'hbb8bba2d),
	.w6(32'hbaea2a4a),
	.w7(32'hbb5e4ab9),
	.w8(32'h36e26dc2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4db077),
	.w1(32'hbc1f8fc3),
	.w2(32'hbc065459),
	.w3(32'hbc153186),
	.w4(32'hbb0e30a4),
	.w5(32'h3a328b7b),
	.w6(32'hbc2a71e2),
	.w7(32'hbb8d6608),
	.w8(32'hbbfc6f36),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91040a),
	.w1(32'hbb3a8e8e),
	.w2(32'h39ce5578),
	.w3(32'hbbe24ace),
	.w4(32'hbb4472ad),
	.w5(32'hba7808da),
	.w6(32'hbba831cf),
	.w7(32'hbacbe403),
	.w8(32'h3a028289),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb512426),
	.w1(32'hbb87e426),
	.w2(32'hbc3dd1b2),
	.w3(32'hb909b58c),
	.w4(32'h3b5f1991),
	.w5(32'hbbc1f994),
	.w6(32'hbbf06a01),
	.w7(32'hbc0516b1),
	.w8(32'hbc252c65),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e27d99),
	.w1(32'hbb1b7b7c),
	.w2(32'hbbc57366),
	.w3(32'hbbb07047),
	.w4(32'hbb3cb34e),
	.w5(32'hbbaa127b),
	.w6(32'hbbdaec70),
	.w7(32'hbb4e341f),
	.w8(32'hbbbf09ff),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc039a72),
	.w1(32'h3b22d833),
	.w2(32'hbbcc5457),
	.w3(32'hbaf99b8f),
	.w4(32'h3af555f4),
	.w5(32'hbb859034),
	.w6(32'hbbbbdcfc),
	.w7(32'h3b1c64a8),
	.w8(32'hbbd107eb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45f390),
	.w1(32'h3c08641d),
	.w2(32'hbac6fe62),
	.w3(32'hbbf988ea),
	.w4(32'h3c7884fd),
	.w5(32'h3bb06be9),
	.w6(32'hbc51b1ff),
	.w7(32'h3bff0c35),
	.w8(32'hbb080137),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefbff9),
	.w1(32'h3b0c324e),
	.w2(32'hbb8ff759),
	.w3(32'hbbef6ebe),
	.w4(32'h3b386828),
	.w5(32'hbb3d70f4),
	.w6(32'hbc2afeda),
	.w7(32'hbb2426b5),
	.w8(32'hbc0805ed),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b6e3f),
	.w1(32'hbb0d695c),
	.w2(32'hbc059e2c),
	.w3(32'hbb84b1cb),
	.w4(32'hba7f5c37),
	.w5(32'hbb9faf7b),
	.w6(32'hbaa107d7),
	.w7(32'h3ad1655a),
	.w8(32'hbbd4c956),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaaef77),
	.w1(32'h3a4554db),
	.w2(32'h3a596c01),
	.w3(32'h390b082c),
	.w4(32'h39c84271),
	.w5(32'hb762b199),
	.w6(32'h38beeea5),
	.w7(32'h3a3260ea),
	.w8(32'h399649d8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21e95f),
	.w1(32'hbbb49194),
	.w2(32'hbc192cd7),
	.w3(32'hbc07256b),
	.w4(32'hba62f9f3),
	.w5(32'hbae51a0e),
	.w6(32'hbb8c3c45),
	.w7(32'h3b2650a6),
	.w8(32'hbb085d80),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb924c798),
	.w1(32'h3a3d6103),
	.w2(32'hbbad2f0c),
	.w3(32'hba5ed466),
	.w4(32'hbae8d172),
	.w5(32'hbbfe03fe),
	.w6(32'hba3a1b88),
	.w7(32'hbac40570),
	.w8(32'hbbd846e0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e648d),
	.w1(32'hba36d7fc),
	.w2(32'hb8dd9c1f),
	.w3(32'hbaad56a7),
	.w4(32'hba4471c1),
	.w5(32'h380149d0),
	.w6(32'hb873d936),
	.w7(32'h3a20a1ef),
	.w8(32'h38c08e26),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb025d35),
	.w1(32'hba913a7d),
	.w2(32'hba24fdfa),
	.w3(32'hbaef999a),
	.w4(32'h39789fd9),
	.w5(32'h378c3af8),
	.w6(32'hbb3bf9dc),
	.w7(32'hba20a149),
	.w8(32'hba34b2d1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cbd5a),
	.w1(32'hba25fbf7),
	.w2(32'hbb869cbd),
	.w3(32'hbbafae2a),
	.w4(32'hbb97feb1),
	.w5(32'hbbddf285),
	.w6(32'hbbeb893b),
	.w7(32'hbbd710fb),
	.w8(32'hbc1762ba),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb409f10),
	.w1(32'h3b297146),
	.w2(32'hbb8582ad),
	.w3(32'hbb8c97eb),
	.w4(32'h3b0ce622),
	.w5(32'hbb1e254c),
	.w6(32'hbb86e7fd),
	.w7(32'hb9bb8f42),
	.w8(32'hbbc7fb3e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc626ca),
	.w1(32'hb781a45a),
	.w2(32'hbb65fb3c),
	.w3(32'hbbf164dd),
	.w4(32'hbae3eb7f),
	.w5(32'hbb199df9),
	.w6(32'hbc1e8ff5),
	.w7(32'hbb9ba17d),
	.w8(32'hbba887aa),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4841f),
	.w1(32'hb90da8ee),
	.w2(32'hb9e881db),
	.w3(32'hbb95916c),
	.w4(32'h3b2b1a5b),
	.w5(32'h3a813c8a),
	.w6(32'hbbb8cfc2),
	.w7(32'hb959255e),
	.w8(32'hbb5bec06),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2389d2),
	.w1(32'h3b470b44),
	.w2(32'hba5c1a24),
	.w3(32'hba917e5e),
	.w4(32'h3b54c848),
	.w5(32'h3a280f7b),
	.w6(32'hbb1e1b01),
	.w7(32'h3a652bb1),
	.w8(32'hbb0e00b3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49374e),
	.w1(32'hbb5d00f1),
	.w2(32'hbba979d8),
	.w3(32'hbac1309f),
	.w4(32'hba098bce),
	.w5(32'hba98c847),
	.w6(32'hb971e113),
	.w7(32'h3a83d7d1),
	.w8(32'hbb4074c3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89c2b1),
	.w1(32'h3abe91a7),
	.w2(32'hb9f43566),
	.w3(32'hba646365),
	.w4(32'h3b066df5),
	.w5(32'hbb0cbf86),
	.w6(32'hbb4bb75b),
	.w7(32'hb988ea9e),
	.w8(32'hbb8604f2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cd53ff),
	.w1(32'hb95a324c),
	.w2(32'h39974968),
	.w3(32'hbaa7db43),
	.w4(32'h39a6b17f),
	.w5(32'h3a8aad82),
	.w6(32'hba192ccf),
	.w7(32'hb9174f48),
	.w8(32'h3a4adc51),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec589c),
	.w1(32'hb928a286),
	.w2(32'hb9b16a1d),
	.w3(32'h39ec5d7d),
	.w4(32'h3a0bf38b),
	.w5(32'h3953d40b),
	.w6(32'hb8ff4bc0),
	.w7(32'h393ed49b),
	.w8(32'h398b47ec),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987698c),
	.w1(32'h3980bb8c),
	.w2(32'h3a621729),
	.w3(32'h3ab6999e),
	.w4(32'h3a2fa5b5),
	.w5(32'h39dec95a),
	.w6(32'h3a6990b2),
	.w7(32'h3ad66feb),
	.w8(32'h3a93d1ef),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa21c9a),
	.w1(32'hb901a731),
	.w2(32'h39570c51),
	.w3(32'h38736efd),
	.w4(32'hb9f0bcf2),
	.w5(32'hb985ed6a),
	.w6(32'h3a0d64a3),
	.w7(32'hb9811a12),
	.w8(32'h3a08fef5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc43c4),
	.w1(32'h3ae09cc5),
	.w2(32'hbb50ccf6),
	.w3(32'hb90578b1),
	.w4(32'h3b93aded),
	.w5(32'hb9a904a0),
	.w6(32'hbb261f37),
	.w7(32'h3b38a3bb),
	.w8(32'hbb258e3c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af7feb),
	.w1(32'hb96368f4),
	.w2(32'hba90e53a),
	.w3(32'hb98030a7),
	.w4(32'h3a227299),
	.w5(32'hb9fc03d8),
	.w6(32'hb98df493),
	.w7(32'hb98f0e26),
	.w8(32'hb93345e1),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a57bc9),
	.w1(32'hbb264e22),
	.w2(32'hbb582dd3),
	.w3(32'hbb6a602f),
	.w4(32'hbb7f07b7),
	.w5(32'hbb512af6),
	.w6(32'hbac3e878),
	.w7(32'hbb7baeb2),
	.w8(32'hbb4dc848),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fe385),
	.w1(32'hbaa6fdef),
	.w2(32'hbb538ef0),
	.w3(32'hbc2504bf),
	.w4(32'h39c17d82),
	.w5(32'hb9efc6e1),
	.w6(32'hbc1d0aa1),
	.w7(32'hb8b2a2a1),
	.w8(32'hbbacc537),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa112d4),
	.w1(32'h391e5009),
	.w2(32'h39733b30),
	.w3(32'h39c0b658),
	.w4(32'h3b287611),
	.w5(32'hba6d96f0),
	.w6(32'hba62ed42),
	.w7(32'h3a5503ed),
	.w8(32'h3a9d3a2a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c252a),
	.w1(32'h398d4231),
	.w2(32'h391697f6),
	.w3(32'hbb20a62f),
	.w4(32'hbac0904d),
	.w5(32'h3a0fc60a),
	.w6(32'hb666e2f7),
	.w7(32'hba2385b0),
	.w8(32'h3a190800),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef266d),
	.w1(32'h3af635db),
	.w2(32'h3aeb8efc),
	.w3(32'h3a05c429),
	.w4(32'hb91a34e4),
	.w5(32'h389cb77e),
	.w6(32'h3a147782),
	.w7(32'h3a14e9d1),
	.w8(32'h3a35126a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3829a971),
	.w1(32'h39e03d83),
	.w2(32'h3956a0a4),
	.w3(32'hbab2d3a4),
	.w4(32'hba4e0d0e),
	.w5(32'hb8dcc79f),
	.w6(32'hbb581adc),
	.w7(32'hbb1b42e0),
	.w8(32'hbaa0ba54),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b065b91),
	.w1(32'hbb8833ad),
	.w2(32'hbb937d2e),
	.w3(32'h3b5630dc),
	.w4(32'hbb0f65b5),
	.w5(32'hbbd7b753),
	.w6(32'h3b3ff601),
	.w7(32'hbb044fdb),
	.w8(32'hbbb51af9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba873dfd),
	.w1(32'hbb791c80),
	.w2(32'hbbd18582),
	.w3(32'hbaf7b5a0),
	.w4(32'hbb1e61f2),
	.w5(32'hbb8ce57c),
	.w6(32'hbb086f85),
	.w7(32'hbb9ca798),
	.w8(32'hbbde702a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384d7448),
	.w1(32'hba0bf014),
	.w2(32'hba5e3ea9),
	.w3(32'h3a01fe6a),
	.w4(32'h3a46e740),
	.w5(32'hb9c7adbd),
	.w6(32'h39b355b0),
	.w7(32'h399bd268),
	.w8(32'hba7933d5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb436a8e),
	.w1(32'hba02f51e),
	.w2(32'h391bcf82),
	.w3(32'hbb06135a),
	.w4(32'hb8e868c1),
	.w5(32'hba749005),
	.w6(32'hbb52dadf),
	.w7(32'hba3bfc55),
	.w8(32'hbace7e50),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd9031),
	.w1(32'h37e092fb),
	.w2(32'hba1269d1),
	.w3(32'hbb1efa88),
	.w4(32'hb83b9d18),
	.w5(32'hbad4111a),
	.w6(32'hbb59977d),
	.w7(32'hb9f240a8),
	.w8(32'hbadd5001),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7fff8),
	.w1(32'h39e6651c),
	.w2(32'hbb4f4add),
	.w3(32'hbaaa7f0f),
	.w4(32'hba1676cd),
	.w5(32'hba4d20f0),
	.w6(32'hbaafacdb),
	.w7(32'hba90fc0c),
	.w8(32'hbadb10a1),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6a549),
	.w1(32'hbb5a612e),
	.w2(32'hbb85ce68),
	.w3(32'hbbb1fc48),
	.w4(32'hba761af6),
	.w5(32'h395144f1),
	.w6(32'hbb796d63),
	.w7(32'hbadacf76),
	.w8(32'hbac30451),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade43cf),
	.w1(32'hbb820138),
	.w2(32'hbbfb7f23),
	.w3(32'hbb49dc98),
	.w4(32'hbb30777e),
	.w5(32'hbbf0240b),
	.w6(32'hbb998c01),
	.w7(32'hbbbd57a5),
	.w8(32'hbc1d6ec3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f19fd),
	.w1(32'h3a946a68),
	.w2(32'hb9c057d5),
	.w3(32'hbb3de2bd),
	.w4(32'h3b3e5518),
	.w5(32'h3a3b9ce8),
	.w6(32'hbb6d134d),
	.w7(32'h3a614a46),
	.w8(32'hbb3aa1bf),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb841647),
	.w1(32'hbb1ae631),
	.w2(32'hbb8e05b9),
	.w3(32'hbb370f73),
	.w4(32'h3b0068e1),
	.w5(32'h38e3a025),
	.w6(32'hbb637a05),
	.w7(32'h39e39c53),
	.w8(32'hbb6ad444),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6989c6),
	.w1(32'hbb51c9da),
	.w2(32'hbb966031),
	.w3(32'hbb96097d),
	.w4(32'hbade0965),
	.w5(32'hbba19371),
	.w6(32'hbac1cc00),
	.w7(32'hba98d106),
	.w8(32'hbb9dfc6c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb995bd8),
	.w1(32'h3a996d4a),
	.w2(32'h3a0e5c92),
	.w3(32'hbb539a15),
	.w4(32'h3b5a0f21),
	.w5(32'h3ac26c15),
	.w6(32'hbbb7fe82),
	.w7(32'h392f725c),
	.w8(32'hbb28856b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39854232),
	.w1(32'h39439790),
	.w2(32'hbb9c97f0),
	.w3(32'hb9975e30),
	.w4(32'h3a08a006),
	.w5(32'hbb27cfea),
	.w6(32'h38c7a43f),
	.w7(32'hb9c5e497),
	.w8(32'hbba44ca1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7eaa0c),
	.w1(32'hba514bba),
	.w2(32'hbae66f13),
	.w3(32'hba1fa422),
	.w4(32'hb9b2c1d7),
	.w5(32'hba703429),
	.w6(32'h3798bd38),
	.w7(32'h3984a9ce),
	.w8(32'hbb01f48a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7e81d),
	.w1(32'h3bcc0d69),
	.w2(32'h3a87048d),
	.w3(32'hbc13fe9a),
	.w4(32'h3b8e5d2d),
	.w5(32'hb94df83c),
	.w6(32'hbc3a2d64),
	.w7(32'h3a83663e),
	.w8(32'hbbb41b75),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1ff6e),
	.w1(32'hb9a802f2),
	.w2(32'hb902529b),
	.w3(32'hbb89495a),
	.w4(32'hb97b58a8),
	.w5(32'hb9ca1360),
	.w6(32'hbbb89894),
	.w7(32'hba99e16a),
	.w8(32'hbb6a6507),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb1754),
	.w1(32'h398df2ee),
	.w2(32'h392311af),
	.w3(32'hb9e44dd8),
	.w4(32'hba9f88e9),
	.w5(32'hb8c59a58),
	.w6(32'h3a3d7db3),
	.w7(32'hba38ddc3),
	.w8(32'h38480711),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39299890),
	.w1(32'h3903c99c),
	.w2(32'hb84f1189),
	.w3(32'h3942079b),
	.w4(32'h3a61e60f),
	.w5(32'h385b7f84),
	.w6(32'hb6d268f3),
	.w7(32'h39270b44),
	.w8(32'h37ab945f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00dfbe),
	.w1(32'hba0397d4),
	.w2(32'hbaa2ce6e),
	.w3(32'hbb0c7f6f),
	.w4(32'hb9a959de),
	.w5(32'hb98a2804),
	.w6(32'hbace6319),
	.w7(32'hb9979d6c),
	.w8(32'hba9636fd),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f73aa),
	.w1(32'hbad014d8),
	.w2(32'hbb32cfc0),
	.w3(32'hbbd45b37),
	.w4(32'h3b23a965),
	.w5(32'h3ab97830),
	.w6(32'hbbfb6c9d),
	.w7(32'h3a88db6e),
	.w8(32'hbb6833a5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ef4d8),
	.w1(32'h3b40082a),
	.w2(32'h393b6a31),
	.w3(32'hbc06d01f),
	.w4(32'hbab7e60b),
	.w5(32'hbad08b6a),
	.w6(32'hbbfe51c0),
	.w7(32'hbb540630),
	.w8(32'hbbd2f30e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba375bbc),
	.w1(32'h3b27fc4b),
	.w2(32'h3ad67747),
	.w3(32'h3b141e8c),
	.w4(32'h3a831181),
	.w5(32'h3a4d80f5),
	.w6(32'h3b0f3843),
	.w7(32'h3a5eb69d),
	.w8(32'h3a69370c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce404e),
	.w1(32'hba68db71),
	.w2(32'hbbb7f889),
	.w3(32'hbafae4fe),
	.w4(32'hba709ef3),
	.w5(32'hbb867ca5),
	.w6(32'hbb472ca6),
	.w7(32'hbb3289c2),
	.w8(32'hbbcc9644),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bce14),
	.w1(32'hb86c4634),
	.w2(32'hbaf41e61),
	.w3(32'hbb4aa615),
	.w4(32'hba898352),
	.w5(32'hba63d8f9),
	.w6(32'hbb85f10d),
	.w7(32'hbb404049),
	.w8(32'hbb99246c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb649961),
	.w1(32'hbb3839ad),
	.w2(32'hbbe3f4d5),
	.w3(32'hbb9ce55f),
	.w4(32'hbb86bade),
	.w5(32'hbbb79d54),
	.w6(32'hbb20b755),
	.w7(32'hbb7fcad2),
	.w8(32'hbb918061),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91790c),
	.w1(32'h3b677c0c),
	.w2(32'hbb6ba06c),
	.w3(32'hbbd51abb),
	.w4(32'h3b95e9dd),
	.w5(32'hbac020d9),
	.w6(32'hbc085094),
	.w7(32'hba8f8118),
	.w8(32'hbba69991),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43dfc5),
	.w1(32'h389fa85c),
	.w2(32'h3a151df2),
	.w3(32'hbb0c42a9),
	.w4(32'h3a9ee4a8),
	.w5(32'hb7cf6c6b),
	.w6(32'hbb797f92),
	.w7(32'h398e8a24),
	.w8(32'hbaa854a2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52730a),
	.w1(32'h3a6d0609),
	.w2(32'h3a246fd7),
	.w3(32'h39060c5e),
	.w4(32'hba6edb84),
	.w5(32'hba6a9cd7),
	.w6(32'hba8a5514),
	.w7(32'hb9e5d57a),
	.w8(32'h39b335d1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f439ef),
	.w1(32'h3b7e17cf),
	.w2(32'hbab5c36e),
	.w3(32'h3b12d8f8),
	.w4(32'h3bdf1060),
	.w5(32'h3adeb55b),
	.w6(32'h3a858437),
	.w7(32'h3b8ad5ed),
	.w8(32'hbaad149f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb984b),
	.w1(32'h3a7549ba),
	.w2(32'hb99939ff),
	.w3(32'hbb8d23c5),
	.w4(32'h3b91aaa8),
	.w5(32'h3951ea55),
	.w6(32'hbc0d9821),
	.w7(32'h38d3c862),
	.w8(32'hbb1036dc),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9abbd),
	.w1(32'h3afa7591),
	.w2(32'hb9871c7b),
	.w3(32'hbb1e94d7),
	.w4(32'h3b677f98),
	.w5(32'h39dfb350),
	.w6(32'hbb3e5b99),
	.w7(32'h3b1b9785),
	.w8(32'hba7ff4ae),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd27f9),
	.w1(32'hbaa63f59),
	.w2(32'hbb05fbc8),
	.w3(32'hba897c94),
	.w4(32'hbb023a6e),
	.w5(32'hbab42206),
	.w6(32'hbab566e6),
	.w7(32'hbb1abbba),
	.w8(32'hbad1d111),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba544e3f),
	.w1(32'hbac76b61),
	.w2(32'hbadbeee0),
	.w3(32'hba3c4c6a),
	.w4(32'hba9ad10e),
	.w5(32'hba8d10b9),
	.w6(32'hba0a0807),
	.w7(32'hba5dc83c),
	.w8(32'hba1dd295),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7abd31),
	.w1(32'hbb6b2a9c),
	.w2(32'hbb902e76),
	.w3(32'hbb41eaf8),
	.w4(32'hbb07d24f),
	.w5(32'hbb77e61a),
	.w6(32'hbb735367),
	.w7(32'hbb3d0109),
	.w8(32'hbba980d9),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987e775),
	.w1(32'hba8698e7),
	.w2(32'hba510e95),
	.w3(32'h3a1547ba),
	.w4(32'h3a4be0fb),
	.w5(32'h39b42185),
	.w6(32'h38b39c13),
	.w7(32'h39e99519),
	.w8(32'h3b0e3755),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d27c58),
	.w1(32'h3b9c675e),
	.w2(32'hba032c4d),
	.w3(32'h3a06903f),
	.w4(32'h3b78e38b),
	.w5(32'hb9ecb2cc),
	.w6(32'h3addb25a),
	.w7(32'h3b3ce7cb),
	.w8(32'hbb1475a5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918b6aa),
	.w1(32'h3a7d791c),
	.w2(32'hb978539a),
	.w3(32'h3a8f4140),
	.w4(32'h3a8c4eb9),
	.w5(32'hb86e7c12),
	.w6(32'h3928c66a),
	.w7(32'hb9d28fdb),
	.w8(32'h390c43ff),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e9cf8),
	.w1(32'hbb07b58e),
	.w2(32'hbbbcbcd1),
	.w3(32'hbb2d94e2),
	.w4(32'hbba0f46f),
	.w5(32'hbc04ddca),
	.w6(32'h3a83a17c),
	.w7(32'hbaeb1615),
	.w8(32'hbbb63a01),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77b62b),
	.w1(32'h3a5b7071),
	.w2(32'h3a932e4b),
	.w3(32'h36e978ae),
	.w4(32'hb9a94841),
	.w5(32'hba43ca06),
	.w6(32'h396e8949),
	.w7(32'h37061697),
	.w8(32'hba965d52),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17a701),
	.w1(32'h394afd20),
	.w2(32'hb9fb2256),
	.w3(32'h38fbb781),
	.w4(32'h3a66d1ee),
	.w5(32'h3a5ee7f7),
	.w6(32'hba947b65),
	.w7(32'hbaeeb0d1),
	.w8(32'h3a254631),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0082e),
	.w1(32'h3b0c1b62),
	.w2(32'hbb00f778),
	.w3(32'hbb0a42eb),
	.w4(32'h3b08f6a4),
	.w5(32'h3aad7431),
	.w6(32'hbb11bc45),
	.w7(32'hbaded18f),
	.w8(32'hbb19632a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45b35a),
	.w1(32'hbae7593b),
	.w2(32'hbc164498),
	.w3(32'hbb0001a5),
	.w4(32'h3ab2a1f4),
	.w5(32'hbc022e43),
	.w6(32'hbbb745f9),
	.w7(32'hbb4b1f92),
	.w8(32'hbc316e46),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf64ef),
	.w1(32'h3b69f0a8),
	.w2(32'h39f20bfd),
	.w3(32'h3ae3360b),
	.w4(32'h3b36fa53),
	.w5(32'hba57f7c3),
	.w6(32'h3976a578),
	.w7(32'h3a8cef12),
	.w8(32'hb9da371c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c6335),
	.w1(32'h3a429540),
	.w2(32'hbb4a5de2),
	.w3(32'hbb733b40),
	.w4(32'h3ac4492d),
	.w5(32'hbb396810),
	.w6(32'hbbb7f482),
	.w7(32'hbad35264),
	.w8(32'hbbe45de1),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1944ea),
	.w1(32'hba93d793),
	.w2(32'hba7c52d0),
	.w3(32'hbb6e0faf),
	.w4(32'hbae0ada6),
	.w5(32'hba37c088),
	.w6(32'hbb325fc2),
	.w7(32'hbb0a272a),
	.w8(32'h3a3f0cee),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba53b0),
	.w1(32'hbacb02b7),
	.w2(32'hbbb1d6ad),
	.w3(32'hbbc9e73e),
	.w4(32'h3a0dcf0e),
	.w5(32'hbba14412),
	.w6(32'hbbf94f05),
	.w7(32'hbb3a7a1f),
	.w8(32'hbc2bd465),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb965067),
	.w1(32'hba635c7d),
	.w2(32'hbbbd6935),
	.w3(32'hbb74f1e9),
	.w4(32'h3a9a01f5),
	.w5(32'hbb26abe1),
	.w6(32'hbb8b2fab),
	.w7(32'hba5713da),
	.w8(32'hbba3f4d7),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2de2d4),
	.w1(32'hbb537681),
	.w2(32'hbbc50958),
	.w3(32'hbb18c4b4),
	.w4(32'hba5cc6ad),
	.w5(32'hbb837a8d),
	.w6(32'hbad4baee),
	.w7(32'hbaa32447),
	.w8(32'hbbb18f24),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4e44d),
	.w1(32'h3a2a1199),
	.w2(32'h39465598),
	.w3(32'h3a2e2505),
	.w4(32'h39e802d8),
	.w5(32'hb9640d78),
	.w6(32'h3a4f7733),
	.w7(32'h3514af68),
	.w8(32'h393b5553),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55c301),
	.w1(32'hbb6396ab),
	.w2(32'hbabb9926),
	.w3(32'hbaec8cc7),
	.w4(32'hb9828897),
	.w5(32'h3a0ce0c7),
	.w6(32'hb9f47471),
	.w7(32'hb9c4cab0),
	.w8(32'hba3f34b2),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6603d),
	.w1(32'h399ab12f),
	.w2(32'h39bcb9a8),
	.w3(32'h35ffc550),
	.w4(32'hba258e42),
	.w5(32'hba24cf09),
	.w6(32'hb92f90a7),
	.w7(32'hb9c73328),
	.w8(32'hb7c6231e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8297287),
	.w1(32'hb9d54a6c),
	.w2(32'hbb13eb72),
	.w3(32'hba917528),
	.w4(32'hb975bd84),
	.w5(32'hba4e19b3),
	.w6(32'hba8ad205),
	.w7(32'hbb028c9c),
	.w8(32'hbb2cccf9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ccd25c),
	.w1(32'h3a2551dd),
	.w2(32'h3a7fbc7a),
	.w3(32'hb9888992),
	.w4(32'h3a58685c),
	.w5(32'hba2f3e98),
	.w6(32'hbafbffc6),
	.w7(32'h39bb8d72),
	.w8(32'hba09479b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b0acf),
	.w1(32'hbb226486),
	.w2(32'hbb916d1c),
	.w3(32'hbbc63a69),
	.w4(32'hbb117fcd),
	.w5(32'hbb0fd091),
	.w6(32'hbbf2dabe),
	.w7(32'hbb5f40e7),
	.w8(32'hbb9efc3b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985ac4a),
	.w1(32'h39a18a37),
	.w2(32'hba6dd749),
	.w3(32'hba2db916),
	.w4(32'hb9d7a471),
	.w5(32'h3a3b6d51),
	.w6(32'h3a113923),
	.w7(32'hb90cbcfd),
	.w8(32'h3aada285),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fc047),
	.w1(32'h3a642f9e),
	.w2(32'h3a865b49),
	.w3(32'h398e09fd),
	.w4(32'h3a226a72),
	.w5(32'h380599e4),
	.w6(32'h3ae55587),
	.w7(32'h3aa8f16d),
	.w8(32'h3a3202fb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b7019),
	.w1(32'h3aa12715),
	.w2(32'h38af2f1b),
	.w3(32'hba28d8a9),
	.w4(32'h3ac9de55),
	.w5(32'h3a8ddac8),
	.w6(32'hba2101c6),
	.w7(32'h3aa0205d),
	.w8(32'h39f7a289),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05e7e4),
	.w1(32'hbb1e9356),
	.w2(32'hbbeca91b),
	.w3(32'hba5912eb),
	.w4(32'hb824c1e2),
	.w5(32'hbb030f00),
	.w6(32'hbb1f8e96),
	.w7(32'hbad79745),
	.w8(32'hbb9edc08),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec91b8),
	.w1(32'h3b24beaf),
	.w2(32'hbaf568b9),
	.w3(32'hbac72868),
	.w4(32'h3ad5e396),
	.w5(32'hbac7e209),
	.w6(32'h3b1500d6),
	.w7(32'h3b8c9ea4),
	.w8(32'hba7772e2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5b957),
	.w1(32'h391c152f),
	.w2(32'h39693866),
	.w3(32'hb9b50408),
	.w4(32'hba5c8c8c),
	.w5(32'hb97762a5),
	.w6(32'hbab27c79),
	.w7(32'hba95b785),
	.w8(32'hba1784a6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b551ab7),
	.w1(32'h3b307bf9),
	.w2(32'hbc0a036f),
	.w3(32'hba9628b0),
	.w4(32'h3beb643e),
	.w5(32'hbb56557a),
	.w6(32'h3c0e9d5f),
	.w7(32'h3c34d208),
	.w8(32'hbb9b22ae),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1588e4),
	.w1(32'h39a110e7),
	.w2(32'hbbf936c9),
	.w3(32'hbc33885f),
	.w4(32'h3bd6b649),
	.w5(32'h39b9d1d4),
	.w6(32'hbc0410e7),
	.w7(32'h3b3ce186),
	.w8(32'hbb2134cc),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac779d1),
	.w1(32'h395ba288),
	.w2(32'hbab57f31),
	.w3(32'h392e62dd),
	.w4(32'hba94393d),
	.w5(32'hbb11bae2),
	.w6(32'h3a6f29e6),
	.w7(32'hb932b4dd),
	.w8(32'hba2b960a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77f2cf),
	.w1(32'h3a172a2f),
	.w2(32'h39bae8fd),
	.w3(32'hba89e3d8),
	.w4(32'hbad366fb),
	.w5(32'hb6d545b2),
	.w6(32'h3a39de67),
	.w7(32'h38edf1c4),
	.w8(32'h3a4695d0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993e94b),
	.w1(32'h3a104e32),
	.w2(32'hb94d87fc),
	.w3(32'hba1e8f35),
	.w4(32'h3982cf81),
	.w5(32'hb846587f),
	.w6(32'hba13ce45),
	.w7(32'hb9956817),
	.w8(32'h3a71c124),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf2516),
	.w1(32'h39835be3),
	.w2(32'h39bf2e85),
	.w3(32'hba03a457),
	.w4(32'h384293ac),
	.w5(32'h39a1dd40),
	.w6(32'h3aaf14c4),
	.w7(32'h3a0c937b),
	.w8(32'h3a23e203),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1531c),
	.w1(32'hba89a7fb),
	.w2(32'hbb6c4187),
	.w3(32'h3907bff1),
	.w4(32'hbb18fb8f),
	.w5(32'hbb850814),
	.w6(32'h3a546b3b),
	.w7(32'hb9fa7cc4),
	.w8(32'hbb8bdd45),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7808e),
	.w1(32'hbb9714a3),
	.w2(32'hbb34f505),
	.w3(32'hbba3475d),
	.w4(32'hba8ee884),
	.w5(32'hbb49ae4f),
	.w6(32'hbba259f7),
	.w7(32'hbb0427e3),
	.w8(32'hbbe1bf1a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5bd39),
	.w1(32'h39149d0d),
	.w2(32'hbb513d4a),
	.w3(32'hbbf955ae),
	.w4(32'h3ab84085),
	.w5(32'h399d3235),
	.w6(32'hbc08c665),
	.w7(32'hbab37069),
	.w8(32'hbb5daaa6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39293148),
	.w1(32'h3a2ceb66),
	.w2(32'hba3855f9),
	.w3(32'hbaa338c0),
	.w4(32'h39fef871),
	.w5(32'hb9729d69),
	.w6(32'hb983abf3),
	.w7(32'hb997d993),
	.w8(32'hba5f4fc3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15b8f3),
	.w1(32'hba0fd89c),
	.w2(32'hbbe615b7),
	.w3(32'hbb509ea4),
	.w4(32'hb996e732),
	.w5(32'hbbb4f742),
	.w6(32'hbbded26b),
	.w7(32'hbb82322d),
	.w8(32'hbc0fb832),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fef58),
	.w1(32'hba2b552e),
	.w2(32'hbb0047a0),
	.w3(32'hba566a92),
	.w4(32'hbb0463ea),
	.w5(32'hbb891f03),
	.w6(32'hbb053d43),
	.w7(32'hbb46aa02),
	.w8(32'hbb7a0b25),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9604d75),
	.w1(32'h399d2c54),
	.w2(32'hb91c39a6),
	.w3(32'h3960524e),
	.w4(32'h39fd769f),
	.w5(32'h39f38952),
	.w6(32'hb8ec309c),
	.w7(32'hba8900df),
	.w8(32'hbac2581a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb305bc6),
	.w1(32'hbb19a489),
	.w2(32'hbb0d4917),
	.w3(32'h39b4c994),
	.w4(32'h3a4a21ac),
	.w5(32'h3ab98889),
	.w6(32'hba36c94a),
	.w7(32'hba3308be),
	.w8(32'h3a87f928),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dac36d),
	.w1(32'hb99efcf9),
	.w2(32'h3951ff45),
	.w3(32'h3a67be4c),
	.w4(32'h3b00cfe6),
	.w5(32'h397e8870),
	.w6(32'h3a0be6f5),
	.w7(32'h3a490ce3),
	.w8(32'h3917d265),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb933999),
	.w1(32'hba6e07a4),
	.w2(32'hbba7810f),
	.w3(32'hbb94189a),
	.w4(32'hba93ac23),
	.w5(32'hbb54b4d6),
	.w6(32'hbb82f96e),
	.w7(32'hbb10b98e),
	.w8(32'hbbc3937b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc178b14),
	.w1(32'h39c0f35a),
	.w2(32'hbaca71f1),
	.w3(32'hbb946082),
	.w4(32'h3bc5ac32),
	.w5(32'h3b38dcda),
	.w6(32'hbc13f148),
	.w7(32'h3b708c2b),
	.w8(32'h39302e36),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bb6be),
	.w1(32'h3a9a9d10),
	.w2(32'hbb38e722),
	.w3(32'hbb27e926),
	.w4(32'h3b63e0b2),
	.w5(32'hba12868e),
	.w6(32'hbb8c54fd),
	.w7(32'hb9052db1),
	.w8(32'hbb90f020),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac85d3d),
	.w1(32'h3b2afaa8),
	.w2(32'h3a4ad636),
	.w3(32'h3a756cd0),
	.w4(32'h3a2d1a0a),
	.w5(32'hbad9633d),
	.w6(32'hb9f9c081),
	.w7(32'hba0e35a6),
	.w8(32'hbb197fa9),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d2c7f),
	.w1(32'hb6023822),
	.w2(32'hbb0f0c55),
	.w3(32'hbbb45ea1),
	.w4(32'h3b49d336),
	.w5(32'hb89aa3fc),
	.w6(32'hbbf59590),
	.w7(32'hba843995),
	.w8(32'hbbadbb0d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb268224),
	.w1(32'hba84aae1),
	.w2(32'hbb7cdacd),
	.w3(32'hbb74a6d2),
	.w4(32'hb903bcb0),
	.w5(32'hbb20b9b3),
	.w6(32'hbb81aeac),
	.w7(32'hbb217c7a),
	.w8(32'hbb6a3a33),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29fdbe),
	.w1(32'h37b67a49),
	.w2(32'hbbb7f954),
	.w3(32'hbc2bacc7),
	.w4(32'hbb9d38dc),
	.w5(32'hbbab5ca7),
	.w6(32'hbc1dabcf),
	.w7(32'hbb4e4966),
	.w8(32'hbc2b8d29),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ae21d),
	.w1(32'hba4e2459),
	.w2(32'hb9468a93),
	.w3(32'h3a673c5b),
	.w4(32'h3a696256),
	.w5(32'h384b6b35),
	.w6(32'h34ee9763),
	.w7(32'h3a32616e),
	.w8(32'hb9042170),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f60d6),
	.w1(32'h3968d629),
	.w2(32'h3a03b64e),
	.w3(32'hb998c446),
	.w4(32'h39e3544c),
	.w5(32'h39d77435),
	.w6(32'hb967872b),
	.w7(32'hb92c3d3a),
	.w8(32'h3acfb79a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84af1b),
	.w1(32'h3ada49f9),
	.w2(32'hbb985e20),
	.w3(32'h3969fb16),
	.w4(32'h3b137585),
	.w5(32'hbb8764b4),
	.w6(32'hbb396528),
	.w7(32'hba0fdc68),
	.w8(32'hbbee6179),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f10f3),
	.w1(32'hb796376a),
	.w2(32'hbc035899),
	.w3(32'hb9d48a66),
	.w4(32'h3b72c112),
	.w5(32'hbc03d499),
	.w6(32'hbb5447c0),
	.w7(32'hba603650),
	.w8(32'hbc40f5cb),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6d6ba),
	.w1(32'hba50402b),
	.w2(32'hbb393885),
	.w3(32'hbb9b1a5b),
	.w4(32'h3b2f90e9),
	.w5(32'h3a528108),
	.w6(32'hbbd23aad),
	.w7(32'hb9bdc912),
	.w8(32'hbb79d13d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad8280),
	.w1(32'hba6fe80e),
	.w2(32'hbaf33414),
	.w3(32'hbb439867),
	.w4(32'hbb91a6cc),
	.w5(32'hbb61d728),
	.w6(32'h3b4fc272),
	.w7(32'h3a4a014e),
	.w8(32'hbae2152d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b4037),
	.w1(32'h39e4612d),
	.w2(32'h3a27b978),
	.w3(32'h38f06756),
	.w4(32'hb8a5e39f),
	.w5(32'h38ad1821),
	.w6(32'hb94e172e),
	.w7(32'hb8294d33),
	.w8(32'h38f030d3),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b1420),
	.w1(32'hba5f685a),
	.w2(32'hb99d5d4d),
	.w3(32'h38f38feb),
	.w4(32'hb712e0ee),
	.w5(32'hb9d490a2),
	.w6(32'h394119ab),
	.w7(32'hb9528aca),
	.w8(32'h3a2fe753),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ef87c),
	.w1(32'h3aaf0517),
	.w2(32'hbbebd1ee),
	.w3(32'hba189e3b),
	.w4(32'hbb025c4e),
	.w5(32'hbc139f6f),
	.w6(32'hba947bca),
	.w7(32'h39ff7e5b),
	.w8(32'hbb9f3b59),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54a8da),
	.w1(32'hbb26fdbd),
	.w2(32'hbbf00b8d),
	.w3(32'hbbc73eb3),
	.w4(32'hbb6dccfb),
	.w5(32'hbbc4c35d),
	.w6(32'hba3b620b),
	.w7(32'hbb563d02),
	.w8(32'hbbd7e24a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba495ae),
	.w1(32'hbbb6eb58),
	.w2(32'hbbba4488),
	.w3(32'hbbac2aee),
	.w4(32'hbbca4191),
	.w5(32'hbb90ac51),
	.w6(32'hbbf3212c),
	.w7(32'hbb96dbd2),
	.w8(32'hbb949da4),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e37db),
	.w1(32'h3b986f00),
	.w2(32'h39735575),
	.w3(32'hbb385e02),
	.w4(32'h3b0fef02),
	.w5(32'h3ad9c6ba),
	.w6(32'hbbf6a1f4),
	.w7(32'hba1fd733),
	.w8(32'hba4d38fb),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc261b6),
	.w1(32'h3a073232),
	.w2(32'hbb9edff6),
	.w3(32'hbb99e66d),
	.w4(32'h3b88cd7e),
	.w5(32'hba0344bb),
	.w6(32'hbbb7ce29),
	.w7(32'h3ab506da),
	.w8(32'hbb509efb),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9e298),
	.w1(32'h391f2b7f),
	.w2(32'h398bf459),
	.w3(32'hba7f8690),
	.w4(32'hba6c80dd),
	.w5(32'h39652752),
	.w6(32'hba010e05),
	.w7(32'hba81a588),
	.w8(32'hb9658851),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38807faa),
	.w1(32'hba0056d3),
	.w2(32'h3978f42a),
	.w3(32'hb9f3587a),
	.w4(32'hbacb6831),
	.w5(32'hba67b2e4),
	.w6(32'hb9d3a173),
	.w7(32'hb904116b),
	.w8(32'hba46f2a2),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa16a1c),
	.w1(32'h39e63074),
	.w2(32'hba34ee13),
	.w3(32'h390c1a0b),
	.w4(32'hba3dbe14),
	.w5(32'hbb19f31f),
	.w6(32'hba350a6c),
	.w7(32'hbabf6b2c),
	.w8(32'hba8a78b9),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a206f),
	.w1(32'hba7960f1),
	.w2(32'hba5d6fd8),
	.w3(32'hb9cf769c),
	.w4(32'hba85bb9e),
	.w5(32'hbb1ad4a6),
	.w6(32'hba18882c),
	.w7(32'hba8e466b),
	.w8(32'hbb89a5a6),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb227f4e),
	.w1(32'hbb244181),
	.w2(32'hbbb0199b),
	.w3(32'h3a8ff5d9),
	.w4(32'hbb469a0e),
	.w5(32'hbbc0abf3),
	.w6(32'hbb03e2bb),
	.w7(32'hbbb3ff79),
	.w8(32'hbb9b6d26),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac6fbe),
	.w1(32'hbb888568),
	.w2(32'hbc0a4827),
	.w3(32'hbb78d9a0),
	.w4(32'hbb21c3fa),
	.w5(32'h3bbd08d5),
	.w6(32'hba47a0de),
	.w7(32'h3a70ea12),
	.w8(32'hbc29a233),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb27042),
	.w1(32'h3bdd2286),
	.w2(32'h3c16db3a),
	.w3(32'h3bfacd74),
	.w4(32'h3c520293),
	.w5(32'h370114b7),
	.w6(32'hbc08f58f),
	.w7(32'h3b4ffcea),
	.w8(32'hbb8fc2da),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7228c),
	.w1(32'hbbbdf229),
	.w2(32'hbb8744a1),
	.w3(32'h3a728b79),
	.w4(32'h3a7ee5e0),
	.w5(32'hb9b09938),
	.w6(32'h3b719d6f),
	.w7(32'hb94722f6),
	.w8(32'hbabfe121),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c3884),
	.w1(32'h39e608f0),
	.w2(32'hbb766e67),
	.w3(32'hbbb7df77),
	.w4(32'hbab30aba),
	.w5(32'hbc3ce21f),
	.w6(32'hbbc767a6),
	.w7(32'hbac61e77),
	.w8(32'hbc078875),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc002462),
	.w1(32'hbb9e5ef1),
	.w2(32'hbb4a71ae),
	.w3(32'hbb2444a1),
	.w4(32'h3adae2c6),
	.w5(32'h3a1a7641),
	.w6(32'h3add5f9e),
	.w7(32'h3b23cbdb),
	.w8(32'hbb2a18ba),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be292e8),
	.w1(32'h3b675344),
	.w2(32'h3c3962dd),
	.w3(32'hbbc7caac),
	.w4(32'hbb0c537a),
	.w5(32'hbb66acaf),
	.w6(32'h3b92ace4),
	.w7(32'h3c1f3815),
	.w8(32'h3a846a90),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f584c),
	.w1(32'hbb817a6f),
	.w2(32'hbba75ed7),
	.w3(32'hbab9ab80),
	.w4(32'hbb20bda6),
	.w5(32'hbb1c9491),
	.w6(32'hbb052107),
	.w7(32'h390558dc),
	.w8(32'hbc0b4194),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba053175),
	.w1(32'h3a3cea3a),
	.w2(32'hbb30a82c),
	.w3(32'h3abc7893),
	.w4(32'hba70708f),
	.w5(32'h3b043edb),
	.w6(32'hb94bbe4f),
	.w7(32'h39ee1633),
	.w8(32'h3887c592),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2220e),
	.w1(32'h3b3ccab6),
	.w2(32'hbb4f250d),
	.w3(32'h3b90d52c),
	.w4(32'h399e8a05),
	.w5(32'hbb9047ae),
	.w6(32'h3beae7ce),
	.w7(32'h3766ae32),
	.w8(32'hbbc6ced9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb994627),
	.w1(32'h3b2b44be),
	.w2(32'h37a31f35),
	.w3(32'h3bfa0680),
	.w4(32'h38f38235),
	.w5(32'hbac7056c),
	.w6(32'h39e558b5),
	.w7(32'hbadc2972),
	.w8(32'hb91b7803),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2c0af),
	.w1(32'hbbcac817),
	.w2(32'hbba94b1b),
	.w3(32'h3acd4d96),
	.w4(32'h3bd83478),
	.w5(32'hba2ad353),
	.w6(32'hbb326c3e),
	.w7(32'h3a8b4268),
	.w8(32'hba010290),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17a5a9),
	.w1(32'hb895d084),
	.w2(32'h38baca4d),
	.w3(32'hbc003789),
	.w4(32'hbbf937e6),
	.w5(32'hbb6748e9),
	.w6(32'hbc13b8fa),
	.w7(32'hbb04a88d),
	.w8(32'hbb030b94),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8bb94),
	.w1(32'hbc3bf49d),
	.w2(32'hbc6b77e6),
	.w3(32'hbb6faeb0),
	.w4(32'hbacaabb3),
	.w5(32'hbc14d077),
	.w6(32'hbba48450),
	.w7(32'hbbc68a53),
	.w8(32'hbc34517a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cab5e),
	.w1(32'hbb7b3120),
	.w2(32'hbc07406b),
	.w3(32'hbad9989e),
	.w4(32'hbb0db25f),
	.w5(32'hbb96c2fb),
	.w6(32'hbb196fd6),
	.w7(32'hbbd0c8b8),
	.w8(32'hbc105554),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba972ce8),
	.w1(32'hbb7986e4),
	.w2(32'hbb9458e9),
	.w3(32'hbbb233f5),
	.w4(32'hbb0fd406),
	.w5(32'hbc383ad1),
	.w6(32'hbbdbfa97),
	.w7(32'hbbaaaadb),
	.w8(32'hbb8b547d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac13237),
	.w1(32'h3ac86d33),
	.w2(32'hbb552a5f),
	.w3(32'hbbdb8284),
	.w4(32'h399b2a65),
	.w5(32'hbab4a0ca),
	.w6(32'hbbc41107),
	.w7(32'hbbbae069),
	.w8(32'h3a9698ae),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cc19a),
	.w1(32'hbbcecf8e),
	.w2(32'hbb6aa3ce),
	.w3(32'hbaf3e837),
	.w4(32'hba5385df),
	.w5(32'h3b604f89),
	.w6(32'hbaa37737),
	.w7(32'hbba1671b),
	.w8(32'h3b10d9b9),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fc5b2),
	.w1(32'hbb6dda57),
	.w2(32'hb9bc28cd),
	.w3(32'h3b899eff),
	.w4(32'h3b817723),
	.w5(32'h3b289e2a),
	.w6(32'h3a2f5bb0),
	.w7(32'h3b6a3b6a),
	.w8(32'hb8a8a038),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8df3b7),
	.w1(32'h3ad02b24),
	.w2(32'h3bfae8a9),
	.w3(32'h3aaccf9b),
	.w4(32'h38cf56fc),
	.w5(32'hba816e7c),
	.w6(32'h3ca8179f),
	.w7(32'h3bad9f69),
	.w8(32'h3b9060aa),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab98d2c),
	.w1(32'h3abdacd1),
	.w2(32'hba0198fd),
	.w3(32'hbb253dfd),
	.w4(32'h3b26791e),
	.w5(32'hbc38809c),
	.w6(32'h3a5664ad),
	.w7(32'h3aa50a21),
	.w8(32'hbc84aac8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f47fe),
	.w1(32'hbb34a713),
	.w2(32'hba2c88c5),
	.w3(32'hbb17feac),
	.w4(32'hbad55559),
	.w5(32'hbba61470),
	.w6(32'hbc0e5bc7),
	.w7(32'hbaf97dd4),
	.w8(32'hb88a9360),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba659b2),
	.w1(32'hbb30e677),
	.w2(32'hbbf0e038),
	.w3(32'hbb24f2d6),
	.w4(32'h3b072467),
	.w5(32'hbb9023b5),
	.w6(32'h3ad52c54),
	.w7(32'hb9907604),
	.w8(32'hbb7eef37),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb202972),
	.w1(32'hba868e13),
	.w2(32'h3a044f3f),
	.w3(32'h39eb36d5),
	.w4(32'hbbde39d7),
	.w5(32'h3a6d1ef7),
	.w6(32'hb9b51bb1),
	.w7(32'hba889d02),
	.w8(32'h3b801286),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc3877),
	.w1(32'hbb8e221f),
	.w2(32'hbb76adf2),
	.w3(32'h3bb86857),
	.w4(32'h3b67a2f3),
	.w5(32'hbb607335),
	.w6(32'h3b223290),
	.w7(32'hbb9b2993),
	.w8(32'hbbdcd5c4),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08471d),
	.w1(32'hbb542b02),
	.w2(32'hbb4e31a1),
	.w3(32'hbb6f08b0),
	.w4(32'hbb9eb7b2),
	.w5(32'hb6d8da5d),
	.w6(32'hbc0d0be1),
	.w7(32'hbb879fa2),
	.w8(32'h3bdca1e5),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63a40d),
	.w1(32'hb9908a98),
	.w2(32'hbb75204a),
	.w3(32'h3b2fc5ae),
	.w4(32'h3aa776f3),
	.w5(32'hbb275de9),
	.w6(32'h3b4f97d7),
	.w7(32'h3aaeb796),
	.w8(32'hbb594a4a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08d513),
	.w1(32'hbc5563f0),
	.w2(32'hbc0e0197),
	.w3(32'hbbff9afa),
	.w4(32'hbbb2ffe7),
	.w5(32'hbb7e4ee5),
	.w6(32'hbb6330c1),
	.w7(32'hbb5f2c5e),
	.w8(32'hbc0a28cd),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc170280),
	.w1(32'hbbdbf95d),
	.w2(32'hbbb387a7),
	.w3(32'h3b3b2182),
	.w4(32'h3b529ec7),
	.w5(32'h3b25f3f4),
	.w6(32'h3aee3943),
	.w7(32'hbad5e391),
	.w8(32'hba8219a0),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94d1af),
	.w1(32'hbb3a5e77),
	.w2(32'h3bc5f657),
	.w3(32'hb9a9045e),
	.w4(32'h3bee9413),
	.w5(32'hba277646),
	.w6(32'hbc3049aa),
	.w7(32'hb8bb0756),
	.w8(32'hbab93637),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule