module layer_10_featuremap_490(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1120a4),
	.w1(32'h3ba293e0),
	.w2(32'hbb1da876),
	.w3(32'hbb3325de),
	.w4(32'h3bcd7590),
	.w5(32'hba024008),
	.w6(32'h3b92ffc8),
	.w7(32'h3b49f381),
	.w8(32'h3b115245),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23bf2d),
	.w1(32'hbb86f36d),
	.w2(32'hb9a718a8),
	.w3(32'hbbab65e4),
	.w4(32'hbbf965ec),
	.w5(32'hbb5dce2a),
	.w6(32'hbb120357),
	.w7(32'hbb64be84),
	.w8(32'h3b601059),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa59f9b),
	.w1(32'hbb3e2e7b),
	.w2(32'hbc0439da),
	.w3(32'h3b01cc85),
	.w4(32'hbbe2ead9),
	.w5(32'hbc01945b),
	.w6(32'h3a9de433),
	.w7(32'hbbd4f239),
	.w8(32'hbc5a5dd6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b7653),
	.w1(32'h3c71ba1e),
	.w2(32'hbaf251c2),
	.w3(32'hbc38f109),
	.w4(32'h3acd6d57),
	.w5(32'h3b4ee117),
	.w6(32'hbc3526aa),
	.w7(32'h3bad8ba6),
	.w8(32'h3bc781cf),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b740772),
	.w1(32'h3a8f13cb),
	.w2(32'h3bceb0db),
	.w3(32'h3c0f1276),
	.w4(32'hba8ae1cb),
	.w5(32'hbbb3437d),
	.w6(32'h3c153b4c),
	.w7(32'hbad1a398),
	.w8(32'hbbb27244),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab47bc4),
	.w1(32'hbbdcc66c),
	.w2(32'hbbff9fca),
	.w3(32'hbbd0b288),
	.w4(32'hbbfac23f),
	.w5(32'hbc176fa2),
	.w6(32'hbbca2e2e),
	.w7(32'hbbe617da),
	.w8(32'h3c39acc5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e8d1c),
	.w1(32'h3b85e198),
	.w2(32'hbbe18bba),
	.w3(32'h3af37a18),
	.w4(32'hbb930537),
	.w5(32'hbb32220c),
	.w6(32'h3b05ff19),
	.w7(32'h3bcf879e),
	.w8(32'h3bdcf156),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a474b),
	.w1(32'h3b4265ad),
	.w2(32'h3a1c0cc0),
	.w3(32'h3aad0d0c),
	.w4(32'h3c1e8212),
	.w5(32'hbb4a06ee),
	.w6(32'h3c0c0478),
	.w7(32'h3b8517d9),
	.w8(32'h3b90b707),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f85655),
	.w1(32'hbadf1398),
	.w2(32'hbb90ebe6),
	.w3(32'hbb19d5cd),
	.w4(32'h37ada520),
	.w5(32'hbae5aec5),
	.w6(32'h3ab85a3a),
	.w7(32'hbb4c4c59),
	.w8(32'h3a40dbce),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac88ef4),
	.w1(32'h3ad10020),
	.w2(32'hb9d95674),
	.w3(32'h3af7b506),
	.w4(32'hbb7a9b70),
	.w5(32'h3b3cfdda),
	.w6(32'hbb2ab769),
	.w7(32'h3963c459),
	.w8(32'h3b93da54),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc60dc0),
	.w1(32'hbb99145d),
	.w2(32'hbb0cc832),
	.w3(32'h3b98e162),
	.w4(32'h3b9cb3d3),
	.w5(32'h3a5a3567),
	.w6(32'h3b439b2d),
	.w7(32'h3b043c04),
	.w8(32'h3b5eccb5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba322a8),
	.w1(32'hbc6005f2),
	.w2(32'hbb0fe5f0),
	.w3(32'hbaf0b656),
	.w4(32'hbb8d4f17),
	.w5(32'h3c51b4a7),
	.w6(32'h3b12ce64),
	.w7(32'h3ad39e16),
	.w8(32'h398832c6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07c870),
	.w1(32'hbb917dc0),
	.w2(32'h3a8af74d),
	.w3(32'h3c3d56f6),
	.w4(32'h3b39ab4c),
	.w5(32'h3cafebf8),
	.w6(32'hbbf3f858),
	.w7(32'h3bfbf8c3),
	.w8(32'h3bd06cf8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58324f),
	.w1(32'hbaeeb69c),
	.w2(32'hbbb8d394),
	.w3(32'h3c112f89),
	.w4(32'hbc015912),
	.w5(32'hbc3bb150),
	.w6(32'hbc16ec54),
	.w7(32'hbacdebaf),
	.w8(32'hbb071f0d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bfac6),
	.w1(32'hbb859cd3),
	.w2(32'hbac4992b),
	.w3(32'hbb3b8a29),
	.w4(32'h3a1b6437),
	.w5(32'hbc9ab70c),
	.w6(32'hb9f95ab3),
	.w7(32'h3b589ba3),
	.w8(32'hbb3626c9),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dcbf1),
	.w1(32'hbbddd9a6),
	.w2(32'h3bb1b7b0),
	.w3(32'hbc3741d1),
	.w4(32'hba3005e0),
	.w5(32'h3a027a4e),
	.w6(32'h3a0df9a9),
	.w7(32'h3b58aa67),
	.w8(32'hbb82e8fd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992680c),
	.w1(32'hba5ed175),
	.w2(32'h3b4e9362),
	.w3(32'hbaf2c2c2),
	.w4(32'hba6ee144),
	.w5(32'hbb19b409),
	.w6(32'h3a04050d),
	.w7(32'h3abf2fde),
	.w8(32'h3b5679b3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ece8c),
	.w1(32'h3c1c9e53),
	.w2(32'hbb6d9415),
	.w3(32'hbbc4f4f0),
	.w4(32'h3bcc4804),
	.w5(32'hbbcbea31),
	.w6(32'h3b80baef),
	.w7(32'hba6d9f8b),
	.w8(32'hba160eaf),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c9972),
	.w1(32'hbbb10164),
	.w2(32'h3b8a6f8e),
	.w3(32'hbc03dd48),
	.w4(32'hbadd9448),
	.w5(32'h3c093c52),
	.w6(32'h3ba577bb),
	.w7(32'h3a76ffab),
	.w8(32'h3b08267b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0657c6),
	.w1(32'hbb4a6561),
	.w2(32'hbbc4732e),
	.w3(32'h3b903eee),
	.w4(32'hbb5ac0e2),
	.w5(32'hbc833a41),
	.w6(32'hbb165db4),
	.w7(32'h3ad6ed3f),
	.w8(32'h3c08beaf),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99de74),
	.w1(32'hbbd3fa9f),
	.w2(32'h3aae33ac),
	.w3(32'hbc024d2f),
	.w4(32'h3befda23),
	.w5(32'h3c775e12),
	.w6(32'hb9cb0dda),
	.w7(32'h3b828811),
	.w8(32'hbb43efde),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badd01a),
	.w1(32'hbafbb596),
	.w2(32'hbbcb8ce3),
	.w3(32'h3b202dd0),
	.w4(32'hbabf376c),
	.w5(32'hbc26032e),
	.w6(32'hbc67b61b),
	.w7(32'hbc1bf0c5),
	.w8(32'hbc571b4f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4df63c),
	.w1(32'hbb00beb7),
	.w2(32'hbb53510e),
	.w3(32'hbc21630b),
	.w4(32'h39bf6390),
	.w5(32'hbc0b5b53),
	.w6(32'hbb3be98c),
	.w7(32'hba3e669f),
	.w8(32'h3b73e918),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c006c40),
	.w1(32'hbbb14371),
	.w2(32'h3a87f6d9),
	.w3(32'h3bdd9ca7),
	.w4(32'h3b2cd2bd),
	.w5(32'h3bf3d053),
	.w6(32'hba553fcc),
	.w7(32'hb61deff6),
	.w8(32'hbb6805ba),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab327e),
	.w1(32'hbb1b9a27),
	.w2(32'hbbf1c647),
	.w3(32'h3af1c2be),
	.w4(32'h3a821dec),
	.w5(32'hbc411f27),
	.w6(32'hbb331346),
	.w7(32'hbbf5f48c),
	.w8(32'hbc38b0d1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1026e3),
	.w1(32'h3b749046),
	.w2(32'h3b35424a),
	.w3(32'hbb3426f0),
	.w4(32'hb9d0f8b2),
	.w5(32'hbaa24c7b),
	.w6(32'hbb6f5b86),
	.w7(32'hbbae8d1e),
	.w8(32'h3a9e212c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c0bd2),
	.w1(32'h3b312f20),
	.w2(32'h3c0a5dc4),
	.w3(32'h3b5ef341),
	.w4(32'h3bdc6842),
	.w5(32'h3af777ae),
	.w6(32'h3c078670),
	.w7(32'h3893e071),
	.w8(32'hbbc8309a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8626f4),
	.w1(32'hbac7f22f),
	.w2(32'hbb8b48e1),
	.w3(32'hbb85f4a0),
	.w4(32'hba1e8468),
	.w5(32'h3acdf50f),
	.w6(32'h3bf4be2d),
	.w7(32'h3b260fc2),
	.w8(32'h3bc28151),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c81ae),
	.w1(32'h3bb74fb1),
	.w2(32'hbbacf2e0),
	.w3(32'h3ba2d247),
	.w4(32'hbb899536),
	.w5(32'h39fd1b95),
	.w6(32'h3c5ec07f),
	.w7(32'h3c0cdd89),
	.w8(32'h3c45caf5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5171e),
	.w1(32'hbb410608),
	.w2(32'h3b25d636),
	.w3(32'h3c163e78),
	.w4(32'h3bd2dbdc),
	.w5(32'h3b9222d6),
	.w6(32'h3a816468),
	.w7(32'h3b9b5b3f),
	.w8(32'hbb1646f1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddae69),
	.w1(32'h3aa8f93e),
	.w2(32'hbb93eaf4),
	.w3(32'h3ad67066),
	.w4(32'hbc0239ab),
	.w5(32'hbb7537e9),
	.w6(32'hbc3ab3d7),
	.w7(32'hbab2bdef),
	.w8(32'h39ee99ca),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac3b14),
	.w1(32'h3b60c830),
	.w2(32'hb911fc31),
	.w3(32'h3ac02384),
	.w4(32'hbba35e0a),
	.w5(32'hbc4c6007),
	.w6(32'h3bb6dbd2),
	.w7(32'hbbbb773b),
	.w8(32'hbc08e137),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ababb),
	.w1(32'hbaab7a9d),
	.w2(32'hbbb76ff8),
	.w3(32'hbc21924e),
	.w4(32'hbbc89bda),
	.w5(32'hbba8c4e1),
	.w6(32'hbb6122f2),
	.w7(32'h3a89006a),
	.w8(32'h38c7aba7),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b513a8e),
	.w1(32'h3bf7329f),
	.w2(32'hbb3bb3e4),
	.w3(32'h3a8c3cad),
	.w4(32'hbac03c72),
	.w5(32'hbc015c52),
	.w6(32'h3bcbf9bc),
	.w7(32'hbb2069c7),
	.w8(32'h3b4f13d4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab409d),
	.w1(32'h3ab1559b),
	.w2(32'hbbd68e17),
	.w3(32'hbb62f556),
	.w4(32'h3855b469),
	.w5(32'hbbfd7701),
	.w6(32'h3c314ff9),
	.w7(32'hbb610553),
	.w8(32'h3a0c2434),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48e995),
	.w1(32'h3b43297c),
	.w2(32'hbb89360c),
	.w3(32'hbaf1d4f6),
	.w4(32'hbbbab586),
	.w5(32'hbbaf4eac),
	.w6(32'h3ae49579),
	.w7(32'h39f3d565),
	.w8(32'h3a1d9b48),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb535f00),
	.w1(32'h3a17fa38),
	.w2(32'h3ad2e545),
	.w3(32'h3b2faee0),
	.w4(32'h3c348f00),
	.w5(32'h3bb8196e),
	.w6(32'h3c0f66c8),
	.w7(32'h3b913ecc),
	.w8(32'h3ba45a55),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba777136),
	.w1(32'hbb76302a),
	.w2(32'hba702554),
	.w3(32'h3af7fedd),
	.w4(32'hbb931785),
	.w5(32'hbb8fb185),
	.w6(32'h3b95b7d6),
	.w7(32'hbad59e11),
	.w8(32'hba77d283),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c406610),
	.w1(32'h3bfce853),
	.w2(32'hbbb4a067),
	.w3(32'h3b059099),
	.w4(32'hbb2b1da1),
	.w5(32'hbc368c5a),
	.w6(32'hbb78c8ba),
	.w7(32'hbc045151),
	.w8(32'hbba70c97),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe11ed0),
	.w1(32'h3b085903),
	.w2(32'hbb4ce2a9),
	.w3(32'hbc1bb6f6),
	.w4(32'hbc0ccaf8),
	.w5(32'hbba9e95f),
	.w6(32'hba665bd9),
	.w7(32'hbace20c2),
	.w8(32'h3b91adbc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bb075),
	.w1(32'h3c33f4c2),
	.w2(32'h3b844162),
	.w3(32'h3b163d2a),
	.w4(32'h3b27a380),
	.w5(32'h381cb5d6),
	.w6(32'h3c0c82e7),
	.w7(32'hbb814627),
	.w8(32'hbbbf427d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace34eb),
	.w1(32'hbbd170c9),
	.w2(32'h3ad7c279),
	.w3(32'hbba38b28),
	.w4(32'h3bb385db),
	.w5(32'h3bb0a498),
	.w6(32'hbbcdea1f),
	.w7(32'hba87e047),
	.w8(32'h3a764d91),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb242b49),
	.w1(32'h3bd935a2),
	.w2(32'h3b3af63f),
	.w3(32'hbbc47962),
	.w4(32'hbb0a5f35),
	.w5(32'hbb4262de),
	.w6(32'hbb5dcdfd),
	.w7(32'hb89d32c1),
	.w8(32'hbba67adc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbaf5a),
	.w1(32'h3c39601f),
	.w2(32'hbaf24474),
	.w3(32'hbc0f3a26),
	.w4(32'hbb257d0b),
	.w5(32'hbb769623),
	.w6(32'hbb55f6b7),
	.w7(32'hba161578),
	.w8(32'h3c1fdc33),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9f2a1),
	.w1(32'hbb533ad2),
	.w2(32'h3bd5b24b),
	.w3(32'h3b93088c),
	.w4(32'h3bcc0030),
	.w5(32'h3c1ef4bb),
	.w6(32'h3c300247),
	.w7(32'h3a464b54),
	.w8(32'h3ab472e4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee42f0),
	.w1(32'hbbb6da49),
	.w2(32'h3c6135b7),
	.w3(32'h3c10e4ca),
	.w4(32'hb90fcd41),
	.w5(32'h3a137c02),
	.w6(32'h3bfd755f),
	.w7(32'h3a26ced7),
	.w8(32'hbc09f050),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba1565),
	.w1(32'hbbb27141),
	.w2(32'h3b754773),
	.w3(32'hba20759e),
	.w4(32'h3ab76e6b),
	.w5(32'h3c5eb29c),
	.w6(32'h3b15848a),
	.w7(32'h3b655d65),
	.w8(32'hb9bddbc4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06a474),
	.w1(32'hbb9d9ea6),
	.w2(32'hbb9a74c2),
	.w3(32'h385ab579),
	.w4(32'hbbf34437),
	.w5(32'hbbbffb99),
	.w6(32'hbb5e2563),
	.w7(32'hbb30b2ed),
	.w8(32'hbae40409),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0fc8a),
	.w1(32'h3c023ce8),
	.w2(32'h3ae19eb5),
	.w3(32'hba2ff33f),
	.w4(32'h3a841d49),
	.w5(32'hbbb4fe6f),
	.w6(32'hba9e206a),
	.w7(32'hbbe53bbd),
	.w8(32'hbb91846e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5eafc0),
	.w1(32'h3bad834e),
	.w2(32'h3aca31cb),
	.w3(32'h39e50548),
	.w4(32'hbb80d683),
	.w5(32'hbb9683bf),
	.w6(32'h3a39037c),
	.w7(32'hba2d8dca),
	.w8(32'hb9fd0869),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac97c9),
	.w1(32'hbba6c082),
	.w2(32'hbae93aea),
	.w3(32'h39947b0e),
	.w4(32'hbc0e7b7c),
	.w5(32'h3c1cc428),
	.w6(32'h3bbbb40a),
	.w7(32'hbb52acfa),
	.w8(32'h3be0196b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c322742),
	.w1(32'hbc2333d4),
	.w2(32'hbbf14a4f),
	.w3(32'h3bd6efdc),
	.w4(32'hbb9742eb),
	.w5(32'hbc5a2ed9),
	.w6(32'hbb826590),
	.w7(32'hbb968a55),
	.w8(32'hbc0ffceb),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb124422),
	.w1(32'hbafb1229),
	.w2(32'hbc046170),
	.w3(32'hb7ea44cd),
	.w4(32'hbbee8a7f),
	.w5(32'hbc134c15),
	.w6(32'h3bc60dca),
	.w7(32'hbb5a1df8),
	.w8(32'h3b82af16),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad156b),
	.w1(32'hba7e98ad),
	.w2(32'h3b06121a),
	.w3(32'hbb7cfb59),
	.w4(32'h3af8e9c8),
	.w5(32'h3b7df74c),
	.w6(32'h39f14a7d),
	.w7(32'h3be540f2),
	.w8(32'h3b00bd7a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90d3ed),
	.w1(32'hbb3fa62b),
	.w2(32'hbbb5652a),
	.w3(32'h3a3349c3),
	.w4(32'hbb67b2fb),
	.w5(32'hbc1a6433),
	.w6(32'h3a79ec9e),
	.w7(32'hbb122409),
	.w8(32'h3a5337be),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3d336),
	.w1(32'hba09fa54),
	.w2(32'h3a023e84),
	.w3(32'hbbb193ea),
	.w4(32'hbbeffb25),
	.w5(32'hbc6de12e),
	.w6(32'h376786ba),
	.w7(32'hbade2354),
	.w8(32'hbbac3933),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0b58f),
	.w1(32'h3ad5cb79),
	.w2(32'h3bb1ec70),
	.w3(32'hbbe1085d),
	.w4(32'h3ac4b51c),
	.w5(32'h3c2c6eef),
	.w6(32'h3bfac13c),
	.w7(32'hba6abae8),
	.w8(32'h3b05e701),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa5af7),
	.w1(32'hba28a395),
	.w2(32'hba8cff34),
	.w3(32'h3ba0e5b6),
	.w4(32'h39497404),
	.w5(32'hbca307f4),
	.w6(32'hbb7614de),
	.w7(32'hbb3158c8),
	.w8(32'hbbdf88a5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eedd6),
	.w1(32'hbb52e71f),
	.w2(32'hbbc41471),
	.w3(32'hbb80ddd9),
	.w4(32'hbb573789),
	.w5(32'hbaeede41),
	.w6(32'hbbbb8f1c),
	.w7(32'hba533226),
	.w8(32'h3a4cbe3a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bbc39),
	.w1(32'h3b9bcc29),
	.w2(32'hba48d423),
	.w3(32'hbb7dc439),
	.w4(32'hbbb366c6),
	.w5(32'hbc46f8af),
	.w6(32'hb999db3f),
	.w7(32'hbaba5638),
	.w8(32'hbb40a1a3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1652a),
	.w1(32'h3bd7310a),
	.w2(32'h3c72b3eb),
	.w3(32'h3ba5378c),
	.w4(32'hbb5581d6),
	.w5(32'hbc8d8102),
	.w6(32'h3a620acd),
	.w7(32'hbc1e7b30),
	.w8(32'h3bb95bd7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad73412),
	.w1(32'h3b23b430),
	.w2(32'hbb7a9688),
	.w3(32'hbc1b87ef),
	.w4(32'h3aa22b28),
	.w5(32'hbc20d9a9),
	.w6(32'h3be7438b),
	.w7(32'hbb5a55fb),
	.w8(32'h3b1c344a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4e351),
	.w1(32'h3b92bd34),
	.w2(32'h3bc83724),
	.w3(32'hbba6875b),
	.w4(32'h3bdb9502),
	.w5(32'h3b1d7466),
	.w6(32'h3c02516f),
	.w7(32'hbac5ad65),
	.w8(32'hbc06c938),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3567b1),
	.w1(32'hbb19f5b0),
	.w2(32'h3c14132d),
	.w3(32'h3a1ff169),
	.w4(32'h3b114f53),
	.w5(32'h3c7076d3),
	.w6(32'hbb489c91),
	.w7(32'hb9f09dbf),
	.w8(32'h3b29cd31),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c093a37),
	.w1(32'hba9040f1),
	.w2(32'h3985bb3b),
	.w3(32'h3bf5912b),
	.w4(32'h3b8d4b0f),
	.w5(32'h3b9758de),
	.w6(32'hbb4cb3ef),
	.w7(32'h3b68edb6),
	.w8(32'h3a6a4e57),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba254b1),
	.w1(32'hbad9eb68),
	.w2(32'hbb88425c),
	.w3(32'h3b968542),
	.w4(32'hbb0f5f2b),
	.w5(32'hbbc02f6d),
	.w6(32'hbb0286a9),
	.w7(32'hbc477b0a),
	.w8(32'hbbed4bb1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45a87d),
	.w1(32'hbb9511f1),
	.w2(32'hbb46d407),
	.w3(32'hbc1b1418),
	.w4(32'hbbe2eba6),
	.w5(32'hb94a1f59),
	.w6(32'hbb837c15),
	.w7(32'hbbe63593),
	.w8(32'h3bd60aea),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b25c8),
	.w1(32'hbafdd9ac),
	.w2(32'h3baad247),
	.w3(32'h3bb784a5),
	.w4(32'h3c10e0db),
	.w5(32'hbb974cf0),
	.w6(32'hbb3bf22b),
	.w7(32'h3b27e522),
	.w8(32'hbb0c4315),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5087a4),
	.w1(32'h3ba56cf1),
	.w2(32'h3b6b16df),
	.w3(32'hbbb240b5),
	.w4(32'hbc0db7b9),
	.w5(32'h3a8e0310),
	.w6(32'h3c08b938),
	.w7(32'hbb12c27c),
	.w8(32'h3bfeb655),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f18ae),
	.w1(32'hb8cde216),
	.w2(32'hbb23fc09),
	.w3(32'h3bfa24fe),
	.w4(32'hbaa7f877),
	.w5(32'hbbce9a11),
	.w6(32'h3a0848a8),
	.w7(32'hbb936db2),
	.w8(32'h3aeecce4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f589e),
	.w1(32'h3a97d9d3),
	.w2(32'hbb154acf),
	.w3(32'h3b493dc3),
	.w4(32'h3b9c16ef),
	.w5(32'hbaa1a9e6),
	.w6(32'hbbdfe4e9),
	.w7(32'h3bf730a1),
	.w8(32'h3ba5d007),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb594410),
	.w1(32'h3b4f157b),
	.w2(32'hbc1de477),
	.w3(32'hbc255dab),
	.w4(32'h38c465ff),
	.w5(32'h3b4ce783),
	.w6(32'hbb76cd71),
	.w7(32'hbc5a9105),
	.w8(32'hbbcc3a61),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba984f3),
	.w1(32'hbaf8a783),
	.w2(32'hba75a807),
	.w3(32'h3a70abd8),
	.w4(32'hbb8129e6),
	.w5(32'h3c939c7d),
	.w6(32'h3b0bd358),
	.w7(32'h3b9e875a),
	.w8(32'h3beffbd7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe25068),
	.w1(32'hbbe7940c),
	.w2(32'hbb8e1a0d),
	.w3(32'h3bb6b989),
	.w4(32'hbad3464c),
	.w5(32'hbc6baf07),
	.w6(32'h3b07b280),
	.w7(32'hbbc329b3),
	.w8(32'hbb105047),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc017ef),
	.w1(32'hbacd6b60),
	.w2(32'h3b3248e5),
	.w3(32'hbbbc46a4),
	.w4(32'h3aa747d6),
	.w5(32'hbc470dbc),
	.w6(32'h3a8d8d28),
	.w7(32'h3c0e7955),
	.w8(32'h3b4a6d5a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f006e),
	.w1(32'h3c1f83a0),
	.w2(32'h3ba20858),
	.w3(32'hbb6cc436),
	.w4(32'h3b72ce1b),
	.w5(32'h3c6dc00f),
	.w6(32'hbc1ca77e),
	.w7(32'hbc2e799f),
	.w8(32'hbb21ac1d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fa05a),
	.w1(32'hbbcbe4b2),
	.w2(32'h3ac98795),
	.w3(32'hbbb5edfa),
	.w4(32'h3bfb9c57),
	.w5(32'hbbc08b23),
	.w6(32'h3a3a1555),
	.w7(32'h3b7ba828),
	.w8(32'h3bf9e598),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13789e),
	.w1(32'h3b86d7db),
	.w2(32'hbc3cb3cc),
	.w3(32'h3b35ed93),
	.w4(32'hbbf8d617),
	.w5(32'hbc1c0076),
	.w6(32'hbaa9406a),
	.w7(32'h3c08e269),
	.w8(32'hbc111f12),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea20d3),
	.w1(32'hbc2b8402),
	.w2(32'hbc28efd0),
	.w3(32'h3b61407b),
	.w4(32'hbc6b1d46),
	.w5(32'hbc82620d),
	.w6(32'hbbafb9f9),
	.w7(32'h3b4d0af2),
	.w8(32'hbbf8251f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7173e2),
	.w1(32'hbc1ca021),
	.w2(32'hbc08a12d),
	.w3(32'hbc5d5210),
	.w4(32'hbb54d627),
	.w5(32'hbcc5226c),
	.w6(32'hbc029dc7),
	.w7(32'hba4fe349),
	.w8(32'hbad32eb2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab059f1),
	.w1(32'h3c394bb1),
	.w2(32'h3bd100bb),
	.w3(32'hbb93a81a),
	.w4(32'h3b20f75b),
	.w5(32'h3b8581d5),
	.w6(32'hbb128a84),
	.w7(32'hbb07adb7),
	.w8(32'h3b93b7c6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68f51a),
	.w1(32'h3a59f453),
	.w2(32'h39b9d570),
	.w3(32'h3c43a150),
	.w4(32'hba643fad),
	.w5(32'h3b8483d4),
	.w6(32'h3c857714),
	.w7(32'hbb90ed96),
	.w8(32'h3a227a1d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb641a68),
	.w1(32'h3acd7674),
	.w2(32'hbb54222c),
	.w3(32'hbbbdc80f),
	.w4(32'hb8fccc92),
	.w5(32'hbc0242bd),
	.w6(32'hbbdc9703),
	.w7(32'hbc33a2d6),
	.w8(32'hbc41cfc6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96b5ae),
	.w1(32'hb9acde8c),
	.w2(32'hbbafd324),
	.w3(32'hbc596454),
	.w4(32'h3b31977a),
	.w5(32'hbb1fb7dd),
	.w6(32'h3a49bd96),
	.w7(32'h3a1264fb),
	.w8(32'h3a84235a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2151de),
	.w1(32'hbb87b581),
	.w2(32'h3b8f8e03),
	.w3(32'hbb3abb42),
	.w4(32'hbc2f46f9),
	.w5(32'h3d356775),
	.w6(32'h3c03a8db),
	.w7(32'hbc0921d7),
	.w8(32'h3c202304),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75dd77),
	.w1(32'h392e187a),
	.w2(32'hbbe31e40),
	.w3(32'hba2390e4),
	.w4(32'h3b8c93cb),
	.w5(32'h3a0ee3de),
	.w6(32'hbb2a2ba4),
	.w7(32'hba3604ae),
	.w8(32'h3a064017),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab87e9b),
	.w1(32'hbc1d33b7),
	.w2(32'hbb12f8c4),
	.w3(32'h3a79e743),
	.w4(32'h3a830e5f),
	.w5(32'h3a494439),
	.w6(32'h3a64d0b5),
	.w7(32'h3baa44c9),
	.w8(32'h3b37c03c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b482562),
	.w1(32'hbbe1f8a3),
	.w2(32'hbc76f695),
	.w3(32'hbb0d6566),
	.w4(32'hbb8c9ac3),
	.w5(32'hbcb291fb),
	.w6(32'h3a9732e3),
	.w7(32'hbb524259),
	.w8(32'h3ab4445a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbace95b),
	.w1(32'hbc214926),
	.w2(32'hba368fc2),
	.w3(32'hbc8bebc4),
	.w4(32'hbba312af),
	.w5(32'hb85d4ac4),
	.w6(32'hbb86fa57),
	.w7(32'h3a815574),
	.w8(32'hbb8e4809),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b654bb3),
	.w1(32'hbb224281),
	.w2(32'hbbd1d036),
	.w3(32'hbbd1b2c8),
	.w4(32'hbb8e6e90),
	.w5(32'h3bcfa37c),
	.w6(32'h3b4f874a),
	.w7(32'h3ad1ddc2),
	.w8(32'h3b2eee9b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc59597),
	.w1(32'h3b19f592),
	.w2(32'hbba84af3),
	.w3(32'hbabde607),
	.w4(32'hbac9b93f),
	.w5(32'h3c39781f),
	.w6(32'hba077a1b),
	.w7(32'h3b0c258c),
	.w8(32'h3bb5b3d8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1be0b5),
	.w1(32'hbbac5170),
	.w2(32'hba9a3622),
	.w3(32'hbc18970c),
	.w4(32'hba74e0dd),
	.w5(32'h3c0a72e0),
	.w6(32'h3a5df69b),
	.w7(32'hb97924ee),
	.w8(32'hba85f145),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43d96d),
	.w1(32'h3bcd7011),
	.w2(32'h3c0e54f2),
	.w3(32'h3b918763),
	.w4(32'h3bf473ff),
	.w5(32'h3cd1691b),
	.w6(32'hba5aa954),
	.w7(32'hb8ae0346),
	.w8(32'h3ca9523e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb890bea4),
	.w1(32'h39dc4265),
	.w2(32'hbbc0c72f),
	.w3(32'h3ab0d519),
	.w4(32'hbae1a47f),
	.w5(32'hbb289214),
	.w6(32'h3c2e81ba),
	.w7(32'hbb147aa8),
	.w8(32'h3bc74388),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ec7b7),
	.w1(32'hbbcfa16f),
	.w2(32'h3ae5dcd6),
	.w3(32'h3b6eace9),
	.w4(32'h3aaa9ed7),
	.w5(32'hbbc6e2b7),
	.w6(32'h3b4a6920),
	.w7(32'hbbb089a3),
	.w8(32'hbc0256f1),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd11f0f),
	.w1(32'h3b88fd29),
	.w2(32'h3c3ef63e),
	.w3(32'hbbd397c4),
	.w4(32'hbb58f906),
	.w5(32'h3c37ab3a),
	.w6(32'hbbe55329),
	.w7(32'hbb802f7e),
	.w8(32'h3cb20569),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa82be),
	.w1(32'hbbf32567),
	.w2(32'hbb142454),
	.w3(32'hbc1a953b),
	.w4(32'hbbfa529b),
	.w5(32'hbb0ddab4),
	.w6(32'h3b7aedff),
	.w7(32'hbc2b430a),
	.w8(32'h3baefa23),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38b572),
	.w1(32'hb94250f7),
	.w2(32'h3bf6179b),
	.w3(32'hbc00a334),
	.w4(32'h3b247bf9),
	.w5(32'h3c6c5fa5),
	.w6(32'hba90a9c8),
	.w7(32'h3b990881),
	.w8(32'h3c229e80),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad94a81),
	.w1(32'hbc08b569),
	.w2(32'hbc09a802),
	.w3(32'h3acdfc29),
	.w4(32'hbbed58ec),
	.w5(32'hbad27926),
	.w6(32'h3bdf9f6e),
	.w7(32'h3b4bd805),
	.w8(32'hbba75343),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadf181),
	.w1(32'hbc3dd85b),
	.w2(32'hbb226436),
	.w3(32'h3b0e0edc),
	.w4(32'h3b8d0c5a),
	.w5(32'hbc366687),
	.w6(32'hb90c81b1),
	.w7(32'hba9a7b27),
	.w8(32'hb975b784),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75d0dd),
	.w1(32'hbb075556),
	.w2(32'hbbbc596a),
	.w3(32'hbb86b8ff),
	.w4(32'h3b9a2ce7),
	.w5(32'hbc3abfc5),
	.w6(32'h39d55657),
	.w7(32'h3a93758f),
	.w8(32'h39d75fa1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f12c04),
	.w1(32'hbc08b27b),
	.w2(32'h3bd00696),
	.w3(32'hbc0c1865),
	.w4(32'hbc4ed36e),
	.w5(32'h3d04f255),
	.w6(32'hbb8f14b7),
	.w7(32'hbc3af36f),
	.w8(32'h3b5a2993),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc401a89),
	.w1(32'hba95fb88),
	.w2(32'hbc9c8f0d),
	.w3(32'hbbab66db),
	.w4(32'h3b816cfa),
	.w5(32'hbcdf44f0),
	.w6(32'hbc3d654b),
	.w7(32'hbc194227),
	.w8(32'hbbc366f2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b6d64),
	.w1(32'h3bcac413),
	.w2(32'hbb2c3384),
	.w3(32'hbc44e304),
	.w4(32'hbb84aeb5),
	.w5(32'h3d3a623b),
	.w6(32'h3a8f3650),
	.w7(32'hbc3e1e91),
	.w8(32'hbadc28fe),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc462990),
	.w1(32'hb9af16a2),
	.w2(32'hbb20f5b0),
	.w3(32'hbaf32321),
	.w4(32'hbb40e6e2),
	.w5(32'h3c28d2b5),
	.w6(32'hbab2f955),
	.w7(32'hbbae31ab),
	.w8(32'hbc053bd4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63e3fb),
	.w1(32'hbb5d3630),
	.w2(32'hbba61b7d),
	.w3(32'hbabd37d0),
	.w4(32'hbb8afc64),
	.w5(32'h3a91fec3),
	.w6(32'hbb42f136),
	.w7(32'hbb842d5b),
	.w8(32'hbbb9c787),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba68646),
	.w1(32'h3be7ad54),
	.w2(32'hba58eba1),
	.w3(32'hbbb15d74),
	.w4(32'h3c24db26),
	.w5(32'hbc5d26ae),
	.w6(32'hbba138a3),
	.w7(32'h3c10143c),
	.w8(32'hbb8ff683),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98bb5b),
	.w1(32'h3b88a5bb),
	.w2(32'hbb492882),
	.w3(32'hbb940e41),
	.w4(32'hbadf571c),
	.w5(32'h3cb647b1),
	.w6(32'hbafe238a),
	.w7(32'h3b407ee0),
	.w8(32'hbad4c2a1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ddcd9),
	.w1(32'h39d1f113),
	.w2(32'h3be4b859),
	.w3(32'h3b983302),
	.w4(32'h39c6d39e),
	.w5(32'h3d3930d9),
	.w6(32'h3b9e3834),
	.w7(32'hbc2da4db),
	.w8(32'hbb874ab7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb74035),
	.w1(32'hbaf49caf),
	.w2(32'hbc123eee),
	.w3(32'h3b87c16e),
	.w4(32'hbaed012b),
	.w5(32'h3d283434),
	.w6(32'h3aa0a7f6),
	.w7(32'hbc322f89),
	.w8(32'h3a3da552),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca027cc),
	.w1(32'hb7ff16d0),
	.w2(32'hbba78954),
	.w3(32'hbc13c778),
	.w4(32'hbad53b0e),
	.w5(32'hb9242187),
	.w6(32'hbc22d830),
	.w7(32'hbb356add),
	.w8(32'hb99ee10a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f4022d),
	.w1(32'hba760c28),
	.w2(32'h3bf876ed),
	.w3(32'hbb96f4ff),
	.w4(32'hbc466349),
	.w5(32'h3c58487f),
	.w6(32'hbb27ff3d),
	.w7(32'hbabffbeb),
	.w8(32'hbc0da7e7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b726e1a),
	.w1(32'hbbd8baea),
	.w2(32'hbb888c4a),
	.w3(32'h3bb23604),
	.w4(32'hbbdbe495),
	.w5(32'hbc283e05),
	.w6(32'h3b18e28a),
	.w7(32'hbc23cfbe),
	.w8(32'h3b875a2f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d53cf),
	.w1(32'hbc3528de),
	.w2(32'hbabf84e6),
	.w3(32'hbc032375),
	.w4(32'hbc2b01f0),
	.w5(32'hbca184f6),
	.w6(32'h3bba368d),
	.w7(32'hbb147848),
	.w8(32'hbbc8142a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc129931),
	.w1(32'hbbc324c8),
	.w2(32'hbbbb6253),
	.w3(32'hbc38fe90),
	.w4(32'h3b1653ed),
	.w5(32'hbc4ae534),
	.w6(32'h39c092a0),
	.w7(32'h3b657da3),
	.w8(32'hbb635b05),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e6276),
	.w1(32'hba828dc5),
	.w2(32'hb9785b51),
	.w3(32'hbb085e3f),
	.w4(32'hba7fdfe3),
	.w5(32'hbb47a1ec),
	.w6(32'h3aa6417d),
	.w7(32'h3aa3ce24),
	.w8(32'hbb251037),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b204027),
	.w1(32'hbb41cf64),
	.w2(32'h3af274ab),
	.w3(32'h3b9830a5),
	.w4(32'h3a3eccf9),
	.w5(32'h3cd11994),
	.w6(32'h3afd2d30),
	.w7(32'hbc117f21),
	.w8(32'h3b8d0825),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e67d6),
	.w1(32'hbb0b5741),
	.w2(32'h3b4eeb14),
	.w3(32'h399fd0c8),
	.w4(32'hbc04c9bc),
	.w5(32'h3a2cb9f3),
	.w6(32'h3b8ac755),
	.w7(32'hbb98fc92),
	.w8(32'h3c3289a6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6eef4e),
	.w1(32'hbbaca635),
	.w2(32'hbc2883a2),
	.w3(32'h3b826b73),
	.w4(32'hbc741439),
	.w5(32'hbc921a91),
	.w6(32'h3b8d4c46),
	.w7(32'hbb6f9ba1),
	.w8(32'hba4221f7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc67945),
	.w1(32'h3b1c62a5),
	.w2(32'h3a5293be),
	.w3(32'hbbe04297),
	.w4(32'hbb92d84e),
	.w5(32'h3c50e4e0),
	.w6(32'hba239ffa),
	.w7(32'hbb2eb443),
	.w8(32'hbb2666a6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a3e40),
	.w1(32'hbb23b26f),
	.w2(32'hb919eb76),
	.w3(32'h3c117a43),
	.w4(32'h3acf10d6),
	.w5(32'h3a99e4c1),
	.w6(32'h3bb4aa05),
	.w7(32'hbb02a8db),
	.w8(32'h3b4fec66),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9b855),
	.w1(32'h3b3db5be),
	.w2(32'h3bf21fab),
	.w3(32'h3b25698b),
	.w4(32'h3b9a7d84),
	.w5(32'h3b102834),
	.w6(32'h3b52f70d),
	.w7(32'hbc002861),
	.w8(32'hba011b08),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d4978),
	.w1(32'hbba597af),
	.w2(32'hbba044f8),
	.w3(32'h3b9162b4),
	.w4(32'h3bc013e1),
	.w5(32'hbc3490ac),
	.w6(32'h3b753f23),
	.w7(32'h3b901747),
	.w8(32'h3b3464e1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83e228),
	.w1(32'h3bc93ede),
	.w2(32'h3c2a5bb7),
	.w3(32'hba8cb8ef),
	.w4(32'hbb40b0cf),
	.w5(32'h3d1c1925),
	.w6(32'h3b0fb8a2),
	.w7(32'hbbc924c9),
	.w8(32'h3bacb133),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b969624),
	.w1(32'h39ca50fa),
	.w2(32'hba86d758),
	.w3(32'h3c5048e2),
	.w4(32'hbaf0817c),
	.w5(32'h3d3f96d2),
	.w6(32'h3c16c388),
	.w7(32'hbc6ab175),
	.w8(32'hbc36499a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52afb4),
	.w1(32'hbb5d571e),
	.w2(32'hbc6788fe),
	.w3(32'h3b3d1b70),
	.w4(32'h3ada6424),
	.w5(32'hbcb6e26c),
	.w6(32'hbb022bf0),
	.w7(32'hbc0738b4),
	.w8(32'hbbc55b1c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ba3a7),
	.w1(32'hba482a1a),
	.w2(32'h3af0518e),
	.w3(32'hbc6ad0fe),
	.w4(32'hbc26433c),
	.w5(32'hbc5594e5),
	.w6(32'hbbe91d24),
	.w7(32'hbb100f3d),
	.w8(32'hbc47cc2d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84cef4),
	.w1(32'h3c644a21),
	.w2(32'h3c02555a),
	.w3(32'hbc3bb5b7),
	.w4(32'h3c6d34db),
	.w5(32'h3b3304f7),
	.w6(32'hbbd9aa84),
	.w7(32'h3ba3512c),
	.w8(32'h3c3a45e5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1b972),
	.w1(32'hba70b731),
	.w2(32'hbb19eacd),
	.w3(32'h3be9898f),
	.w4(32'h3b12c69b),
	.w5(32'h39a525ca),
	.w6(32'h3c21bb79),
	.w7(32'h3b195975),
	.w8(32'h3b9d0e51),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a282806),
	.w1(32'hbc01d3c0),
	.w2(32'hbc8bfda1),
	.w3(32'h394e2a69),
	.w4(32'hbc30d31d),
	.w5(32'hbbc0e3c6),
	.w6(32'hbb03c7d6),
	.w7(32'hbb3c6be1),
	.w8(32'hbc04be56),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fc1e5),
	.w1(32'h3b9f33e2),
	.w2(32'h3c0d9349),
	.w3(32'h3bb0d803),
	.w4(32'h3bb7eb92),
	.w5(32'h3d269fa4),
	.w6(32'h3b5ca013),
	.w7(32'hbb11be80),
	.w8(32'h3b98c0f4),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe85cde),
	.w1(32'hbc3b6cb9),
	.w2(32'hbc0a1fd7),
	.w3(32'hbb7a820a),
	.w4(32'hbc293210),
	.w5(32'hbc89debd),
	.w6(32'h3b48410c),
	.w7(32'hbc2a8638),
	.w8(32'hbb813b15),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e9067),
	.w1(32'hbbd9838a),
	.w2(32'h3b588d3b),
	.w3(32'hbc08457d),
	.w4(32'hbbc1be6d),
	.w5(32'h3d0cda14),
	.w6(32'hbb8193c5),
	.w7(32'hbba18827),
	.w8(32'h3abf3aed),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30ec01),
	.w1(32'h3ba01f22),
	.w2(32'h3babf72a),
	.w3(32'h3bb4ff8f),
	.w4(32'hbb2ce932),
	.w5(32'hbc6c83ee),
	.w6(32'h3b83eaa3),
	.w7(32'h3a6c8b32),
	.w8(32'hbb97fe6f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b353768),
	.w1(32'hbadfd28e),
	.w2(32'h3b918b41),
	.w3(32'hbb20c577),
	.w4(32'hbb8b17eb),
	.w5(32'hbc768ba9),
	.w6(32'hbb158021),
	.w7(32'h3b205e61),
	.w8(32'h3c3bbbef),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7d42e),
	.w1(32'hbc0aebe4),
	.w2(32'hbc8b4507),
	.w3(32'hbbc53f97),
	.w4(32'hbb8d63a6),
	.w5(32'hbccd7859),
	.w6(32'hbb2fbc9c),
	.w7(32'h3c00771f),
	.w8(32'hbbe352fd),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14366b),
	.w1(32'h3b603b84),
	.w2(32'h3ae16344),
	.w3(32'hbc0c0525),
	.w4(32'hbbb6b6f4),
	.w5(32'h3c5b18c7),
	.w6(32'hbc03b298),
	.w7(32'hbb1f3426),
	.w8(32'hbb034542),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53936d),
	.w1(32'hbba0b4ee),
	.w2(32'hbc1d1cd3),
	.w3(32'h3ba3fc80),
	.w4(32'h3a8fae01),
	.w5(32'hbc41ee0c),
	.w6(32'h3b03b6c8),
	.w7(32'hbbfea21c),
	.w8(32'hbc802570),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46956f),
	.w1(32'h3bfccc0d),
	.w2(32'h3ca342d5),
	.w3(32'hbb961dff),
	.w4(32'hbc6708bd),
	.w5(32'h3cf855e7),
	.w6(32'hbbdf1d98),
	.w7(32'hbc0dd60a),
	.w8(32'hbc13a792),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9baa462),
	.w1(32'h3aaaca15),
	.w2(32'h3c010c8d),
	.w3(32'h3cbfb031),
	.w4(32'h3b5b0604),
	.w5(32'h3be1443b),
	.w6(32'hb9b87b87),
	.w7(32'h39e8087c),
	.w8(32'hba406f07),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91d4cb),
	.w1(32'hbc0a5fab),
	.w2(32'hbbdfaaaf),
	.w3(32'h3b908ee2),
	.w4(32'hbb8ef033),
	.w5(32'hbcae1cb6),
	.w6(32'hbc06ea88),
	.w7(32'h3bddd408),
	.w8(32'hbc78f2be),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3aac6),
	.w1(32'h3b770491),
	.w2(32'h3a14a6d4),
	.w3(32'hbbb8b51c),
	.w4(32'h3c228074),
	.w5(32'h3d657d86),
	.w6(32'h3bacf5b5),
	.w7(32'hbc3f6c69),
	.w8(32'h3c3dddb0),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc167f38),
	.w1(32'h3aa3c1dd),
	.w2(32'h3bef2cf1),
	.w3(32'hbc247e00),
	.w4(32'hbbef99bd),
	.w5(32'h3d291b90),
	.w6(32'h39992125),
	.w7(32'hbc5c5fd3),
	.w8(32'hbb011607),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd72d7),
	.w1(32'h37ae3e01),
	.w2(32'h3ae0389d),
	.w3(32'h3c25a51b),
	.w4(32'h3aac5946),
	.w5(32'h3b19ab39),
	.w6(32'h3ab40068),
	.w7(32'h3a346586),
	.w8(32'hbb9c86a0),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b253800),
	.w1(32'h399be5bf),
	.w2(32'hbb3ca709),
	.w3(32'h3a37d14b),
	.w4(32'hbc2dc920),
	.w5(32'hbc28152c),
	.w6(32'hbbe59f15),
	.w7(32'h3abce3a1),
	.w8(32'hbbc8acc7),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf23500),
	.w1(32'h3a182458),
	.w2(32'h3ba36015),
	.w3(32'hbb2791f7),
	.w4(32'h3b14770b),
	.w5(32'hbbcddd95),
	.w6(32'hbc0094ef),
	.w7(32'h3ace505e),
	.w8(32'h3b95ffb6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba290a),
	.w1(32'hba5095e3),
	.w2(32'h3c2db00e),
	.w3(32'hbbe66b61),
	.w4(32'hbc356d08),
	.w5(32'h3c92506d),
	.w6(32'hbbf6bd98),
	.w7(32'hbc19294a),
	.w8(32'hbc058db0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23a243),
	.w1(32'h3c0f81db),
	.w2(32'h3b9ad9ae),
	.w3(32'h3c16423b),
	.w4(32'h38e90bbc),
	.w5(32'h3a9d9d89),
	.w6(32'hbafb87d8),
	.w7(32'hbacfc822),
	.w8(32'hbb4564a7),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb255727),
	.w1(32'h3c197b61),
	.w2(32'h3b189dce),
	.w3(32'hbafbdfe5),
	.w4(32'hbaa538fe),
	.w5(32'h3c05c275),
	.w6(32'h382ac289),
	.w7(32'hb9d2ef38),
	.w8(32'h3acc8625),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57150e),
	.w1(32'hbb9c83ff),
	.w2(32'hbba08cfc),
	.w3(32'h3bd65244),
	.w4(32'hbaa87595),
	.w5(32'h3aaad801),
	.w6(32'h39ecd267),
	.w7(32'hbaa9ee46),
	.w8(32'hba72b1a7),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8b10d),
	.w1(32'h3b88c058),
	.w2(32'h3b31bb0e),
	.w3(32'hbbf22e4e),
	.w4(32'h3c2c38b4),
	.w5(32'h3b8fa0bc),
	.w6(32'hbb9a6e44),
	.w7(32'hbb801e4c),
	.w8(32'h3b4db52e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf81b7),
	.w1(32'h3a6075aa),
	.w2(32'h3bd5ab43),
	.w3(32'h3be4a594),
	.w4(32'h37da5e4b),
	.w5(32'h3a31a937),
	.w6(32'hb97bd3c6),
	.w7(32'hbbc025c2),
	.w8(32'hbb6a3fe2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb71464),
	.w1(32'h3b904769),
	.w2(32'hbb4ec874),
	.w3(32'h39446ceb),
	.w4(32'h3bbe559d),
	.w5(32'h3a12af63),
	.w6(32'hb9c09e61),
	.w7(32'h3accf72f),
	.w8(32'hbaf29ee5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb882894),
	.w1(32'h3b31c9e9),
	.w2(32'hba3bfee3),
	.w3(32'hbb95fd0d),
	.w4(32'h3b406835),
	.w5(32'hbba42412),
	.w6(32'hb9bc29a3),
	.w7(32'h3ac2b770),
	.w8(32'h3bd483a7),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7b5a7),
	.w1(32'hbb442812),
	.w2(32'h3bbe1684),
	.w3(32'h3c438f55),
	.w4(32'hbc0c3633),
	.w5(32'hbc1f64ed),
	.w6(32'h3be6a847),
	.w7(32'hbc2c0443),
	.w8(32'h3ab11df2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5b1c2),
	.w1(32'h3b139228),
	.w2(32'hbbdb94f4),
	.w3(32'hbc3e6aeb),
	.w4(32'h3ad9f830),
	.w5(32'hbbb5c683),
	.w6(32'hbb9563c9),
	.w7(32'h3bd63ee7),
	.w8(32'h3af05f72),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72ea93),
	.w1(32'h3ba7dd17),
	.w2(32'hbb042a79),
	.w3(32'hbb36c758),
	.w4(32'h3c1892c2),
	.w5(32'hbc2e1080),
	.w6(32'hbba1895a),
	.w7(32'h3a180ac2),
	.w8(32'hb9c67fbd),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10c869),
	.w1(32'hbaf24be2),
	.w2(32'hbb4fa9e6),
	.w3(32'hba72c6fc),
	.w4(32'h3b04ca4e),
	.w5(32'h39e86c46),
	.w6(32'hbb749eaf),
	.w7(32'h3b4a58c1),
	.w8(32'h3b1342dc),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe907c3),
	.w1(32'h3b6ec838),
	.w2(32'hb96ccf36),
	.w3(32'hbbfe6d7b),
	.w4(32'h3ab543ea),
	.w5(32'h3a5809f1),
	.w6(32'hbc01832c),
	.w7(32'h3b201522),
	.w8(32'h3bfe2165),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03f89f),
	.w1(32'hba84ad8e),
	.w2(32'h3a8fdd2b),
	.w3(32'h3b79f06c),
	.w4(32'hbb9fe545),
	.w5(32'h3c95df91),
	.w6(32'h3961953d),
	.w7(32'h38f90393),
	.w8(32'h3abcf945),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb373cb3),
	.w1(32'hb9ee9a1a),
	.w2(32'hbb19a06c),
	.w3(32'h3b9af9ad),
	.w4(32'h3b2b92d0),
	.w5(32'hbbaf6d63),
	.w6(32'h3b9399df),
	.w7(32'hb93de157),
	.w8(32'hbb3d8a4e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb44455),
	.w1(32'hbb2b92e1),
	.w2(32'hbbdc32d2),
	.w3(32'hbb225664),
	.w4(32'h37f85c33),
	.w5(32'hbc784b06),
	.w6(32'h3baf1cc3),
	.w7(32'hbadbd4e2),
	.w8(32'h3c0e30f9),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08da86),
	.w1(32'h3a55ee5f),
	.w2(32'h3c00da7e),
	.w3(32'h3ab945b5),
	.w4(32'hbb165447),
	.w5(32'h3bdb584f),
	.w6(32'h3aca0c0a),
	.w7(32'hbb7ca2f0),
	.w8(32'hba23abcf),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae98aeb),
	.w1(32'hbaa81c50),
	.w2(32'hbb1463b6),
	.w3(32'hbba92d89),
	.w4(32'hbb23ffaf),
	.w5(32'hbca24dbc),
	.w6(32'h3b8ca78c),
	.w7(32'h3b0810be),
	.w8(32'hbb5ec884),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a6114),
	.w1(32'hbb3f7a09),
	.w2(32'h3c35f9c1),
	.w3(32'hbb9f6ba9),
	.w4(32'hbbd8498e),
	.w5(32'h3ccb2d95),
	.w6(32'hbb14358b),
	.w7(32'hba30bcb1),
	.w8(32'h3bafce01),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5274db),
	.w1(32'h39c2027a),
	.w2(32'hbbd2fea0),
	.w3(32'h3c666c70),
	.w4(32'hbc245522),
	.w5(32'hbc0b05dc),
	.w6(32'h3c44ba0c),
	.w7(32'h3add26b5),
	.w8(32'hbc489965),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5489c3),
	.w1(32'h3978ac31),
	.w2(32'h3a54f36f),
	.w3(32'h3b89a558),
	.w4(32'hbba0c0e2),
	.w5(32'h3c7afe00),
	.w6(32'h3b8c0163),
	.w7(32'hbbaf69eb),
	.w8(32'hbb831492),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab98e29),
	.w1(32'hbbe36432),
	.w2(32'hbbc4496f),
	.w3(32'h3c16a74d),
	.w4(32'hbb9261b7),
	.w5(32'hbc380c13),
	.w6(32'h399bcfb8),
	.w7(32'hbbb26383),
	.w8(32'hbc1f48d7),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f5d00),
	.w1(32'hbbb8ca37),
	.w2(32'hbc80d257),
	.w3(32'h3abdc438),
	.w4(32'h3c565d34),
	.w5(32'h39218582),
	.w6(32'hbb37cb68),
	.w7(32'hbbfbef24),
	.w8(32'h39b8fb10),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb68050),
	.w1(32'h3b20e0be),
	.w2(32'h3c04b4da),
	.w3(32'hbc102344),
	.w4(32'hbb8dbc6d),
	.w5(32'h3c0745b1),
	.w6(32'h3af22a24),
	.w7(32'hbbaeb1b1),
	.w8(32'hbac28643),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a219b51),
	.w1(32'hbbbab296),
	.w2(32'hbc1c19a0),
	.w3(32'h3beab16d),
	.w4(32'hbc14f1fd),
	.w5(32'hbc865f9a),
	.w6(32'h3ba0dd80),
	.w7(32'hbbe30c32),
	.w8(32'hbc0e4865),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83501d),
	.w1(32'h3b5ac0f6),
	.w2(32'h3a1285ed),
	.w3(32'hbc957913),
	.w4(32'h3b4ab342),
	.w5(32'hbc13f6b3),
	.w6(32'hbbb8e364),
	.w7(32'h3bcb9f82),
	.w8(32'h3b874a23),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d3c8c),
	.w1(32'hbad3094b),
	.w2(32'h3b34a08e),
	.w3(32'h3b1ee39e),
	.w4(32'hbb339dfd),
	.w5(32'h3b603b26),
	.w6(32'h3b6756eb),
	.w7(32'hbbb78e41),
	.w8(32'h3b9876a1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe307c5),
	.w1(32'h3b454f8f),
	.w2(32'hbbb660df),
	.w3(32'hbb8083b9),
	.w4(32'h3b0e5617),
	.w5(32'h3b3875bb),
	.w6(32'hbad5f3c6),
	.w7(32'h3b4b7f73),
	.w8(32'h3b992726),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e939b),
	.w1(32'hba865f77),
	.w2(32'hbb592f6b),
	.w3(32'hba7c0fda),
	.w4(32'h3baca245),
	.w5(32'h3aec2328),
	.w6(32'hbbcebbcb),
	.w7(32'h3a7114e8),
	.w8(32'hbb7fe262),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20a213),
	.w1(32'hbb1489e9),
	.w2(32'hba859032),
	.w3(32'hbb844bde),
	.w4(32'hbbe87d9c),
	.w5(32'hbab5a3fa),
	.w6(32'h3a9a4424),
	.w7(32'h3a97609d),
	.w8(32'hbb384f2c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f296b),
	.w1(32'h3c2bb1b7),
	.w2(32'h3c0e7fda),
	.w3(32'hbb20b57e),
	.w4(32'h3c6df714),
	.w5(32'h3ced54d9),
	.w6(32'h3a272e82),
	.w7(32'h3be134a1),
	.w8(32'h3c138f39),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b960af0),
	.w1(32'hbbe3a048),
	.w2(32'hbc841ec8),
	.w3(32'h3c4dd0c0),
	.w4(32'hb996ad3b),
	.w5(32'hbc5bde44),
	.w6(32'h3c0b67be),
	.w7(32'h3b671654),
	.w8(32'hbc1c76df),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6645fb),
	.w1(32'h3a87a827),
	.w2(32'hb9c42c01),
	.w3(32'hbbb438c9),
	.w4(32'hbafa1908),
	.w5(32'hbab1538f),
	.w6(32'hbc0364c5),
	.w7(32'h3b4692e7),
	.w8(32'hba5053f3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7167ec),
	.w1(32'h3b13926c),
	.w2(32'h3be0cd93),
	.w3(32'h3bc70fab),
	.w4(32'h3bab79b1),
	.w5(32'h3acc1cc1),
	.w6(32'hbb6a5f40),
	.w7(32'hbb172a91),
	.w8(32'h3bf22a12),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73e8d6),
	.w1(32'h3b4fbe5e),
	.w2(32'hbbe6a471),
	.w3(32'h39bad7e9),
	.w4(32'h3a44de61),
	.w5(32'hbc2bafcc),
	.w6(32'h3abd606b),
	.w7(32'h3b862c07),
	.w8(32'hbb1e5e95),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5eddb),
	.w1(32'hbc0c1086),
	.w2(32'hbc3e4200),
	.w3(32'h3bdc4d87),
	.w4(32'hbc5872b9),
	.w5(32'hbc825907),
	.w6(32'h3b5908e3),
	.w7(32'h3a7168a1),
	.w8(32'hbc21f42b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fdc37),
	.w1(32'hbad847ca),
	.w2(32'h3a86ccdc),
	.w3(32'hbc0ac1a8),
	.w4(32'hbb9ef357),
	.w5(32'h389a23bd),
	.w6(32'hbbec7e49),
	.w7(32'hbb744da6),
	.w8(32'hbc2e10dc),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc020583),
	.w1(32'hbacd8446),
	.w2(32'h3a25820b),
	.w3(32'hbb94839c),
	.w4(32'hbc1e0a4b),
	.w5(32'h3c871ae4),
	.w6(32'hba899aec),
	.w7(32'h39c53892),
	.w8(32'hba18c81e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc07cb6),
	.w1(32'hbb18d8e6),
	.w2(32'h3b653364),
	.w3(32'hbbd9c470),
	.w4(32'hb9cda22b),
	.w5(32'hbc04f9bb),
	.w6(32'hbb2f1abd),
	.w7(32'h3b8e4da4),
	.w8(32'hbb6e9d15),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a1b13),
	.w1(32'h3acad66e),
	.w2(32'hb93ea32d),
	.w3(32'hba759b49),
	.w4(32'hbc126529),
	.w5(32'hbbe8e632),
	.w6(32'h39a363e9),
	.w7(32'hba92d5fe),
	.w8(32'hbc10cdad),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a10d4),
	.w1(32'h3b331501),
	.w2(32'hbbf3aff3),
	.w3(32'hba997c83),
	.w4(32'h3bccdef8),
	.w5(32'hbc537804),
	.w6(32'hbc2aaee8),
	.w7(32'h3bc98d17),
	.w8(32'hbc1ec966),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ad5e9),
	.w1(32'hba610ee5),
	.w2(32'hbc149367),
	.w3(32'h3a72e8da),
	.w4(32'hbbb8cc7e),
	.w5(32'hbb892b2b),
	.w6(32'hbb9ab6d1),
	.w7(32'h3ba74eb8),
	.w8(32'hbbcc7c4d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb068982),
	.w1(32'hba7536dc),
	.w2(32'hbbda5eed),
	.w3(32'h3b610415),
	.w4(32'hbbb42717),
	.w5(32'hbb28214a),
	.w6(32'h3b3210fc),
	.w7(32'h3b26592e),
	.w8(32'hbb9b9ed9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0466c6),
	.w1(32'h3abb11ab),
	.w2(32'h3bae7236),
	.w3(32'hbb1a8860),
	.w4(32'hbc133e79),
	.w5(32'h3d3e827b),
	.w6(32'hb9fd1417),
	.w7(32'hbc01bb91),
	.w8(32'h3bd24bc5),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf737db),
	.w1(32'hbb271291),
	.w2(32'hbc429c78),
	.w3(32'h3b441678),
	.w4(32'h3b45b1d3),
	.w5(32'hbbd0aa24),
	.w6(32'h3c03f12e),
	.w7(32'h391e7a68),
	.w8(32'hbb21d203),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10671c),
	.w1(32'h3bb3fd8f),
	.w2(32'hbb174e8d),
	.w3(32'hbc3978dd),
	.w4(32'h3b61252e),
	.w5(32'hbb491ec1),
	.w6(32'hba6b6237),
	.w7(32'h3bdf8fe3),
	.w8(32'h393c9d35),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f83e3),
	.w1(32'h3c0be4af),
	.w2(32'h3b45291b),
	.w3(32'hbb67f824),
	.w4(32'h3bd5d432),
	.w5(32'hbbf2f0c2),
	.w6(32'hbb7d6f3c),
	.w7(32'h3ae5b77a),
	.w8(32'hbb3b4b15),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd901bb),
	.w1(32'h3c518ada),
	.w2(32'h3c45ed24),
	.w3(32'hba96b1f4),
	.w4(32'h3bcc4394),
	.w5(32'h3cd78b23),
	.w6(32'hbb2da827),
	.w7(32'hbbc90cb0),
	.w8(32'h3c22ea4b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e14df),
	.w1(32'h39e207ac),
	.w2(32'hbc187ec1),
	.w3(32'h3c2a648d),
	.w4(32'h3bde02d0),
	.w5(32'h3bba9c70),
	.w6(32'h3c563e07),
	.w7(32'h3b709bbe),
	.w8(32'h3b851f13),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b4fb3),
	.w1(32'h3b9069ac),
	.w2(32'hbb9fc844),
	.w3(32'hbc0cd332),
	.w4(32'h3a780e80),
	.w5(32'h3b6ef62a),
	.w6(32'h37a96477),
	.w7(32'h3c0707e7),
	.w8(32'h3b12f0eb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c3ec0),
	.w1(32'hbc009b51),
	.w2(32'h3a552f77),
	.w3(32'hbca36d27),
	.w4(32'h3af5c8f7),
	.w5(32'hbae63fb6),
	.w6(32'hbbb3bf57),
	.w7(32'h3c4baf4b),
	.w8(32'hbad144a8),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b952d),
	.w1(32'h3b453383),
	.w2(32'h3ae1c563),
	.w3(32'hba66997c),
	.w4(32'h3c185c59),
	.w5(32'h3a1f3043),
	.w6(32'h3a161a5e),
	.w7(32'h3c0f1895),
	.w8(32'hb91304fd),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb676a98),
	.w1(32'hba11d88b),
	.w2(32'hbb16ffe6),
	.w3(32'hbb1f4168),
	.w4(32'hbb5c8a91),
	.w5(32'hbb04cd8c),
	.w6(32'h3a400c9c),
	.w7(32'hbaa45016),
	.w8(32'hbb5171cf),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27a1c0),
	.w1(32'hbb06a4cf),
	.w2(32'hbb57c0d1),
	.w3(32'h382c0446),
	.w4(32'h3ae355a2),
	.w5(32'h3c2ddcab),
	.w6(32'hbab36e99),
	.w7(32'h3bbd21fa),
	.w8(32'h3ac66bac),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedb6ba),
	.w1(32'h3b62461e),
	.w2(32'hbb8e7b81),
	.w3(32'hbaf47300),
	.w4(32'h3ae29ab5),
	.w5(32'hbba9c7a0),
	.w6(32'h3af2f8b8),
	.w7(32'h3b3b4138),
	.w8(32'hba83190a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba02425),
	.w1(32'h3ae43cc0),
	.w2(32'hbb9aa635),
	.w3(32'hbc1c1ce4),
	.w4(32'h3984c2c0),
	.w5(32'hbc1351b6),
	.w6(32'hbbd4b915),
	.w7(32'hba5263d4),
	.w8(32'hbab15ffc),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d726f6),
	.w1(32'h3a545c28),
	.w2(32'hba8966e7),
	.w3(32'h3c039efc),
	.w4(32'hbb0322c8),
	.w5(32'hbac19b15),
	.w6(32'h3bbd1fbf),
	.w7(32'hbad3c8b6),
	.w8(32'hbaaba665),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0a021),
	.w1(32'h3b45909d),
	.w2(32'hbb2164df),
	.w3(32'hbb1aaf96),
	.w4(32'hba62515f),
	.w5(32'hbbea15bd),
	.w6(32'h3b5643a5),
	.w7(32'hbb4aeba0),
	.w8(32'hbb63216f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946670b),
	.w1(32'hbbc234e2),
	.w2(32'hbba179b5),
	.w3(32'h3b166949),
	.w4(32'hbb314ae2),
	.w5(32'hbaf04930),
	.w6(32'hbb261d98),
	.w7(32'hbb384ecc),
	.w8(32'hba8fbf36),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad120a),
	.w1(32'h3b9ebcbb),
	.w2(32'hbb495db5),
	.w3(32'h398d5c28),
	.w4(32'h3b60c4a5),
	.w5(32'h3a61dd53),
	.w6(32'hbb9254cc),
	.w7(32'h3b3e9774),
	.w8(32'h3abc9218),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb596db7),
	.w1(32'h3aa28857),
	.w2(32'hbb22c0c4),
	.w3(32'h3b5e3d8f),
	.w4(32'h39fe65b5),
	.w5(32'h3b78c81a),
	.w6(32'h3b1a13e1),
	.w7(32'hbb0c3d25),
	.w8(32'hbb23ea55),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd87853),
	.w1(32'hbb281742),
	.w2(32'hba874ece),
	.w3(32'h3bcbaac3),
	.w4(32'hbb6de163),
	.w5(32'hbb6aa977),
	.w6(32'h3b7c0109),
	.w7(32'hbb87a588),
	.w8(32'h3af577f0),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983738c),
	.w1(32'h3b2ea8e2),
	.w2(32'h3b90e1c4),
	.w3(32'hbbabd95f),
	.w4(32'h3c51b44a),
	.w5(32'h3b4f94d9),
	.w6(32'h3ab94dda),
	.w7(32'h3c4575cc),
	.w8(32'h3bc2f678),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8804a0),
	.w1(32'hb9db888e),
	.w2(32'h3abf0bc0),
	.w3(32'h3c052e5d),
	.w4(32'hbaec9d59),
	.w5(32'h390dfabb),
	.w6(32'h3bc166a8),
	.w7(32'h3a839493),
	.w8(32'h3a96ed63),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2a152),
	.w1(32'hbb3cc56f),
	.w2(32'h3a4a3660),
	.w3(32'hba1d3c3d),
	.w4(32'h3b592c7e),
	.w5(32'h3bbde7ae),
	.w6(32'h3a869047),
	.w7(32'h3b163727),
	.w8(32'hbb4793a5),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a0073),
	.w1(32'h3bb9dd9f),
	.w2(32'h372bf351),
	.w3(32'hbb912906),
	.w4(32'h3b8c4d50),
	.w5(32'hbb193363),
	.w6(32'hbb8c4b10),
	.w7(32'h39f79a11),
	.w8(32'h388018a0),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba27697),
	.w1(32'h3ac9dc36),
	.w2(32'hbb2b3ef9),
	.w3(32'h3b4fe2c1),
	.w4(32'h39a1b2bf),
	.w5(32'hbb38eb92),
	.w6(32'h3ae4644f),
	.w7(32'h3b9ad6ce),
	.w8(32'h3a934510),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf5a27),
	.w1(32'hbb45046e),
	.w2(32'hba936fc4),
	.w3(32'h3ba5f5df),
	.w4(32'h3b08f196),
	.w5(32'h3ab68b9e),
	.w6(32'h3b8244b7),
	.w7(32'hbb9117fd),
	.w8(32'hbc01d816),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5a3ed),
	.w1(32'hbaf17add),
	.w2(32'hbac4891e),
	.w3(32'hbbc88d32),
	.w4(32'hbb5079f4),
	.w5(32'hb9f9681a),
	.w6(32'hbab87162),
	.w7(32'h3aacb48b),
	.w8(32'h3a957325),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13e9e0),
	.w1(32'hba55b6be),
	.w2(32'h3a805bc4),
	.w3(32'h3b38f56c),
	.w4(32'hbbcf7486),
	.w5(32'h3ba50e51),
	.w6(32'h3ad030f7),
	.w7(32'h3affd8d2),
	.w8(32'hbb6f1549),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad63d59),
	.w1(32'hbb08f168),
	.w2(32'h3b1c9086),
	.w3(32'hb9ebf18b),
	.w4(32'hba739cd1),
	.w5(32'h39f10b1e),
	.w6(32'h37db2873),
	.w7(32'hbaf639fb),
	.w8(32'hbb33aac1),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac57e5c),
	.w1(32'hbad92764),
	.w2(32'h3ab1e8b4),
	.w3(32'h3b849b42),
	.w4(32'hbb70b2cf),
	.w5(32'h3a0912d3),
	.w6(32'hbb1e0eca),
	.w7(32'hbb55a039),
	.w8(32'hba744faa),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66ff52),
	.w1(32'hbaca153d),
	.w2(32'hbb26686b),
	.w3(32'hbb48eba9),
	.w4(32'hbba72642),
	.w5(32'hbbd079ce),
	.w6(32'hbb3c1c62),
	.w7(32'hbb8cc75b),
	.w8(32'hbc08e66f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc125439),
	.w1(32'hba37c828),
	.w2(32'h3af2cdaf),
	.w3(32'hbb829c1d),
	.w4(32'hbb294fe8),
	.w5(32'h3b015704),
	.w6(32'hbc10303f),
	.w7(32'h3b277bb2),
	.w8(32'h3b7ba1ae),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd3f58),
	.w1(32'hbaf31f91),
	.w2(32'h3b4e25a5),
	.w3(32'hbb3f9117),
	.w4(32'hbb453e80),
	.w5(32'h3b11c19d),
	.w6(32'h3bbe8a87),
	.w7(32'hbb4e11a8),
	.w8(32'hba25164d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b405578),
	.w1(32'h3ad6a80f),
	.w2(32'hbb459ea9),
	.w3(32'hbb4ddb30),
	.w4(32'h3bd97bd9),
	.w5(32'hbae7c6eb),
	.w6(32'hbb872299),
	.w7(32'h3b3c1c5e),
	.w8(32'h3b8fdef9),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e8f22),
	.w1(32'h3b382bf7),
	.w2(32'h3b71eb8e),
	.w3(32'hb9650fe0),
	.w4(32'hbb1f6ee9),
	.w5(32'hbba9b7b0),
	.w6(32'h3ab13312),
	.w7(32'hbb710dd7),
	.w8(32'h3ad55fa8),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7834c),
	.w1(32'h3bcb0e13),
	.w2(32'h3b163790),
	.w3(32'hbb9a603f),
	.w4(32'h3b38cee3),
	.w5(32'hbabd70d8),
	.w6(32'h3a226587),
	.w7(32'h3b86a03d),
	.w8(32'h3b4613b1),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0423a),
	.w1(32'h3b1d41e1),
	.w2(32'hbb067002),
	.w3(32'h3be68f3b),
	.w4(32'h3aebd574),
	.w5(32'hbb56fc74),
	.w6(32'h3be013f9),
	.w7(32'h3ae6bbad),
	.w8(32'hbb8cda6c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2799b4),
	.w1(32'hbb5a66bf),
	.w2(32'h3b3c93a1),
	.w3(32'h3a227234),
	.w4(32'h3823c692),
	.w5(32'hb9ac9365),
	.w6(32'h3a6860de),
	.w7(32'hbb65db4b),
	.w8(32'h3ab01225),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b869cc9),
	.w1(32'hba961a6d),
	.w2(32'h3b742e0e),
	.w3(32'h3b9916e0),
	.w4(32'h392fb395),
	.w5(32'h3ab8df1b),
	.w6(32'h3b54f9b1),
	.w7(32'h3b2da781),
	.w8(32'h3acad4de),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62e487),
	.w1(32'h3bf66e0f),
	.w2(32'h3bbe590e),
	.w3(32'hbb76bdec),
	.w4(32'hba8aa200),
	.w5(32'hbaa2b556),
	.w6(32'hbb2559c9),
	.w7(32'h39a3aae6),
	.w8(32'hbb11240a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49eaa2),
	.w1(32'h3b13feec),
	.w2(32'h3a481e25),
	.w3(32'hb996fe5c),
	.w4(32'h3b2f6233),
	.w5(32'hbb0e9aba),
	.w6(32'hbb509098),
	.w7(32'hb9a9fab3),
	.w8(32'h3a91b076),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fb9e0),
	.w1(32'hba7c6805),
	.w2(32'hbbb1352e),
	.w3(32'h3b1f7dbc),
	.w4(32'h39d95fc9),
	.w5(32'hbbc3bba7),
	.w6(32'h3b36949a),
	.w7(32'hbacda6ef),
	.w8(32'hbb6c37fd),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0661a7),
	.w1(32'hbc081bfb),
	.w2(32'hba9d2816),
	.w3(32'hb9b55cf9),
	.w4(32'h3a580da8),
	.w5(32'h3c7a068b),
	.w6(32'h3a0f24d4),
	.w7(32'h3b4c27b0),
	.w8(32'hbb12d1d8),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe27118),
	.w1(32'h3b795004),
	.w2(32'hbb48663d),
	.w3(32'hbab80fd8),
	.w4(32'h39a29f3f),
	.w5(32'hba4c582b),
	.w6(32'hbabfd557),
	.w7(32'h3b04ba0e),
	.w8(32'hbb4c4f05),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8915c),
	.w1(32'h3a32acb2),
	.w2(32'h3afdcc4b),
	.w3(32'h3ba0c414),
	.w4(32'h3a8ff348),
	.w5(32'h3b3884f9),
	.w6(32'h3b08c90e),
	.w7(32'h3ab360f7),
	.w8(32'h3ba78608),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd7415),
	.w1(32'h3b267aed),
	.w2(32'h3baed744),
	.w3(32'h3b989aee),
	.w4(32'h3b9f2694),
	.w5(32'h3be8f267),
	.w6(32'h3a678faa),
	.w7(32'h3ad5cce5),
	.w8(32'h3b95b478),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8726f4),
	.w1(32'h3943bdbf),
	.w2(32'hbba15434),
	.w3(32'h3b38634d),
	.w4(32'hbaab0a06),
	.w5(32'hbbb1d65d),
	.w6(32'h3b6eca2d),
	.w7(32'hba676ff7),
	.w8(32'hbb6d058a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba72401),
	.w1(32'hbad6e2b6),
	.w2(32'h388f63dd),
	.w3(32'h3ac3dace),
	.w4(32'hbb37f135),
	.w5(32'hbb3de951),
	.w6(32'h3b029a7f),
	.w7(32'h3b2a2b5e),
	.w8(32'hbab51521),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c3a46),
	.w1(32'h3baec843),
	.w2(32'h3af7c74a),
	.w3(32'hbabafcf0),
	.w4(32'h3bac9cd4),
	.w5(32'hbab7a260),
	.w6(32'h3b08cd5c),
	.w7(32'h3b886a2e),
	.w8(32'h3b8028c5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eb2b1),
	.w1(32'h3adc0bb1),
	.w2(32'h3a0ac19d),
	.w3(32'h3bf5edf9),
	.w4(32'h3ac6c841),
	.w5(32'hbb409668),
	.w6(32'h3bb8e9ae),
	.w7(32'hba348664),
	.w8(32'h3bd39e11),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58175a),
	.w1(32'hbaca99ae),
	.w2(32'hbb8b2891),
	.w3(32'h3ba3fbb8),
	.w4(32'hba450ade),
	.w5(32'hbbd0959b),
	.w6(32'h3b01c74c),
	.w7(32'h3a8a51b2),
	.w8(32'h3a262bd6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b07c2),
	.w1(32'hbb3aa812),
	.w2(32'hba986093),
	.w3(32'hba04847a),
	.w4(32'h3b8fd0dc),
	.w5(32'hbb9a017b),
	.w6(32'h3ac82be2),
	.w7(32'hbb0e54c0),
	.w8(32'hbb97fe5d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c0a64),
	.w1(32'hbbbd0866),
	.w2(32'h3b0aac68),
	.w3(32'hbbd390e7),
	.w4(32'hba612130),
	.w5(32'h3b256bf9),
	.w6(32'hbb988bd2),
	.w7(32'hbb666a28),
	.w8(32'hba15b468),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeaeb2),
	.w1(32'h3c3fffb9),
	.w2(32'hbbc3c968),
	.w3(32'hbb45ef7a),
	.w4(32'h3c3c19f4),
	.w5(32'hbc0acd64),
	.w6(32'hba8cb9da),
	.w7(32'h3b8ae101),
	.w8(32'hba7410d2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1900aa),
	.w1(32'hbb912966),
	.w2(32'hbc09d3ea),
	.w3(32'h3c9c54da),
	.w4(32'hbb758c3d),
	.w5(32'hbb2865a3),
	.w6(32'h3c21a4a3),
	.w7(32'hbc0022ea),
	.w8(32'hbbecae6c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7949d),
	.w1(32'hbb670ffe),
	.w2(32'hbb48df99),
	.w3(32'hbba473da),
	.w4(32'hbb63f9cb),
	.w5(32'hbb085df8),
	.w6(32'hbbf05743),
	.w7(32'hbb81db1a),
	.w8(32'hbb157ebc),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb975e2e),
	.w1(32'h3a9eb7e8),
	.w2(32'hb8d904c6),
	.w3(32'hbae781ae),
	.w4(32'h3be80b7e),
	.w5(32'h3b16ae6d),
	.w6(32'hbb34d59b),
	.w7(32'h3b869952),
	.w8(32'h3ba3ca17),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75907a),
	.w1(32'hbb484afb),
	.w2(32'hbb180915),
	.w3(32'h3accdf6c),
	.w4(32'hbc01592f),
	.w5(32'hbbb54bb0),
	.w6(32'hb94d3e07),
	.w7(32'hbbb7436a),
	.w8(32'hba154611),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db88c),
	.w1(32'h3b60adb5),
	.w2(32'h3b9ca73b),
	.w3(32'h3a71dc2e),
	.w4(32'h3a158723),
	.w5(32'h39dd1a84),
	.w6(32'hbb3a851b),
	.w7(32'h3ba628b8),
	.w8(32'h3ba37f31),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e2af6),
	.w1(32'hbb367428),
	.w2(32'h3c1429cf),
	.w3(32'h3b2c24df),
	.w4(32'h3b82c764),
	.w5(32'h3c30e798),
	.w6(32'h3baba862),
	.w7(32'h3a389f18),
	.w8(32'h3b4f7ecd),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb124acf),
	.w1(32'hba8f2bed),
	.w2(32'h38a23a72),
	.w3(32'hbc0dd889),
	.w4(32'h39495649),
	.w5(32'h39a9beae),
	.w6(32'hbbddef52),
	.w7(32'h39a56d6e),
	.w8(32'hbae4546c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a1c80),
	.w1(32'hbb525c0d),
	.w2(32'h3b9f58b6),
	.w3(32'h3b9ae57a),
	.w4(32'h3acbf6d8),
	.w5(32'hbba907b7),
	.w6(32'hbbaf341e),
	.w7(32'hbb4fa4e3),
	.w8(32'hbbc4b3ed),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22699c),
	.w1(32'hbaedb079),
	.w2(32'hbab9ca46),
	.w3(32'hbbfe29d9),
	.w4(32'hbab2b938),
	.w5(32'h3a8aa55b),
	.w6(32'hbb519591),
	.w7(32'h38f1f3fb),
	.w8(32'hbb8b88e0),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace721f),
	.w1(32'h3a2d24c4),
	.w2(32'h3b6765ee),
	.w3(32'hbb66e860),
	.w4(32'h3b9504e6),
	.w5(32'hbad97d30),
	.w6(32'hbacb5ba2),
	.w7(32'hbadaf194),
	.w8(32'hbb3765fb),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13366d),
	.w1(32'h3b1aa6da),
	.w2(32'h3a02c30d),
	.w3(32'h3b7f29cb),
	.w4(32'h3a015fe5),
	.w5(32'hba872119),
	.w6(32'h3aebeeba),
	.w7(32'h3b903077),
	.w8(32'h3b928bed),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af61782),
	.w1(32'h3a38721c),
	.w2(32'hbb16c53a),
	.w3(32'h3bd02036),
	.w4(32'hbb192d20),
	.w5(32'h3adbc2c7),
	.w6(32'h3ad82b8a),
	.w7(32'hbb388a78),
	.w8(32'h3ad292e0),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34230f),
	.w1(32'hba78f773),
	.w2(32'hb9c1f316),
	.w3(32'h3be1a6f7),
	.w4(32'hbbf2fbff),
	.w5(32'hba43ce2c),
	.w6(32'h3b96295d),
	.w7(32'hbb9ab4fd),
	.w8(32'hbb9865af),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af45498),
	.w1(32'hbb2530d1),
	.w2(32'hba42cb78),
	.w3(32'hbb980ed0),
	.w4(32'hbba49850),
	.w5(32'hbae8be86),
	.w6(32'hbba4ae3b),
	.w7(32'hbb56428b),
	.w8(32'hbaf280db),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule