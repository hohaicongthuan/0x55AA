module layer_8_featuremap_111(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e821e),
	.w1(32'hbb27e369),
	.w2(32'h3be790a9),
	.w3(32'hbbcb2595),
	.w4(32'hb93195b9),
	.w5(32'hbb36f7aa),
	.w6(32'hbbe81b86),
	.w7(32'h3ac22be9),
	.w8(32'hbc13c956),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfed332),
	.w1(32'h39d5479c),
	.w2(32'h3c0ab9b7),
	.w3(32'h3a5bb3cf),
	.w4(32'h3c60b4e0),
	.w5(32'h3c2ee9e9),
	.w6(32'hbac34771),
	.w7(32'h3c424817),
	.w8(32'hba8fd50a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23c8dd),
	.w1(32'hbbe372aa),
	.w2(32'h3bd0afb0),
	.w3(32'hbace9fdb),
	.w4(32'hb7d49ab7),
	.w5(32'h3c3a334c),
	.w6(32'hbb500ee4),
	.w7(32'h3c40178f),
	.w8(32'h3b98a09a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c830918),
	.w1(32'hbbb54741),
	.w2(32'hbc9cf4a3),
	.w3(32'h38b6b18f),
	.w4(32'h3bb81334),
	.w5(32'h3ab87db5),
	.w6(32'hbb51afba),
	.w7(32'hbc715fb1),
	.w8(32'h3b629cd6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc992812),
	.w1(32'h39e6c6e4),
	.w2(32'h3b29218b),
	.w3(32'h3b7d89bb),
	.w4(32'h3c74975a),
	.w5(32'h3b615115),
	.w6(32'h39b9a2cb),
	.w7(32'h3a0d3f70),
	.w8(32'h3ad18d00),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5735a),
	.w1(32'h3b805647),
	.w2(32'h3a49032c),
	.w3(32'hbad00a7a),
	.w4(32'h3bef4b02),
	.w5(32'h3a8831c7),
	.w6(32'hbc0baa29),
	.w7(32'hbc1fbb45),
	.w8(32'hbb89a0a4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e626e),
	.w1(32'hbb8d9c35),
	.w2(32'h3bc07359),
	.w3(32'h3aefde5c),
	.w4(32'h3bc10fbb),
	.w5(32'hbb327831),
	.w6(32'h3b2248c1),
	.w7(32'hba6a6504),
	.w8(32'hbb8f996e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb981dc7),
	.w1(32'h3ade39dd),
	.w2(32'h3c321016),
	.w3(32'h3b83b7e0),
	.w4(32'h3c695ca5),
	.w5(32'h3bfbca86),
	.w6(32'h3bbce2bb),
	.w7(32'h3c35c814),
	.w8(32'h3a4859c7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ea97d),
	.w1(32'hbb9ce575),
	.w2(32'h3b8076e1),
	.w3(32'hbab413f3),
	.w4(32'h3bf4d65e),
	.w5(32'h3bfa0da2),
	.w6(32'hbb815b5b),
	.w7(32'hbb551dfe),
	.w8(32'hbbff0e1f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3214de),
	.w1(32'h3b8b044b),
	.w2(32'hbc59732f),
	.w3(32'h3aaf6543),
	.w4(32'h3b8b0fdf),
	.w5(32'h3b810ac2),
	.w6(32'hbb25e700),
	.w7(32'hbc9934d2),
	.w8(32'hbc17b424),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6c095),
	.w1(32'hbc127020),
	.w2(32'hbcc0f902),
	.w3(32'hb9f84c90),
	.w4(32'hbc4ac8a1),
	.w5(32'h3af69866),
	.w6(32'hbba0893a),
	.w7(32'hbbd04cbb),
	.w8(32'hbc457ed0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3053a),
	.w1(32'hbc8a8e55),
	.w2(32'h3bf3a91d),
	.w3(32'hbbfdd3ac),
	.w4(32'h3c111c71),
	.w5(32'h3ab5411e),
	.w6(32'hbb0fed01),
	.w7(32'hbab690fb),
	.w8(32'hbb6e84a1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7c18a),
	.w1(32'hb93e8f54),
	.w2(32'h3a6ce2b9),
	.w3(32'h3ba191a8),
	.w4(32'h3bafa420),
	.w5(32'h3bf50ecf),
	.w6(32'h3afd40da),
	.w7(32'h3bed9453),
	.w8(32'h3c964971),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a7a93),
	.w1(32'hbaa2f28b),
	.w2(32'h3a88f23a),
	.w3(32'h3a6cff22),
	.w4(32'h3a894d5d),
	.w5(32'hbb0c63d9),
	.w6(32'h3c2e881d),
	.w7(32'h3b972479),
	.w8(32'hbad3d2d8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff539f),
	.w1(32'h3b39a284),
	.w2(32'h3aec551a),
	.w3(32'h3b07c6a8),
	.w4(32'h3b08eff0),
	.w5(32'h396f1878),
	.w6(32'h3b30137b),
	.w7(32'h3b84d1ea),
	.w8(32'h3aaba49c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d2e20),
	.w1(32'h3b994fa3),
	.w2(32'h3a61760d),
	.w3(32'h3b746d76),
	.w4(32'h39fb94b8),
	.w5(32'h3a0c1ee0),
	.w6(32'h3b9c58ed),
	.w7(32'hbb03cf77),
	.w8(32'h3bc72e39),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e4882),
	.w1(32'h3bc29ada),
	.w2(32'h3b2dcea3),
	.w3(32'hb8e99dc3),
	.w4(32'h3bd29d33),
	.w5(32'hbb0a6465),
	.w6(32'h3ac02a82),
	.w7(32'h3b9729a2),
	.w8(32'hbb6d716e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a0508),
	.w1(32'hbb9a143e),
	.w2(32'h3aa6ecf1),
	.w3(32'hbadfa4f2),
	.w4(32'h3b6f37a2),
	.w5(32'hbbdccd56),
	.w6(32'hbbbf3ee3),
	.w7(32'h3b5c3803),
	.w8(32'hbc06a6d0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55dc80),
	.w1(32'hbc97df30),
	.w2(32'hbc5b5dfd),
	.w3(32'hbc916619),
	.w4(32'hbc74d02a),
	.w5(32'hbc79ac15),
	.w6(32'hbc1f8262),
	.w7(32'hbbbeeeae),
	.w8(32'hbba862b4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb298123),
	.w1(32'hbbb2d225),
	.w2(32'hbc12ffd2),
	.w3(32'hbbf3bbfd),
	.w4(32'hbc76520f),
	.w5(32'h3a2abf9d),
	.w6(32'h3b4e155b),
	.w7(32'h3c294068),
	.w8(32'h3c7158d4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb5421),
	.w1(32'hbb4ca6d9),
	.w2(32'hbc3753f7),
	.w3(32'hba68b148),
	.w4(32'hb9bb946c),
	.w5(32'h3ba3f5c1),
	.w6(32'h3a312bc9),
	.w7(32'hbc9cdd0e),
	.w8(32'hbc0d5f78),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc023304),
	.w1(32'h3c747957),
	.w2(32'h3a0f1921),
	.w3(32'h3c8ae1cd),
	.w4(32'hbba1c28b),
	.w5(32'hbb12334b),
	.w6(32'h3be3e949),
	.w7(32'hbb42f10e),
	.w8(32'hbb9f33b8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b88f7),
	.w1(32'h3b34c600),
	.w2(32'h3bcc074f),
	.w3(32'h3c3a74af),
	.w4(32'h3c116e7b),
	.w5(32'h3c72dc4c),
	.w6(32'h3c8fd420),
	.w7(32'h3cc26a13),
	.w8(32'h3cd628da),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a64fa8),
	.w1(32'h3bae58c6),
	.w2(32'h3c393f4e),
	.w3(32'hbb5e9383),
	.w4(32'h3bfa8752),
	.w5(32'h3c5eb2c9),
	.w6(32'h3b8fc6cb),
	.w7(32'h3c7741dc),
	.w8(32'h3c8b5c0f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07c1ce),
	.w1(32'hb8b199cb),
	.w2(32'hbbcf3171),
	.w3(32'hbb194fc1),
	.w4(32'hbaf010eb),
	.w5(32'hbc18ebed),
	.w6(32'hbb3841bc),
	.w7(32'hbc7d9733),
	.w8(32'hbcae2586),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59f63c),
	.w1(32'h3b917607),
	.w2(32'h3b1c45d0),
	.w3(32'h3c1b90f5),
	.w4(32'hbb7fd65c),
	.w5(32'h398993c3),
	.w6(32'h3be61d88),
	.w7(32'h3b1941fb),
	.w8(32'hbb3f45b2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdcc3b),
	.w1(32'h3cb0f82c),
	.w2(32'hbb7014b9),
	.w3(32'h3c49c597),
	.w4(32'hbb010d76),
	.w5(32'hba931190),
	.w6(32'h3b53cf66),
	.w7(32'hbbf5e44d),
	.w8(32'hbc3df90f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9627bb),
	.w1(32'hbbbe8a2f),
	.w2(32'h3bdc0974),
	.w3(32'hbc25735b),
	.w4(32'hbd36fe7b),
	.w5(32'hbd789372),
	.w6(32'hbd5ddfb7),
	.w7(32'hbceb882b),
	.w8(32'hbca26b89),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc707991),
	.w1(32'hbc3b901c),
	.w2(32'h3ab0e3bb),
	.w3(32'hbc0899d8),
	.w4(32'hbb3551c2),
	.w5(32'hba98c49f),
	.w6(32'hba77464b),
	.w7(32'h3beb009a),
	.w8(32'h3c0bbd20),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba98ce9),
	.w1(32'hbb066b21),
	.w2(32'hbb9fb8a6),
	.w3(32'hbbcfaf9b),
	.w4(32'h3c53a7f3),
	.w5(32'h3cbd43ad),
	.w6(32'h3abfbcd2),
	.w7(32'h3ca486d2),
	.w8(32'h3c5c8753),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94932b),
	.w1(32'hbd08a746),
	.w2(32'h3b64132b),
	.w3(32'hbb4b0912),
	.w4(32'h3b296561),
	.w5(32'h3b9f8488),
	.w6(32'hbc2b7bcf),
	.w7(32'h3aca88b6),
	.w8(32'h3bb0ff5f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fe92a),
	.w1(32'h3b6a0a41),
	.w2(32'hbaa347e9),
	.w3(32'h3c0652fb),
	.w4(32'hbc116f91),
	.w5(32'h3b2a1fce),
	.w6(32'h3c19a231),
	.w7(32'hbbd4a904),
	.w8(32'h3c9f4df2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92dbbb),
	.w1(32'hbb966f70),
	.w2(32'hbbbe7ee9),
	.w3(32'h3b718caa),
	.w4(32'h3c99c504),
	.w5(32'h3d08980e),
	.w6(32'h3c35da13),
	.w7(32'h3c7bf950),
	.w8(32'h3ce746dd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1a2d3),
	.w1(32'h3b6ef46b),
	.w2(32'hbb1475d1),
	.w3(32'h39e2fbae),
	.w4(32'h3b81b35e),
	.w5(32'hbc01978c),
	.w6(32'h3c13148c),
	.w7(32'h3bd8293a),
	.w8(32'hbc2926dd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc81847),
	.w1(32'h3c2113e1),
	.w2(32'h3c7f83af),
	.w3(32'hbb54d227),
	.w4(32'h3c04ac42),
	.w5(32'h3c627e76),
	.w6(32'hbb12bf1a),
	.w7(32'h3c3e2ee8),
	.w8(32'h3c8618c0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dc2ce),
	.w1(32'hb99acc0e),
	.w2(32'h3b03938d),
	.w3(32'h3b574e40),
	.w4(32'h3c00292f),
	.w5(32'h3c94a868),
	.w6(32'h3b436ae2),
	.w7(32'h3c1f3ca7),
	.w8(32'h3c7f1870),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd5bd1),
	.w1(32'h3bd8178e),
	.w2(32'hbc08a893),
	.w3(32'h3c0764b5),
	.w4(32'h3aed5de4),
	.w5(32'h3bd5fd27),
	.w6(32'h3ca45db5),
	.w7(32'hbc0f850d),
	.w8(32'h38133bfa),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac77bde),
	.w1(32'h3b5d1607),
	.w2(32'h3c8c8ce4),
	.w3(32'h3c394843),
	.w4(32'h3c21c47e),
	.w5(32'h3bc2792c),
	.w6(32'h3bb56f1f),
	.w7(32'h3c870011),
	.w8(32'h3c4660ed),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd7278),
	.w1(32'h3b1b69be),
	.w2(32'hba7045ef),
	.w3(32'h3ba21053),
	.w4(32'h3a1289f8),
	.w5(32'hbbb1252b),
	.w6(32'h3babae04),
	.w7(32'hbb158c7e),
	.w8(32'h38ebbed1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ece02),
	.w1(32'hb9a0656e),
	.w2(32'h3baef490),
	.w3(32'hbb2fc9ce),
	.w4(32'h3b37493d),
	.w5(32'h3b79c5b3),
	.w6(32'h3ad1aee1),
	.w7(32'h3aedf8ce),
	.w8(32'h3b57bd51),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b3a15),
	.w1(32'h3c42a460),
	.w2(32'h3bd6e1af),
	.w3(32'h3bb7ea40),
	.w4(32'hb9578828),
	.w5(32'h3be3be3c),
	.w6(32'h3b2b6810),
	.w7(32'h3c055bf1),
	.w8(32'h3c55865c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd7421),
	.w1(32'h3ac3452f),
	.w2(32'hbb251d0b),
	.w3(32'h398d3746),
	.w4(32'h3ba83c1b),
	.w5(32'h3c20d44b),
	.w6(32'hbb2f092c),
	.w7(32'hbc00c86e),
	.w8(32'hbad3d7b7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02be8e),
	.w1(32'h3b8e8102),
	.w2(32'h3b5ba3e2),
	.w3(32'h3b771544),
	.w4(32'h3bbfe1e5),
	.w5(32'h3c8f6fe6),
	.w6(32'hbb39c287),
	.w7(32'h3cbe16e9),
	.w8(32'h3d09b71b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a1f9e),
	.w1(32'hbbf01419),
	.w2(32'hbafb26ec),
	.w3(32'hbaa78103),
	.w4(32'hb91e941e),
	.w5(32'h3a824e0b),
	.w6(32'h3c481df8),
	.w7(32'h3b945bcc),
	.w8(32'h3c5719d7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b148396),
	.w1(32'hbbc01f1b),
	.w2(32'hbad48c04),
	.w3(32'hbb866fa1),
	.w4(32'hbb9737bf),
	.w5(32'hbc57d635),
	.w6(32'h3bc1dc48),
	.w7(32'hbb1f3f0c),
	.w8(32'hbc3e5631),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44b157),
	.w1(32'hbba81b78),
	.w2(32'hb9c3ab19),
	.w3(32'hbab11651),
	.w4(32'hbb28fcc0),
	.w5(32'h3ca16af2),
	.w6(32'hbbaba6ad),
	.w7(32'h3bd55699),
	.w8(32'h3ce99510),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92dc34),
	.w1(32'hbb974194),
	.w2(32'hbb414a4d),
	.w3(32'h3b974b89),
	.w4(32'hbbd60e43),
	.w5(32'h3bb3b871),
	.w6(32'h3bbf7a94),
	.w7(32'hba49ace1),
	.w8(32'h3bce48fd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa6023),
	.w1(32'h3b5b83c8),
	.w2(32'h3b1ab18e),
	.w3(32'h3c2266b5),
	.w4(32'h3b5f4420),
	.w5(32'h3c091439),
	.w6(32'h3c283c17),
	.w7(32'h3c8370d8),
	.w8(32'h3c6f4097),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a3d47),
	.w1(32'hbbae2a10),
	.w2(32'hbc8e97d3),
	.w3(32'h3b947761),
	.w4(32'hbbd935df),
	.w5(32'hbc2a5239),
	.w6(32'h3b1f808e),
	.w7(32'hbca6e4ed),
	.w8(32'hbcb358b6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc307167),
	.w1(32'hbbd608c8),
	.w2(32'hbc8395b5),
	.w3(32'hbc2884d6),
	.w4(32'hbc673163),
	.w5(32'hbcc54dd3),
	.w6(32'hbc6849c3),
	.w7(32'hbc94b9c9),
	.w8(32'hbccf5c80),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24e0a5),
	.w1(32'h396628a4),
	.w2(32'hba886be9),
	.w3(32'hb9f5d78f),
	.w4(32'h3c02a5cb),
	.w5(32'h3c245ef4),
	.w6(32'hbbdb7017),
	.w7(32'h3bb4971e),
	.w8(32'h3c32ce8f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48e025),
	.w1(32'hbb2bec29),
	.w2(32'hbbf0443a),
	.w3(32'hbcbc7258),
	.w4(32'hbc0bc2cc),
	.w5(32'hbbf64d91),
	.w6(32'hbbf95593),
	.w7(32'hbbafb36a),
	.w8(32'hbb8c0b7e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb951573),
	.w1(32'hbc005641),
	.w2(32'hba5e018c),
	.w3(32'hbbd7fe44),
	.w4(32'h3a7f38bd),
	.w5(32'hbbe6b06b),
	.w6(32'hbae2644b),
	.w7(32'h3bbff751),
	.w8(32'h3c15791f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe7840),
	.w1(32'hbc4efe0e),
	.w2(32'hbb27c5a8),
	.w3(32'hbc657824),
	.w4(32'hbb01b783),
	.w5(32'hbadb3477),
	.w6(32'hbb8485f2),
	.w7(32'h3ba26b19),
	.w8(32'h3bf0d38e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c0458),
	.w1(32'hbacf60d9),
	.w2(32'hbbcc1814),
	.w3(32'hb9a5366a),
	.w4(32'h3ba3e3eb),
	.w5(32'h3a92a85f),
	.w6(32'h3b56c4e1),
	.w7(32'h3a3cb961),
	.w8(32'hbb8d41fb),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc451ff4),
	.w1(32'hbc4f5c92),
	.w2(32'hba27faff),
	.w3(32'hb9008e80),
	.w4(32'hbc054819),
	.w5(32'hbbd95686),
	.w6(32'hbc37325b),
	.w7(32'h3bfd882e),
	.w8(32'h3bcbb20f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb224ae0),
	.w1(32'h3ace6542),
	.w2(32'h3bc26b23),
	.w3(32'hbb51d8a2),
	.w4(32'h3af7c13a),
	.w5(32'h3aa773e0),
	.w6(32'h3b88ddd0),
	.w7(32'h3ba1bb1d),
	.w8(32'h3b8c98eb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11ebcf),
	.w1(32'h3c2db355),
	.w2(32'h3b768137),
	.w3(32'h3baf4001),
	.w4(32'hbc277265),
	.w5(32'hbbd2fb4b),
	.w6(32'h3bbb3b68),
	.w7(32'h3b4b1746),
	.w8(32'h39ff46f1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc292cbf),
	.w1(32'hbb4510cc),
	.w2(32'hbb137f01),
	.w3(32'hbb53c3c2),
	.w4(32'h3a3fef25),
	.w5(32'h3a50eb3b),
	.w6(32'h3b931b90),
	.w7(32'h3b8566a9),
	.w8(32'h3c122975),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bada634),
	.w1(32'hba21b522),
	.w2(32'h3acf4220),
	.w3(32'h39ea6410),
	.w4(32'hbd263cb8),
	.w5(32'hbc7b8b47),
	.w6(32'h3bc06c36),
	.w7(32'hbcdc8bce),
	.w8(32'h3c1c2446),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8dd1e),
	.w1(32'h3cec797d),
	.w2(32'h3bed95e7),
	.w3(32'hbb28705c),
	.w4(32'hbc395265),
	.w5(32'hbba1c769),
	.w6(32'h3c5e2579),
	.w7(32'h3bb6ba3a),
	.w8(32'h3bf42bbc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be48136),
	.w1(32'h3ab4bd77),
	.w2(32'h3c09be9c),
	.w3(32'hbc40af21),
	.w4(32'h3bca09ec),
	.w5(32'h39e8094c),
	.w6(32'h3b48a70f),
	.w7(32'h3b3c3074),
	.w8(32'hbbf6609b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967bf6),
	.w1(32'h3bc9723c),
	.w2(32'h3b9926a0),
	.w3(32'h3b08e63c),
	.w4(32'hbb4fdf51),
	.w5(32'hbabc9276),
	.w6(32'h3950f095),
	.w7(32'h3bd0d15a),
	.w8(32'h3c3135be),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb23ce),
	.w1(32'hba369cd8),
	.w2(32'hbb0de07c),
	.w3(32'hbbfa1378),
	.w4(32'hb7112523),
	.w5(32'h3a69e2eb),
	.w6(32'hba300eb4),
	.w7(32'h3b73c60e),
	.w8(32'h3c2d837a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08a34d),
	.w1(32'hbb8cca59),
	.w2(32'h3c2aefab),
	.w3(32'h38013869),
	.w4(32'h3b44ba78),
	.w5(32'h3bd7b4e5),
	.w6(32'h3c08a9fb),
	.w7(32'hbab2675a),
	.w8(32'h3b626eef),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1464c0),
	.w1(32'h3c15b7d0),
	.w2(32'h3c2eb459),
	.w3(32'h3bb01b91),
	.w4(32'h3c68e07d),
	.w5(32'hbb0d4b5d),
	.w6(32'h3af1e297),
	.w7(32'h3c981597),
	.w8(32'hbaa4ce37),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe59632),
	.w1(32'h3c34c28c),
	.w2(32'hbb15828c),
	.w3(32'h3c09d203),
	.w4(32'h3bad5f53),
	.w5(32'h3af6746a),
	.w6(32'h3c38df07),
	.w7(32'h3bb2a1c1),
	.w8(32'h3b97bea2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95e155),
	.w1(32'hbbf09cae),
	.w2(32'hbbb53970),
	.w3(32'hbbd91878),
	.w4(32'h3b15c1aa),
	.w5(32'h3c61df56),
	.w6(32'hbba64e3f),
	.w7(32'hbbdfb1ac),
	.w8(32'h3c7f8444),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd30739),
	.w1(32'hbbbc7994),
	.w2(32'hbbda8c16),
	.w3(32'hbc041b0b),
	.w4(32'hbc02538d),
	.w5(32'hbc573161),
	.w6(32'hb9fd8986),
	.w7(32'hbc5cdd95),
	.w8(32'hbb620851),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcac738),
	.w1(32'hbbf36d87),
	.w2(32'hbb6e289c),
	.w3(32'hbc2beb48),
	.w4(32'hba8726ff),
	.w5(32'h3a9ab71b),
	.w6(32'hbc001bb8),
	.w7(32'hbac2edcf),
	.w8(32'hbaae16b0),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94087c),
	.w1(32'hbbfbd011),
	.w2(32'hbbecd5bb),
	.w3(32'hbc049e02),
	.w4(32'hbbc0ce5d),
	.w5(32'hbc0676e9),
	.w6(32'hbb77a6e3),
	.w7(32'hbc1cb8d2),
	.w8(32'hbbc88229),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb609d52),
	.w1(32'hbb670ba7),
	.w2(32'hbc54138e),
	.w3(32'hbc813791),
	.w4(32'hbac02b34),
	.w5(32'hbbd3329a),
	.w6(32'hbb8d87a4),
	.w7(32'hba9b6231),
	.w8(32'hbc3e71a6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fde76),
	.w1(32'hbb24c592),
	.w2(32'hbb3d11c9),
	.w3(32'hbb31e2c1),
	.w4(32'h39696d50),
	.w5(32'h3b562d8f),
	.w6(32'hbb896b78),
	.w7(32'hbc889a52),
	.w8(32'hbbffa168),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6a2b4),
	.w1(32'hbc1109b9),
	.w2(32'hbc47aa1a),
	.w3(32'h3acb97ef),
	.w4(32'h3b4cbc2f),
	.w5(32'h3a955594),
	.w6(32'hbb491979),
	.w7(32'h3b11047b),
	.w8(32'h3c922f5a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e5615),
	.w1(32'hbc52f160),
	.w2(32'hbbaf9d4c),
	.w3(32'hbc4f9687),
	.w4(32'hbb552db9),
	.w5(32'h3a7fbe2a),
	.w6(32'hbbb05e6f),
	.w7(32'hbbc2548a),
	.w8(32'hbb663127),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb226f6),
	.w1(32'hbb2818f9),
	.w2(32'hbbcf9fe9),
	.w3(32'h3b452fb0),
	.w4(32'hbb11e097),
	.w5(32'hbbc1d668),
	.w6(32'hbb899267),
	.w7(32'hbb7e10c7),
	.w8(32'hbbf2b47f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26e885),
	.w1(32'hbb8bd386),
	.w2(32'h3ad7b032),
	.w3(32'hba3da223),
	.w4(32'h3a802505),
	.w5(32'hbb37edb5),
	.w6(32'hb91a0331),
	.w7(32'h3b232405),
	.w8(32'h3be43a48),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb73b7b),
	.w1(32'h3b2fa440),
	.w2(32'h3a95a1ea),
	.w3(32'hba462aa7),
	.w4(32'hbad0d9d2),
	.w5(32'hbb9334c3),
	.w6(32'h399a01ab),
	.w7(32'h3b4a736e),
	.w8(32'h3b066eca),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae104c),
	.w1(32'hbb0c49d7),
	.w2(32'h3b9ed574),
	.w3(32'h3988963f),
	.w4(32'h39854de5),
	.w5(32'h3b33cd40),
	.w6(32'h3afa59e6),
	.w7(32'h3bdb896b),
	.w8(32'h3bcf394c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b180296),
	.w1(32'hba9cbded),
	.w2(32'hbbef70a7),
	.w3(32'h3b981e61),
	.w4(32'h3b830155),
	.w5(32'h3b09bafc),
	.w6(32'h3b30dcbe),
	.w7(32'hb9d03308),
	.w8(32'h3ccd9bbb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b6fec),
	.w1(32'hbb4e1e8a),
	.w2(32'h3bf1789e),
	.w3(32'hbbd6f788),
	.w4(32'hba0a535c),
	.w5(32'h3a625093),
	.w6(32'h3c483acc),
	.w7(32'hbbd5740a),
	.w8(32'h3a1a8bca),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dd4c7),
	.w1(32'h3b35df88),
	.w2(32'hbac2f629),
	.w3(32'hb9c6343a),
	.w4(32'hbc515bcf),
	.w5(32'hbcb7062d),
	.w6(32'h3a414c87),
	.w7(32'hbbf31428),
	.w8(32'hbca7cbc8),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73ae47),
	.w1(32'h3c3e08aa),
	.w2(32'hbb2d3630),
	.w3(32'hbc05ba79),
	.w4(32'h3a9877ff),
	.w5(32'h3bc59158),
	.w6(32'h3ae6226a),
	.w7(32'hbb6710a5),
	.w8(32'h3b7a6624),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fddd1),
	.w1(32'hbb3d124e),
	.w2(32'h3ad55bbf),
	.w3(32'h3a251c8b),
	.w4(32'hbb2c5b7d),
	.w5(32'hbc1a84c4),
	.w6(32'h3b5e80e6),
	.w7(32'h3cc574f5),
	.w8(32'h3b53a4bd),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c154e02),
	.w1(32'h3b9335c6),
	.w2(32'h3b549980),
	.w3(32'h3c2c26ce),
	.w4(32'h3bd46a3b),
	.w5(32'h3ce21809),
	.w6(32'hbcc58ef0),
	.w7(32'hbc86bbe5),
	.w8(32'h3bed64af),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c0dee),
	.w1(32'h3c2d29a1),
	.w2(32'hbb61a39c),
	.w3(32'h3cb204c0),
	.w4(32'hbc550425),
	.w5(32'hbc8add12),
	.w6(32'hbb281646),
	.w7(32'h3b65f106),
	.w8(32'hbc55aeb4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13113f),
	.w1(32'hbb96b284),
	.w2(32'hbbeda4b8),
	.w3(32'hbc942e58),
	.w4(32'hbb33eeac),
	.w5(32'h3bc27a5c),
	.w6(32'hbb2d0373),
	.w7(32'hbbd59fb4),
	.w8(32'h3baf7058),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafb800),
	.w1(32'h3bf120de),
	.w2(32'h3b8c6d1a),
	.w3(32'h3bdbf8b9),
	.w4(32'hbb4f5150),
	.w5(32'hbc074ac8),
	.w6(32'hbba098bd),
	.w7(32'h3aeec0cc),
	.w8(32'hbb870339),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba706e7c),
	.w1(32'hbb8b9d42),
	.w2(32'h3ba0b094),
	.w3(32'hbb129227),
	.w4(32'h3b3a0273),
	.w5(32'h3b8c0f43),
	.w6(32'hbadbf256),
	.w7(32'hbb792c75),
	.w8(32'hbb85f355),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be29cd6),
	.w1(32'h3b8dfe89),
	.w2(32'h3c9062fb),
	.w3(32'h3b35691b),
	.w4(32'hbba286f6),
	.w5(32'h3c80e7b1),
	.w6(32'hba2a887d),
	.w7(32'hbc847e8a),
	.w8(32'hbd2d82ed),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b8682),
	.w1(32'hbc617f4b),
	.w2(32'hbbeffc5e),
	.w3(32'h3c35ec90),
	.w4(32'hbb930629),
	.w5(32'hbc681033),
	.w6(32'hbd155033),
	.w7(32'h3c84e3dc),
	.w8(32'h3ba5603e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89b26c),
	.w1(32'h3a90d501),
	.w2(32'hbc810116),
	.w3(32'h3cb0a74b),
	.w4(32'h3b6eef43),
	.w5(32'h3ce507ca),
	.w6(32'h3ba456a3),
	.w7(32'h3c3af3f3),
	.w8(32'h3c9e6eb3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc0a98),
	.w1(32'hbb7b6c3a),
	.w2(32'h3b9ba61f),
	.w3(32'h3c8fed8e),
	.w4(32'h3c3af9de),
	.w5(32'hbac1447c),
	.w6(32'hbbb9ea88),
	.w7(32'hbbf11a68),
	.w8(32'hbc8a6168),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6399b8),
	.w1(32'hbbb44e35),
	.w2(32'hbb3aa0d8),
	.w3(32'h3c3360b7),
	.w4(32'hbb90f0ec),
	.w5(32'hbc8c10dd),
	.w6(32'hbb75d129),
	.w7(32'h3d045773),
	.w8(32'h3cf0c7c7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c170bb2),
	.w1(32'h3a43e09a),
	.w2(32'h3b4dd1d4),
	.w3(32'hbcfacf8c),
	.w4(32'h3b507a48),
	.w5(32'h3b90398e),
	.w6(32'hbc556889),
	.w7(32'h3c055860),
	.w8(32'h3c0d6ad0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb114588),
	.w1(32'hbb63e0b7),
	.w2(32'hbc770b8b),
	.w3(32'hbb1388bf),
	.w4(32'h3aabac58),
	.w5(32'h3c0bc311),
	.w6(32'h390ebfa9),
	.w7(32'h3c220d2c),
	.w8(32'h3d34888a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d9193),
	.w1(32'h3c444ea7),
	.w2(32'h3b8525b3),
	.w3(32'hbc3c31b7),
	.w4(32'h3c27f39f),
	.w5(32'hbbab32c4),
	.w6(32'h3ca3fcd1),
	.w7(32'h3cf636fe),
	.w8(32'h3b11c2fd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60e5c2),
	.w1(32'hbbdee257),
	.w2(32'h3c360de3),
	.w3(32'hbb924175),
	.w4(32'h3be422da),
	.w5(32'h3c4f9dd3),
	.w6(32'hbc2a867d),
	.w7(32'hbc35806c),
	.w8(32'hbc531ec9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8663cd),
	.w1(32'h378c3c56),
	.w2(32'h3b7e94dd),
	.w3(32'h3bb7b14a),
	.w4(32'h3c400eee),
	.w5(32'h3c516e21),
	.w6(32'h3b5acbb0),
	.w7(32'h3b9f6512),
	.w8(32'h3c086632),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be54b18),
	.w1(32'h3bbfeefa),
	.w2(32'hba0f29cd),
	.w3(32'h3c235c13),
	.w4(32'hbc2e3b35),
	.w5(32'hbb13092c),
	.w6(32'h3be99ed8),
	.w7(32'h3c1e8149),
	.w8(32'hba8f9ab5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc3359),
	.w1(32'h3c0249b1),
	.w2(32'hbc265550),
	.w3(32'hbba6fd55),
	.w4(32'hbc23f54c),
	.w5(32'hbc46e543),
	.w6(32'h3bc5df99),
	.w7(32'hbc0b97bc),
	.w8(32'h3c202af7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca91c7c),
	.w1(32'hbc8c2b9e),
	.w2(32'hbb7e4917),
	.w3(32'hbc29086d),
	.w4(32'h3b9a0c1b),
	.w5(32'h3ba89d38),
	.w6(32'h3c796cec),
	.w7(32'hbc227b1c),
	.w8(32'hbbcdea15),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cdce0),
	.w1(32'h3b373b5b),
	.w2(32'hbbc9f5a8),
	.w3(32'hbb67876b),
	.w4(32'h3b003a71),
	.w5(32'hbba3e340),
	.w6(32'hbb8e1931),
	.w7(32'hbc59b9a3),
	.w8(32'hbc76aad5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb99dbf),
	.w1(32'hbc0c1998),
	.w2(32'h3b2ff40e),
	.w3(32'hbb3b1b8a),
	.w4(32'hb9c6bda4),
	.w5(32'hbbd3e5ed),
	.w6(32'hbc303cf6),
	.w7(32'h3b2fd514),
	.w8(32'hba80c3c0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae663ca),
	.w1(32'h3b8a1f74),
	.w2(32'hbbd7e77d),
	.w3(32'hbc03089b),
	.w4(32'h3aff72e3),
	.w5(32'hbc252df7),
	.w6(32'hbbad4044),
	.w7(32'h39b3587e),
	.w8(32'h3b5422d6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85ca42),
	.w1(32'hbc0cec9d),
	.w2(32'hbbe36228),
	.w3(32'hbc5d161e),
	.w4(32'hbcb4fd87),
	.w5(32'h3c063784),
	.w6(32'hbc2ae17d),
	.w7(32'h3c68d093),
	.w8(32'hbc135c4d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97a074),
	.w1(32'hbc11304a),
	.w2(32'hbc85619f),
	.w3(32'h3d0ba190),
	.w4(32'h3ca4df1a),
	.w5(32'h3c1951aa),
	.w6(32'hbc6d996a),
	.w7(32'hbbbe16dc),
	.w8(32'h3cc1bebf),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2c213),
	.w1(32'h3b6fb421),
	.w2(32'h3b9ec901),
	.w3(32'hbc26d4cf),
	.w4(32'h3b6b261d),
	.w5(32'h390c9fa5),
	.w6(32'h3ca33302),
	.w7(32'h3c26bdf7),
	.w8(32'h3c274884),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6b909),
	.w1(32'h3b96f1af),
	.w2(32'h3b7f7d26),
	.w3(32'h3b0e9f1c),
	.w4(32'h399cb365),
	.w5(32'hbb288f9f),
	.w6(32'h3b43b3af),
	.w7(32'hbb8697d7),
	.w8(32'hbbaa0d08),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e0164),
	.w1(32'h38929045),
	.w2(32'hbc72151b),
	.w3(32'h3c621d96),
	.w4(32'hbc0c3fb1),
	.w5(32'hbbe0847f),
	.w6(32'h3baeb696),
	.w7(32'h3c84737a),
	.w8(32'h3c8e9f6e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef2b31),
	.w1(32'h3c1532b8),
	.w2(32'h3c2f0c21),
	.w3(32'hbc919da8),
	.w4(32'hba287ed5),
	.w5(32'hba552c89),
	.w6(32'h3c7e61c2),
	.w7(32'hbbc498e2),
	.w8(32'hbc9cb87b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b797d8b),
	.w1(32'h3bd16b0d),
	.w2(32'h3bd058d1),
	.w3(32'hba5d0193),
	.w4(32'hbb390a65),
	.w5(32'hbb8fabf4),
	.w6(32'hbbb578e1),
	.w7(32'h3a5449cb),
	.w8(32'hbadfa671),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19ce45),
	.w1(32'hbb59d7e4),
	.w2(32'h3c3e2bab),
	.w3(32'hbb8b7f43),
	.w4(32'hbc54cf8a),
	.w5(32'hbcbd99db),
	.w6(32'h3a72cf58),
	.w7(32'h3c1e4976),
	.w8(32'hbc89c4d3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ed471),
	.w1(32'hbbd421c7),
	.w2(32'hbbf5feb9),
	.w3(32'hbbf62773),
	.w4(32'hbc917d7f),
	.w5(32'hbcb9c769),
	.w6(32'hbc91769b),
	.w7(32'hbc35b3fb),
	.w8(32'hbc79b070),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc301884),
	.w1(32'hbc2b1fb2),
	.w2(32'hbb080629),
	.w3(32'hbc426710),
	.w4(32'hbc23f8e5),
	.w5(32'h3c33514d),
	.w6(32'hbbe60436),
	.w7(32'hbc8980d1),
	.w8(32'hbcd9f972),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b831593),
	.w1(32'hbb19f5a3),
	.w2(32'hbb9c83d3),
	.w3(32'h3a1dbe75),
	.w4(32'h3bf06fb7),
	.w5(32'h3bda866a),
	.w6(32'hbc957dfc),
	.w7(32'hbc11be40),
	.w8(32'hbb9f989c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b001fca),
	.w1(32'h3a680d7f),
	.w2(32'h3b38b75d),
	.w3(32'h3bc7b9b9),
	.w4(32'h398c5cd5),
	.w5(32'h3a1b674e),
	.w6(32'hb8b6ed0f),
	.w7(32'h3b861955),
	.w8(32'hbc6251e3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6cc75),
	.w1(32'h3be677b0),
	.w2(32'h3b34b530),
	.w3(32'hbb7848c7),
	.w4(32'hbae13929),
	.w5(32'hbb57d287),
	.w6(32'hbbe3756a),
	.w7(32'h3bcf8db6),
	.w8(32'h3bcbfb27),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944a3dd),
	.w1(32'hbabd325f),
	.w2(32'hbc06b6cb),
	.w3(32'h3ad091c6),
	.w4(32'hbbcc1678),
	.w5(32'hbb3377b4),
	.w6(32'h3b8464fe),
	.w7(32'hbb87ab9e),
	.w8(32'hbc6d31cd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac9183),
	.w1(32'hbbc1449b),
	.w2(32'hbae82072),
	.w3(32'h3bb3d863),
	.w4(32'hbc16a4fc),
	.w5(32'hbc6569cb),
	.w6(32'hba35cd84),
	.w7(32'hbbe22041),
	.w8(32'hbbf28ef8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390215d1),
	.w1(32'hbb8ade68),
	.w2(32'h3a971ead),
	.w3(32'hbb836e15),
	.w4(32'h3b1fb00d),
	.w5(32'h3c04e0a2),
	.w6(32'h3a5a6884),
	.w7(32'h3bbcc6d6),
	.w8(32'h3ba56bed),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3327c3),
	.w1(32'h3a88be12),
	.w2(32'hb94f8c7c),
	.w3(32'h3c1b27a3),
	.w4(32'h3c18f8f8),
	.w5(32'h3c3d9f07),
	.w6(32'hbb022d88),
	.w7(32'h3b1bca55),
	.w8(32'h3c88071c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b389ce6),
	.w1(32'h3bde32cf),
	.w2(32'h39c590b6),
	.w3(32'h3ae78b36),
	.w4(32'hb9ded04a),
	.w5(32'hbb3e6bc8),
	.w6(32'h3a965392),
	.w7(32'h3b923403),
	.w8(32'h3b887828),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba56a00),
	.w1(32'h3abcd40e),
	.w2(32'h3bc2e1be),
	.w3(32'h3b6061e3),
	.w4(32'h3ba03745),
	.w5(32'h3d25b8e9),
	.w6(32'h3b2fe12c),
	.w7(32'hbd6407c6),
	.w8(32'hbcbeaf38),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec4d5d),
	.w1(32'h3a300172),
	.w2(32'hb991a1de),
	.w3(32'h3cca920f),
	.w4(32'h391c7434),
	.w5(32'h3c8de2e8),
	.w6(32'h3c3b9593),
	.w7(32'hbbad30aa),
	.w8(32'hbc923909),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8a04f),
	.w1(32'h3c49725f),
	.w2(32'hbb59712c),
	.w3(32'h3cc006a9),
	.w4(32'hba02b62c),
	.w5(32'h3ae2e174),
	.w6(32'hbbeb0ab8),
	.w7(32'hbb88caaa),
	.w8(32'hbaddc4c1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7a3b9),
	.w1(32'hbb08c0d2),
	.w2(32'h3bd7f57a),
	.w3(32'h3b226e6a),
	.w4(32'h3bdf9f89),
	.w5(32'hbba9441f),
	.w6(32'h3ad8bfdb),
	.w7(32'hba95107d),
	.w8(32'hbb32620e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf97ba),
	.w1(32'h3acd3dd7),
	.w2(32'h3981fdba),
	.w3(32'hbc4690b8),
	.w4(32'h3bf3de6d),
	.w5(32'hbb0a2123),
	.w6(32'hbb311ba3),
	.w7(32'h3a2e74d6),
	.w8(32'hbc0f19ee),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule