module layer_10_featuremap_197(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f384ea),
	.w1(32'hb98c4eeb),
	.w2(32'h3a5d454b),
	.w3(32'h392ba35b),
	.w4(32'h38a4a77e),
	.w5(32'h36d03d69),
	.w6(32'hb9e78949),
	.w7(32'h38d759ff),
	.w8(32'hba766415),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fd3f2),
	.w1(32'h3b9659bf),
	.w2(32'h3b3b74d5),
	.w3(32'h3bc4263a),
	.w4(32'h3b0488e9),
	.w5(32'h3ad51aa0),
	.w6(32'h3af0117e),
	.w7(32'hbb52f54c),
	.w8(32'hbb79a812),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6a635),
	.w1(32'h3a91ad5f),
	.w2(32'h3a85f528),
	.w3(32'h381a079f),
	.w4(32'h3a2de73e),
	.w5(32'h39f1def7),
	.w6(32'h39e8534d),
	.w7(32'h39a57175),
	.w8(32'h3951cebe),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5fc2e),
	.w1(32'h3a136ac4),
	.w2(32'hb99f5a4d),
	.w3(32'h39c2f641),
	.w4(32'hbb1179c9),
	.w5(32'hbaf8c86c),
	.w6(32'h3a48b6b5),
	.w7(32'h39cea30b),
	.w8(32'hb932a90d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1615b0),
	.w1(32'hba35804f),
	.w2(32'hba4f8840),
	.w3(32'hba6d6db6),
	.w4(32'hb9d4f829),
	.w5(32'hba253e76),
	.w6(32'h3a34ff12),
	.w7(32'h3b02ee3f),
	.w8(32'h3af302e4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999f692),
	.w1(32'h3a1e2c8a),
	.w2(32'h3a83823b),
	.w3(32'hba161369),
	.w4(32'h3a04c9a8),
	.w5(32'h3a3af178),
	.w6(32'h3a621a41),
	.w7(32'h3a2bfb35),
	.w8(32'h39c69830),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98bf77),
	.w1(32'hba6554c5),
	.w2(32'h3b9b0531),
	.w3(32'hbb534709),
	.w4(32'hbafa1947),
	.w5(32'hbba32d16),
	.w6(32'hbbb92ef1),
	.w7(32'hbafc072a),
	.w8(32'hbb8b53c3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56fedc),
	.w1(32'hbad92bc7),
	.w2(32'hbc344d30),
	.w3(32'hbc8cd3fe),
	.w4(32'hbbc71b63),
	.w5(32'hbbbdc926),
	.w6(32'h3bb05f98),
	.w7(32'h39c12566),
	.w8(32'h3c073bf2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a014035),
	.w1(32'h38fa7082),
	.w2(32'hba18f8d4),
	.w3(32'h3aa6c18d),
	.w4(32'h3a7deb9f),
	.w5(32'h3956e0c0),
	.w6(32'h3a441548),
	.w7(32'h3a2b3fee),
	.w8(32'h39d5ee29),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf26516),
	.w1(32'hbb011e0a),
	.w2(32'hbb2127b3),
	.w3(32'hbbe83812),
	.w4(32'hbb4515b7),
	.w5(32'hbbb0f073),
	.w6(32'hbb4339a0),
	.w7(32'hbabc10fe),
	.w8(32'hbb64fe79),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d15cf6),
	.w1(32'hbadf841e),
	.w2(32'hbb169dd9),
	.w3(32'hba203180),
	.w4(32'hba5a9ada),
	.w5(32'hb96296fd),
	.w6(32'hbaa1997c),
	.w7(32'hbaa89542),
	.w8(32'hbb0c7598),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc477e),
	.w1(32'h3a93bb6f),
	.w2(32'h3c206dbb),
	.w3(32'hb949a19e),
	.w4(32'h3b5754af),
	.w5(32'h3a474761),
	.w6(32'h3abb2fcc),
	.w7(32'h3b30c3f2),
	.w8(32'h3bf94d99),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76a277),
	.w1(32'hbc12126f),
	.w2(32'hbbaf09dc),
	.w3(32'hbc1a927a),
	.w4(32'hbbd7599b),
	.w5(32'hbbb0e85e),
	.w6(32'h3a9ba677),
	.w7(32'h3bbfe711),
	.w8(32'h3b2c6283),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6e196),
	.w1(32'h3b0bfa1e),
	.w2(32'hba44c8aa),
	.w3(32'hbb0c3e80),
	.w4(32'hbaf33fb3),
	.w5(32'hbb539e2b),
	.w6(32'hbad8dd48),
	.w7(32'hba3d3576),
	.w8(32'hbb0ee532),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd9f67),
	.w1(32'hba9dc6b1),
	.w2(32'hbb843508),
	.w3(32'h3b5b8740),
	.w4(32'h3a65fe5f),
	.w5(32'h3a849e17),
	.w6(32'hba695cd7),
	.w7(32'hbab81e41),
	.w8(32'h399629d9),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9304b8f),
	.w1(32'h3b934f66),
	.w2(32'h39551839),
	.w3(32'h3b0f07b3),
	.w4(32'h3ac18894),
	.w5(32'hb925b81b),
	.w6(32'h3b53d68e),
	.w7(32'h3ab20157),
	.w8(32'h3a29e312),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933f828),
	.w1(32'hb9205674),
	.w2(32'h39a219fd),
	.w3(32'hba0d47ec),
	.w4(32'hba4bcf54),
	.w5(32'h39f3d878),
	.w6(32'hb9955324),
	.w7(32'hba6bac53),
	.w8(32'hbabb5561),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b01bf),
	.w1(32'hbb3f5f09),
	.w2(32'hb9a2c025),
	.w3(32'hbb9e0607),
	.w4(32'hbba779e8),
	.w5(32'hbbbd1234),
	.w6(32'h3b5d8202),
	.w7(32'h3bf97cc4),
	.w8(32'h3be34d75),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc101e00),
	.w1(32'hbb2f6b8f),
	.w2(32'hb98349d2),
	.w3(32'hbbac1f62),
	.w4(32'hbb78db89),
	.w5(32'hbb4dfa2e),
	.w6(32'h3b678611),
	.w7(32'h3b99e984),
	.w8(32'h3b638de7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377c6193),
	.w1(32'h39f0a8f5),
	.w2(32'h391bcf25),
	.w3(32'hb8acd141),
	.w4(32'h39b5bf73),
	.w5(32'h39990c49),
	.w6(32'h39e401a0),
	.w7(32'hb898c51f),
	.w8(32'h394fad1c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9918459),
	.w1(32'hb8cfa731),
	.w2(32'h37c60313),
	.w3(32'hb9bd9ee5),
	.w4(32'hba07e15f),
	.w5(32'hba3e8b4f),
	.w6(32'hb896f323),
	.w7(32'hba4ba3f0),
	.w8(32'hb9c985cc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7ce5c),
	.w1(32'h3ad58c60),
	.w2(32'h3ab0a511),
	.w3(32'h3b19e685),
	.w4(32'h3aa53790),
	.w5(32'h3b71fc32),
	.w6(32'h3aa5f283),
	.w7(32'hba95ca95),
	.w8(32'hb897195a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e1534),
	.w1(32'hbb1ff17d),
	.w2(32'hbadfe62b),
	.w3(32'h3b6cec48),
	.w4(32'h3c1c56c7),
	.w5(32'h3b9edc13),
	.w6(32'h3b6d248a),
	.w7(32'h3b2c4277),
	.w8(32'h3ba43d8b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc6b3a),
	.w1(32'h3a1aac18),
	.w2(32'h39cee504),
	.w3(32'h3b1d53ad),
	.w4(32'h3a94d3ae),
	.w5(32'hba1f1006),
	.w6(32'h3b6be3ad),
	.w7(32'h3b3b9291),
	.w8(32'h3b379efc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e4ff8),
	.w1(32'h3c0c33ea),
	.w2(32'h3b30ab3f),
	.w3(32'h3c590bd7),
	.w4(32'h3b03c8a8),
	.w5(32'h3b1bad51),
	.w6(32'h3b188d7b),
	.w7(32'hbbdba102),
	.w8(32'hbb89224a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae2c44),
	.w1(32'h3b35cbab),
	.w2(32'h3af6ce47),
	.w3(32'hbaa9bef1),
	.w4(32'h3a96d542),
	.w5(32'h3a8b685f),
	.w6(32'hba1ae652),
	.w7(32'hb9fda12f),
	.w8(32'hb9e3b8e6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a427ccb),
	.w1(32'h39dcc876),
	.w2(32'h38a7b59c),
	.w3(32'h3a4837e7),
	.w4(32'h39ad2e50),
	.w5(32'h39a26f04),
	.w6(32'h38d0c6da),
	.w7(32'hb9c4fa51),
	.w8(32'hb7057861),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34a1ef),
	.w1(32'hb9f643db),
	.w2(32'hbaf995ad),
	.w3(32'h3b5fa1c7),
	.w4(32'hbc29b940),
	.w5(32'hbc23365b),
	.w6(32'h3a90b1f5),
	.w7(32'hbc34870d),
	.w8(32'hbc37570d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03ec45),
	.w1(32'h39a84c6f),
	.w2(32'h387d77d1),
	.w3(32'h3a72b014),
	.w4(32'h3ae06c1f),
	.w5(32'h3b039ff3),
	.w6(32'h3aac1137),
	.w7(32'h3a0a06ef),
	.w8(32'h3b065b37),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ae948),
	.w1(32'h3beb5c10),
	.w2(32'h3b25d1b4),
	.w3(32'h3ba4a9fc),
	.w4(32'hbc1410f1),
	.w5(32'hbc069a0b),
	.w6(32'h3abd53ff),
	.w7(32'hbc131cb9),
	.w8(32'hbc4639b4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385b4828),
	.w1(32'hb9792b93),
	.w2(32'hb82711c8),
	.w3(32'hb8b6ab35),
	.w4(32'hb9abc0be),
	.w5(32'hb96aa530),
	.w6(32'hb8e6869b),
	.w7(32'hb9e2e86a),
	.w8(32'hb9b46630),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e14c9b),
	.w1(32'hb9a93827),
	.w2(32'hb9be0b8a),
	.w3(32'hb9b0ecfa),
	.w4(32'hba06befe),
	.w5(32'hb8edfc89),
	.w6(32'hb9e0f30b),
	.w7(32'hb9e299e7),
	.w8(32'hb943fe81),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab27418),
	.w1(32'h3a1fc3f4),
	.w2(32'hba7c3c96),
	.w3(32'hbaefc89a),
	.w4(32'hb9d6ae55),
	.w5(32'hbb462118),
	.w6(32'h3aa8f3b6),
	.w7(32'h3a9d1b28),
	.w8(32'h3aa71222),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36d98c),
	.w1(32'h3b72a986),
	.w2(32'h3b040869),
	.w3(32'h39b10abe),
	.w4(32'h3b021439),
	.w5(32'h3b87f3a3),
	.w6(32'h3b0d7b99),
	.w7(32'hba39d890),
	.w8(32'h3a1ad254),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae55d1e),
	.w1(32'h3a8c196c),
	.w2(32'h3adfe2b4),
	.w3(32'hba4e1e76),
	.w4(32'hba752c75),
	.w5(32'h388c3abc),
	.w6(32'hbadfde5a),
	.w7(32'hbaa82150),
	.w8(32'hbaa9126d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe65bae),
	.w1(32'hbafb4483),
	.w2(32'h3af17cc8),
	.w3(32'hbb88ff29),
	.w4(32'hba05bff3),
	.w5(32'hbae02e6f),
	.w6(32'hbab41726),
	.w7(32'h3aae8ad6),
	.w8(32'h3b265388),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c44b7),
	.w1(32'hbc91bd1b),
	.w2(32'h3bc4b863),
	.w3(32'hbb350e29),
	.w4(32'h3bb851c8),
	.w5(32'h3c9c87b0),
	.w6(32'h3a2a0b40),
	.w7(32'hbb125bc3),
	.w8(32'h3c84ad60),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97eb12),
	.w1(32'h3b2c42e3),
	.w2(32'h3b933b64),
	.w3(32'h3c05f8f2),
	.w4(32'hba414e75),
	.w5(32'h3c0ae4c1),
	.w6(32'hbadfdce6),
	.w7(32'hbc52a690),
	.w8(32'hbb8b64ec),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbea44c),
	.w1(32'h3bad4857),
	.w2(32'h3a3a5c9c),
	.w3(32'h3c3e4c6b),
	.w4(32'hbbb6ca36),
	.w5(32'hbbad8a85),
	.w6(32'h3b93d5ec),
	.w7(32'hbc654172),
	.w8(32'hbc6e69fb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8429e3),
	.w1(32'h3a8aac3b),
	.w2(32'h3a6766e1),
	.w3(32'h3973e538),
	.w4(32'hba9f59ba),
	.w5(32'h39d6146d),
	.w6(32'hbabba5f9),
	.w7(32'hbb3bc6c4),
	.w8(32'hba32a174),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913d552),
	.w1(32'hbac667bf),
	.w2(32'hbaba3b38),
	.w3(32'hb97d53dc),
	.w4(32'hba8956bd),
	.w5(32'hbabbd8d1),
	.w6(32'hba600990),
	.w7(32'hba07a4c2),
	.w8(32'h3a4b98fc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c3a7e),
	.w1(32'h38cc435d),
	.w2(32'hb930728b),
	.w3(32'hb7cce01c),
	.w4(32'h39c950a0),
	.w5(32'h3a6665cb),
	.w6(32'h3a486551),
	.w7(32'h3a41cdd0),
	.w8(32'h3938e633),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa537f2),
	.w1(32'h3ac88f4d),
	.w2(32'h3b593b2e),
	.w3(32'h3aa1634f),
	.w4(32'h3b075910),
	.w5(32'h3b3922ca),
	.w6(32'h377fcebb),
	.w7(32'h3acabd64),
	.w8(32'h3b1a245b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a9de1),
	.w1(32'hbb0298d7),
	.w2(32'hbbbad68c),
	.w3(32'hbb76cd05),
	.w4(32'hb92da87e),
	.w5(32'hbbd9f5bf),
	.w6(32'h3b560d94),
	.w7(32'h3c09f2b7),
	.w8(32'hbb836267),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b941a07),
	.w1(32'hba81a1b7),
	.w2(32'hba01c19e),
	.w3(32'h3bdac006),
	.w4(32'h39069c7c),
	.w5(32'h3b02c274),
	.w6(32'h3b5bef30),
	.w7(32'hb993192a),
	.w8(32'h3a9b30bb),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb860ce10),
	.w1(32'hbb07a94d),
	.w2(32'h39a948cd),
	.w3(32'h3b936e6f),
	.w4(32'h3b1b0cc7),
	.w5(32'h3a9fc36a),
	.w6(32'h3ba6a3df),
	.w7(32'h3b8ec9f5),
	.w8(32'h3b6de888),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38f953),
	.w1(32'hb9c8ca2a),
	.w2(32'h383e98d4),
	.w3(32'h3b3ced24),
	.w4(32'hba484b82),
	.w5(32'h3aad3ac6),
	.w6(32'h3b6f9a44),
	.w7(32'h3b4930b7),
	.w8(32'h3b8fbbed),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbb67f8),
	.w1(32'hbc05169d),
	.w2(32'hba9029fa),
	.w3(32'hbc84b8c0),
	.w4(32'hbc05d9bf),
	.w5(32'hbbb1bc0a),
	.w6(32'h3b45d6c6),
	.w7(32'h3c1d24b8),
	.w8(32'h3c0c884e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9af7c9),
	.w1(32'h3a07fcda),
	.w2(32'h3831c8e1),
	.w3(32'hb96a0093),
	.w4(32'h39c9e7c8),
	.w5(32'h3a245c40),
	.w6(32'h39301236),
	.w7(32'hb810d45f),
	.w8(32'h394ff6e8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb057426),
	.w1(32'hba071043),
	.w2(32'hba2f9eed),
	.w3(32'hba887632),
	.w4(32'hb9a7bceb),
	.w5(32'hba4c151e),
	.w6(32'h3844bbfa),
	.w7(32'h39d16a20),
	.w8(32'hb999b4e9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a102bda),
	.w1(32'h3a28040a),
	.w2(32'hb9b9b759),
	.w3(32'h3a355c68),
	.w4(32'h3a8dcfc5),
	.w5(32'h39170b24),
	.w6(32'hb94f0a07),
	.w7(32'h398f6e57),
	.w8(32'h38af9d7a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc06f2),
	.w1(32'hb9bb3df3),
	.w2(32'hbbcf0daf),
	.w3(32'h3b652599),
	.w4(32'hbb1cc334),
	.w5(32'hbb90b3fc),
	.w6(32'h3ab0deb2),
	.w7(32'h3b3c8d9c),
	.w8(32'hbab3427d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2468e6),
	.w1(32'h3a88224b),
	.w2(32'h3a50f2f1),
	.w3(32'hbb34633d),
	.w4(32'h3a9a4a32),
	.w5(32'h39efbc6f),
	.w6(32'h3ad4e3bd),
	.w7(32'h3a8186b7),
	.w8(32'h3a9e4e6b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79e506),
	.w1(32'hbc1aeba4),
	.w2(32'hbb5a5b0d),
	.w3(32'hbc5064e9),
	.w4(32'hbba91b3b),
	.w5(32'hbbba5ac4),
	.w6(32'h3b8ffdbf),
	.w7(32'h3c103a26),
	.w8(32'h3b92d8a3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fd7a0),
	.w1(32'h3abb55c0),
	.w2(32'h39a34fb4),
	.w3(32'h3a7c40e0),
	.w4(32'h3aefe906),
	.w5(32'h39bb2065),
	.w6(32'h3b5d435f),
	.w7(32'h3b4e644b),
	.w8(32'h3a3d3f06),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1703de),
	.w1(32'hba478f8b),
	.w2(32'hbaa826d2),
	.w3(32'hb841fa89),
	.w4(32'hbaaaadde),
	.w5(32'hbb2129f4),
	.w6(32'hba001160),
	.w7(32'hba1942d8),
	.w8(32'h3a17c50c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bf86fb),
	.w1(32'h3a7a2ec6),
	.w2(32'h3a21e732),
	.w3(32'hba08c3b5),
	.w4(32'h398c835a),
	.w5(32'h3a423179),
	.w6(32'h3a13b197),
	.w7(32'hb936e40b),
	.w8(32'h3a1a054a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4c3dd),
	.w1(32'hb9ed9306),
	.w2(32'h39d16396),
	.w3(32'h3ad0c193),
	.w4(32'hb987082b),
	.w5(32'hb984e29f),
	.w6(32'h395a7aa0),
	.w7(32'hb9251b84),
	.w8(32'hb98af042),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1023d),
	.w1(32'h3a1fe80e),
	.w2(32'h3a976dd8),
	.w3(32'h3a45e688),
	.w4(32'h39acea5a),
	.w5(32'h3a83aebe),
	.w6(32'hb88e3378),
	.w7(32'h38e1aa4d),
	.w8(32'h38d4275d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22d3a2),
	.w1(32'h3a219086),
	.w2(32'h3a98b6a2),
	.w3(32'h39381427),
	.w4(32'h39a17c12),
	.w5(32'h3a0f4315),
	.w6(32'h39aac7e0),
	.w7(32'hb8bbf292),
	.w8(32'h3a16ff2e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74f7b0),
	.w1(32'h3a806c17),
	.w2(32'h3b18b7b9),
	.w3(32'hb9ced438),
	.w4(32'h3b1ae80b),
	.w5(32'hb9bee568),
	.w6(32'h3ba02e63),
	.w7(32'h3bc8ad61),
	.w8(32'h3b7e2d64),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb796444),
	.w1(32'h3b139219),
	.w2(32'hbb32e094),
	.w3(32'h3b8ad430),
	.w4(32'hbaaabc27),
	.w5(32'hbb119d3a),
	.w6(32'h3a635a04),
	.w7(32'h3a0eff09),
	.w8(32'hb992621e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba347587),
	.w1(32'h398a2874),
	.w2(32'hba5f2dbd),
	.w3(32'hba600c38),
	.w4(32'h39be91e2),
	.w5(32'hb823142b),
	.w6(32'hb885491d),
	.w7(32'hba40b3bb),
	.w8(32'h3b0293b3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15a56e),
	.w1(32'h38197314),
	.w2(32'hb987beff),
	.w3(32'h38ec4d2b),
	.w4(32'h3980db9c),
	.w5(32'h39b0722b),
	.w6(32'hba2a762d),
	.w7(32'hba38b2bd),
	.w8(32'hba2ac120),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c03b59),
	.w1(32'h399243e9),
	.w2(32'hb9c50d8f),
	.w3(32'h3a543100),
	.w4(32'h393aa363),
	.w5(32'hba123f84),
	.w6(32'hb912d0fb),
	.w7(32'hba1a6ca0),
	.w8(32'hba46800f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba711d4e),
	.w1(32'hba6ced55),
	.w2(32'hb9d083db),
	.w3(32'hb9c78f4d),
	.w4(32'hba34298f),
	.w5(32'h39cef588),
	.w6(32'h39ab319f),
	.w7(32'hb97b29b8),
	.w8(32'hba81f698),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de4446),
	.w1(32'h3b5da09d),
	.w2(32'h3c01d111),
	.w3(32'hbb0a105d),
	.w4(32'h3af61212),
	.w5(32'h3b4744cc),
	.w6(32'h3ab06142),
	.w7(32'h3bad59a8),
	.w8(32'h3acf4ea4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdcb26),
	.w1(32'h3b5a6d8b),
	.w2(32'h3abe941a),
	.w3(32'h3b9221ac),
	.w4(32'h3aab4546),
	.w5(32'hbb95e547),
	.w6(32'h3c159af5),
	.w7(32'h3c5f697d),
	.w8(32'h3c2f9daf),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26ff40),
	.w1(32'h3b6a8c59),
	.w2(32'h3afdc2d6),
	.w3(32'h3c368652),
	.w4(32'h3bd10f96),
	.w5(32'h3b915f65),
	.w6(32'h3bbf912f),
	.w7(32'h3bf1fd1c),
	.w8(32'h3c03260c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca44a79),
	.w1(32'h3c0aa8e7),
	.w2(32'hb9933240),
	.w3(32'h3c73ef42),
	.w4(32'hb8bff880),
	.w5(32'h3a70f52e),
	.w6(32'h3b37384b),
	.w7(32'hbbe4150a),
	.w8(32'hbbab7bd3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c5cb2),
	.w1(32'hba1e1761),
	.w2(32'hb97e9a93),
	.w3(32'hb9c39ea0),
	.w4(32'hb9e05bf1),
	.w5(32'h39b0534e),
	.w6(32'hba5a7429),
	.w7(32'hba3c1f32),
	.w8(32'hba4c0bd9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a7eef),
	.w1(32'hb99ff3e6),
	.w2(32'h39d6d7ab),
	.w3(32'hb784ff8d),
	.w4(32'hb9c11652),
	.w5(32'h399b5a6d),
	.w6(32'h371e0558),
	.w7(32'h388d1d93),
	.w8(32'h38c009a5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944e433),
	.w1(32'hb8dd6981),
	.w2(32'hb97d1284),
	.w3(32'h39a9495c),
	.w4(32'hb928c0a3),
	.w5(32'hb98c5921),
	.w6(32'h395b40e2),
	.w7(32'h38fa7ae5),
	.w8(32'h39dd98a5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0de042),
	.w1(32'hbabc44e1),
	.w2(32'h39496f0d),
	.w3(32'hbae60245),
	.w4(32'hbaaaaf2b),
	.w5(32'hb9a6b0ab),
	.w6(32'h3a3a907a),
	.w7(32'h39f1eb9f),
	.w8(32'h3a962ab0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcdbc1),
	.w1(32'h380b3027),
	.w2(32'hb99936ee),
	.w3(32'hb9e2a057),
	.w4(32'hb930eaae),
	.w5(32'hb95c3d9f),
	.w6(32'hb8998eff),
	.w7(32'h37cb8cf5),
	.w8(32'hba2604c4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a7028),
	.w1(32'hbbe33fd1),
	.w2(32'hba9d956f),
	.w3(32'hbbd07e1b),
	.w4(32'hbacafc34),
	.w5(32'h3a5684ec),
	.w6(32'hb9ec7535),
	.w7(32'h3ac0d9e5),
	.w8(32'h3b251892),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaf70d),
	.w1(32'hbc044f8b),
	.w2(32'hbb17b3e4),
	.w3(32'hbc1b76fc),
	.w4(32'hbb14432f),
	.w5(32'h3a61a875),
	.w6(32'hbad6d877),
	.w7(32'h3b11daea),
	.w8(32'h3c3687c4),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4aced),
	.w1(32'hb94282dc),
	.w2(32'hba5e9aec),
	.w3(32'h39ff9356),
	.w4(32'hbb97d9bc),
	.w5(32'hbaf2726d),
	.w6(32'h3b86eca2),
	.w7(32'hb88d0987),
	.w8(32'h3a818711),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56e54f),
	.w1(32'h39dc360c),
	.w2(32'hb7e17f55),
	.w3(32'h3b2e26bc),
	.w4(32'h3aca5b0e),
	.w5(32'hba7d59ea),
	.w6(32'h3b54ca46),
	.w7(32'h3aeb4c3d),
	.w8(32'hba0dd931),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb66327),
	.w1(32'hbb1c937f),
	.w2(32'h3bb03a57),
	.w3(32'hbbc36a75),
	.w4(32'hb9cfa441),
	.w5(32'h3ac8cd94),
	.w6(32'hbb346101),
	.w7(32'hb9334341),
	.w8(32'hba0c46db),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34a030),
	.w1(32'hbadb0b13),
	.w2(32'hbb85ca22),
	.w3(32'h3b3585f5),
	.w4(32'hba9e2ff0),
	.w5(32'hbb05aa2a),
	.w6(32'h3a86ebbf),
	.w7(32'hba2eb1a4),
	.w8(32'hbad83e97),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf177be),
	.w1(32'hbaec2d87),
	.w2(32'hb9d5a09b),
	.w3(32'hbbb6c004),
	.w4(32'hbafc25f6),
	.w5(32'hba0b9631),
	.w6(32'h3a813c77),
	.w7(32'h3b48e2c3),
	.w8(32'h3af8be93),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a160217),
	.w1(32'h399afd63),
	.w2(32'h388820fc),
	.w3(32'h3a365342),
	.w4(32'h38428a7b),
	.w5(32'hba08e8e0),
	.w6(32'h3a073fdc),
	.w7(32'h39c0db29),
	.w8(32'h39f75322),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f96911),
	.w1(32'h39fd5f8b),
	.w2(32'h3a8be888),
	.w3(32'hb9c3cf22),
	.w4(32'h39b9266c),
	.w5(32'h39fa51b7),
	.w6(32'h394f38b7),
	.w7(32'h39ac2eb4),
	.w8(32'hb7cbcbe8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba49cd),
	.w1(32'hbaa3ecbb),
	.w2(32'hba07eb84),
	.w3(32'h3a2bf216),
	.w4(32'h3ac74517),
	.w5(32'h3a9de406),
	.w6(32'h39e0d363),
	.w7(32'h39acc7fe),
	.w8(32'h3a0387ff),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce3c89),
	.w1(32'h3a008979),
	.w2(32'h3a3d7abd),
	.w3(32'h3a69a2d7),
	.w4(32'hbab5a398),
	.w5(32'hb9d257be),
	.w6(32'h397088dd),
	.w7(32'hba5bfb62),
	.w8(32'hb923a3d1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c133f51),
	.w1(32'h3a9d2088),
	.w2(32'h3b4d949f),
	.w3(32'h3baff621),
	.w4(32'h3b1fd1d7),
	.w5(32'h3bba7d49),
	.w6(32'h3b156d38),
	.w7(32'hbabaa7c9),
	.w8(32'h3a215cd8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a774f83),
	.w1(32'hba139db1),
	.w2(32'h3a4d8d46),
	.w3(32'h39c85058),
	.w4(32'hba874051),
	.w5(32'hb7f27888),
	.w6(32'hb9c44baf),
	.w7(32'hb9f8073d),
	.w8(32'h3a20ac59),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4086ca),
	.w1(32'h388076bf),
	.w2(32'hba3becf2),
	.w3(32'h3b878f89),
	.w4(32'h3b05b95e),
	.w5(32'hba881fcf),
	.w6(32'h3b6c834d),
	.w7(32'h3b3199ee),
	.w8(32'hb7d4d20f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09319c),
	.w1(32'hbb706094),
	.w2(32'h39bab4b8),
	.w3(32'hbbe95316),
	.w4(32'hbb91650b),
	.w5(32'hbaa69f72),
	.w6(32'h3a2cb25d),
	.w7(32'h3af5f8b9),
	.w8(32'h3bbb4e48),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf87e10),
	.w1(32'h3902a431),
	.w2(32'hba55abcd),
	.w3(32'h3b30972a),
	.w4(32'hbb57e8e4),
	.w5(32'hbaf3dfa1),
	.w6(32'h3adcf1d2),
	.w7(32'hbbc19c5d),
	.w8(32'hbb4fa412),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ad1ad),
	.w1(32'hbbcf358d),
	.w2(32'h3b2d53cf),
	.w3(32'hbc09ca35),
	.w4(32'h3be85ab0),
	.w5(32'h3c1eac2f),
	.w6(32'hbb91d93e),
	.w7(32'h3b7e87fa),
	.w8(32'h3bb81716),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7f336),
	.w1(32'h3b40ee8c),
	.w2(32'h3ad3449f),
	.w3(32'h3bca259c),
	.w4(32'h3a208219),
	.w5(32'hbaea9a79),
	.w6(32'h3b609b3b),
	.w7(32'hbb4c7ac0),
	.w8(32'hbb3b143f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba825a5),
	.w1(32'hbac9c464),
	.w2(32'hb9f5fc69),
	.w3(32'h3bac9c12),
	.w4(32'h3ba99280),
	.w5(32'h3a55808d),
	.w6(32'h3beac698),
	.w7(32'h3c07883e),
	.w8(32'h3bd3f631),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb352d4),
	.w1(32'h3bd415ff),
	.w2(32'h3b834a12),
	.w3(32'h3bb2581a),
	.w4(32'h3b98e8ea),
	.w5(32'h3ab11407),
	.w6(32'h3be389c3),
	.w7(32'h3ba69a1e),
	.w8(32'h3aba3451),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59803d),
	.w1(32'h3b8012d1),
	.w2(32'h3a166926),
	.w3(32'h3a629f38),
	.w4(32'hbbcee575),
	.w5(32'hbb80791c),
	.w6(32'hb8051ed6),
	.w7(32'hbbf3e4e9),
	.w8(32'hbbbd04ee),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71efab),
	.w1(32'h398a3617),
	.w2(32'h3a66d6ff),
	.w3(32'h3a675f2b),
	.w4(32'h3a4efcf8),
	.w5(32'h3a0570a0),
	.w6(32'h3a7a3c71),
	.w7(32'h3aacb052),
	.w8(32'hb978d165),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd33eab),
	.w1(32'h3a304ece),
	.w2(32'hba494b7e),
	.w3(32'hba9e3831),
	.w4(32'h3a4c7877),
	.w5(32'hbb70d94f),
	.w6(32'h3be422c6),
	.w7(32'h3bce7f0d),
	.w8(32'h3b347bdc),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40c8a0),
	.w1(32'hbb0922c4),
	.w2(32'h3b9df209),
	.w3(32'hbb0e5ea1),
	.w4(32'h3bbb0995),
	.w5(32'h3c0ed364),
	.w6(32'h3be28d49),
	.w7(32'h3bfcd03c),
	.w8(32'h3bf2a7ab),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eea4d),
	.w1(32'hbc4797e4),
	.w2(32'hbba169cd),
	.w3(32'hbba8009d),
	.w4(32'h3b76e8d8),
	.w5(32'h3b540c9c),
	.w6(32'hbbf75ef9),
	.w7(32'hbba3e388),
	.w8(32'h3c4132bc),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4014a),
	.w1(32'h37830774),
	.w2(32'h3ba145c7),
	.w3(32'h3ba6b271),
	.w4(32'h3b85d9bb),
	.w5(32'h3bd78780),
	.w6(32'hbb5f1230),
	.w7(32'hbbf19d4e),
	.w8(32'hbafee92b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb904c6),
	.w1(32'hba303dab),
	.w2(32'hbb20fec8),
	.w3(32'h3bdb76c3),
	.w4(32'hba9fe034),
	.w5(32'hbb4ced79),
	.w6(32'h3a839994),
	.w7(32'hbb2e2ba9),
	.w8(32'hbb9241b7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50641c),
	.w1(32'hbafd43f5),
	.w2(32'h3bf8390c),
	.w3(32'hbb21c633),
	.w4(32'h3c4a56b5),
	.w5(32'h3c103c57),
	.w6(32'h3b0ef9d9),
	.w7(32'h3c28dc05),
	.w8(32'h3c3e85f3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0e9e3),
	.w1(32'h398d080e),
	.w2(32'h3ac8fcfa),
	.w3(32'h399bc63a),
	.w4(32'h3a5e856d),
	.w5(32'h3b0dbdc8),
	.w6(32'h3a4bcd00),
	.w7(32'h3b1d76a3),
	.w8(32'h3aebbab0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8974bd),
	.w1(32'hbc8c0736),
	.w2(32'hbbe65435),
	.w3(32'hbc42c02c),
	.w4(32'hba9beb8f),
	.w5(32'h3b923b61),
	.w6(32'h3b95b1d2),
	.w7(32'h3b88ad86),
	.w8(32'h3c01bed1),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59e689),
	.w1(32'hbbee8551),
	.w2(32'hba3e2af0),
	.w3(32'h3af5517f),
	.w4(32'hbab790a6),
	.w5(32'hb998034f),
	.w6(32'hba372762),
	.w7(32'hba632b84),
	.w8(32'h3a8ebf06),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be40c5),
	.w1(32'h3a9c38d0),
	.w2(32'h3a9807a4),
	.w3(32'hb90d5e0c),
	.w4(32'h3a00e6ca),
	.w5(32'h3a785d44),
	.w6(32'h3ab59268),
	.w7(32'h3a7b21c4),
	.w8(32'h3a87821b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bfc94),
	.w1(32'h3a4560e0),
	.w2(32'hba1c1d14),
	.w3(32'h3b897541),
	.w4(32'h3a534f54),
	.w5(32'h3a953de3),
	.w6(32'hba57a288),
	.w7(32'h3957da38),
	.w8(32'h38d4b857),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd93d9f),
	.w1(32'hba6b5425),
	.w2(32'h39461f9e),
	.w3(32'hbb9f0d01),
	.w4(32'hbb23749b),
	.w5(32'hbb83d90d),
	.w6(32'h3a9d5d61),
	.w7(32'h3b402812),
	.w8(32'h3a682d76),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce867c),
	.w1(32'h3b73115f),
	.w2(32'h3ac771c8),
	.w3(32'h3ba7752f),
	.w4(32'h38162b90),
	.w5(32'hb8a0d056),
	.w6(32'h3b23a895),
	.w7(32'hbb162ee4),
	.w8(32'hbae27e52),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c055168),
	.w1(32'h391d94d4),
	.w2(32'hbb60c1c2),
	.w3(32'h3b85ce96),
	.w4(32'hbaf98991),
	.w5(32'hbb772a8d),
	.w6(32'h3a9bb00c),
	.w7(32'hbbdf1751),
	.w8(32'hbb9e2fe1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cd57c),
	.w1(32'hb96dd294),
	.w2(32'hb98d1dbf),
	.w3(32'h3b0f1077),
	.w4(32'h3a0c4536),
	.w5(32'hbaa6302e),
	.w6(32'h39d26300),
	.w7(32'hbaa0a2b4),
	.w8(32'hbad30112),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4d721),
	.w1(32'h3b2d4cc6),
	.w2(32'h3bc96edf),
	.w3(32'hbaaa934a),
	.w4(32'h3b3d7284),
	.w5(32'h3b87e659),
	.w6(32'h3b6ef820),
	.w7(32'h3bcccc57),
	.w8(32'h3c3ced9c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35867f),
	.w1(32'h3aa411a6),
	.w2(32'hb9cb0e60),
	.w3(32'hbb16024f),
	.w4(32'h3adeeaa6),
	.w5(32'h3a93ba7c),
	.w6(32'h3ae0dc96),
	.w7(32'h3a62a69f),
	.w8(32'hbac4771e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c02b3),
	.w1(32'hb96641f5),
	.w2(32'hbaadfc8c),
	.w3(32'h3b4dfb0f),
	.w4(32'h3a0df5ab),
	.w5(32'hba901e1e),
	.w6(32'h3ae6f125),
	.w7(32'h3a296748),
	.w8(32'h3a10bcb5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987ec3f),
	.w1(32'h3a1bc2ea),
	.w2(32'h39d02c0d),
	.w3(32'hba77d0c5),
	.w4(32'h391c2b2b),
	.w5(32'h39185d21),
	.w6(32'h39f546da),
	.w7(32'hb9192f65),
	.w8(32'h3a559fc5),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2964a0),
	.w1(32'hb7600bb3),
	.w2(32'h3a8f1c84),
	.w3(32'h3a806cf2),
	.w4(32'hb983e9d1),
	.w5(32'h3a9cfae3),
	.w6(32'h3a68fee8),
	.w7(32'h398a675b),
	.w8(32'h39e1ac7d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395aca82),
	.w1(32'hb741a320),
	.w2(32'h3919874b),
	.w3(32'h39cec16a),
	.w4(32'h37accd82),
	.w5(32'h396d3f77),
	.w6(32'h39ff6695),
	.w7(32'h38d14326),
	.w8(32'h39ea4054),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e355ba),
	.w1(32'hba1b5d29),
	.w2(32'hba36a6e4),
	.w3(32'h3a9c2b82),
	.w4(32'h3a738834),
	.w5(32'h3a871d23),
	.w6(32'h388506ae),
	.w7(32'h39b05fd8),
	.w8(32'hb836ce13),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f76d6),
	.w1(32'h3ab48bf9),
	.w2(32'hba08be85),
	.w3(32'h3b86f584),
	.w4(32'h3b3da389),
	.w5(32'h38189a68),
	.w6(32'h3b55ebf8),
	.w7(32'h3b1737bc),
	.w8(32'h3a4fbb32),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8a0c2),
	.w1(32'hb9abd1ba),
	.w2(32'hba0a8847),
	.w3(32'hb9f434b0),
	.w4(32'hb8e94229),
	.w5(32'hb94fba39),
	.w6(32'h3a194654),
	.w7(32'h3913fb9d),
	.w8(32'hb9cf6c0d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d87fe),
	.w1(32'hbb4f95a6),
	.w2(32'h3981968a),
	.w3(32'hbb88d4de),
	.w4(32'h39805492),
	.w5(32'hb82a5690),
	.w6(32'hba9fef49),
	.w7(32'h3b77b118),
	.w8(32'h3b615965),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c610b68),
	.w1(32'h3c0bc71f),
	.w2(32'h3b63ce41),
	.w3(32'h3bc9bffe),
	.w4(32'hbab5a1ae),
	.w5(32'hb994bb97),
	.w6(32'hbaef14e5),
	.w7(32'hbc0f7409),
	.w8(32'hbc1c3577),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10912d),
	.w1(32'hba88a57c),
	.w2(32'hb99886aa),
	.w3(32'h3966324f),
	.w4(32'h386eb8a4),
	.w5(32'h380841b0),
	.w6(32'hb6909a5f),
	.w7(32'h396b32f0),
	.w8(32'hb88eb124),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3443336e),
	.w1(32'h3a47683d),
	.w2(32'h3a4323b4),
	.w3(32'hb95566cf),
	.w4(32'h39f908cf),
	.w5(32'h3a95dc06),
	.w6(32'h3a317cb8),
	.w7(32'hb944297b),
	.w8(32'hb994bf82),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b604c),
	.w1(32'h371b6013),
	.w2(32'hb98b4508),
	.w3(32'h39633394),
	.w4(32'hb884e086),
	.w5(32'hb99f13e3),
	.w6(32'h393453f0),
	.w7(32'hba09a4ab),
	.w8(32'hb96a3d83),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54f55f),
	.w1(32'h39c186ee),
	.w2(32'h39b8d3fa),
	.w3(32'hb97dc9a0),
	.w4(32'h37582ff3),
	.w5(32'hb987243b),
	.w6(32'h3a45e3d9),
	.w7(32'h3a1f78e7),
	.w8(32'h39b56255),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd941c),
	.w1(32'hba909180),
	.w2(32'h3b6d5fe1),
	.w3(32'hbb4d602e),
	.w4(32'hbb0b6142),
	.w5(32'hbc3e0ae0),
	.w6(32'hbba2ab64),
	.w7(32'h3b6c6e43),
	.w8(32'h3bc7a7b3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd12fc1),
	.w1(32'hba9238f3),
	.w2(32'h3a01b32c),
	.w3(32'hbbba5735),
	.w4(32'hbb2e318d),
	.w5(32'hbbc381e2),
	.w6(32'h3ae3d9cb),
	.w7(32'h3b89bfc9),
	.w8(32'h3a8df6d3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4ddab),
	.w1(32'hba67bf00),
	.w2(32'h3a07a531),
	.w3(32'hbaa31620),
	.w4(32'h3956f73c),
	.w5(32'h39cf5583),
	.w6(32'h39e1bb4c),
	.w7(32'h3a83efd0),
	.w8(32'h3a3753e3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5816a),
	.w1(32'hba7f6328),
	.w2(32'h3a65af59),
	.w3(32'h39dbf64c),
	.w4(32'h3abd4cfb),
	.w5(32'h39bc4548),
	.w6(32'h3af42633),
	.w7(32'h3b32d448),
	.w8(32'h3b75503d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eb14c),
	.w1(32'h3974b1a7),
	.w2(32'h3a4fb32a),
	.w3(32'h3acfd27e),
	.w4(32'hb9dbaa70),
	.w5(32'h39941d74),
	.w6(32'h3ae1ae87),
	.w7(32'hba440640),
	.w8(32'h3940ecf9),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bf3e8a),
	.w1(32'h3a53359a),
	.w2(32'hb9e8253c),
	.w3(32'h3a480ff6),
	.w4(32'h39d1257a),
	.w5(32'hba4389b0),
	.w6(32'h3b09478f),
	.w7(32'h3ac22d2f),
	.w8(32'h3ab415f4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6aeec),
	.w1(32'h3b205b36),
	.w2(32'h3a5fa477),
	.w3(32'h3bd625d3),
	.w4(32'h3b108594),
	.w5(32'h3b15eb65),
	.w6(32'h3b98e30f),
	.w7(32'hb9ead161),
	.w8(32'hba7af700),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77633a),
	.w1(32'hbb849fbc),
	.w2(32'h3aa67eb3),
	.w3(32'hbc1081e9),
	.w4(32'hbab49a86),
	.w5(32'hbae67f16),
	.w6(32'hbae2773f),
	.w7(32'h3bc3441b),
	.w8(32'h3b3690bc),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2aafb),
	.w1(32'h3abd7850),
	.w2(32'hb9e3d87c),
	.w3(32'h3ada874f),
	.w4(32'hbafb0b75),
	.w5(32'hbb2208da),
	.w6(32'hba9dbd1f),
	.w7(32'hbba8437c),
	.w8(32'hbb8aabfc),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc51d08),
	.w1(32'h3ad6c858),
	.w2(32'h3a8bd63a),
	.w3(32'hbb05d3cb),
	.w4(32'h3b2151b4),
	.w5(32'h3b073950),
	.w6(32'h3a15254d),
	.w7(32'h3b3f02f3),
	.w8(32'h3aee72eb),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34709e),
	.w1(32'hbb7e5623),
	.w2(32'h3997ff18),
	.w3(32'hbb648bd1),
	.w4(32'h3b55959a),
	.w5(32'h3a849fd3),
	.w6(32'h3af318fe),
	.w7(32'h3bac3113),
	.w8(32'h3b30d4bd),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f0333),
	.w1(32'h38f158e2),
	.w2(32'h3ad79d6c),
	.w3(32'h3bb73cbc),
	.w4(32'h3b220946),
	.w5(32'h3b934068),
	.w6(32'h3af4cc94),
	.w7(32'h3a9970ea),
	.w8(32'h3b9792bd),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89f82f),
	.w1(32'hbab8ee42),
	.w2(32'h3a9cce53),
	.w3(32'hbb02b0be),
	.w4(32'h3b139d02),
	.w5(32'h3a997502),
	.w6(32'h3aa82a07),
	.w7(32'h3b54bbeb),
	.w8(32'h3a43a8ba),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb845ad81),
	.w1(32'hb94f1c75),
	.w2(32'hb9b50121),
	.w3(32'hb9812e18),
	.w4(32'hb9c36155),
	.w5(32'hb9b52130),
	.w6(32'h39f4c959),
	.w7(32'hb8e832c6),
	.w8(32'h3814943d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c791fb0),
	.w1(32'h3b8b0364),
	.w2(32'h3ba8e88c),
	.w3(32'h3baed7f4),
	.w4(32'hbbe62f4b),
	.w5(32'hbbb955ca),
	.w6(32'h3acc0515),
	.w7(32'hbc39aacc),
	.w8(32'hbc280884),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40323f),
	.w1(32'h3a85ad59),
	.w2(32'h3b0228a6),
	.w3(32'h3b163e73),
	.w4(32'h3afd2769),
	.w5(32'h3b06a118),
	.w6(32'hb9041586),
	.w7(32'h3ab5fce6),
	.w8(32'h3b312056),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388ab384),
	.w1(32'hb7af04c2),
	.w2(32'h393a2c4f),
	.w3(32'hba2cc25c),
	.w4(32'hb78df4e7),
	.w5(32'h39339dcc),
	.w6(32'hb961f7b3),
	.w7(32'h38e1979f),
	.w8(32'h39b58bfb),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b388c),
	.w1(32'h38e83b5c),
	.w2(32'h39b14912),
	.w3(32'h38c565ed),
	.w4(32'h392450bd),
	.w5(32'h398fa386),
	.w6(32'h39060622),
	.w7(32'hb8febcb4),
	.w8(32'h38efd054),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb042f33),
	.w1(32'hbb279199),
	.w2(32'h399f8d8a),
	.w3(32'hba995b9b),
	.w4(32'hba3550a8),
	.w5(32'h3a643f60),
	.w6(32'h3a37cd84),
	.w7(32'h3aa60b91),
	.w8(32'h3b093689),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be999e2),
	.w1(32'h3a8fd23b),
	.w2(32'h3b2d7630),
	.w3(32'h3b7872d1),
	.w4(32'hba2b6e06),
	.w5(32'h3b7ddb6b),
	.w6(32'h3a0d61ba),
	.w7(32'hbb31242c),
	.w8(32'h3995d574),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05bbfd),
	.w1(32'hbbc9d712),
	.w2(32'hbad616b8),
	.w3(32'hbbc46bf2),
	.w4(32'hbbf2872a),
	.w5(32'hbb9bf8b1),
	.w6(32'h3b2e1616),
	.w7(32'h38b364a5),
	.w8(32'h3a53290a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f39e88),
	.w1(32'hb92f84e4),
	.w2(32'hb92117af),
	.w3(32'h3589d11f),
	.w4(32'hb9143530),
	.w5(32'hb93bc30e),
	.w6(32'h387ccea5),
	.w7(32'h388ebbaf),
	.w8(32'h39072b29),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64f8ac),
	.w1(32'hbaeef718),
	.w2(32'hba298efd),
	.w3(32'hbb7a40da),
	.w4(32'hbadecab3),
	.w5(32'hbb45f8e8),
	.w6(32'h3aa9f200),
	.w7(32'h3ac0ebc5),
	.w8(32'hbaf25877),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80a38a),
	.w1(32'h39cf066e),
	.w2(32'hba2ea4f0),
	.w3(32'hb9361885),
	.w4(32'hba727c4f),
	.w5(32'hbb5e6ed2),
	.w6(32'h3a4f8fd7),
	.w7(32'h3919be02),
	.w8(32'hbb049a92),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49e28e),
	.w1(32'hbb7db42b),
	.w2(32'h39f3ac5a),
	.w3(32'hbbb151dd),
	.w4(32'h3b74d2e6),
	.w5(32'h3b91c888),
	.w6(32'hba0d20e6),
	.w7(32'h3bf186c7),
	.w8(32'h3bfc17a2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b40b8),
	.w1(32'hba2d6718),
	.w2(32'hbb07c96a),
	.w3(32'h3bc1c3df),
	.w4(32'hbba62a62),
	.w5(32'h3a3e6854),
	.w6(32'h3b8640b7),
	.w7(32'hbbd675cf),
	.w8(32'hbc026128),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc21fa2),
	.w1(32'h3b2368dc),
	.w2(32'h3ab51495),
	.w3(32'h3b76039f),
	.w4(32'h3acbec87),
	.w5(32'h3b005a13),
	.w6(32'h3a8b7327),
	.w7(32'hbac92e58),
	.w8(32'hbb0bd041),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c5b1e),
	.w1(32'h3901fb7c),
	.w2(32'h3ab97c1c),
	.w3(32'h3a6452a7),
	.w4(32'h3abf20c9),
	.w5(32'h3b008b35),
	.w6(32'h3aba2e19),
	.w7(32'h3abcc7a9),
	.w8(32'h3b1453b1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03365a),
	.w1(32'hb9b1c554),
	.w2(32'h3a815f54),
	.w3(32'h3b544fee),
	.w4(32'h39d2dc19),
	.w5(32'h3af626ff),
	.w6(32'h3b0a69ec),
	.w7(32'h3aaebebf),
	.w8(32'h3b31397b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8752a),
	.w1(32'h3b219dab),
	.w2(32'h3b64bdfd),
	.w3(32'h3be37866),
	.w4(32'h3b2ecd3b),
	.w5(32'h3bb8f8e2),
	.w6(32'h3be2afdd),
	.w7(32'h3abca617),
	.w8(32'h3b1fc84e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd44514),
	.w1(32'h3b37133b),
	.w2(32'h3b04a1e3),
	.w3(32'h3b66e11c),
	.w4(32'h394b1bfc),
	.w5(32'h3ae64dde),
	.w6(32'h3a91cf49),
	.w7(32'hbb469a3d),
	.w8(32'hbaaa216b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e876e),
	.w1(32'hbaf4a2bb),
	.w2(32'h39582628),
	.w3(32'hbb0e4178),
	.w4(32'h3a225bb8),
	.w5(32'h3a918d14),
	.w6(32'h38843030),
	.w7(32'h3af7d888),
	.w8(32'h3ad7d3fc),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7ef8d),
	.w1(32'h38ea91ee),
	.w2(32'h39333aa7),
	.w3(32'h3a46705a),
	.w4(32'h3a130ede),
	.w5(32'h39fae3d4),
	.w6(32'h3a2fd793),
	.w7(32'h395e486e),
	.w8(32'hb8f4189b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe956ae),
	.w1(32'hba217e1a),
	.w2(32'h3b1fee99),
	.w3(32'hbb99fe0d),
	.w4(32'h3a809ea7),
	.w5(32'h3a321c8b),
	.w6(32'hb910d6ac),
	.w7(32'h3b4cab6a),
	.w8(32'h3b60a5e4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96506a),
	.w1(32'hba9a9a58),
	.w2(32'h3a933409),
	.w3(32'hb9e1934e),
	.w4(32'hb6dd33aa),
	.w5(32'h3aafc7f4),
	.w6(32'hba32b7e3),
	.w7(32'hba621069),
	.w8(32'h3a2c1b63),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a720d3e),
	.w1(32'h3b232dc7),
	.w2(32'h3ad7ab12),
	.w3(32'h3b743626),
	.w4(32'h3a214504),
	.w5(32'hba4d830a),
	.w6(32'h3ad9f6d9),
	.w7(32'h3a1f8374),
	.w8(32'hb9625aee),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900ef58),
	.w1(32'h38bf2361),
	.w2(32'h3987e9a1),
	.w3(32'hb999943f),
	.w4(32'hb93c7841),
	.w5(32'h398a2cc5),
	.w6(32'hb96aab36),
	.w7(32'h38b71384),
	.w8(32'h39850bb6),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe36ec),
	.w1(32'h3bba15f9),
	.w2(32'h3ba6d434),
	.w3(32'h3b2c883b),
	.w4(32'hba8a0852),
	.w5(32'hbbcaf1d6),
	.w6(32'h3bae26df),
	.w7(32'h3b50f21c),
	.w8(32'hba983cda),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d66f54),
	.w1(32'hb71a68e1),
	.w2(32'h38a1a04d),
	.w3(32'hb915a38e),
	.w4(32'hb7e7f323),
	.w5(32'h38459e88),
	.w6(32'hb8df62bf),
	.w7(32'h395454b7),
	.w8(32'h38923135),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39937968),
	.w1(32'hb9492fae),
	.w2(32'hba1c7e6d),
	.w3(32'h3a188e96),
	.w4(32'hb932671b),
	.w5(32'hba12f549),
	.w6(32'h3a19cbeb),
	.w7(32'hb8838629),
	.w8(32'hba08a3be),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92238d),
	.w1(32'h3a718991),
	.w2(32'hba14e0cb),
	.w3(32'h3b828c78),
	.w4(32'h3add986d),
	.w5(32'h3b1b4fdc),
	.w6(32'h3a8edbae),
	.w7(32'h3a07ba1d),
	.w8(32'h3ac05173),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcebfe9),
	.w1(32'h39f7c5b7),
	.w2(32'h3b36bc74),
	.w3(32'hbb8e3dc5),
	.w4(32'h38cae07d),
	.w5(32'h394ec684),
	.w6(32'hbb12a753),
	.w7(32'h3b7636c5),
	.w8(32'h3bc7713a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc8922),
	.w1(32'h39803bff),
	.w2(32'h3a3be35e),
	.w3(32'h3a67978d),
	.w4(32'hb8d65a27),
	.w5(32'h39ece31a),
	.w6(32'h38f4b939),
	.w7(32'hb95573c2),
	.w8(32'hb8207e34),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83339f),
	.w1(32'h3b3a924a),
	.w2(32'hba80202b),
	.w3(32'h3a86ee6d),
	.w4(32'hbaf8bac6),
	.w5(32'hbb9f7012),
	.w6(32'h3a8b07d0),
	.w7(32'hbb06f902),
	.w8(32'hbba18c39),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18e447),
	.w1(32'hb9fe3d34),
	.w2(32'hbb0b85cb),
	.w3(32'h3a1e9aa6),
	.w4(32'hbb87336f),
	.w5(32'hbb183127),
	.w6(32'h3889587b),
	.w7(32'hbb27ab16),
	.w8(32'hbb7d926f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd768b),
	.w1(32'hba8bead1),
	.w2(32'hbb0df220),
	.w3(32'h3bcd8325),
	.w4(32'hb7f5fa92),
	.w5(32'hbb863b0f),
	.w6(32'h3c0ddf7a),
	.w7(32'h3c178a22),
	.w8(32'h3b507d05),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf90883),
	.w1(32'hba2889ab),
	.w2(32'hba8064ac),
	.w3(32'h395d63cd),
	.w4(32'h3a964e71),
	.w5(32'h3b05c671),
	.w6(32'h3aff1de4),
	.w7(32'h3adf6a99),
	.w8(32'h3b1eebf5),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099502),
	.w1(32'hbafdd917),
	.w2(32'hb98004a6),
	.w3(32'hbb94453c),
	.w4(32'hb9cac98d),
	.w5(32'hbb5a0a46),
	.w6(32'h3b23f7a0),
	.w7(32'h3b9b104a),
	.w8(32'h3aaeba65),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8daedd1),
	.w1(32'h3a2420e4),
	.w2(32'h3a6069e0),
	.w3(32'hb9ff06f1),
	.w4(32'h3a5fff6a),
	.w5(32'h3aa1f9eb),
	.w6(32'hb9e020a9),
	.w7(32'h3997a887),
	.w8(32'h3a92e893),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12d8aa),
	.w1(32'h3b43378a),
	.w2(32'h3a608094),
	.w3(32'h3b3da1be),
	.w4(32'h3ada1cec),
	.w5(32'hba181580),
	.w6(32'h3b53da72),
	.w7(32'h3ab27a11),
	.w8(32'hbaf671b5),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c6c367),
	.w1(32'hb65004f4),
	.w2(32'h3809adec),
	.w3(32'h38c67bf9),
	.w4(32'hb6fd2558),
	.w5(32'hb7266460),
	.w6(32'h38f39332),
	.w7(32'h390bd16e),
	.w8(32'h391129d6),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6de72e),
	.w1(32'h38ab8ac6),
	.w2(32'h39cd7397),
	.w3(32'h3a85cd08),
	.w4(32'h396959d2),
	.w5(32'h3a682f76),
	.w6(32'h3ab3b857),
	.w7(32'hb835fbd6),
	.w8(32'h3a7a92c9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae95ccd),
	.w1(32'h3a897804),
	.w2(32'h390411af),
	.w3(32'h3ac5ce1b),
	.w4(32'hb913d4ff),
	.w5(32'h38da27e8),
	.w6(32'h38efb035),
	.w7(32'hbaa484bf),
	.w8(32'hba68bc81),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec779a),
	.w1(32'h3abaae92),
	.w2(32'h3a59e679),
	.w3(32'h392b2e0d),
	.w4(32'hbaf0dced),
	.w5(32'hbaed6553),
	.w6(32'h3ac174bf),
	.w7(32'hb812b369),
	.w8(32'hba8cc952),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39075bf7),
	.w1(32'hb93c8b15),
	.w2(32'hb8fbce0f),
	.w3(32'h380c6f6b),
	.w4(32'hb9a43c2a),
	.w5(32'hb92820cf),
	.w6(32'hb802f181),
	.w7(32'hb8c9a951),
	.w8(32'hb88417a7),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9730288),
	.w1(32'hb91cd604),
	.w2(32'h381b44dc),
	.w3(32'hb99c50c0),
	.w4(32'h38beee90),
	.w5(32'h38ce53ff),
	.w6(32'hb925fcc0),
	.w7(32'h37636ae1),
	.w8(32'hb5af781d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b074ca9),
	.w1(32'h3b191f92),
	.w2(32'h3a68aaef),
	.w3(32'h3b522f13),
	.w4(32'h3b1af445),
	.w5(32'h3b0a0bf8),
	.w6(32'h3ad3870a),
	.w7(32'h3af6c920),
	.w8(32'h3a8947cd),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f1bac),
	.w1(32'hbb188f32),
	.w2(32'h3a76ddc0),
	.w3(32'h3bd905f3),
	.w4(32'h3a991b12),
	.w5(32'h3acca491),
	.w6(32'h3bb3a35c),
	.w7(32'h3a78e742),
	.w8(32'h39d49237),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d1e72),
	.w1(32'hbbbee600),
	.w2(32'h3a4d6235),
	.w3(32'hbbf3f456),
	.w4(32'hba9a36ea),
	.w5(32'h3be53efc),
	.w6(32'hbb381138),
	.w7(32'h395e35aa),
	.w8(32'h3be3d72e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992bba4),
	.w1(32'hba93137f),
	.w2(32'hba67ef2b),
	.w3(32'h36e6641e),
	.w4(32'hba244fdb),
	.w5(32'hba8721f6),
	.w6(32'h3a56076c),
	.w7(32'h38aa7c6c),
	.w8(32'hb9d0ffc9),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa49ed),
	.w1(32'hbc0d3ec7),
	.w2(32'hbaa73a10),
	.w3(32'hbba7aa8c),
	.w4(32'hba6ad144),
	.w5(32'hbb22181c),
	.w6(32'h3bff8af4),
	.w7(32'h3c9e74e5),
	.w8(32'h3c8f3249),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e998f),
	.w1(32'h3b99cb44),
	.w2(32'h3b27ec67),
	.w3(32'h3c20924f),
	.w4(32'hb9f3190e),
	.w5(32'h3b518ef3),
	.w6(32'h3bfd95f7),
	.w7(32'hb9aac9cc),
	.w8(32'hbb979320),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86382c),
	.w1(32'hbb324554),
	.w2(32'h3a5c0aa1),
	.w3(32'hbb024124),
	.w4(32'h38cb373c),
	.w5(32'h3a987e05),
	.w6(32'hba980a3d),
	.w7(32'hbae391ad),
	.w8(32'hba54cdd0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4cc57),
	.w1(32'hb9090b20),
	.w2(32'h3828f763),
	.w3(32'hb8f03711),
	.w4(32'h38b45a59),
	.w5(32'hb8f2613e),
	.w6(32'hb9079464),
	.w7(32'hb8ada38a),
	.w8(32'hb7cf5f1e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3911ab1f),
	.w1(32'hb9940543),
	.w2(32'hb9afb741),
	.w3(32'h39991159),
	.w4(32'hb889ac47),
	.w5(32'hb9a9f11d),
	.w6(32'h3852b4d5),
	.w7(32'h37b8108c),
	.w8(32'hb9b03f50),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7657950),
	.w1(32'hb92ff036),
	.w2(32'h388895b8),
	.w3(32'hb74320ea),
	.w4(32'hb9345fc9),
	.w5(32'hb8e13881),
	.w6(32'hb872b38f),
	.w7(32'hb7320436),
	.w8(32'hb85d6399),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e05ed),
	.w1(32'hb71eed48),
	.w2(32'h3b579bab),
	.w3(32'hbaec8109),
	.w4(32'hb9e245e5),
	.w5(32'hbad05119),
	.w6(32'hbaba1451),
	.w7(32'h38e6add6),
	.w8(32'h3917ec5b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d60a7a),
	.w1(32'hb8b6c254),
	.w2(32'h3a329ca9),
	.w3(32'h3ac8dc70),
	.w4(32'h3aa092dd),
	.w5(32'h3ab8e03b),
	.w6(32'h3ad78a0e),
	.w7(32'hb9f12ae7),
	.w8(32'h3a6adf6c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf52427),
	.w1(32'h39b487bc),
	.w2(32'hbab3f3f8),
	.w3(32'h3b2bfd72),
	.w4(32'hbb545c90),
	.w5(32'hbae3861f),
	.w6(32'h3922e000),
	.w7(32'hbbb304ba),
	.w8(32'hbb5cb38f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a832eca),
	.w1(32'hb976c5e3),
	.w2(32'hb9fd58a6),
	.w3(32'h3ae7d068),
	.w4(32'h39d59f20),
	.w5(32'h399c3f87),
	.w6(32'h3a82a4c6),
	.w7(32'h3a4c59ac),
	.w8(32'h3a3de081),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc191f40),
	.w1(32'hb9e4c11e),
	.w2(32'hb9ed6ffa),
	.w3(32'hbb909175),
	.w4(32'hba1e3c07),
	.w5(32'hbb599868),
	.w6(32'h3b8f8b69),
	.w7(32'h3bc7eab0),
	.w8(32'h3b33ff94),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70ee76),
	.w1(32'hbbcaa333),
	.w2(32'hbb3a43a5),
	.w3(32'hbb07d9c8),
	.w4(32'hba417e15),
	.w5(32'h3a82fe1b),
	.w6(32'hba5c2c51),
	.w7(32'hb983bf20),
	.w8(32'h3a9b4b3e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84974a4),
	.w1(32'hb90c3197),
	.w2(32'h37cf52e7),
	.w3(32'hb85a02d1),
	.w4(32'hb8efb002),
	.w5(32'hb8506bd9),
	.w6(32'hb895694b),
	.w7(32'h370a052e),
	.w8(32'h38d9f928),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb097b8e),
	.w1(32'hb89dca18),
	.w2(32'h390fe1c1),
	.w3(32'h3a2fd981),
	.w4(32'h3b2b831b),
	.w5(32'hba883727),
	.w6(32'h3bbe39ff),
	.w7(32'h3b7cbebb),
	.w8(32'h3a9809a5),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cf6407),
	.w1(32'hb8a9b982),
	.w2(32'h38105d6b),
	.w3(32'h3698d309),
	.w4(32'hb54a8bca),
	.w5(32'h38e3009e),
	.w6(32'h3700736c),
	.w7(32'hb61b229e),
	.w8(32'h38bd4178),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39080243),
	.w1(32'h3b354cdd),
	.w2(32'h3b2b0366),
	.w3(32'hb93e1fb4),
	.w4(32'h3aec2914),
	.w5(32'h397e0830),
	.w6(32'h3b47b21e),
	.w7(32'h3b868f4d),
	.w8(32'h3ad5b586),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a9dc5),
	.w1(32'h3b6a10e9),
	.w2(32'h3b1e9a69),
	.w3(32'h3c0ab04e),
	.w4(32'h3b8f6c49),
	.w5(32'h3c0c6edd),
	.w6(32'h3b246107),
	.w7(32'hba959743),
	.w8(32'h3b0205a1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91ece6),
	.w1(32'h3ac8eb0c),
	.w2(32'h396e11e4),
	.w3(32'h3b93f73d),
	.w4(32'h3ab42c7a),
	.w5(32'h3aa83938),
	.w6(32'h3b891b85),
	.w7(32'h3a65752f),
	.w8(32'h3ac0fb70),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3d5da),
	.w1(32'hb790b780),
	.w2(32'h38f9d001),
	.w3(32'h3a0bc5c4),
	.w4(32'h39c445e5),
	.w5(32'h39a3608e),
	.w6(32'hba1cffe6),
	.w7(32'hb9fbb12f),
	.w8(32'hba1bb9f0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cf767),
	.w1(32'h3b5f8cb0),
	.w2(32'hba50dba1),
	.w3(32'h3bcf89f7),
	.w4(32'h39e9e504),
	.w5(32'hba4d9293),
	.w6(32'h3b8a2439),
	.w7(32'hba90c586),
	.w8(32'hbb14b468),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6944a),
	.w1(32'hbb060259),
	.w2(32'hba3853d2),
	.w3(32'hbb6fb5d0),
	.w4(32'hba3c8f0f),
	.w5(32'hbb042588),
	.w6(32'hbaa0fdbf),
	.w7(32'h3aba96ad),
	.w8(32'h3a0b1fe8),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25fe90),
	.w1(32'hbb80e8cd),
	.w2(32'hba9b5b48),
	.w3(32'hbbfba565),
	.w4(32'hbbe7936e),
	.w5(32'hbb60b7b2),
	.w6(32'h3ad5f3de),
	.w7(32'h3b779da4),
	.w8(32'h3b759d16),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a09903),
	.w1(32'h37eeac8f),
	.w2(32'h399b6c49),
	.w3(32'h396fd112),
	.w4(32'hb7ea505b),
	.w5(32'h39596de3),
	.w6(32'h391382c0),
	.w7(32'h398db2f0),
	.w8(32'h395e0680),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399645b4),
	.w1(32'h388944d8),
	.w2(32'h38eef6e9),
	.w3(32'h3934b182),
	.w4(32'hb83855de),
	.w5(32'h38f32ff6),
	.w6(32'h3a0828d7),
	.w7(32'h389d64ea),
	.w8(32'h3898f249),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba974d7),
	.w1(32'hbb83ba0d),
	.w2(32'h3b2fdc08),
	.w3(32'h3a565996),
	.w4(32'hb79e80e8),
	.w5(32'h3b40e8e3),
	.w6(32'h3b121661),
	.w7(32'h3c12626a),
	.w8(32'h3c16cc52),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd1458),
	.w1(32'h391ae3d2),
	.w2(32'h3ac399e2),
	.w3(32'h3a0b21bc),
	.w4(32'h3b5615c8),
	.w5(32'h3b05568c),
	.w6(32'hb9d74325),
	.w7(32'h3bd46d74),
	.w8(32'h3bc73d99),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7f193),
	.w1(32'h3aa8ee40),
	.w2(32'h39e96c60),
	.w3(32'h3bbc478b),
	.w4(32'h3b0bd798),
	.w5(32'h3a93958d),
	.w6(32'h3b8515af),
	.w7(32'h3adb6c09),
	.w8(32'h3af7a282),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bf809),
	.w1(32'h3a579d40),
	.w2(32'h3c20e317),
	.w3(32'hbb822ce5),
	.w4(32'h3bb15cee),
	.w5(32'h3c0a2f79),
	.w6(32'hba12ef53),
	.w7(32'h3bae47f4),
	.w8(32'h3ae31036),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4aa49),
	.w1(32'h39e4bc10),
	.w2(32'h396ded2c),
	.w3(32'h392ae6ca),
	.w4(32'hb8746ac0),
	.w5(32'hb8d41edd),
	.w6(32'hba465bef),
	.w7(32'hb98401d5),
	.w8(32'h384f6876),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2aedee),
	.w1(32'h38d2d42c),
	.w2(32'h3a260b1e),
	.w3(32'hbb0c39b6),
	.w4(32'hb9ec3bff),
	.w5(32'hb8c90bf8),
	.w6(32'hb9423af9),
	.w7(32'h389a665c),
	.w8(32'h39ca9c59),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b9103),
	.w1(32'hbc546af3),
	.w2(32'h3ba3610d),
	.w3(32'hbbc3b512),
	.w4(32'hbb5f66ef),
	.w5(32'h3bef13c5),
	.w6(32'hbba1093b),
	.w7(32'hbaf06a64),
	.w8(32'h3bcf456f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9077e7),
	.w1(32'hbbd5613b),
	.w2(32'h3989b51a),
	.w3(32'hbc033a91),
	.w4(32'hbb3e4028),
	.w5(32'hb9cfba5e),
	.w6(32'h3b9db6d8),
	.w7(32'h3c32e95e),
	.w8(32'h3c394f95),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a1261),
	.w1(32'hbb26134b),
	.w2(32'h3b662338),
	.w3(32'hbbd3a08f),
	.w4(32'h3b3a6d66),
	.w5(32'h3ac97fd4),
	.w6(32'hbac0636a),
	.w7(32'h3bc5b257),
	.w8(32'h3bb7ac94),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1ce33),
	.w1(32'h3b4490ed),
	.w2(32'h3b397aa8),
	.w3(32'h3b899336),
	.w4(32'hba8c0854),
	.w5(32'h3a9c1e76),
	.w6(32'h3a173ab8),
	.w7(32'hbb893795),
	.w8(32'hbacbc251),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf30796),
	.w1(32'h3b13a25b),
	.w2(32'hba515dfb),
	.w3(32'h3b6393fa),
	.w4(32'hbab0d4f5),
	.w5(32'h3ac78ace),
	.w6(32'h38826d68),
	.w7(32'hbbb451e6),
	.w8(32'hbb5054a0),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae6cc6),
	.w1(32'hb7878b2d),
	.w2(32'h37aba0b5),
	.w3(32'h397309f2),
	.w4(32'h36cb9f00),
	.w5(32'h3816a718),
	.w6(32'hb919c5b1),
	.w7(32'hb93d367c),
	.w8(32'hb926a27e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bcf2b4),
	.w1(32'hb89ab37b),
	.w2(32'hb8d53dc1),
	.w3(32'hb69aaaca),
	.w4(32'hb8a2688e),
	.w5(32'h37749c83),
	.w6(32'h369eb9bf),
	.w7(32'h38e74600),
	.w8(32'h3844e06d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d2dbe),
	.w1(32'h3b84941b),
	.w2(32'h3b9de0dd),
	.w3(32'hbb4998ca),
	.w4(32'hbb3534bd),
	.w5(32'hbb4f839e),
	.w6(32'h3941a79a),
	.w7(32'h3b08bc90),
	.w8(32'h3ad51599),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8659bc9),
	.w1(32'hb9406073),
	.w2(32'hb95e441e),
	.w3(32'hb95e22bb),
	.w4(32'h36a08d11),
	.w5(32'hb7b58a52),
	.w6(32'hb96e8b2f),
	.w7(32'hb918885a),
	.w8(32'h38032e60),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa5671),
	.w1(32'hbaaaa598),
	.w2(32'h39a594a0),
	.w3(32'hbb2a1307),
	.w4(32'hbb852d91),
	.w5(32'hbb4c1390),
	.w6(32'hbabc847e),
	.w7(32'hbb36adb0),
	.w8(32'hbae519be),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ae1f0),
	.w1(32'h3aad0327),
	.w2(32'h3ab42956),
	.w3(32'h3b24693e),
	.w4(32'h3b521b97),
	.w5(32'h3a13470e),
	.w6(32'hba182f4d),
	.w7(32'h3b58d275),
	.w8(32'h3b8d504d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adde91f),
	.w1(32'h3a5040e4),
	.w2(32'hb98f9e15),
	.w3(32'h3ad4d17d),
	.w4(32'h3a06ed11),
	.w5(32'hb930ded7),
	.w6(32'h3aa2788d),
	.w7(32'h3a438b84),
	.w8(32'h3a42f5e4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a425fd),
	.w1(32'hb815b6dc),
	.w2(32'hb9fb4650),
	.w3(32'h390e74f8),
	.w4(32'hb977fc83),
	.w5(32'hb9a04b72),
	.w6(32'h389c5545),
	.w7(32'hb898e70f),
	.w8(32'hb94e13b4),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c229f),
	.w1(32'hbb4ef946),
	.w2(32'h3b241296),
	.w3(32'hbc5d58d7),
	.w4(32'hbb1bae8b),
	.w5(32'hbad97333),
	.w6(32'hbbe9cfc6),
	.w7(32'h3bf89e90),
	.w8(32'h3c244b93),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac0431),
	.w1(32'hba019f28),
	.w2(32'h3a5e7cb5),
	.w3(32'hbb23e737),
	.w4(32'h39f96ed7),
	.w5(32'hba6f19d8),
	.w6(32'h3a941b37),
	.w7(32'h3b637d58),
	.w8(32'h3b0f745d),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73bab67),
	.w1(32'h390de4d5),
	.w2(32'h394a211f),
	.w3(32'h38a95b86),
	.w4(32'h39948f94),
	.w5(32'h3928f6fb),
	.w6(32'h37ed942c),
	.w7(32'h3912b3c4),
	.w8(32'h38e66f19),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ac14b),
	.w1(32'hbb9d391b),
	.w2(32'hba54ff93),
	.w3(32'hbbdfc511),
	.w4(32'hbb071495),
	.w5(32'hbaac3009),
	.w6(32'hbb15f9ce),
	.w7(32'h3ae06760),
	.w8(32'h3b13e2ef),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb8ea5),
	.w1(32'h3994a755),
	.w2(32'h39a303f4),
	.w3(32'h39948670),
	.w4(32'h39534961),
	.w5(32'h39037cd5),
	.w6(32'hb8f14aa7),
	.w7(32'hb8e1664e),
	.w8(32'hb9095013),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991e0f3),
	.w1(32'h392a4cd2),
	.w2(32'h39843b58),
	.w3(32'hb8a77aef),
	.w4(32'h3817ab1e),
	.w5(32'h398e1940),
	.w6(32'h37927571),
	.w7(32'h3a29b981),
	.w8(32'h3a622d36),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c2ccf2),
	.w1(32'h38200685),
	.w2(32'h37975c03),
	.w3(32'hb8902d37),
	.w4(32'h38a22be1),
	.w5(32'h38396319),
	.w6(32'h39684654),
	.w7(32'h39281489),
	.w8(32'h395b3aef),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395200e8),
	.w1(32'hb9278a44),
	.w2(32'h38e3221a),
	.w3(32'h39418fb4),
	.w4(32'hb8eeee8b),
	.w5(32'hb8224fd7),
	.w6(32'hb8ce88aa),
	.w7(32'hb7cfbf4c),
	.w8(32'hb8cc96bb),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29a82f),
	.w1(32'h3aad446b),
	.w2(32'h3b2dff8b),
	.w3(32'h3abbed81),
	.w4(32'hba4c51c1),
	.w5(32'h3ae7986c),
	.w6(32'h3a27eab7),
	.w7(32'hba902b7a),
	.w8(32'h3b00b489),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6965c0),
	.w1(32'h39fb7094),
	.w2(32'hbb510d38),
	.w3(32'hba659ae1),
	.w4(32'h3a6606b9),
	.w5(32'hbb1a9130),
	.w6(32'h3af742fb),
	.w7(32'h3a1b360c),
	.w8(32'hbb3f6ff5),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19b76d),
	.w1(32'hbbac6942),
	.w2(32'hbb2170b1),
	.w3(32'hbb617103),
	.w4(32'hb98287a5),
	.w5(32'hbb0318e6),
	.w6(32'h3ab2149a),
	.w7(32'h3b89bc69),
	.w8(32'h3aeea050),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc137c4e),
	.w1(32'hbb3cd600),
	.w2(32'h3a93276b),
	.w3(32'hbbbde031),
	.w4(32'hbb0bec4a),
	.w5(32'hbb0eb98c),
	.w6(32'h39d34874),
	.w7(32'h3b140af4),
	.w8(32'h39abc188),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f5b47),
	.w1(32'h3949074c),
	.w2(32'h3917590f),
	.w3(32'h39274227),
	.w4(32'h38498464),
	.w5(32'h38995eaa),
	.w6(32'h399f62ff),
	.w7(32'h3968ce1b),
	.w8(32'h394f8b5b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f1f64),
	.w1(32'h3a42c99e),
	.w2(32'hb8b0fcef),
	.w3(32'hb987a8c5),
	.w4(32'hb8b49e2a),
	.w5(32'hba4f4e85),
	.w6(32'h3a2b1fcd),
	.w7(32'h39eb1a5f),
	.w8(32'h392a678b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38745c83),
	.w1(32'hb90128bf),
	.w2(32'hb7e07b0c),
	.w3(32'h37a3fcbd),
	.w4(32'hb8869df5),
	.w5(32'hb7a8ccab),
	.w6(32'hb8855fa3),
	.w7(32'h370ce226),
	.w8(32'h388bb8f3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38162562),
	.w1(32'hb8cdfe4d),
	.w2(32'hb86e314d),
	.w3(32'h38d4eeed),
	.w4(32'hb6f46d6b),
	.w5(32'h37cab641),
	.w6(32'h38cb8341),
	.w7(32'h393d818c),
	.w8(32'h39406ff2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57e9bc),
	.w1(32'h3b408a3a),
	.w2(32'hb8e58dae),
	.w3(32'h3b666f24),
	.w4(32'h3b01a195),
	.w5(32'hbb4deb14),
	.w6(32'h3beb8b2e),
	.w7(32'h3b9b6f7d),
	.w8(32'h3ab42768),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3d9fa),
	.w1(32'hba14eaab),
	.w2(32'hb9842a4f),
	.w3(32'hba150d1d),
	.w4(32'hba10a990),
	.w5(32'hb93d3c06),
	.w6(32'hb9efabb4),
	.w7(32'hba0b0e3a),
	.w8(32'hba05a59a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6b2bb),
	.w1(32'h38f5c1d8),
	.w2(32'h39a94d0e),
	.w3(32'h3ab95a54),
	.w4(32'h3a5be5a2),
	.w5(32'h39f38d0b),
	.w6(32'h39f22d70),
	.w7(32'h3a22fcb0),
	.w8(32'h39879982),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5cb94),
	.w1(32'hba8843fa),
	.w2(32'hbac49d55),
	.w3(32'hb9a80b92),
	.w4(32'hba547f63),
	.w5(32'hb98ee3d0),
	.w6(32'h3a47f9ef),
	.w7(32'hba3b0cc8),
	.w8(32'hba03178e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92b15eb),
	.w1(32'hb852634a),
	.w2(32'hb7c68774),
	.w3(32'hb8cadca7),
	.w4(32'hb8239196),
	.w5(32'hb8ab3e79),
	.w6(32'h38e5dd85),
	.w7(32'h38efb9c6),
	.w8(32'h384220a5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b6455),
	.w1(32'h39d50da2),
	.w2(32'h3a014989),
	.w3(32'hb9e9fd4b),
	.w4(32'hb8d143fd),
	.w5(32'hba1c24cb),
	.w6(32'h3ab9ba83),
	.w7(32'h3b093fcc),
	.w8(32'h3aa24e6c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db7a4d),
	.w1(32'h395d932c),
	.w2(32'h361ef61e),
	.w3(32'h3989735c),
	.w4(32'hb7b4f6be),
	.w5(32'hb9558cb6),
	.w6(32'h3a06d8fd),
	.w7(32'h3912db19),
	.w8(32'hb6b7c09c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae721e7),
	.w1(32'h3b636941),
	.w2(32'hbb5f45cc),
	.w3(32'h3bae5a6e),
	.w4(32'h3a1494ba),
	.w5(32'hbb0d9141),
	.w6(32'h3bb8e882),
	.w7(32'h3b3fd47d),
	.w8(32'hbb1b0ff4),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93555ed),
	.w1(32'hb8a9ee8c),
	.w2(32'hb923a893),
	.w3(32'hba044856),
	.w4(32'hb9bf86c4),
	.w5(32'hba14d916),
	.w6(32'hb65fa35f),
	.w7(32'h3973c25a),
	.w8(32'hb92cb7f7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3afe27),
	.w1(32'hbc0522aa),
	.w2(32'hbb7fca4f),
	.w3(32'h3b92722d),
	.w4(32'h3b754788),
	.w5(32'h3a958cf1),
	.w6(32'h3b8504a1),
	.w7(32'h3bb2b754),
	.w8(32'h3b7e6d01),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule