module layer_10_featuremap_76(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1a6a7),
	.w1(32'hbc2fa7be),
	.w2(32'h3c2145ae),
	.w3(32'h3ba211da),
	.w4(32'h3b1c508b),
	.w5(32'hbbc68195),
	.w6(32'hbc69daaf),
	.w7(32'hbbeed694),
	.w8(32'hbc47fd9c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b291de8),
	.w1(32'hbb98c967),
	.w2(32'hbb7d7b14),
	.w3(32'h3c1b36b6),
	.w4(32'h3bf7529b),
	.w5(32'h3c8f1cef),
	.w6(32'h3aad8a8f),
	.w7(32'h3a637742),
	.w8(32'h3b939aa3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6eb123),
	.w1(32'hbba2fef8),
	.w2(32'h3c358186),
	.w3(32'h3c895258),
	.w4(32'hbc29e6a9),
	.w5(32'hbb81ba12),
	.w6(32'h3c683de3),
	.w7(32'h3bd3b4d4),
	.w8(32'h3c0e91cd),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6919ca),
	.w1(32'h3ba0922c),
	.w2(32'hbb9dcccd),
	.w3(32'h3bc3821c),
	.w4(32'h3c5c1dcf),
	.w5(32'h3b0e5395),
	.w6(32'h3bc2be4d),
	.w7(32'h39e5eba4),
	.w8(32'h3b8f517f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb776a0c),
	.w1(32'hbbcecb11),
	.w2(32'h3b8a7131),
	.w3(32'hbb520198),
	.w4(32'hbaec1916),
	.w5(32'h3c0350c3),
	.w6(32'h3bd8662a),
	.w7(32'hbb41c221),
	.w8(32'h3c447f2c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b8432),
	.w1(32'h3bb3ac7d),
	.w2(32'hbb6ebf7f),
	.w3(32'hbb82d745),
	.w4(32'h39e29278),
	.w5(32'h3ae60c3c),
	.w6(32'h3c602819),
	.w7(32'h3b4ce8ae),
	.w8(32'hba68096b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc668b4),
	.w1(32'hbb832f63),
	.w2(32'hbc1d7651),
	.w3(32'hbb2292c5),
	.w4(32'hb980190d),
	.w5(32'hbbc28075),
	.w6(32'hbb30b79a),
	.w7(32'h3a5d36f5),
	.w8(32'h3ba85b39),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42d0e3),
	.w1(32'hbbeda9a6),
	.w2(32'hbbf375b8),
	.w3(32'hbc892365),
	.w4(32'hbca67b01),
	.w5(32'hbce3e439),
	.w6(32'hbad0bd45),
	.w7(32'h39bde4d8),
	.w8(32'hbc43a7ec),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9841f2),
	.w1(32'hbb4ff713),
	.w2(32'hba54608c),
	.w3(32'hbcbf33aa),
	.w4(32'hbb881abc),
	.w5(32'hbb08494f),
	.w6(32'hbcd42f25),
	.w7(32'hbc3d525b),
	.w8(32'h3aed2cce),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e5c034),
	.w1(32'h3bc39cab),
	.w2(32'hb9731318),
	.w3(32'h3b172888),
	.w4(32'h3bd70113),
	.w5(32'h3bae8ca8),
	.w6(32'h3b94c602),
	.w7(32'h3bf7ba2d),
	.w8(32'h3bcc6e94),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd9f51),
	.w1(32'hb9f71940),
	.w2(32'h3bbaffd3),
	.w3(32'h3ad0d07d),
	.w4(32'hbaf78ae6),
	.w5(32'h3c180beb),
	.w6(32'h3c04ab80),
	.w7(32'h3ba349b9),
	.w8(32'h3b42c6ad),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6907f4),
	.w1(32'h3b17127a),
	.w2(32'h3b43e384),
	.w3(32'h3ccab6ea),
	.w4(32'h3c3ff019),
	.w5(32'h3ad98e12),
	.w6(32'h3ac88f39),
	.w7(32'h3c084e3e),
	.w8(32'h3b87e47e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11be85),
	.w1(32'h3adbb4b9),
	.w2(32'hbafa12b4),
	.w3(32'h3af55f32),
	.w4(32'h3b681d28),
	.w5(32'h3bc6e278),
	.w6(32'h3b58fa9c),
	.w7(32'h3ae6883e),
	.w8(32'h3c2e12c3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb10423),
	.w1(32'h3ba815bb),
	.w2(32'h3be21cca),
	.w3(32'h3c06216e),
	.w4(32'hba84f27d),
	.w5(32'h3b9a9a47),
	.w6(32'h3acc5d26),
	.w7(32'h3c166282),
	.w8(32'h3c6763d8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cebafda),
	.w1(32'h3d1da309),
	.w2(32'hbc82a06a),
	.w3(32'hbbd1ffaa),
	.w4(32'h3ce69b52),
	.w5(32'h3b8c6d5d),
	.w6(32'h3c592970),
	.w7(32'h3b31a45c),
	.w8(32'h3c41c4df),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6e69f),
	.w1(32'hbc011890),
	.w2(32'hba8ba7d2),
	.w3(32'hbc5d8370),
	.w4(32'hbc8e495c),
	.w5(32'h3b95274b),
	.w6(32'h3c264662),
	.w7(32'h3b08d8a6),
	.w8(32'h3bff4985),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb985437),
	.w1(32'hbb7ef130),
	.w2(32'hbbe45f3a),
	.w3(32'hbae1774a),
	.w4(32'hbb88df92),
	.w5(32'hbc125324),
	.w6(32'h3bb08d90),
	.w7(32'h3b0f0819),
	.w8(32'hbb6137a9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9e6b5),
	.w1(32'h3bbfa299),
	.w2(32'h3b3fa7dc),
	.w3(32'hbc543a49),
	.w4(32'h39a6fc36),
	.w5(32'hba428571),
	.w6(32'hbc337fea),
	.w7(32'hb97808a8),
	.w8(32'h3bdae2be),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af658e7),
	.w1(32'hbb10ba3d),
	.w2(32'h3bcc0ca9),
	.w3(32'hb9b25160),
	.w4(32'h3b347514),
	.w5(32'hbb5f425b),
	.w6(32'h3b04b0a4),
	.w7(32'h3b4b1c35),
	.w8(32'h3c8863a4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2c8c88),
	.w1(32'h3cad1c40),
	.w2(32'h3a3aa480),
	.w3(32'h3c6b431f),
	.w4(32'h3d13feae),
	.w5(32'h3a012c4a),
	.w6(32'h3bb95c8e),
	.w7(32'h3aba7baa),
	.w8(32'h3c0e6a42),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67f804),
	.w1(32'h3b85493d),
	.w2(32'hb9e2777a),
	.w3(32'h3b30ebc8),
	.w4(32'h3b8b54f9),
	.w5(32'hbb87f85c),
	.w6(32'h3a5d9ce2),
	.w7(32'h3b1ae446),
	.w8(32'h3c202c3a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf237a),
	.w1(32'hba6add5d),
	.w2(32'hbb6adb31),
	.w3(32'h3ac708d4),
	.w4(32'h3c0e4a2c),
	.w5(32'hbc6bf074),
	.w6(32'hbbd43683),
	.w7(32'h3b03f848),
	.w8(32'h3ba305d5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9743e8),
	.w1(32'hbc415ec3),
	.w2(32'hbacbc5fe),
	.w3(32'hbce403b2),
	.w4(32'hbc887279),
	.w5(32'h3a1e6734),
	.w6(32'hbc603c1e),
	.w7(32'hbca0251d),
	.w8(32'hbb052097),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94d531),
	.w1(32'hbb5aab5b),
	.w2(32'hba01660d),
	.w3(32'h3a0fa6ba),
	.w4(32'h3a809364),
	.w5(32'h3b31bd15),
	.w6(32'hbaeeea33),
	.w7(32'h393230c1),
	.w8(32'h3bd4d18f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60e172),
	.w1(32'hbb059067),
	.w2(32'h3c8b9e05),
	.w3(32'h3bd7d4a7),
	.w4(32'h3c442c2b),
	.w5(32'hbac9a090),
	.w6(32'h3b069a16),
	.w7(32'h3c2e73bb),
	.w8(32'h3c1f1e09),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce8e01b),
	.w1(32'h3c3ffcfe),
	.w2(32'h3c5e6c04),
	.w3(32'h3ab61985),
	.w4(32'h3ca0d0bb),
	.w5(32'h3c65828a),
	.w6(32'h3bd8794a),
	.w7(32'hb7fe7b12),
	.w8(32'h3b847c3b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c028789),
	.w1(32'h3bbe60cb),
	.w2(32'h3ae99c93),
	.w3(32'h3c76930c),
	.w4(32'h3c34661c),
	.w5(32'h3b38cb34),
	.w6(32'h3bb34e04),
	.w7(32'h3bdb1cdc),
	.w8(32'h3a923eea),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc2a07),
	.w1(32'h3a8cd59c),
	.w2(32'hbbd1ac45),
	.w3(32'h3b901466),
	.w4(32'h3b4a0b0f),
	.w5(32'hbb845754),
	.w6(32'h3a347388),
	.w7(32'h388688c7),
	.w8(32'hbc07079c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ccb65),
	.w1(32'hbc19fc4b),
	.w2(32'hbb843a03),
	.w3(32'h3b9249d3),
	.w4(32'hba84e9a4),
	.w5(32'h3ba7c87f),
	.w6(32'hba26124c),
	.w7(32'hbb80f44e),
	.w8(32'h3b91b586),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc684fc6),
	.w1(32'hbbd13a1d),
	.w2(32'hbad1bcb5),
	.w3(32'h39e0f169),
	.w4(32'hbc95e510),
	.w5(32'h3aa34c3a),
	.w6(32'h3c58c4fc),
	.w7(32'hbba35831),
	.w8(32'hba659b76),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f933ac),
	.w1(32'h39eb968a),
	.w2(32'hbac2044f),
	.w3(32'hba813bed),
	.w4(32'hb9990c8e),
	.w5(32'hbb65458a),
	.w6(32'hbaf006f4),
	.w7(32'hbb74a4ff),
	.w8(32'h3c60ac42),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8924bb),
	.w1(32'h3bacf191),
	.w2(32'hbbb4e202),
	.w3(32'hbc547dbb),
	.w4(32'hbb611bc1),
	.w5(32'hbbbbe160),
	.w6(32'hbc55d850),
	.w7(32'hbc90646e),
	.w8(32'hbb914a5f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9dd25),
	.w1(32'h38f1a42e),
	.w2(32'hbaf00ba3),
	.w3(32'hbb37cc36),
	.w4(32'hbb9b5559),
	.w5(32'h399b80e9),
	.w6(32'hbb9c6def),
	.w7(32'h3ab6638d),
	.w8(32'hba321099),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98181c1),
	.w1(32'hba632e85),
	.w2(32'hbbcd701e),
	.w3(32'hb9e335cc),
	.w4(32'hb9bb15a6),
	.w5(32'hbb6a01cb),
	.w6(32'h3a2bfd67),
	.w7(32'hba14fbea),
	.w8(32'h3ab3b89a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3985c8),
	.w1(32'hbb929541),
	.w2(32'hbbbd0491),
	.w3(32'hbcb26fb3),
	.w4(32'hbc8a03ec),
	.w5(32'hbb6b370e),
	.w6(32'hbc4ce344),
	.w7(32'hbcbeeafa),
	.w8(32'h3a1035a7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca881c),
	.w1(32'hb9b76634),
	.w2(32'hbb75f906),
	.w3(32'hbb938b44),
	.w4(32'hbab514f1),
	.w5(32'hbc0f7df1),
	.w6(32'hbb5d088f),
	.w7(32'hbadd6f88),
	.w8(32'hbb0336d2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b095af2),
	.w1(32'h3a191a07),
	.w2(32'hbc620c38),
	.w3(32'hbc473e24),
	.w4(32'hbb07c29c),
	.w5(32'hbbc8b9a9),
	.w6(32'hbc7166e6),
	.w7(32'hbc55e64c),
	.w8(32'hbc1f02e3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc63d3f),
	.w1(32'hbc1bba25),
	.w2(32'h3c4b253d),
	.w3(32'h3b5fecd1),
	.w4(32'h3ab16123),
	.w5(32'h3c432ecd),
	.w6(32'h3b552b22),
	.w7(32'h3afecfbc),
	.w8(32'h3c024c53),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5e17f),
	.w1(32'h39b429d7),
	.w2(32'hba0253cb),
	.w3(32'h3c1492fd),
	.w4(32'h3ab7cb82),
	.w5(32'h3bb13337),
	.w6(32'h3c88fdf7),
	.w7(32'h3ae3e95d),
	.w8(32'h3c01f456),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc819b),
	.w1(32'hbbbe2d94),
	.w2(32'h3a76b140),
	.w3(32'h3b8e66d3),
	.w4(32'hbb1ca5b6),
	.w5(32'hb9d11106),
	.w6(32'h3bd2fc24),
	.w7(32'hbac82724),
	.w8(32'h3bc3ab0d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba853f06),
	.w1(32'h3c216896),
	.w2(32'hbb4ec0ba),
	.w3(32'hb9f567c0),
	.w4(32'h3c172742),
	.w5(32'hbb4038af),
	.w6(32'h3b42d9a9),
	.w7(32'h3bfe0465),
	.w8(32'h3b5fa19e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0411b),
	.w1(32'hb7cbaee1),
	.w2(32'h3b1833d8),
	.w3(32'hbb457c6a),
	.w4(32'hbba05b1a),
	.w5(32'hbac1abd8),
	.w6(32'h3b4ae129),
	.w7(32'hbc22ddd9),
	.w8(32'h3b6dd233),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe46b59),
	.w1(32'hbb48d660),
	.w2(32'hbbd1c5d0),
	.w3(32'hbc3da600),
	.w4(32'hbc4a2d1b),
	.w5(32'hbbdc197a),
	.w6(32'hbb31fc3e),
	.w7(32'hbbec4a5a),
	.w8(32'hbb29bdaa),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1147df),
	.w1(32'hbac20267),
	.w2(32'hbae986fb),
	.w3(32'h3a0b07a2),
	.w4(32'h3b460963),
	.w5(32'h3a1cac0e),
	.w6(32'h3aa41111),
	.w7(32'h3b7652bf),
	.w8(32'h39066d1c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0688a3),
	.w1(32'hbb239b3f),
	.w2(32'hb9d9f952),
	.w3(32'h3b429d96),
	.w4(32'h3ad5f2ba),
	.w5(32'h39647425),
	.w6(32'h3ccc679a),
	.w7(32'h3c59d515),
	.w8(32'hbb24b407),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9891f2),
	.w1(32'h3ba09eef),
	.w2(32'hbc2be44c),
	.w3(32'h3bc8a076),
	.w4(32'h3c0e7251),
	.w5(32'hbb1df83f),
	.w6(32'h3bd03ae0),
	.w7(32'h3bafbc27),
	.w8(32'hbc0a93fb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61a534),
	.w1(32'h3b687f34),
	.w2(32'h397f91be),
	.w3(32'h3acfd65b),
	.w4(32'h3bed42cf),
	.w5(32'h3b9e24d9),
	.w6(32'hbba12c3a),
	.w7(32'h3c7c97dd),
	.w8(32'h3bbd74ad),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb975738),
	.w1(32'hbbdb7617),
	.w2(32'hbba5f965),
	.w3(32'h3b996877),
	.w4(32'h3932ac92),
	.w5(32'hbb0c3d6d),
	.w6(32'h3b3f877d),
	.w7(32'hbb105c0e),
	.w8(32'hba5b03a1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cc937),
	.w1(32'hbae49e62),
	.w2(32'h3ab03bf5),
	.w3(32'h3b06c012),
	.w4(32'h3b353989),
	.w5(32'hbbfee94f),
	.w6(32'h3b802134),
	.w7(32'h3b933df8),
	.w8(32'hbac16a3c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a53b0),
	.w1(32'hbb0aa9de),
	.w2(32'hbc8ce752),
	.w3(32'hbbe0a4b2),
	.w4(32'h3c0cd746),
	.w5(32'hbc8126d4),
	.w6(32'hba765ab7),
	.w7(32'hbb23bce3),
	.w8(32'hbcb1eb4a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce479e6),
	.w1(32'hbc97d37c),
	.w2(32'hbc1211d3),
	.w3(32'hbd179bec),
	.w4(32'hbcf7a2f2),
	.w5(32'hbc8c4e4e),
	.w6(32'hbce9dd21),
	.w7(32'hbcc0555d),
	.w8(32'hbb70c8da),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc341ce9),
	.w1(32'h3b2d69c2),
	.w2(32'hbba2f5b0),
	.w3(32'hbcc5a068),
	.w4(32'hbbd39229),
	.w5(32'hbc0c3bbc),
	.w6(32'hbc6c1c91),
	.w7(32'hbb5e14a1),
	.w8(32'hbc47af67),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc790858),
	.w1(32'hbc45f3a4),
	.w2(32'h3bd91993),
	.w3(32'hbca27e60),
	.w4(32'hbc2299eb),
	.w5(32'h3a9a88c2),
	.w6(32'hbcdb1c95),
	.w7(32'hbc333b89),
	.w8(32'h3b62e189),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5992b),
	.w1(32'h3c25ea6b),
	.w2(32'h3bfd2836),
	.w3(32'hba6fbcdf),
	.w4(32'h3b5f1b32),
	.w5(32'h3bc10d27),
	.w6(32'hbbc5d36d),
	.w7(32'hbb8a54c2),
	.w8(32'h3bfcce3b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc51375),
	.w1(32'h3b3d3007),
	.w2(32'hbb18fb3c),
	.w3(32'hbc062b52),
	.w4(32'hbc6968d2),
	.w5(32'hba87ff4b),
	.w6(32'h3b28e6ec),
	.w7(32'hbc092d60),
	.w8(32'h3b8204e1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1588c8),
	.w1(32'h3c0a6caa),
	.w2(32'hba2a16fb),
	.w3(32'hbb9eb755),
	.w4(32'hbaa0a2cf),
	.w5(32'h3a949852),
	.w6(32'hbc3a37c3),
	.w7(32'hb6ca191b),
	.w8(32'h3b96fab5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcc260),
	.w1(32'hbc8356d9),
	.w2(32'hbaa5fbaf),
	.w3(32'h3c1fc237),
	.w4(32'h3b7e1b15),
	.w5(32'hbb63d53c),
	.w6(32'h3aafe42b),
	.w7(32'h3c254c9b),
	.w8(32'hbbc92bcb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf26f55),
	.w1(32'hbbd630b9),
	.w2(32'h3a547ae5),
	.w3(32'hbb76962b),
	.w4(32'h39ef66ec),
	.w5(32'hbb187737),
	.w6(32'hbb3bb3be),
	.w7(32'hbad8d479),
	.w8(32'h3b93d2f5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d2b02),
	.w1(32'hbb4ce23e),
	.w2(32'h3c19bbc3),
	.w3(32'hba995d51),
	.w4(32'h390e152b),
	.w5(32'h3b3b3dd5),
	.w6(32'h3beee93a),
	.w7(32'h3c1656c1),
	.w8(32'h3ab4d69e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bcb9f),
	.w1(32'h3b521c50),
	.w2(32'hbb93fcc9),
	.w3(32'hb8004c94),
	.w4(32'h3ab2fd68),
	.w5(32'hbb503034),
	.w6(32'h3b1a5e95),
	.w7(32'h3a39800e),
	.w8(32'h3b8ae523),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83bda7),
	.w1(32'h3bc05ffb),
	.w2(32'h3bd8bb51),
	.w3(32'hbb811236),
	.w4(32'h3ae37584),
	.w5(32'hba0525c9),
	.w6(32'hbba062ba),
	.w7(32'hbb5a1f95),
	.w8(32'hbb946bfc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92a92c),
	.w1(32'h3bcb0abe),
	.w2(32'hba51f6f9),
	.w3(32'h3cfbe276),
	.w4(32'h3cdaa552),
	.w5(32'h3b0abd86),
	.w6(32'h3c52d14d),
	.w7(32'h3cd7518f),
	.w8(32'hbb94aa26),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87a573),
	.w1(32'hbb8fef80),
	.w2(32'hbaae5a2e),
	.w3(32'h3bffe3c2),
	.w4(32'h3b6c93b0),
	.w5(32'h3aedf7b8),
	.w6(32'h3c1fad9c),
	.w7(32'h3bd5153f),
	.w8(32'h3c4d9877),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b434715),
	.w1(32'h3befacb1),
	.w2(32'h3bb88367),
	.w3(32'h3968054d),
	.w4(32'h3aa40bc9),
	.w5(32'h3bcb230f),
	.w6(32'h3ba3db1c),
	.w7(32'h3a118d1a),
	.w8(32'h3bf7853d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc38025),
	.w1(32'h3c15bea5),
	.w2(32'h3b912006),
	.w3(32'h3ae31b50),
	.w4(32'h3bd1dbf8),
	.w5(32'h3a7ee14d),
	.w6(32'hbc2c1e9e),
	.w7(32'hbb089b4f),
	.w8(32'h3b09edc0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa26ead),
	.w1(32'hbbbedad2),
	.w2(32'hbc283742),
	.w3(32'h3b8fc5b8),
	.w4(32'hb9da5fe1),
	.w5(32'hbc2a695b),
	.w6(32'h3c01a12a),
	.w7(32'h3b75576b),
	.w8(32'hbc12adce),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e34b0),
	.w1(32'hbc01f0b6),
	.w2(32'hbc750d71),
	.w3(32'hb9365921),
	.w4(32'hba1173d9),
	.w5(32'hbc3759b2),
	.w6(32'hbb997fe4),
	.w7(32'hbb0a6b94),
	.w8(32'hbb6831e6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98376c),
	.w1(32'h3a9afb0e),
	.w2(32'h3b2ba86c),
	.w3(32'hbcef0edc),
	.w4(32'hbc34dc64),
	.w5(32'h3baba114),
	.w6(32'hbcceb6dc),
	.w7(32'hbc815517),
	.w8(32'h3ba5132c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bacf4),
	.w1(32'h3b80efd3),
	.w2(32'h3c2a4609),
	.w3(32'h3b9a8560),
	.w4(32'h3b66bb50),
	.w5(32'h3c1b4be4),
	.w6(32'h3bc1b770),
	.w7(32'h3ba9a88e),
	.w8(32'h3c33cfc7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d3f72),
	.w1(32'h3c094eb6),
	.w2(32'hbc773538),
	.w3(32'h3c9f9f77),
	.w4(32'h3c0ba4f9),
	.w5(32'hbb2644c3),
	.w6(32'h3cb107a5),
	.w7(32'h3c5a91cb),
	.w8(32'hbb90905c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ec154),
	.w1(32'hbc6ee42a),
	.w2(32'h3c0415dc),
	.w3(32'h3b69a613),
	.w4(32'hbb6a0623),
	.w5(32'h3b8ddcdd),
	.w6(32'hbb8d1ba9),
	.w7(32'hba197371),
	.w8(32'hbb7d2928),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83df96),
	.w1(32'hbbce2b96),
	.w2(32'hbcdbd457),
	.w3(32'h3bd5c225),
	.w4(32'hbb8070e6),
	.w5(32'hbcd7dfea),
	.w6(32'h39ed46a7),
	.w7(32'h3a2a5dcb),
	.w8(32'hbc5d3543),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9102bd),
	.w1(32'h3b37ac37),
	.w2(32'hbb609025),
	.w3(32'hbd17c19b),
	.w4(32'hbc5cc9d2),
	.w5(32'h3b44597e),
	.w6(32'hbcda5c47),
	.w7(32'hbca7b1a9),
	.w8(32'h3b50ce83),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1ed88),
	.w1(32'hbba0a835),
	.w2(32'hbb243dab),
	.w3(32'hba2302e4),
	.w4(32'hbb1d9df6),
	.w5(32'h3abc164c),
	.w6(32'h3bd736e8),
	.w7(32'h3ae071e5),
	.w8(32'h3b6b0f6f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1803ca),
	.w1(32'h3b156d5b),
	.w2(32'hbc05049f),
	.w3(32'h3a7e8280),
	.w4(32'h3b46dd5c),
	.w5(32'hbc0ae24c),
	.w6(32'h3a2b7677),
	.w7(32'h38e0539a),
	.w8(32'hbbe931ee),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd98e2d),
	.w1(32'hbb43302a),
	.w2(32'hbbd23847),
	.w3(32'hbc80713d),
	.w4(32'hbbeae816),
	.w5(32'hbc296fc2),
	.w6(32'hbc264aa6),
	.w7(32'hbc3bd365),
	.w8(32'hbc1ef379),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bacce),
	.w1(32'hbc070112),
	.w2(32'hbc24bd93),
	.w3(32'hbcbedb18),
	.w4(32'hbc3cf0e0),
	.w5(32'hbca76471),
	.w6(32'hbc70c243),
	.w7(32'hbc379360),
	.w8(32'hbc18fd10),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f37e4),
	.w1(32'hbbedcb25),
	.w2(32'h3c1f5e3b),
	.w3(32'hbd36fda8),
	.w4(32'hbcbad289),
	.w5(32'h3bf8d705),
	.w6(32'hbcd08d28),
	.w7(32'hbd03ebd3),
	.w8(32'hb9bc4847),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbddf9c),
	.w1(32'hba508942),
	.w2(32'h3b812e4b),
	.w3(32'h3c8c56bf),
	.w4(32'h3c20f4a5),
	.w5(32'h3b0cec32),
	.w6(32'h3c50b550),
	.w7(32'h3c8165bb),
	.w8(32'h3a9dca9d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b610d13),
	.w1(32'h3afa9aef),
	.w2(32'h3b20ee70),
	.w3(32'h3bd43c3b),
	.w4(32'h3b6def16),
	.w5(32'h3afd3c93),
	.w6(32'h3b40e716),
	.w7(32'h3aa4e394),
	.w8(32'h3b845a5d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94587a),
	.w1(32'hbada3718),
	.w2(32'h3b1bd89b),
	.w3(32'hbb04962c),
	.w4(32'hbb12c7b4),
	.w5(32'h3b4e4842),
	.w6(32'hbb8f5887),
	.w7(32'hbb4e46e4),
	.w8(32'h3b744194),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf6a33),
	.w1(32'h3ba10446),
	.w2(32'hbc01c5af),
	.w3(32'h3be08812),
	.w4(32'h3bc5d864),
	.w5(32'hbbeb67cc),
	.w6(32'h3b6ea4af),
	.w7(32'hba83c006),
	.w8(32'hbadf192b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ecaec),
	.w1(32'h3b8401c3),
	.w2(32'h3bb3fc48),
	.w3(32'hbc81b4ec),
	.w4(32'hbba1cef6),
	.w5(32'hbad746ac),
	.w6(32'hbc9374a2),
	.w7(32'hbc7c6d7f),
	.w8(32'hbc4cf730),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd25351),
	.w1(32'h3befd102),
	.w2(32'hbb98aa24),
	.w3(32'h3c131d14),
	.w4(32'h3c399135),
	.w5(32'hbc96ca19),
	.w6(32'h3b58d10d),
	.w7(32'h3c394ada),
	.w8(32'hbbc82cee),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c2185),
	.w1(32'h3a43fdd7),
	.w2(32'hba01eb49),
	.w3(32'hbbb23754),
	.w4(32'h3bf8aac4),
	.w5(32'hbc4127b5),
	.w6(32'hbc42be62),
	.w7(32'h3b9ae7fb),
	.w8(32'hbbb38a71),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31223d),
	.w1(32'h3c163d5b),
	.w2(32'hba636b6c),
	.w3(32'hba109601),
	.w4(32'h3c4e58fa),
	.w5(32'hbb9f3b46),
	.w6(32'hbc7afea0),
	.w7(32'h3b936f5c),
	.w8(32'hbb17d506),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb124df2),
	.w1(32'h3b3f47ba),
	.w2(32'h3b680292),
	.w3(32'hba68faca),
	.w4(32'h3baaa181),
	.w5(32'h3a8f44be),
	.w6(32'hbaea2821),
	.w7(32'h3b412b03),
	.w8(32'h3b0ae66e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae445b),
	.w1(32'h3b97fb9d),
	.w2(32'hbc867694),
	.w3(32'hba471c29),
	.w4(32'h3b0182ce),
	.w5(32'hbc8c8381),
	.w6(32'hb823eda2),
	.w7(32'h3a84954c),
	.w8(32'hbc7d19b1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd2aac4),
	.w1(32'hbc0ab10c),
	.w2(32'hbad23b60),
	.w3(32'hbd016e77),
	.w4(32'hbcca9f6f),
	.w5(32'h3a0dd78d),
	.w6(32'hbccd69e5),
	.w7(32'hbc91f6eb),
	.w8(32'h3bb74db3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b573276),
	.w1(32'h3c45c1c1),
	.w2(32'hbb94bf0b),
	.w3(32'hbc14ea4d),
	.w4(32'h3b11f635),
	.w5(32'hbb98d626),
	.w6(32'hbc234836),
	.w7(32'hbc250889),
	.w8(32'h3b68672c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ababbc9),
	.w1(32'hbb04337b),
	.w2(32'hba7b11eb),
	.w3(32'h3bbb261c),
	.w4(32'h3acb7a9a),
	.w5(32'hbb862efd),
	.w6(32'h3c0379c5),
	.w7(32'h3b405b4c),
	.w8(32'hbc284cca),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5228a),
	.w1(32'hbc0c7118),
	.w2(32'h3afa1c16),
	.w3(32'h3bd918b0),
	.w4(32'h3aee3af0),
	.w5(32'h3b03d8af),
	.w6(32'hbbd46c0b),
	.w7(32'hbba8bc59),
	.w8(32'h39b94828),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b703dd9),
	.w1(32'hb94bd49a),
	.w2(32'hbb5fe78b),
	.w3(32'h3bba589f),
	.w4(32'h3b5acc0e),
	.w5(32'hbbac509c),
	.w6(32'h3bd5575e),
	.w7(32'h3c0334de),
	.w8(32'hbb879b11),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12bab2),
	.w1(32'hbad3620e),
	.w2(32'h3bbd3aef),
	.w3(32'hbac3e058),
	.w4(32'hba7a644c),
	.w5(32'h3c0026d7),
	.w6(32'hbb94b016),
	.w7(32'hbb6b23af),
	.w8(32'h3adc7050),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6ec10),
	.w1(32'h3b9647a8),
	.w2(32'hbc388d74),
	.w3(32'h3b5ecef1),
	.w4(32'h3c007be2),
	.w5(32'hbbbaf1d6),
	.w6(32'h3c13a7d5),
	.w7(32'h3be4e07a),
	.w8(32'h3a35a867),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7a01f),
	.w1(32'hbb47a20f),
	.w2(32'hbb3da0a3),
	.w3(32'hbab97410),
	.w4(32'hbb9f5c28),
	.w5(32'h38d5b97b),
	.w6(32'hbbb1326e),
	.w7(32'hbaddecfb),
	.w8(32'h3abe51fe),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39344dbf),
	.w1(32'h3a847c83),
	.w2(32'h3c5761ea),
	.w3(32'hbc8e913a),
	.w4(32'hbbb738d2),
	.w5(32'h3b9921bc),
	.w6(32'hbbb942c6),
	.w7(32'hbc23fbd3),
	.w8(32'hba7b85e1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb62221),
	.w1(32'h3b85ef7d),
	.w2(32'hbc228bb0),
	.w3(32'h3d2c3739),
	.w4(32'h3cf27fd4),
	.w5(32'hbc591e8f),
	.w6(32'h3cbf898a),
	.w7(32'h3d106415),
	.w8(32'hbb1952e6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8432f7),
	.w1(32'hb8c21efd),
	.w2(32'hbba5bc2e),
	.w3(32'hbd0a325f),
	.w4(32'hbc98362a),
	.w5(32'h3b7eedac),
	.w6(32'hbd07a06b),
	.w7(32'hbccddec7),
	.w8(32'hbb5867b2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38b8a8),
	.w1(32'h3b87abd2),
	.w2(32'hbb9cdb78),
	.w3(32'h3b83fbe1),
	.w4(32'h3c5c7c82),
	.w5(32'hbb4d9b59),
	.w6(32'hbb083782),
	.w7(32'h3c043881),
	.w8(32'h3c2ec362),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07da2c),
	.w1(32'h3b8bb5ba),
	.w2(32'hbaecc860),
	.w3(32'hbcf1d434),
	.w4(32'hbc874cc7),
	.w5(32'hbb60e4f1),
	.w6(32'hbc5ff8a4),
	.w7(32'hbcce0a5f),
	.w8(32'h3c8b758d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a357859),
	.w1(32'h3c667d19),
	.w2(32'hbb89227f),
	.w3(32'hbcddacfd),
	.w4(32'hbc9b6e3d),
	.w5(32'h3af29e9b),
	.w6(32'hbc2d46e8),
	.w7(32'hbcdd51db),
	.w8(32'h3b51ce2f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06d3bc),
	.w1(32'h3b843e96),
	.w2(32'hbb14cbd9),
	.w3(32'hba1a06f9),
	.w4(32'h3b4d6394),
	.w5(32'hbb03ef3f),
	.w6(32'h3b78eb82),
	.w7(32'h394b7667),
	.w8(32'h3c404945),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13a897),
	.w1(32'h3c3f7824),
	.w2(32'h3b964805),
	.w3(32'hbc0dbb88),
	.w4(32'h3b3e0917),
	.w5(32'hb953fcbe),
	.w6(32'hba7fe45b),
	.w7(32'h3bb27698),
	.w8(32'h3ab839cb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a5218),
	.w1(32'h3c47d26e),
	.w2(32'h3bb59906),
	.w3(32'h3b7b2ea8),
	.w4(32'h3c5b70c1),
	.w5(32'h3a01672b),
	.w6(32'hbb89996b),
	.w7(32'h3ba02120),
	.w8(32'h3ba64da7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babcd5c),
	.w1(32'h3c1af6ba),
	.w2(32'h3b32ec54),
	.w3(32'h3b134550),
	.w4(32'h3c1f6294),
	.w5(32'hba831d49),
	.w6(32'hbb4123fa),
	.w7(32'h3bb194b1),
	.w8(32'hb9b6ab09),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7695a5),
	.w1(32'h3886d1be),
	.w2(32'h3b2238f9),
	.w3(32'h3bd363b7),
	.w4(32'h3bf4e12e),
	.w5(32'h3b0dbc7a),
	.w6(32'h3ada1de2),
	.w7(32'h3be83483),
	.w8(32'hbbdce199),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcad5c3),
	.w1(32'hba816bee),
	.w2(32'h3ac81fb9),
	.w3(32'h3c7a28da),
	.w4(32'h3c6a0eef),
	.w5(32'hbc14ffe8),
	.w6(32'h3ad5c30d),
	.w7(32'h3c65ab78),
	.w8(32'hbc80958b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a521531),
	.w1(32'hbbe689d3),
	.w2(32'h3ade47df),
	.w3(32'hbb6391a8),
	.w4(32'h3b101e14),
	.w5(32'h3c02ceec),
	.w6(32'hbbbf32cc),
	.w7(32'h3c28c937),
	.w8(32'h3c47a6de),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97246a),
	.w1(32'h3aeb02e1),
	.w2(32'h3c0e42b1),
	.w3(32'hbb5fd1ac),
	.w4(32'hbbee395c),
	.w5(32'h3c562c3a),
	.w6(32'h39a2f760),
	.w7(32'hbb8a25f7),
	.w8(32'h3b6d10c2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee7dc2),
	.w1(32'h3bad2407),
	.w2(32'hbbdf14c1),
	.w3(32'h3ceb61b0),
	.w4(32'h3c476df8),
	.w5(32'hbb977701),
	.w6(32'h3cd271bb),
	.w7(32'h3c75c6f4),
	.w8(32'h3b2c866f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae98b3),
	.w1(32'h3b508aaa),
	.w2(32'hbc194418),
	.w3(32'h39af8d05),
	.w4(32'h3b95543a),
	.w5(32'hbbcd04b4),
	.w6(32'hbafbedfe),
	.w7(32'h3bbc64b7),
	.w8(32'hb9c53641),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaca15),
	.w1(32'hbb9b4017),
	.w2(32'h3c436245),
	.w3(32'hbbc4bd3c),
	.w4(32'hbc3d120d),
	.w5(32'h3c58a641),
	.w6(32'hbc229487),
	.w7(32'hbc5c9220),
	.w8(32'h3bc4db26),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dbed4),
	.w1(32'h3ba4d737),
	.w2(32'hbc324c76),
	.w3(32'h3ca216eb),
	.w4(32'h3c0bb520),
	.w5(32'hbc019ba9),
	.w6(32'h3c8df182),
	.w7(32'h3c90ab42),
	.w8(32'h3b40f426),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf25fe),
	.w1(32'hbb9d17b5),
	.w2(32'h3a96f731),
	.w3(32'hbc23422a),
	.w4(32'hbc28d2e7),
	.w5(32'hbb14dd73),
	.w6(32'hb9cfcfeb),
	.w7(32'hbbe37a9d),
	.w8(32'hbb938067),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b1d9f),
	.w1(32'h38378b09),
	.w2(32'hbc36dc3f),
	.w3(32'h3b9a483e),
	.w4(32'h3b425c30),
	.w5(32'hbc17cf3b),
	.w6(32'h3b6668db),
	.w7(32'h3b1b9c8e),
	.w8(32'hbc3eb97a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0add35),
	.w1(32'h3aa6a40e),
	.w2(32'h3be8dec4),
	.w3(32'hbab5e8a9),
	.w4(32'hbb00e3b4),
	.w5(32'hb99a65d4),
	.w6(32'hbbe909a1),
	.w7(32'hbb96b5c4),
	.w8(32'h3c0477fb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e9e8a),
	.w1(32'h3b64eaf0),
	.w2(32'hbc32b765),
	.w3(32'hbb0e7203),
	.w4(32'hbb4e49f4),
	.w5(32'hbc21f2aa),
	.w6(32'h3bd132c7),
	.w7(32'h3bc60da1),
	.w8(32'h3bd2aca6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a8152),
	.w1(32'h3bf6c830),
	.w2(32'hbbb718cd),
	.w3(32'hbd048c95),
	.w4(32'hbc9afe2c),
	.w5(32'hbbff5c57),
	.w6(32'hbc81ec76),
	.w7(32'hbcc57521),
	.w8(32'h3c6642d7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc17c6c),
	.w1(32'h3c31e120),
	.w2(32'hbb3d95b4),
	.w3(32'hbceb9c16),
	.w4(32'hbc5fa52f),
	.w5(32'hbbc31e3e),
	.w6(32'hbc48bdab),
	.w7(32'hbd09f39d),
	.w8(32'hba40d6ac),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb782de),
	.w1(32'hbc344c66),
	.w2(32'h3aaae006),
	.w3(32'h3b57965d),
	.w4(32'hbaad8e68),
	.w5(32'h3b3953a5),
	.w6(32'h3c009f48),
	.w7(32'h3b97d86e),
	.w8(32'h3b7490e2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13161f),
	.w1(32'h3b802a76),
	.w2(32'hbb87ff17),
	.w3(32'h3b39849c),
	.w4(32'h3a9c3eed),
	.w5(32'hba9fb532),
	.w6(32'h3b0146a1),
	.w7(32'h3b2cd549),
	.w8(32'hba0f5006),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d8b2a),
	.w1(32'h3a0b1c8c),
	.w2(32'hba62480b),
	.w3(32'hbbc0b14b),
	.w4(32'hbad34532),
	.w5(32'h3b0669b1),
	.w6(32'hbb42d064),
	.w7(32'hbae68fd0),
	.w8(32'h3b9e33cd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc734805),
	.w1(32'hba095088),
	.w2(32'h3ba3d8b3),
	.w3(32'hbbd744c2),
	.w4(32'hbbbbdb55),
	.w5(32'h3b940545),
	.w6(32'h3b92a28f),
	.w7(32'hbbb94206),
	.w8(32'h3b811fd7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8b2b5),
	.w1(32'h3b9d7613),
	.w2(32'hbcaff436),
	.w3(32'h3ba90cc5),
	.w4(32'h3ba34c30),
	.w5(32'hbc9a5766),
	.w6(32'h3b571e1f),
	.w7(32'h3b93d311),
	.w8(32'hbc1a7edd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb57b58),
	.w1(32'hbc0099bb),
	.w2(32'hbcf79d3e),
	.w3(32'hbd1644b6),
	.w4(32'hbc79acc6),
	.w5(32'hbc650356),
	.w6(32'hbca89ed6),
	.w7(32'hbc911759),
	.w8(32'hbb72429b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40dcd5),
	.w1(32'h3b585f3c),
	.w2(32'hbcc69337),
	.w3(32'hbcde6ed3),
	.w4(32'hbb62d788),
	.w5(32'hbcbf9c46),
	.w6(32'hbca1c416),
	.w7(32'hbc975932),
	.w8(32'hbc8ae2b3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba54ad),
	.w1(32'h3baa9698),
	.w2(32'h3c5f97f5),
	.w3(32'hbd3b009f),
	.w4(32'hbc633b27),
	.w5(32'h3c060716),
	.w6(32'hbd1eeb4e),
	.w7(32'hbca0e2ca),
	.w8(32'hb9363573),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c903842),
	.w1(32'hbb25d194),
	.w2(32'hbaf77e52),
	.w3(32'h3c3c0643),
	.w4(32'h3c1db2f7),
	.w5(32'hbb8c4742),
	.w6(32'h3a8047c1),
	.w7(32'h3c3a1a78),
	.w8(32'h3a1de183),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc16a41),
	.w1(32'hbc5f78c4),
	.w2(32'hbb19dc7d),
	.w3(32'h3c6c6d4d),
	.w4(32'h3c3f6f4d),
	.w5(32'h3ab798cb),
	.w6(32'hbc078954),
	.w7(32'h3b7d3d57),
	.w8(32'h39f4271c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11072e),
	.w1(32'hbb0de886),
	.w2(32'h3ab818f4),
	.w3(32'h3ae24a5e),
	.w4(32'hbbb4ecee),
	.w5(32'hbaf4f312),
	.w6(32'h3ad7d847),
	.w7(32'hbbe5f916),
	.w8(32'hbbad3a60),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50ea97),
	.w1(32'h3a43e32c),
	.w2(32'hbc23f46c),
	.w3(32'hbca033bb),
	.w4(32'hbc92f88f),
	.w5(32'hbc895b25),
	.w6(32'hbbeed280),
	.w7(32'hbc4a6dcb),
	.w8(32'hbb378788),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3edc3),
	.w1(32'hbbb25a52),
	.w2(32'hbc06e655),
	.w3(32'hbcfbde59),
	.w4(32'hbc3b4aa1),
	.w5(32'hbc8d7d38),
	.w6(32'hbc890af7),
	.w7(32'hbcc1524b),
	.w8(32'hbbee28f7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29ac19),
	.w1(32'h3c04854e),
	.w2(32'hb67e0535),
	.w3(32'hbc701af7),
	.w4(32'hbbe23e52),
	.w5(32'h390aca6a),
	.w6(32'hbbd94852),
	.w7(32'h3b4f1377),
	.w8(32'h3b7d17a2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962ae09),
	.w1(32'h3bc282bd),
	.w2(32'h39cc8270),
	.w3(32'hb8352b83),
	.w4(32'h3bac5bf5),
	.w5(32'h3970a1e9),
	.w6(32'hbb01b604),
	.w7(32'hbae089a3),
	.w8(32'h3b8c150b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4275b),
	.w1(32'hb7844f5a),
	.w2(32'h3c0b0205),
	.w3(32'hbbb64c2e),
	.w4(32'hbbbab37d),
	.w5(32'h377b238f),
	.w6(32'hba032b3d),
	.w7(32'hbb9489b1),
	.w8(32'h3b19e31b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be95613),
	.w1(32'hbb8600ac),
	.w2(32'h3c030e7d),
	.w3(32'h3c4f169d),
	.w4(32'hba2f8105),
	.w5(32'h3a8f4793),
	.w6(32'h3c60f469),
	.w7(32'h3bcb62e4),
	.w8(32'hbae2dfbf),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85cd21),
	.w1(32'h3b55b3af),
	.w2(32'h3a37b34f),
	.w3(32'h3b0f154b),
	.w4(32'hb7b5ff26),
	.w5(32'h3afda98a),
	.w6(32'h398959d5),
	.w7(32'h3a7a0189),
	.w8(32'h3addfb7d),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcb88c),
	.w1(32'h3b17dace),
	.w2(32'hba4b5114),
	.w3(32'h3acd5756),
	.w4(32'h3b305743),
	.w5(32'hbbd48c4b),
	.w6(32'h3b1741ef),
	.w7(32'h3ad6bc06),
	.w8(32'hbad60336),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3baa31),
	.w1(32'h3b2c10e8),
	.w2(32'h3a6aa267),
	.w3(32'hbc691ce5),
	.w4(32'hbc365481),
	.w5(32'h3a0edf64),
	.w6(32'hbc88c60d),
	.w7(32'hbc75590b),
	.w8(32'hba718e6a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4d05d),
	.w1(32'h39c479b0),
	.w2(32'hbb98c090),
	.w3(32'h3b5631e7),
	.w4(32'h3b086228),
	.w5(32'h39f8d925),
	.w6(32'h3b0ff1e3),
	.w7(32'h3b269b6f),
	.w8(32'hbb67cf79),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb883f35),
	.w1(32'hbb5fd275),
	.w2(32'h3c08b0e4),
	.w3(32'hb9da2ae0),
	.w4(32'h3b6bc212),
	.w5(32'h3c38738b),
	.w6(32'hbb218e92),
	.w7(32'h3b958c70),
	.w8(32'h3c929fe5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb145f),
	.w1(32'hbabb2662),
	.w2(32'h3b9015a6),
	.w3(32'hbc052e05),
	.w4(32'hbcc69e4e),
	.w5(32'hbb4c116d),
	.w6(32'h3b28414c),
	.w7(32'hbc331f94),
	.w8(32'h3bbc67fe),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b167824),
	.w1(32'hb9c9292c),
	.w2(32'h3a8c92b1),
	.w3(32'h3a0dbe93),
	.w4(32'hbbad6488),
	.w5(32'h39d65bb3),
	.w6(32'h3ba0bd8a),
	.w7(32'h3b7ff04c),
	.w8(32'hb9663b0c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25e72d),
	.w1(32'h3aee9eb3),
	.w2(32'h3beca9c9),
	.w3(32'h3b38fe51),
	.w4(32'h3b0cc511),
	.w5(32'h3c22c2cf),
	.w6(32'h38e3d32e),
	.w7(32'hba097688),
	.w8(32'h3c705028),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5936cb),
	.w1(32'h3b8cc719),
	.w2(32'hba38041e),
	.w3(32'h3bd52958),
	.w4(32'h3ad33ba2),
	.w5(32'hbbb42cbb),
	.w6(32'h3c180868),
	.w7(32'h3a672e7d),
	.w8(32'hbc12a275),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd18c4f),
	.w1(32'hbb7e68da),
	.w2(32'h3bcb50bc),
	.w3(32'hbb9e4088),
	.w4(32'h385c21d5),
	.w5(32'h3b8bf590),
	.w6(32'hbb1c3164),
	.w7(32'hbb51fa86),
	.w8(32'hbb98eca4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c9978),
	.w1(32'h3b49d315),
	.w2(32'hbb3dded1),
	.w3(32'h3c737a45),
	.w4(32'h3c5ac715),
	.w5(32'h3abdaddb),
	.w6(32'h3be6045f),
	.w7(32'h3c93c242),
	.w8(32'h3bc83c45),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f27d8),
	.w1(32'h3b379bfb),
	.w2(32'h3c612cc3),
	.w3(32'hbbaffbcf),
	.w4(32'h3b2becf9),
	.w5(32'h3c348383),
	.w6(32'hba2c1724),
	.w7(32'h3b513266),
	.w8(32'hbb13557c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5c9d4),
	.w1(32'h3baf15ca),
	.w2(32'h3bb8e724),
	.w3(32'h3d0be501),
	.w4(32'h3cef148b),
	.w5(32'hb9e51d8e),
	.w6(32'h3cc8d4e9),
	.w7(32'h3d049751),
	.w8(32'hbb1a067c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02ee61),
	.w1(32'h3aa2d132),
	.w2(32'h3b1754ad),
	.w3(32'h3c503605),
	.w4(32'h3c044024),
	.w5(32'h3baf99fd),
	.w6(32'h3bd056f4),
	.w7(32'h3bc7641d),
	.w8(32'h3b5c4d8d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad35490),
	.w1(32'h3b8050e1),
	.w2(32'h3b01ff27),
	.w3(32'h3aca5a1d),
	.w4(32'h3a7b81b9),
	.w5(32'hb9f3b49e),
	.w6(32'h3b4bfc9c),
	.w7(32'h3b38c26b),
	.w8(32'hba75b8f1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc59ae),
	.w1(32'h3b67fdf4),
	.w2(32'h3bedf04c),
	.w3(32'h3bb6368f),
	.w4(32'h3ae4fd20),
	.w5(32'hbb43f632),
	.w6(32'h3b792994),
	.w7(32'h3ae92bbc),
	.w8(32'hbbf3e77d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a161d),
	.w1(32'hbb9de685),
	.w2(32'hbbae8dec),
	.w3(32'hba264b61),
	.w4(32'h3af5113a),
	.w5(32'hbc8a428d),
	.w6(32'hbbdd6bcd),
	.w7(32'hbb92cf61),
	.w8(32'hbb9dd397),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe760fb),
	.w1(32'hbc24439b),
	.w2(32'h3a997679),
	.w3(32'hbcc28f6b),
	.w4(32'hbc47d8d9),
	.w5(32'hba01c0c8),
	.w6(32'hbcab7fcc),
	.w7(32'hbc81e76b),
	.w8(32'hba94f902),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbdccb),
	.w1(32'h3b15c45d),
	.w2(32'hba24f323),
	.w3(32'hbad02cba),
	.w4(32'h3926ecc0),
	.w5(32'hbb0e8793),
	.w6(32'hbaf12743),
	.w7(32'hb8bfe6bd),
	.w8(32'hbadf00c8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9440b7),
	.w1(32'hbb88f811),
	.w2(32'hbb12cc90),
	.w3(32'hbba90118),
	.w4(32'hbbcd82c3),
	.w5(32'h3a370a8b),
	.w6(32'hbbd22eab),
	.w7(32'hbbf7975c),
	.w8(32'hba80f58d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb992d71),
	.w1(32'hbabe169a),
	.w2(32'h3ab5f4f6),
	.w3(32'hbb9eb1b8),
	.w4(32'hbbde0f6a),
	.w5(32'h3b6df539),
	.w6(32'h39a6d7ec),
	.w7(32'h3a520295),
	.w8(32'h3bcf03f4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a571c2f),
	.w1(32'h3abf37da),
	.w2(32'h39fe82a7),
	.w3(32'h3b8efda3),
	.w4(32'h3b8b87b2),
	.w5(32'hbb03ddc4),
	.w6(32'h3be864fe),
	.w7(32'h3be3318a),
	.w8(32'h3b1b4c1c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7f780),
	.w1(32'h39cb8ebe),
	.w2(32'hbaa8e0e7),
	.w3(32'hba37d00d),
	.w4(32'h39b11fea),
	.w5(32'hba451255),
	.w6(32'hba1637d7),
	.w7(32'h3b380c35),
	.w8(32'h3b0ab468),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7900d),
	.w1(32'h3c00e113),
	.w2(32'hbc14a858),
	.w3(32'h3b33a15b),
	.w4(32'h3bb269f2),
	.w5(32'hbbbe5ed4),
	.w6(32'h3b665b4c),
	.w7(32'h3b284a54),
	.w8(32'h3b41b7bd),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e3b54),
	.w1(32'hbc32c196),
	.w2(32'h3b8634dc),
	.w3(32'hbbc56bd0),
	.w4(32'hbbd2abc0),
	.w5(32'h3be478e7),
	.w6(32'h3b3f97c3),
	.w7(32'h3aa6005a),
	.w8(32'hbb694545),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cd21f),
	.w1(32'h3ba62509),
	.w2(32'h3a845d60),
	.w3(32'h3a0dc5d2),
	.w4(32'h3b12ccfb),
	.w5(32'hba139f9c),
	.w6(32'hba9cb28b),
	.w7(32'h3a841f4f),
	.w8(32'h3a7231b9),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9404a9d),
	.w1(32'hba3abd4d),
	.w2(32'h3bd506a2),
	.w3(32'hbab334b2),
	.w4(32'hbac94ab9),
	.w5(32'h3b13483d),
	.w6(32'hba8f5484),
	.w7(32'hbab4fba6),
	.w8(32'h3ad2ae8c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0170c6),
	.w1(32'h3bb6ec9d),
	.w2(32'hbbc527b0),
	.w3(32'h3b33525a),
	.w4(32'h38ee408f),
	.w5(32'hbb4457f2),
	.w6(32'hbb3753ee),
	.w7(32'h3b211beb),
	.w8(32'h3baf73dd),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25c77c),
	.w1(32'hbc0a1ce8),
	.w2(32'hba32376c),
	.w3(32'hbbfb55a9),
	.w4(32'hbbdd7965),
	.w5(32'hbb38da46),
	.w6(32'h3a61b649),
	.w7(32'h3b1dca77),
	.w8(32'hbbbac4a5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcde99f),
	.w1(32'hbbd388ed),
	.w2(32'hb9cc4567),
	.w3(32'hbbcf81f6),
	.w4(32'hbb703a73),
	.w5(32'hbae23d9b),
	.w6(32'hbbad0b1c),
	.w7(32'hbbd33b66),
	.w8(32'h3b3d8c37),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb187a25),
	.w1(32'hbaae8651),
	.w2(32'h39252c26),
	.w3(32'hbaad69df),
	.w4(32'h3a8f5b14),
	.w5(32'h3a1c7efa),
	.w6(32'hbb56b2a9),
	.w7(32'h3b3bd7f9),
	.w8(32'hba77ccd0),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b322ec9),
	.w1(32'h39f0e28a),
	.w2(32'hbb0275e4),
	.w3(32'h3a831383),
	.w4(32'h3a85827f),
	.w5(32'hbb900cb2),
	.w6(32'h3ae51ab9),
	.w7(32'hb9912c8b),
	.w8(32'hb99bbff9),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4f41e),
	.w1(32'hbb36da0f),
	.w2(32'hbb1247d2),
	.w3(32'hbbb8780f),
	.w4(32'hbaf13dae),
	.w5(32'hbbd7f4aa),
	.w6(32'hbb2266cb),
	.w7(32'hba589e20),
	.w8(32'hb9c71a57),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadefe2f),
	.w1(32'h3a956063),
	.w2(32'h3bc51d27),
	.w3(32'h3a9bd946),
	.w4(32'hbb13b557),
	.w5(32'hb9a3a1c3),
	.w6(32'h3997aed9),
	.w7(32'h3a14a406),
	.w8(32'hbc00385b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e86ab),
	.w1(32'h3c4d2f52),
	.w2(32'h38a2f7cd),
	.w3(32'h3b313381),
	.w4(32'h3b423475),
	.w5(32'h3b09b451),
	.w6(32'hbbf1643e),
	.w7(32'hbbbb44c1),
	.w8(32'h3aa39cc7),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e9a3f),
	.w1(32'hbc069f44),
	.w2(32'hbbb1e5ae),
	.w3(32'hbbebe213),
	.w4(32'hbbf0adf2),
	.w5(32'hbbe1fc6d),
	.w6(32'h3b2efa3f),
	.w7(32'hbbefe32c),
	.w8(32'h3bea5db5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef4a25),
	.w1(32'h3b500cdb),
	.w2(32'h3a10f796),
	.w3(32'hbbb45f44),
	.w4(32'hbb4c37f5),
	.w5(32'h3aef33d6),
	.w6(32'hbb1771eb),
	.w7(32'hbba49962),
	.w8(32'h3a63d2db),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b211066),
	.w1(32'hbb5b566b),
	.w2(32'hbb82c7f3),
	.w3(32'h3b4fe962),
	.w4(32'h3ac10546),
	.w5(32'hbb0000e4),
	.w6(32'h3b4e3f95),
	.w7(32'h3b0f0620),
	.w8(32'hbbcc9167),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78d920),
	.w1(32'h3ae17109),
	.w2(32'h3b2ee4b0),
	.w3(32'h3a3d0dc0),
	.w4(32'h39e8ebb6),
	.w5(32'h3ae84560),
	.w6(32'hbb43bc83),
	.w7(32'hbb07aa9b),
	.w8(32'h3a940851),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad320f2),
	.w1(32'h3a9ab2d3),
	.w2(32'hbbe4b357),
	.w3(32'h36ff89ae),
	.w4(32'hb95afc5c),
	.w5(32'hbbdae326),
	.w6(32'hbaac3b45),
	.w7(32'h39cd29db),
	.w8(32'hba859e38),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a6846),
	.w1(32'h3bb11eb0),
	.w2(32'h3ae53fd7),
	.w3(32'hbba581a9),
	.w4(32'h3a5e3401),
	.w5(32'hbb577b0b),
	.w6(32'h3baeb5c5),
	.w7(32'hb892bc19),
	.w8(32'h3b004c45),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd405b),
	.w1(32'h3b159eca),
	.w2(32'h3b7e12ef),
	.w3(32'h3b3a6024),
	.w4(32'h3b3de7ba),
	.w5(32'h3b00d5e8),
	.w6(32'h3c000ba2),
	.w7(32'hba3eb9da),
	.w8(32'hbafcfff2),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd044f8),
	.w1(32'hbb98da30),
	.w2(32'hba84088e),
	.w3(32'h3ba1d23b),
	.w4(32'hbb9c02de),
	.w5(32'hbaeca4a3),
	.w6(32'hb9bd9a2a),
	.w7(32'hb9b3d049),
	.w8(32'hbb6f496d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79746f),
	.w1(32'hba147438),
	.w2(32'h3b6280b5),
	.w3(32'hbb530024),
	.w4(32'h35ce4953),
	.w5(32'h3aba6a36),
	.w6(32'hbb1e8f7c),
	.w7(32'hbb1291f3),
	.w8(32'h3a9f2867),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c031003),
	.w1(32'h3b8b8a00),
	.w2(32'hbbb39cc0),
	.w3(32'hbab211e1),
	.w4(32'hbb027971),
	.w5(32'hbae9145d),
	.w6(32'h3a2f275a),
	.w7(32'hba331501),
	.w8(32'h3b19289c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb886098),
	.w1(32'hbb0e3c57),
	.w2(32'h3bc2e3ee),
	.w3(32'hba7eb53e),
	.w4(32'hbbdf5d06),
	.w5(32'h3c009c58),
	.w6(32'hbb9d13e8),
	.w7(32'h3a5db882),
	.w8(32'h3b1543f5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be428d0),
	.w1(32'h3c23ef55),
	.w2(32'h39423c1d),
	.w3(32'h3c188895),
	.w4(32'h3ba72f28),
	.w5(32'h3b013a08),
	.w6(32'h3adf0b8e),
	.w7(32'hbaa6d183),
	.w8(32'h3bb5b766),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a007ef),
	.w1(32'h3bbecb61),
	.w2(32'h39d92466),
	.w3(32'hba533e36),
	.w4(32'hbb36e589),
	.w5(32'h3aa2c4af),
	.w6(32'hbb162358),
	.w7(32'hbb0ed3d8),
	.w8(32'h3abf9158),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8da00fc),
	.w1(32'hba87a07c),
	.w2(32'hbaba38f8),
	.w3(32'h3b09ecfb),
	.w4(32'h3a2c69c7),
	.w5(32'hbad1d6dd),
	.w6(32'h3b11c549),
	.w7(32'hba7d7015),
	.w8(32'hbb83b1bb),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ddbda),
	.w1(32'hbb721af8),
	.w2(32'hba9242a0),
	.w3(32'hbb4d0c38),
	.w4(32'hbb76424a),
	.w5(32'hba9f81e3),
	.w6(32'hbb295e0a),
	.w7(32'hbb9476ba),
	.w8(32'hbb07bd90),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94316c),
	.w1(32'h3bd33e25),
	.w2(32'h3aa6d7b1),
	.w3(32'hbb5222c2),
	.w4(32'h3a47911e),
	.w5(32'hbaebad10),
	.w6(32'hbb03d84b),
	.w7(32'h38d425ca),
	.w8(32'h399a5f30),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5ad12),
	.w1(32'hbb6ee6a9),
	.w2(32'h3b98076c),
	.w3(32'hbb515a3d),
	.w4(32'hbb698f5a),
	.w5(32'h3b1ec374),
	.w6(32'h3a8621b4),
	.w7(32'hba8c08af),
	.w8(32'hb99a4873),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34a331),
	.w1(32'h3b2b8841),
	.w2(32'hbb4f0532),
	.w3(32'h3b9c7c26),
	.w4(32'hbb069539),
	.w5(32'hbb231c82),
	.w6(32'h3b7d02ce),
	.w7(32'h3974a27d),
	.w8(32'hbae831ed),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60cf05),
	.w1(32'hbb0e5bef),
	.w2(32'hba920a9d),
	.w3(32'hbb9ab68a),
	.w4(32'hbb43af76),
	.w5(32'hbba02e73),
	.w6(32'hbb868bbc),
	.w7(32'hbb14380c),
	.w8(32'h39ffebce),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82368df),
	.w1(32'h3aa292d7),
	.w2(32'h3b885f92),
	.w3(32'hbb4eb58b),
	.w4(32'hbac89a8a),
	.w5(32'hbc0659b6),
	.w6(32'h3ac02dc6),
	.w7(32'h3b0c9389),
	.w8(32'hbb2adc47),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fbdcdc),
	.w1(32'h39bae518),
	.w2(32'h3a7c5371),
	.w3(32'hbbab5644),
	.w4(32'hbbaf8b70),
	.w5(32'h38c0fe6a),
	.w6(32'hbac32e3b),
	.w7(32'hba656bb2),
	.w8(32'h3a83403f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a904d34),
	.w1(32'h3a2a58bb),
	.w2(32'h3c26334c),
	.w3(32'hb8783864),
	.w4(32'hba9c2b08),
	.w5(32'h3ba654a2),
	.w6(32'h3ae91ed4),
	.w7(32'h38d32179),
	.w8(32'hba7fbd90),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52e307),
	.w1(32'h3c7a5908),
	.w2(32'hbb9cc63f),
	.w3(32'h3bda781e),
	.w4(32'h3bd1ede4),
	.w5(32'hbb1fae99),
	.w6(32'hbae39ec8),
	.w7(32'hbaa12351),
	.w8(32'hba8ee69b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39188e83),
	.w1(32'h3b0c1713),
	.w2(32'hbacd96b4),
	.w3(32'h39c95bd8),
	.w4(32'hba94dd5f),
	.w5(32'hbb3984e6),
	.w6(32'h3af73a4f),
	.w7(32'hba9697ce),
	.w8(32'hbb9354e6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae63fff),
	.w1(32'h3a593f4e),
	.w2(32'h3b712a4f),
	.w3(32'hbb952893),
	.w4(32'hbb70a20b),
	.w5(32'h3b9c4aa4),
	.w6(32'hbb0caee8),
	.w7(32'hbb4e2f8b),
	.w8(32'h3ba81f4f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b784c78),
	.w1(32'h3b88a36f),
	.w2(32'h3be37105),
	.w3(32'h3b986777),
	.w4(32'h3bb79002),
	.w5(32'h3c005d34),
	.w6(32'h3b9e19e3),
	.w7(32'h3b970469),
	.w8(32'h3b980ac8),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c074e63),
	.w1(32'h3b87ef81),
	.w2(32'h39d7e1e1),
	.w3(32'h3bbf1afd),
	.w4(32'h3ab6e3ab),
	.w5(32'h3aca2bc6),
	.w6(32'hb9344565),
	.w7(32'hbac8ef3d),
	.w8(32'h3a807d41),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16f6cb),
	.w1(32'hba6938e5),
	.w2(32'hbba59b41),
	.w3(32'h3b3625f4),
	.w4(32'hbb84495d),
	.w5(32'hbb2496dd),
	.w6(32'h3a6135c5),
	.w7(32'hbb74ab88),
	.w8(32'hbb236552),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa54be3),
	.w1(32'h392db858),
	.w2(32'h3a9ffcf8),
	.w3(32'hb897142c),
	.w4(32'hba20d639),
	.w5(32'h3ab4386c),
	.w6(32'h3b25ef2a),
	.w7(32'hbb0a8b62),
	.w8(32'h3a63aa93),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1870a1),
	.w1(32'h3964a579),
	.w2(32'h3ad3222b),
	.w3(32'hbaea6828),
	.w4(32'hba4b6dd0),
	.w5(32'h3a92400e),
	.w6(32'hbb0b9c87),
	.w7(32'hbb7d4c61),
	.w8(32'hbacf4e45),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac78cf0),
	.w1(32'h3a63f253),
	.w2(32'hbb346131),
	.w3(32'h3a713afc),
	.w4(32'hba1cb26c),
	.w5(32'hbbcb98e8),
	.w6(32'hbb0de61a),
	.w7(32'hbb1e9c51),
	.w8(32'hbba5d0e4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34c7c7),
	.w1(32'hbb965d73),
	.w2(32'h3acc09e7),
	.w3(32'hbb81da0e),
	.w4(32'hbbcf5b4c),
	.w5(32'h3a9eb0e2),
	.w6(32'hbb6f33f4),
	.w7(32'hbbccc63b),
	.w8(32'hbb5544fd),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7356ff),
	.w1(32'hbbe3e37e),
	.w2(32'h3b1dc6a8),
	.w3(32'hbb3bc63f),
	.w4(32'hbbc0878c),
	.w5(32'h3a8e0548),
	.w6(32'hbb7022b2),
	.w7(32'hbbf636f9),
	.w8(32'hbacbfe6f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6016ea),
	.w1(32'h399e78f2),
	.w2(32'hbbf791f4),
	.w3(32'hbbca2266),
	.w4(32'hbaa36beb),
	.w5(32'hbbccdb57),
	.w6(32'hba3943da),
	.w7(32'hbac1981d),
	.w8(32'hbb2a5ae4),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f73ae),
	.w1(32'hbb16d2e6),
	.w2(32'h3aa9a927),
	.w3(32'hbb8f5e29),
	.w4(32'hbae7531c),
	.w5(32'h3aa949e0),
	.w6(32'hbb3fa1d7),
	.w7(32'hbab05379),
	.w8(32'hba8d8c38),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b592357),
	.w1(32'h3b4621e9),
	.w2(32'hba7a4512),
	.w3(32'h3b2eb81b),
	.w4(32'h3aeb942c),
	.w5(32'h3b37ff78),
	.w6(32'h3b06694e),
	.w7(32'hb91ed6c2),
	.w8(32'h399824d8),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70d654),
	.w1(32'h3babac77),
	.w2(32'h3b72dcfb),
	.w3(32'h3bb7f043),
	.w4(32'h3b99007d),
	.w5(32'h3a8d09fc),
	.w6(32'h3b16f0d9),
	.w7(32'h39b98a96),
	.w8(32'hbb199ac7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba13e9),
	.w1(32'h3c221e79),
	.w2(32'hbb95a39e),
	.w3(32'h3b2f63e8),
	.w4(32'h3bb54129),
	.w5(32'hbbe37881),
	.w6(32'hbaf0b828),
	.w7(32'h37812d60),
	.w8(32'hbbb0a843),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b3fc4),
	.w1(32'hbaff7a6c),
	.w2(32'hbb93f8a3),
	.w3(32'hb994b744),
	.w4(32'h3aab02f2),
	.w5(32'hbacab0f4),
	.w6(32'h3ab0db4e),
	.w7(32'h3b614683),
	.w8(32'hbaf78728),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b2e542),
	.w1(32'h3b41cbcb),
	.w2(32'h3ae0e3d6),
	.w3(32'h3b73030f),
	.w4(32'h3b57114b),
	.w5(32'h3ac41d2a),
	.w6(32'h3b4c76aa),
	.w7(32'h3b1a41e5),
	.w8(32'h3b85423c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad44e1),
	.w1(32'hbb193adf),
	.w2(32'hbbb3cf69),
	.w3(32'h3b7f7fed),
	.w4(32'hbb19eea9),
	.w5(32'hbb9150cf),
	.w6(32'hb9075c1d),
	.w7(32'h3b344fba),
	.w8(32'h38852997),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadd2d8),
	.w1(32'hbbd03f1f),
	.w2(32'hbb226a58),
	.w3(32'hbacb3ba9),
	.w4(32'hbbeedc97),
	.w5(32'hba3c70fc),
	.w6(32'hbb630e23),
	.w7(32'hbc02cf66),
	.w8(32'hbac78591),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21bb6f),
	.w1(32'hbae58a97),
	.w2(32'h3c05490c),
	.w3(32'hb998a26d),
	.w4(32'hba3e4854),
	.w5(32'h3bfeeb69),
	.w6(32'hbacda953),
	.w7(32'hbb0a6788),
	.w8(32'h3bb4cf66),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c8179),
	.w1(32'h3c217b85),
	.w2(32'h3b052a58),
	.w3(32'h3c2b5cdd),
	.w4(32'h3c166ee1),
	.w5(32'hbb7974e2),
	.w6(32'h3c146951),
	.w7(32'h3baaf5b4),
	.w8(32'h3b16202c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baec839),
	.w1(32'h3be3138f),
	.w2(32'h39c006fe),
	.w3(32'h3b335f4c),
	.w4(32'h3b18af1d),
	.w5(32'h3b3d2d55),
	.w6(32'h3beaff1f),
	.w7(32'h3a89519b),
	.w8(32'h3b1d33da),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9c3c8),
	.w1(32'h3bc873f6),
	.w2(32'h3c12910d),
	.w3(32'h3b60e64b),
	.w4(32'hbb016cc2),
	.w5(32'h3bdca36d),
	.w6(32'h3b04f127),
	.w7(32'hbb21dbe8),
	.w8(32'h3bffdc48),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c136807),
	.w1(32'h3b256cd9),
	.w2(32'h3bb554c7),
	.w3(32'h3abe3e2a),
	.w4(32'hbb2bf5ba),
	.w5(32'h3bedd1f4),
	.w6(32'h3b3e3f9d),
	.w7(32'h3b300632),
	.w8(32'h3c0cef63),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55585e),
	.w1(32'hbb0c0d1b),
	.w2(32'hbab65534),
	.w3(32'hbacf9850),
	.w4(32'h3aafb061),
	.w5(32'hba4cbb04),
	.w6(32'h3b173174),
	.w7(32'h3bedc3b0),
	.w8(32'hba04c494),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba640071),
	.w1(32'hbb44dcb4),
	.w2(32'h3c3d10b4),
	.w3(32'h39e24951),
	.w4(32'hbaf9812d),
	.w5(32'h3bec6205),
	.w6(32'h3ab9f398),
	.w7(32'hbb394084),
	.w8(32'hba87410d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bab77),
	.w1(32'h3c62d37d),
	.w2(32'hba0442c5),
	.w3(32'h3c1b7094),
	.w4(32'h3c27ddb6),
	.w5(32'hba91573e),
	.w6(32'h3a49cefb),
	.w7(32'h3a0b80ae),
	.w8(32'hbb8b85cf),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8b2c6),
	.w1(32'hbb4cafcb),
	.w2(32'h3a9d5647),
	.w3(32'hbafb1e32),
	.w4(32'hbb621d74),
	.w5(32'h3b10c38e),
	.w6(32'hbb62be18),
	.w7(32'hbb77bcba),
	.w8(32'hb95f41e2),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b06116),
	.w1(32'h3b161780),
	.w2(32'hbadbe036),
	.w3(32'h39a9de17),
	.w4(32'h3a4995f7),
	.w5(32'hbae03af8),
	.w6(32'h3c053133),
	.w7(32'h3b70eb94),
	.w8(32'hb84c85e5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1be52d),
	.w1(32'h3b30ea81),
	.w2(32'h3bda8f31),
	.w3(32'hb98b7f82),
	.w4(32'hbb8787b7),
	.w5(32'hba1b9567),
	.w6(32'hbb28cd70),
	.w7(32'hbac6a472),
	.w8(32'h3b86d3d5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b484a05),
	.w1(32'h3aa47dee),
	.w2(32'h3b81be17),
	.w3(32'h3bbb4f73),
	.w4(32'h390f388f),
	.w5(32'hba2fde80),
	.w6(32'h3ae3f793),
	.w7(32'h3b9d0791),
	.w8(32'hb9168b12),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c057f22),
	.w1(32'h3afdbfd8),
	.w2(32'h3a407178),
	.w3(32'h3b886b0c),
	.w4(32'hb8b1c934),
	.w5(32'h3b4e58c2),
	.w6(32'hba14bf22),
	.w7(32'h3bb280fd),
	.w8(32'hba511a1d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8008e8),
	.w1(32'h3bc6ffed),
	.w2(32'hbba2973b),
	.w3(32'hba2e3fa2),
	.w4(32'h3ab59f90),
	.w5(32'hbbbe953b),
	.w6(32'hbb842347),
	.w7(32'h3a17a955),
	.w8(32'hbb713d47),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fb6b9),
	.w1(32'hbb62bf65),
	.w2(32'hbbaf3100),
	.w3(32'hbbcc2349),
	.w4(32'hbb89bc79),
	.w5(32'hbb2ee3d5),
	.w6(32'hbb7d0d39),
	.w7(32'hbb611bb3),
	.w8(32'hbbdef759),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f5bf4),
	.w1(32'hba09c555),
	.w2(32'hbad6e3f8),
	.w3(32'hbb2200df),
	.w4(32'hb964401e),
	.w5(32'hba623523),
	.w6(32'hbb99413e),
	.w7(32'h3a2d51ab),
	.w8(32'hbaddea55),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95766e),
	.w1(32'h3b96007f),
	.w2(32'hbaa9ad1e),
	.w3(32'hb9283134),
	.w4(32'h3ac13d45),
	.w5(32'h3b4da96c),
	.w6(32'hbaab47bd),
	.w7(32'hb8afefd1),
	.w8(32'h3b51272e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb621b),
	.w1(32'h3bbcce3a),
	.w2(32'h398314ee),
	.w3(32'h3b8c94b8),
	.w4(32'h3b661312),
	.w5(32'hbaca35f6),
	.w6(32'h3b8f65a3),
	.w7(32'h3aa2cb63),
	.w8(32'hba95cb92),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fde0a),
	.w1(32'h39f3fe83),
	.w2(32'h3b1aa5da),
	.w3(32'h390fbba6),
	.w4(32'hbb2e7307),
	.w5(32'h3af1251c),
	.w6(32'hba9c3d32),
	.w7(32'hbb2217fe),
	.w8(32'hba10ca69),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6f78e),
	.w1(32'h3a18f04e),
	.w2(32'hba179a65),
	.w3(32'h3b2e41e3),
	.w4(32'h36d654a4),
	.w5(32'h3a84b82c),
	.w6(32'hba3a1acf),
	.w7(32'hbbccff7a),
	.w8(32'hba8dcb71),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cf02b),
	.w1(32'hb8985ef6),
	.w2(32'hbb9e56a7),
	.w3(32'h3abe0eeb),
	.w4(32'hba32fad8),
	.w5(32'hbb8c408d),
	.w6(32'hbb278491),
	.w7(32'hbbb33c98),
	.w8(32'hbbe58584),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ff181),
	.w1(32'h3b83cb73),
	.w2(32'h3aabd424),
	.w3(32'hbb6bb563),
	.w4(32'hb95adbda),
	.w5(32'h3b7c7a5b),
	.w6(32'hbb679cca),
	.w7(32'hba68885b),
	.w8(32'h3ab4ed1b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1506dd),
	.w1(32'h3b44d0ec),
	.w2(32'hbbb40e8e),
	.w3(32'h3b201b6f),
	.w4(32'h3ad1dbb1),
	.w5(32'hbb762c0d),
	.w6(32'h3b4badd6),
	.w7(32'h3ab54597),
	.w8(32'hbb8b9576),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3293a4),
	.w1(32'hba5872f5),
	.w2(32'hbb612641),
	.w3(32'hbaa82b32),
	.w4(32'hba0ae838),
	.w5(32'h3a0804f2),
	.w6(32'hbb45bc97),
	.w7(32'hb9d6849c),
	.w8(32'hbb21502c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab94835),
	.w1(32'hba8f6444),
	.w2(32'h3a02e8d7),
	.w3(32'hbbb488b9),
	.w4(32'hbbd80fd3),
	.w5(32'h3a9048e4),
	.w6(32'hbb8ca521),
	.w7(32'hbad68456),
	.w8(32'h3b8d6a1f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bf2af),
	.w1(32'h3b30681a),
	.w2(32'hbb3fe49f),
	.w3(32'hbb391c69),
	.w4(32'hbbdded25),
	.w5(32'hbabef6b2),
	.w6(32'hbb2ae2d4),
	.w7(32'hbb3b61bc),
	.w8(32'hba3fa5bd),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ff68c),
	.w1(32'h3c7d778b),
	.w2(32'hba973035),
	.w3(32'h3bced29c),
	.w4(32'h3c3e52dc),
	.w5(32'h3ad991bf),
	.w6(32'h3bc50600),
	.w7(32'h3c28f023),
	.w8(32'hb83cb807),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980772a),
	.w1(32'h3b50e20b),
	.w2(32'h3a80ee24),
	.w3(32'h3b7c5daa),
	.w4(32'hb9a2279c),
	.w5(32'h3bbbb87e),
	.w6(32'h39e92ceb),
	.w7(32'h3b53fc4c),
	.w8(32'h3b0cce97),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b485c),
	.w1(32'h3b017037),
	.w2(32'hbbcb0816),
	.w3(32'hba3833ac),
	.w4(32'h3bbda088),
	.w5(32'hbb8eae6d),
	.w6(32'h3af777ea),
	.w7(32'h3b8721a9),
	.w8(32'hbb8cbb7b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb940b7b),
	.w1(32'hb9b461f0),
	.w2(32'h3c2b2299),
	.w3(32'hbb9d6915),
	.w4(32'hbadb2dc4),
	.w5(32'h3b3db921),
	.w6(32'hbb935e89),
	.w7(32'hbb1ec9df),
	.w8(32'h3ac3b122),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc235e),
	.w1(32'h3ad3700d),
	.w2(32'hbbf36a28),
	.w3(32'h3aacae55),
	.w4(32'hba898cd2),
	.w5(32'hbbb60e2c),
	.w6(32'h3ae441ee),
	.w7(32'hba12fc21),
	.w8(32'hbb8d5d13),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56944c),
	.w1(32'h3a54ed38),
	.w2(32'h393f55e3),
	.w3(32'hbb90b475),
	.w4(32'hbb21da2a),
	.w5(32'h3b7ca4de),
	.w6(32'hbb0ea327),
	.w7(32'hbadcf3c8),
	.w8(32'hbb808d87),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f183f),
	.w1(32'h3a6ed95a),
	.w2(32'hbb8a5a3d),
	.w3(32'h3b0001e4),
	.w4(32'h3aa3ff93),
	.w5(32'hbb43729b),
	.w6(32'hbb431155),
	.w7(32'h38b520df),
	.w8(32'hba2c8854),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb960a976),
	.w1(32'hbb009f2d),
	.w2(32'hbb21cbe0),
	.w3(32'hbb13805c),
	.w4(32'hbb618274),
	.w5(32'hbad775a1),
	.w6(32'hbb1345ab),
	.w7(32'hbb2d2b5e),
	.w8(32'h3acfa123),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab82890),
	.w1(32'hbb41f0ee),
	.w2(32'hbaaf3b20),
	.w3(32'hb8c6025c),
	.w4(32'hba92e948),
	.w5(32'h39c59d9c),
	.w6(32'hba6f8ec9),
	.w7(32'hb9307f06),
	.w8(32'h3b356a23),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e642d),
	.w1(32'hbb7208de),
	.w2(32'h399f1832),
	.w3(32'hb8d9a0cd),
	.w4(32'hba562e78),
	.w5(32'h3a85dce4),
	.w6(32'h3b3bca95),
	.w7(32'h3afa3ffc),
	.w8(32'h3b14aa5b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c03ff),
	.w1(32'hba7cf6c3),
	.w2(32'hbb3b4aa3),
	.w3(32'h3aed3996),
	.w4(32'h3a8fdacf),
	.w5(32'hbba699a9),
	.w6(32'h3b7d380c),
	.w7(32'h3ad3646b),
	.w8(32'hbbbc0277),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a5c78),
	.w1(32'h3b3288a3),
	.w2(32'hbaf2e2ec),
	.w3(32'hbb83a9dd),
	.w4(32'h3bc9e313),
	.w5(32'hb94c12af),
	.w6(32'h3b02adb5),
	.w7(32'h3ab30760),
	.w8(32'hb9cd92e2),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad1649),
	.w1(32'hb9371453),
	.w2(32'h3b8b6450),
	.w3(32'hb8c02fd9),
	.w4(32'hba319a52),
	.w5(32'h3a877629),
	.w6(32'hbacf68e3),
	.w7(32'hbb3b934b),
	.w8(32'hbb3c0179),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03ec9b),
	.w1(32'h3c02995d),
	.w2(32'h3a0b92e9),
	.w3(32'h3b2f7aee),
	.w4(32'h3bb7d853),
	.w5(32'hba0f9eb7),
	.w6(32'h3c1265fa),
	.w7(32'h3b427c84),
	.w8(32'h3b0393a2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb173ada),
	.w1(32'hbaf83d46),
	.w2(32'hba577cd2),
	.w3(32'h3bd9e43f),
	.w4(32'hbaaecead),
	.w5(32'hbbb8fcea),
	.w6(32'h3c4dad6f),
	.w7(32'hbb666a16),
	.w8(32'hbb812948),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa776b7),
	.w1(32'hbb7b4962),
	.w2(32'hbb1d8918),
	.w3(32'hbb523755),
	.w4(32'hbb990118),
	.w5(32'hba59c34d),
	.w6(32'h3ba1625f),
	.w7(32'hbb835f4d),
	.w8(32'hbaf803ea),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule