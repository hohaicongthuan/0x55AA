module layer_10_featuremap_13(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b153751),
	.w1(32'h3a5cfe67),
	.w2(32'hbb55df68),
	.w3(32'hbbb0b9bb),
	.w4(32'hbc1adae0),
	.w5(32'hba1ad4a5),
	.w6(32'hbc359c59),
	.w7(32'hbb5a6f75),
	.w8(32'hbc184efc),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97c4a7),
	.w1(32'h3af1a5d5),
	.w2(32'hbc279478),
	.w3(32'h3c8c3cb1),
	.w4(32'h3cfc95e1),
	.w5(32'h3c56f72a),
	.w6(32'hbc5afde4),
	.w7(32'hbbf4ec29),
	.w8(32'hba827cc1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e455b),
	.w1(32'hbba5ae61),
	.w2(32'h3b667e56),
	.w3(32'h3c33956a),
	.w4(32'h3c8b3fe2),
	.w5(32'hbb3a2d1e),
	.w6(32'hbb7f56bb),
	.w7(32'hbb5f8cc2),
	.w8(32'hbc3711b2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8848d6),
	.w1(32'h3b80dbaf),
	.w2(32'hbc6aacdb),
	.w3(32'hbc456dbc),
	.w4(32'hbc1de98f),
	.w5(32'h3af66bc5),
	.w6(32'hbbc060e6),
	.w7(32'hbb0bc6fc),
	.w8(32'hbca3a670),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd34495),
	.w1(32'h3b9833d6),
	.w2(32'h3c2bab83),
	.w3(32'hbbf25d03),
	.w4(32'hbcbe9577),
	.w5(32'hbb10e5dc),
	.w6(32'hbccb8d55),
	.w7(32'hbc778ef0),
	.w8(32'hbb102c36),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c37f9),
	.w1(32'hbad7d066),
	.w2(32'hbb9c07d6),
	.w3(32'hbbc7e5f7),
	.w4(32'hbb181220),
	.w5(32'hbb9b815d),
	.w6(32'h3b55a8c7),
	.w7(32'h3c334b85),
	.w8(32'hb9be0120),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb229a0e),
	.w1(32'h3a15c7d1),
	.w2(32'hbc0b8677),
	.w3(32'hbb857572),
	.w4(32'h3b11b90d),
	.w5(32'h3c103a3a),
	.w6(32'hbab5c371),
	.w7(32'h3b04a7d1),
	.w8(32'h3b385449),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ce267),
	.w1(32'hbbf955b6),
	.w2(32'h3b18c317),
	.w3(32'h3c881f54),
	.w4(32'h3c6805ec),
	.w5(32'hbbd14e29),
	.w6(32'hbbdb62ed),
	.w7(32'hbc089861),
	.w8(32'h3bf5e0f5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b47c9),
	.w1(32'h3b3ae122),
	.w2(32'hbbb896dc),
	.w3(32'hbafb71e2),
	.w4(32'hbbd05d54),
	.w5(32'hbb5b21d3),
	.w6(32'h3bbc1df3),
	.w7(32'hbaacb3da),
	.w8(32'h39431075),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8621e4),
	.w1(32'hbc8c0f8a),
	.w2(32'h39a53e88),
	.w3(32'hbbf7472d),
	.w4(32'hbbe6bfee),
	.w5(32'hbac562bd),
	.w6(32'hbb789040),
	.w7(32'hbbebc5bd),
	.w8(32'hbb665876),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb391f94),
	.w1(32'hba4bb2d2),
	.w2(32'h3bb32c6c),
	.w3(32'hbb53c79b),
	.w4(32'hba10ca61),
	.w5(32'hbbd793c0),
	.w6(32'hbb899607),
	.w7(32'hbb1bf630),
	.w8(32'hbc209bcf),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f43b1),
	.w1(32'h3a0c6242),
	.w2(32'h3b0360a3),
	.w3(32'hbc00e197),
	.w4(32'hbc6a4caf),
	.w5(32'h3c10a70d),
	.w6(32'hbc32d2e1),
	.w7(32'h3b4c1e21),
	.w8(32'h3bf7be0e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea90ef),
	.w1(32'hbabd60ba),
	.w2(32'hbaa1a97d),
	.w3(32'hba61ca13),
	.w4(32'h3aee2241),
	.w5(32'hbb06834a),
	.w6(32'hba685095),
	.w7(32'h3ab9edb5),
	.w8(32'hbbab4a8e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c2e1c),
	.w1(32'hbc0794e1),
	.w2(32'hbc3530e9),
	.w3(32'h3b187493),
	.w4(32'hbaaa848f),
	.w5(32'h3bec72fa),
	.w6(32'h3c25025b),
	.w7(32'h3b8c52cc),
	.w8(32'hbc8934a8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfb461),
	.w1(32'h3c2caad9),
	.w2(32'hbc0486c8),
	.w3(32'h3ba3694f),
	.w4(32'hbb1fea76),
	.w5(32'hbb3d1e37),
	.w6(32'hbc19fce3),
	.w7(32'hbc9c1e59),
	.w8(32'h3adf92e4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae893d4),
	.w1(32'h38155bbb),
	.w2(32'h3aa0159a),
	.w3(32'h3bbbe9c1),
	.w4(32'h3bdc6b67),
	.w5(32'hbb8e62a0),
	.w6(32'h3941e66b),
	.w7(32'hbab9c6a8),
	.w8(32'hbb8fa229),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f124e),
	.w1(32'h3a33f455),
	.w2(32'hb9dbd208),
	.w3(32'hbaa34fbb),
	.w4(32'h3aa553a8),
	.w5(32'hbb44f6c3),
	.w6(32'hbad61b05),
	.w7(32'h3a1dd1a7),
	.w8(32'hbb8d169c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc2d75),
	.w1(32'hbbd80de2),
	.w2(32'h3ba171ff),
	.w3(32'hbb5ec797),
	.w4(32'h3b1a6492),
	.w5(32'h3ad5fbe5),
	.w6(32'hbc1d7835),
	.w7(32'h39c596f8),
	.w8(32'hba17c2f0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba83c40),
	.w1(32'hbb89fdc4),
	.w2(32'h3a97d85e),
	.w3(32'h3b8bbb73),
	.w4(32'hba3a0b4f),
	.w5(32'hbc797c65),
	.w6(32'hbaa3782f),
	.w7(32'h3a257f1f),
	.w8(32'hbadd7b1e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90a61b),
	.w1(32'h35cfbe9f),
	.w2(32'h3b0b6ef8),
	.w3(32'hbc4a7460),
	.w4(32'hbc2cbc8f),
	.w5(32'hbb8933a6),
	.w6(32'hbc05f18b),
	.w7(32'hbc2670ba),
	.w8(32'h3b2d2140),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24d99c),
	.w1(32'h3b2602a4),
	.w2(32'h3c1058f1),
	.w3(32'hbbdbc382),
	.w4(32'hb9f6693b),
	.w5(32'hbc10d598),
	.w6(32'h3a531e64),
	.w7(32'h3c187b99),
	.w8(32'h3bf81ccc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b6c74),
	.w1(32'h3bc7236d),
	.w2(32'h3ba83f21),
	.w3(32'hbc2c8916),
	.w4(32'hbc87acf1),
	.w5(32'hbb3bebda),
	.w6(32'h3bbf84fd),
	.w7(32'h3b89dc2c),
	.w8(32'h3b241fae),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d6def),
	.w1(32'h3af4e7f2),
	.w2(32'h3c6c4575),
	.w3(32'h3ad57c9f),
	.w4(32'hbbcc7135),
	.w5(32'h3c11ad25),
	.w6(32'hba2cb7d6),
	.w7(32'h3a29a68e),
	.w8(32'h3b214d26),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ab8e6),
	.w1(32'hbab70f47),
	.w2(32'hbb9c725b),
	.w3(32'h3a53e71c),
	.w4(32'hba940c1d),
	.w5(32'hbb895a55),
	.w6(32'hbb6b9b15),
	.w7(32'hbb68bb39),
	.w8(32'hbc05e7cc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b061429),
	.w1(32'hbc1a27ff),
	.w2(32'h39b2756f),
	.w3(32'h3a7de01b),
	.w4(32'hbbe19e79),
	.w5(32'hbc2524a0),
	.w6(32'h3bf4d46b),
	.w7(32'h38b9b1fa),
	.w8(32'hbc7cd057),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4937e),
	.w1(32'h3b24bb2e),
	.w2(32'hba0ce76b),
	.w3(32'h3b2b0874),
	.w4(32'h39540182),
	.w5(32'hbc36bbde),
	.w6(32'hbc4a22cc),
	.w7(32'hbc55498f),
	.w8(32'h3c09625e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2fd03),
	.w1(32'h3b6e7401),
	.w2(32'hbafec905),
	.w3(32'hbb2d0d62),
	.w4(32'hbbb240aa),
	.w5(32'hbb331134),
	.w6(32'hbc4bdbe7),
	.w7(32'hbc19bfe0),
	.w8(32'hba8c7dd2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb154609),
	.w1(32'h38d93a8a),
	.w2(32'h3c230968),
	.w3(32'h3b089720),
	.w4(32'h3ad99f2f),
	.w5(32'h3b65d8bc),
	.w6(32'h3b2ebfef),
	.w7(32'h3beae3dc),
	.w8(32'h3b9f1944),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ceb81),
	.w1(32'h3bc83090),
	.w2(32'hbb0f326f),
	.w3(32'h390994da),
	.w4(32'h3c0bce83),
	.w5(32'hbbbf468a),
	.w6(32'h3b8280c0),
	.w7(32'h3bb58f8a),
	.w8(32'h3b889318),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb698ab8),
	.w1(32'h398cbb69),
	.w2(32'hbb8bab02),
	.w3(32'hbc227fdc),
	.w4(32'hbc81300b),
	.w5(32'hbb51e9cb),
	.w6(32'hbb5fafba),
	.w7(32'hbc63a86e),
	.w8(32'h393c50e8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ffc59),
	.w1(32'hbb358206),
	.w2(32'h3ad4d0e3),
	.w3(32'hbb755fd0),
	.w4(32'h3a21a959),
	.w5(32'hbb97327f),
	.w6(32'h3a435498),
	.w7(32'h3a5b8cff),
	.w8(32'h3b507984),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b460d2e),
	.w1(32'hb7e6dfbb),
	.w2(32'hbac727f0),
	.w3(32'hbb8a9fa4),
	.w4(32'hbb38e70b),
	.w5(32'hbbf9e84c),
	.w6(32'hba11a02c),
	.w7(32'hb9240dd1),
	.w8(32'h3a52c756),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1b816),
	.w1(32'hb89daca9),
	.w2(32'h3a49870a),
	.w3(32'hbc3df841),
	.w4(32'hbc07e43c),
	.w5(32'h3b13c97b),
	.w6(32'hbb81b4aa),
	.w7(32'hbc0e8500),
	.w8(32'hba84e859),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b9b24),
	.w1(32'hbb449b0b),
	.w2(32'h3a9732f8),
	.w3(32'hbb91c991),
	.w4(32'hbab4c8a1),
	.w5(32'hbb311aaa),
	.w6(32'hbb66b118),
	.w7(32'hbb15964f),
	.w8(32'hbb8402e5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6dfad),
	.w1(32'h3b72909f),
	.w2(32'hba8088e0),
	.w3(32'h3947a62b),
	.w4(32'h3c1115a0),
	.w5(32'hbb6ecdd6),
	.w6(32'hbb3bd410),
	.w7(32'h3b5e76bb),
	.w8(32'hbbbc3233),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3fa0a),
	.w1(32'hbacd105d),
	.w2(32'h3c2f9d34),
	.w3(32'hbc113302),
	.w4(32'hbc19e81f),
	.w5(32'hbc2bc629),
	.w6(32'hbc6784bd),
	.w7(32'hbc4c7fa1),
	.w8(32'hbcdd5199),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be913f8),
	.w1(32'hbb97ba7d),
	.w2(32'h3c7382de),
	.w3(32'hbc6a783b),
	.w4(32'hbca7122e),
	.w5(32'h3c647e5a),
	.w6(32'hbd1cdf09),
	.w7(32'hbcacfd8d),
	.w8(32'h3c6c9f7d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74a373),
	.w1(32'hbb2df450),
	.w2(32'hbb9e773a),
	.w3(32'hb9dc8ae3),
	.w4(32'h392274c9),
	.w5(32'h3b3f8024),
	.w6(32'h3be984d1),
	.w7(32'h3b80aed0),
	.w8(32'h3c702f85),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f27c8),
	.w1(32'hbbd7df27),
	.w2(32'h3c43530a),
	.w3(32'hbc3ea320),
	.w4(32'hbba856fe),
	.w5(32'h3c35d370),
	.w6(32'h3c2c1b01),
	.w7(32'h3c471174),
	.w8(32'h3c30a7e2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2f454),
	.w1(32'hbc43682b),
	.w2(32'hbaa8e40b),
	.w3(32'h3a6f5acd),
	.w4(32'hbc4304a2),
	.w5(32'hb9d25100),
	.w6(32'h3bddc64e),
	.w7(32'hbaaa360a),
	.w8(32'h3b6330d4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea940e),
	.w1(32'hbc0cb02d),
	.w2(32'hbc1481a8),
	.w3(32'hbbbb006f),
	.w4(32'hbbd5875b),
	.w5(32'hbbd88362),
	.w6(32'hbb821b9f),
	.w7(32'hbb92755f),
	.w8(32'h3b895a9b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef6b81),
	.w1(32'hb9d7b9f8),
	.w2(32'h3bd9db8b),
	.w3(32'hbc725ed4),
	.w4(32'hbc41c5d5),
	.w5(32'h3ace20ea),
	.w6(32'hbbdcd4e4),
	.w7(32'hbc18b4be),
	.w8(32'h3b541040),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba898bfb),
	.w1(32'hbb88f27d),
	.w2(32'h3b393c01),
	.w3(32'hb9e2cb0d),
	.w4(32'hbc2bee10),
	.w5(32'h3abb0dba),
	.w6(32'hbbcad566),
	.w7(32'hbc395533),
	.w8(32'hbab93d4e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe343f),
	.w1(32'h3bcf5104),
	.w2(32'h3b5bfa73),
	.w3(32'h3b39dd44),
	.w4(32'h3b6b5a20),
	.w5(32'h3bbf2acd),
	.w6(32'hbb9be322),
	.w7(32'hbadb32de),
	.w8(32'h3af92b21),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba907221),
	.w1(32'h3b235ad0),
	.w2(32'h3bcea738),
	.w3(32'hbabf166d),
	.w4(32'hbc1e9135),
	.w5(32'hba02e6d7),
	.w6(32'hbb7b01d4),
	.w7(32'hbc6d160e),
	.w8(32'h3c10526d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c046d63),
	.w1(32'h3c8a6cc9),
	.w2(32'h3bb39e19),
	.w3(32'h3c4ca0d3),
	.w4(32'h3c87ff3a),
	.w5(32'h3a82c423),
	.w6(32'h3c6c2ed1),
	.w7(32'h396af03b),
	.w8(32'hbaf753e7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba608c0),
	.w1(32'h3c070446),
	.w2(32'hbaa3d3c9),
	.w3(32'h3c01b968),
	.w4(32'h3b19076f),
	.w5(32'hbb9a7248),
	.w6(32'hbb507435),
	.w7(32'hbc3c36cd),
	.w8(32'hbc2199b2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbf794),
	.w1(32'h3c31abbc),
	.w2(32'h3c11cb0d),
	.w3(32'hbc4fadbc),
	.w4(32'h3ba1d0d0),
	.w5(32'h3bf0b754),
	.w6(32'hbcb5e48a),
	.w7(32'hbc8562c0),
	.w8(32'h3bbf3988),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b400149),
	.w1(32'h39488946),
	.w2(32'hb9d6ceb9),
	.w3(32'h39d768e4),
	.w4(32'hbbb86273),
	.w5(32'h3b92b68f),
	.w6(32'hba1c7488),
	.w7(32'hbb6cb6ee),
	.w8(32'h3a8f4007),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9a355),
	.w1(32'h3ab40184),
	.w2(32'hbab4e7d3),
	.w3(32'h3c217dc9),
	.w4(32'h3ba94181),
	.w5(32'h3b975fb1),
	.w6(32'h3c89399f),
	.w7(32'h3be63c75),
	.w8(32'hbc10aaa9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f375a),
	.w1(32'h3c92a44c),
	.w2(32'h3c433ffc),
	.w3(32'hba31352f),
	.w4(32'h3bb55dc5),
	.w5(32'h3b140e43),
	.w6(32'hbb80d76e),
	.w7(32'h3ac770d5),
	.w8(32'h3ad070ef),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40d7b6),
	.w1(32'hb921c6be),
	.w2(32'h3b76006b),
	.w3(32'hbad1d8a5),
	.w4(32'hbbd639dc),
	.w5(32'h3b2deadc),
	.w6(32'hbc1174fc),
	.w7(32'hbad021c2),
	.w8(32'hbb2490ab),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd67850),
	.w1(32'h3c83afd8),
	.w2(32'h3ac23286),
	.w3(32'h3bf3c03e),
	.w4(32'h3c0f2df6),
	.w5(32'hbb840271),
	.w6(32'hbbe396ab),
	.w7(32'hbb069891),
	.w8(32'h3b066219),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a6d02),
	.w1(32'hbb08747f),
	.w2(32'hba6586f9),
	.w3(32'hbc10f10c),
	.w4(32'hbafb080c),
	.w5(32'hbc0c4f3e),
	.w6(32'hbb61f8ec),
	.w7(32'h3aa36247),
	.w8(32'hbc1ace23),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f3692),
	.w1(32'hbbd78176),
	.w2(32'hba479b0c),
	.w3(32'hbccb60bc),
	.w4(32'hbd0310b6),
	.w5(32'hbbe71345),
	.w6(32'hbcc98d07),
	.w7(32'hbc4c3719),
	.w8(32'h3bd653d2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb0cde),
	.w1(32'hbc040d4b),
	.w2(32'h3b96f237),
	.w3(32'hbc2cdc0b),
	.w4(32'hbc30a020),
	.w5(32'h3c65d235),
	.w6(32'h3c1daa2d),
	.w7(32'hba52881c),
	.w8(32'h3c3b8e76),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f4699),
	.w1(32'hba5171e8),
	.w2(32'h3b9edf76),
	.w3(32'hbb74a9ad),
	.w4(32'hbb8912e3),
	.w5(32'h3a07ae46),
	.w6(32'hbab4860a),
	.w7(32'hbbf666be),
	.w8(32'h3b049a5a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fd943),
	.w1(32'h3bc0f337),
	.w2(32'hbb168098),
	.w3(32'h377254ac),
	.w4(32'h3ba7d3ea),
	.w5(32'hbb9e896e),
	.w6(32'h3a7193c5),
	.w7(32'h3ab65fb6),
	.w8(32'h3c1ff7f3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb749e88),
	.w1(32'hbba6ae4a),
	.w2(32'h3af1fe3a),
	.w3(32'hbbf59ab4),
	.w4(32'hbbe00d2d),
	.w5(32'h3a9256bc),
	.w6(32'h3c18c040),
	.w7(32'h3c11ab6d),
	.w8(32'h3a8d528e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf856c),
	.w1(32'h3af040fe),
	.w2(32'h3c2c0b0a),
	.w3(32'hbad5d5c7),
	.w4(32'hbb029bc6),
	.w5(32'h3bf49b8e),
	.w6(32'h3b063e89),
	.w7(32'h3b4eb28a),
	.w8(32'h3c405860),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5247d9),
	.w1(32'h3c23ccf7),
	.w2(32'hbb9431cd),
	.w3(32'h3c562b35),
	.w4(32'h3c5cef85),
	.w5(32'hbae27da7),
	.w6(32'h3c869183),
	.w7(32'h3c0a668a),
	.w8(32'h3b62c0cc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385fb0aa),
	.w1(32'hbc057010),
	.w2(32'h3bb4f5b5),
	.w3(32'h3bc5fc1d),
	.w4(32'hbb9ad134),
	.w5(32'h3b956f06),
	.w6(32'h3b87da6d),
	.w7(32'hbc514c37),
	.w8(32'hbb8d02d4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b221670),
	.w1(32'h39c2491d),
	.w2(32'h3bbf7a0b),
	.w3(32'h3c00d370),
	.w4(32'h3b1505cd),
	.w5(32'h3b80a218),
	.w6(32'hbb5b9e72),
	.w7(32'hba81dfa0),
	.w8(32'h3c08c01c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12fe06),
	.w1(32'h3bb6705f),
	.w2(32'hbb001128),
	.w3(32'h3bb0a443),
	.w4(32'h3b1e0c19),
	.w5(32'hbb296205),
	.w6(32'h3c256bcb),
	.w7(32'h3b9aab98),
	.w8(32'hbb5f27f2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11c35f),
	.w1(32'h3b9b11ed),
	.w2(32'h39e928ba),
	.w3(32'hbb5d912d),
	.w4(32'hba3e5c7b),
	.w5(32'hbb526dd0),
	.w6(32'hbc0946da),
	.w7(32'hbb0c28cd),
	.w8(32'hba702d15),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d0a04),
	.w1(32'h3c0a6c87),
	.w2(32'h3bdea2b8),
	.w3(32'hbb04bb0d),
	.w4(32'h3b95294d),
	.w5(32'h3c0535d8),
	.w6(32'h3adb46e0),
	.w7(32'h3c0a5591),
	.w8(32'h3b4999e7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f8ab9),
	.w1(32'h3c7ddb55),
	.w2(32'h3b97dc0b),
	.w3(32'h3c88e5ba),
	.w4(32'h3cb213d9),
	.w5(32'hbb5ede34),
	.w6(32'h3c2cab10),
	.w7(32'h3c88d19b),
	.w8(32'hbbed8ca8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb723d93),
	.w1(32'h3ac51973),
	.w2(32'h3b7519c3),
	.w3(32'hbc67cdea),
	.w4(32'hbc174c60),
	.w5(32'h3b9de0b9),
	.w6(32'hbce045d7),
	.w7(32'hbcb91fa2),
	.w8(32'hbb88c5d0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d6417),
	.w1(32'h3bf84110),
	.w2(32'hb94f5126),
	.w3(32'h3c1d924a),
	.w4(32'h3c384c60),
	.w5(32'hba2661d3),
	.w6(32'hbae657e4),
	.w7(32'hbb850510),
	.w8(32'h3a51d1be),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6c6da),
	.w1(32'hbbe6c247),
	.w2(32'hbbad0a8c),
	.w3(32'h3b0befa1),
	.w4(32'hb94d4fc9),
	.w5(32'hbbb860dc),
	.w6(32'h3c5cf806),
	.w7(32'h3c036862),
	.w8(32'hbc1a0ffd),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0bedd),
	.w1(32'hbba0fefa),
	.w2(32'hbbe0825d),
	.w3(32'hbba331a8),
	.w4(32'hbbfb6df7),
	.w5(32'hbc0d0e8f),
	.w6(32'hbc6ed949),
	.w7(32'hbc41833a),
	.w8(32'hba744c88),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ce487),
	.w1(32'hbbbfac38),
	.w2(32'h3c1b20a6),
	.w3(32'hbc03200f),
	.w4(32'hba8774b5),
	.w5(32'h3ba76fef),
	.w6(32'hbad99646),
	.w7(32'hba6f219a),
	.w8(32'hbb76a1c7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a1ce7),
	.w1(32'h3a3436a0),
	.w2(32'hbc15f7b3),
	.w3(32'hbc5eeee5),
	.w4(32'hbc3ffc11),
	.w5(32'hbb58501a),
	.w6(32'hbcd063a1),
	.w7(32'hbcc30cc2),
	.w8(32'h3b389de2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c166b),
	.w1(32'h3ba45b80),
	.w2(32'h3c1e1a4b),
	.w3(32'h3c513107),
	.w4(32'h3c7f7d39),
	.w5(32'h3bb2a423),
	.w6(32'h3cb61c24),
	.w7(32'h3cd166cd),
	.w8(32'h3bfc1386),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6115d),
	.w1(32'h3b6fb3f2),
	.w2(32'h3a3d299a),
	.w3(32'hb94690ac),
	.w4(32'hba9c7449),
	.w5(32'hbc0808d0),
	.w6(32'h3b00cc3a),
	.w7(32'h38054418),
	.w8(32'hbc2f3b4b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9352da),
	.w1(32'hbb154641),
	.w2(32'h3af5f32d),
	.w3(32'hbc77a82c),
	.w4(32'hbc82df7f),
	.w5(32'hbb59d568),
	.w6(32'hbcf8be3d),
	.w7(32'hbcc22504),
	.w8(32'hbb802b68),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0700f2),
	.w1(32'h39eb3c76),
	.w2(32'h3b3aa237),
	.w3(32'hbaedda27),
	.w4(32'h3c0481ec),
	.w5(32'hbb894fd7),
	.w6(32'hbc627026),
	.w7(32'hbb172d3a),
	.w8(32'hbbc7a29c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc004085),
	.w1(32'hbba592d5),
	.w2(32'hbb83b535),
	.w3(32'hbc585324),
	.w4(32'hbb17c3dc),
	.w5(32'hbbcaa280),
	.w6(32'hbc2acbbc),
	.w7(32'hbb386209),
	.w8(32'hbb45bfee),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc01432),
	.w1(32'h39ad52fb),
	.w2(32'hbb7a6096),
	.w3(32'hbc70e740),
	.w4(32'hbc4409fc),
	.w5(32'hbbe2a15a),
	.w6(32'hbcb14ec5),
	.w7(32'hbcc80729),
	.w8(32'hbb678f5f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8778a1),
	.w1(32'hba18fb55),
	.w2(32'hbb1cb824),
	.w3(32'hbbaba538),
	.w4(32'hb8a05694),
	.w5(32'h3959f178),
	.w6(32'hbaa11db5),
	.w7(32'h3ba25697),
	.w8(32'h3abe0c5f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ccde2),
	.w1(32'hbad973d0),
	.w2(32'hbc28823c),
	.w3(32'hbc03d2e7),
	.w4(32'hbba8d14f),
	.w5(32'hbc5dda0b),
	.w6(32'hbb53242c),
	.w7(32'hbab5cde3),
	.w8(32'hbc5b2f67),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52c7c0),
	.w1(32'hbb8f6e13),
	.w2(32'h3c2d5574),
	.w3(32'hbc3ef7ec),
	.w4(32'hbaaaf68d),
	.w5(32'h3b948fcf),
	.w6(32'hbc508cfa),
	.w7(32'hbae1988c),
	.w8(32'hbc29cc36),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42dce3),
	.w1(32'h3c52cf70),
	.w2(32'h3ad603b1),
	.w3(32'h3a60992f),
	.w4(32'h3c00b164),
	.w5(32'h3af86b8c),
	.w6(32'hbc4b050a),
	.w7(32'h3b13f70c),
	.w8(32'hbb107021),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad159ae),
	.w1(32'hbb117689),
	.w2(32'hba5d4cd7),
	.w3(32'hbb277b08),
	.w4(32'hbbdb0973),
	.w5(32'hbb9ab8f4),
	.w6(32'hbc949c77),
	.w7(32'hbc9c3d47),
	.w8(32'hbab66122),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6994af),
	.w1(32'hb8c7e404),
	.w2(32'h3bf99876),
	.w3(32'hbba534b4),
	.w4(32'hbbdca266),
	.w5(32'h3b361677),
	.w6(32'hbc23c7da),
	.w7(32'hbc258b75),
	.w8(32'hbbb45d22),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd60075),
	.w1(32'hbb09c831),
	.w2(32'hba952bdb),
	.w3(32'hbc34005b),
	.w4(32'hbbf7bab0),
	.w5(32'hbb420d23),
	.w6(32'hbca14474),
	.w7(32'hbc0a6edd),
	.w8(32'hbb5a1926),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb28d18),
	.w1(32'hbbd8df69),
	.w2(32'hbb34fb7e),
	.w3(32'hbba33f7f),
	.w4(32'hbb8b4965),
	.w5(32'hbb9e10ab),
	.w6(32'hbb726029),
	.w7(32'hbb8abd73),
	.w8(32'hbb8259eb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d9c64),
	.w1(32'hbb17c118),
	.w2(32'hbbcb2ee2),
	.w3(32'hbb759893),
	.w4(32'hbad9a3af),
	.w5(32'hbb1a9c89),
	.w6(32'hbb98e05a),
	.w7(32'hb9ebb71f),
	.w8(32'hbb679ded),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bba0b),
	.w1(32'h3bd9a6e2),
	.w2(32'hba319af0),
	.w3(32'h3c0144e5),
	.w4(32'h3c079aac),
	.w5(32'hbc4aafe5),
	.w6(32'h3b5595ea),
	.w7(32'h3b789f46),
	.w8(32'hbc0b43a6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bb399),
	.w1(32'h3a21375f),
	.w2(32'h3c819cc0),
	.w3(32'hbcae74fc),
	.w4(32'hbc522346),
	.w5(32'h3c8c3fcd),
	.w6(32'hbc9a66fb),
	.w7(32'hbbd17c2e),
	.w8(32'h3ba97b91),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0afb74),
	.w1(32'h3bdb0e5b),
	.w2(32'h3cd86f40),
	.w3(32'h3c4a2ea8),
	.w4(32'h3b9bec88),
	.w5(32'h3d01ef76),
	.w6(32'h3b2c0640),
	.w7(32'hbb9a20d6),
	.w8(32'h3d0797b1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf1fa6c),
	.w1(32'h3ce2dbdf),
	.w2(32'hbbf60b93),
	.w3(32'h3d142ba0),
	.w4(32'h3d07196d),
	.w5(32'hbc29dc4c),
	.w6(32'h3d22783b),
	.w7(32'h3d0f9107),
	.w8(32'hbbe35ed3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1489a1),
	.w1(32'hbc6660ac),
	.w2(32'h3ac24837),
	.w3(32'hbc436e36),
	.w4(32'hbc6f3869),
	.w5(32'h391c43be),
	.w6(32'hbbe8d32d),
	.w7(32'hbbf4cc14),
	.w8(32'hbaf3f856),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be26277),
	.w1(32'h3be374d8),
	.w2(32'h3ab1c7af),
	.w3(32'h3bc815de),
	.w4(32'h3bf5b2be),
	.w5(32'h3bad4a2e),
	.w6(32'h3b2289e1),
	.w7(32'h3b6fe959),
	.w8(32'hbb87784a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0eb01),
	.w1(32'h3bfed6af),
	.w2(32'hbc739540),
	.w3(32'h3c191ac1),
	.w4(32'h3c512026),
	.w5(32'hbae2cff9),
	.w6(32'hbaa67f3a),
	.w7(32'h3c05789f),
	.w8(32'h3c848c9a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81bcea),
	.w1(32'hbb2b3031),
	.w2(32'hbb29aa01),
	.w3(32'h3c52e12a),
	.w4(32'h3c853c1d),
	.w5(32'hbc2f32c2),
	.w6(32'h3d27f852),
	.w7(32'h3ccee2ee),
	.w8(32'hbc319a19),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb395aa8),
	.w1(32'hbaf00191),
	.w2(32'h3b236225),
	.w3(32'hbc0f995f),
	.w4(32'hbc45a343),
	.w5(32'h3b71bc6e),
	.w6(32'hbc91a0cd),
	.w7(32'hbc84a939),
	.w8(32'h3acbc59d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed6cae),
	.w1(32'hbb07e9ac),
	.w2(32'h3b9742b6),
	.w3(32'hbb42341b),
	.w4(32'h39a2f0ca),
	.w5(32'hbb30609a),
	.w6(32'hbc3d9575),
	.w7(32'hbc0eac63),
	.w8(32'h3ac13b5a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f4336),
	.w1(32'h3b685d33),
	.w2(32'hbacd7ab5),
	.w3(32'hb86db118),
	.w4(32'h3c20a82e),
	.w5(32'h3b91c64d),
	.w6(32'h3bd59575),
	.w7(32'h3c165da9),
	.w8(32'h3bcf5c43),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d5cdf),
	.w1(32'h3c091914),
	.w2(32'h3b475f1a),
	.w3(32'h3b78daad),
	.w4(32'hbaa18a70),
	.w5(32'h3be53546),
	.w6(32'h3bade1cc),
	.w7(32'hbb2bb933),
	.w8(32'h3c15f623),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb73229),
	.w1(32'h3ac797e7),
	.w2(32'h3a901055),
	.w3(32'h3c1f84b4),
	.w4(32'hbb5f26cf),
	.w5(32'h3ad2ad6a),
	.w6(32'h3c1a561a),
	.w7(32'h3b6e67c9),
	.w8(32'h3a46bf0a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb309b),
	.w1(32'h3aa0c0d6),
	.w2(32'hba057f39),
	.w3(32'hbb57b4f3),
	.w4(32'hba525b07),
	.w5(32'h3b0a0186),
	.w6(32'h3b8c534a),
	.w7(32'h3bbc9a23),
	.w8(32'hbbd243e0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84a505),
	.w1(32'h3b73b51b),
	.w2(32'h3b62fd6a),
	.w3(32'h39c7f2ac),
	.w4(32'hbb5b0c5e),
	.w5(32'h3b137c95),
	.w6(32'hbba1c87e),
	.w7(32'hbbbdde79),
	.w8(32'h39abc916),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce224e),
	.w1(32'h3ada80f6),
	.w2(32'h3c6302bc),
	.w3(32'h3a58424c),
	.w4(32'hbb1d9c09),
	.w5(32'h3b11eef1),
	.w6(32'hbbc5ee7c),
	.w7(32'hbb468a37),
	.w8(32'hbc6fcd51),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d443d),
	.w1(32'h3c7763b5),
	.w2(32'h3ad72e72),
	.w3(32'h3c20f82a),
	.w4(32'hb9f31d45),
	.w5(32'h3a2b584f),
	.w6(32'hbc90fc40),
	.w7(32'hbc9b0f33),
	.w8(32'hbbdffaaf),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc9723),
	.w1(32'h39e1a0bd),
	.w2(32'hbc2863d5),
	.w3(32'hbbcf1bfc),
	.w4(32'hbb7cccf2),
	.w5(32'hbc580719),
	.w6(32'hbbb0b9f4),
	.w7(32'hbbc9dc18),
	.w8(32'hbc72a6ee),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1949d8),
	.w1(32'hbb86767a),
	.w2(32'hbbb56203),
	.w3(32'hbc6fec6a),
	.w4(32'hbb942de4),
	.w5(32'h3b1edbc0),
	.w6(32'hbc7fafe7),
	.w7(32'hbbc03441),
	.w8(32'h3c17ac59),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3941d6ba),
	.w1(32'h39a767d8),
	.w2(32'h3baf4556),
	.w3(32'h3a4b7640),
	.w4(32'hb9cba708),
	.w5(32'h3c3a4e88),
	.w6(32'h3b40fdc1),
	.w7(32'h3ae4dcb8),
	.w8(32'h3b3ba78d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8d37d),
	.w1(32'hbb43a79e),
	.w2(32'h3bc9bf06),
	.w3(32'hbba20a2a),
	.w4(32'hbc0ebca1),
	.w5(32'h3b4e809f),
	.w6(32'hbc23d2d1),
	.w7(32'hbc7416ec),
	.w8(32'h3b99b8ef),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24a32f),
	.w1(32'hbb99f5b6),
	.w2(32'hbb418fe2),
	.w3(32'h3b2c3cf3),
	.w4(32'hbbff36eb),
	.w5(32'hbbcb18f4),
	.w6(32'hbb705c80),
	.w7(32'hbbd743a3),
	.w8(32'hbb12d24b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1df519),
	.w1(32'h3acfe347),
	.w2(32'h3c1befc6),
	.w3(32'hbbdf4112),
	.w4(32'hbc566ba2),
	.w5(32'h3bf98495),
	.w6(32'hbca2ac27),
	.w7(32'hbc83130a),
	.w8(32'h3bd8c032),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1713ff),
	.w1(32'h3a8d1458),
	.w2(32'hbba07a8f),
	.w3(32'h3c4f3a75),
	.w4(32'h3b86ec6d),
	.w5(32'hb9b0d287),
	.w6(32'h3c0f8afb),
	.w7(32'hbb1b8a38),
	.w8(32'h39e80296),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe56a43),
	.w1(32'hb8a3f592),
	.w2(32'hbbf24e7e),
	.w3(32'h3c4a47ac),
	.w4(32'h3c893b9f),
	.w5(32'h3c361cfb),
	.w6(32'h39c42488),
	.w7(32'h3bd054bb),
	.w8(32'h3c42038e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd18f00),
	.w1(32'hbc378dfa),
	.w2(32'hbc1eda1a),
	.w3(32'h3b4708c5),
	.w4(32'hbb87017f),
	.w5(32'h3b1eea06),
	.w6(32'h3c2466a7),
	.w7(32'hbba4791d),
	.w8(32'h3bdf96f2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c3c49),
	.w1(32'hbb0a202c),
	.w2(32'hbb234607),
	.w3(32'h3c170126),
	.w4(32'h3c1b0385),
	.w5(32'h3b3b2f09),
	.w6(32'h3c7de275),
	.w7(32'h3c35030e),
	.w8(32'h3b7c0b1b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac44288),
	.w1(32'hbb18053e),
	.w2(32'h3c99eefe),
	.w3(32'h3bbcc36f),
	.w4(32'h3b72941c),
	.w5(32'h3ba7d3c5),
	.w6(32'h3c357d8c),
	.w7(32'h3c039ced),
	.w8(32'h3bdf39cb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c675069),
	.w1(32'h3c0e2670),
	.w2(32'h3b0cfd9b),
	.w3(32'h3ad3af67),
	.w4(32'hba61e1ad),
	.w5(32'hba81f00a),
	.w6(32'h3ac3567c),
	.w7(32'h39c1a599),
	.w8(32'h3c064081),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5553fb),
	.w1(32'h3af5ffbe),
	.w2(32'h3b8cf8af),
	.w3(32'hbb60c2bb),
	.w4(32'h3a8c22ba),
	.w5(32'h3aafc645),
	.w6(32'h3be87316),
	.w7(32'h3bca04fa),
	.w8(32'hbb72569d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3262b),
	.w1(32'hba31f559),
	.w2(32'h3c1d47eb),
	.w3(32'hbbb826db),
	.w4(32'hbc0c9c4e),
	.w5(32'hbad900c9),
	.w6(32'hba7914f3),
	.w7(32'h3b8eb103),
	.w8(32'h3b5215e0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe7f41),
	.w1(32'h3b341b9c),
	.w2(32'h3c50b0f3),
	.w3(32'hba5d0506),
	.w4(32'hbba0a2a9),
	.w5(32'h3c3474f1),
	.w6(32'h3ba4099d),
	.w7(32'h3b8592bf),
	.w8(32'hbaf11083),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd236a7),
	.w1(32'h3af9ecf8),
	.w2(32'hbb99250d),
	.w3(32'h3c451b22),
	.w4(32'h3c003168),
	.w5(32'hbae4ed11),
	.w6(32'h3af667cc),
	.w7(32'hbb27ce73),
	.w8(32'hb985aba2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf2a66),
	.w1(32'hbb896b6e),
	.w2(32'h3b338646),
	.w3(32'hbbaafc21),
	.w4(32'hbb659030),
	.w5(32'hbb34e518),
	.w6(32'hbb185dd7),
	.w7(32'hba9dd6e1),
	.w8(32'hbb3a1322),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac9907),
	.w1(32'hbbdfd235),
	.w2(32'hbc3bced5),
	.w3(32'hbc0485c2),
	.w4(32'hbc22e60d),
	.w5(32'hbc8fbd81),
	.w6(32'hbbab8a6c),
	.w7(32'hbc1ae44e),
	.w8(32'hbbaa5240),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43a6c8),
	.w1(32'h3c287ce6),
	.w2(32'hbb8f9402),
	.w3(32'h3b3f83d5),
	.w4(32'h3b2dcee2),
	.w5(32'hba97e68b),
	.w6(32'h3c0499a1),
	.w7(32'hba260e9d),
	.w8(32'h3bb35e23),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d33ad),
	.w1(32'hbaeb418c),
	.w2(32'h3c21043a),
	.w3(32'hbac170fb),
	.w4(32'h3b47dc40),
	.w5(32'h3bb71807),
	.w6(32'h3c03f077),
	.w7(32'h3c18d27f),
	.w8(32'hbb425255),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cc198),
	.w1(32'h3c60c216),
	.w2(32'h3bf84166),
	.w3(32'h3c094ee9),
	.w4(32'h3c976e6f),
	.w5(32'h3b4e0582),
	.w6(32'hbb7347b0),
	.w7(32'h39865f48),
	.w8(32'hbc12557c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3b7d6),
	.w1(32'h3b2e1e54),
	.w2(32'h3c2dea20),
	.w3(32'hbb2277ed),
	.w4(32'hbb1cd37e),
	.w5(32'hbbbf3534),
	.w6(32'hbc7b2f7b),
	.w7(32'hbc9195f5),
	.w8(32'hbc41b99b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8d2a2),
	.w1(32'hbac6f52a),
	.w2(32'hb8ce4d24),
	.w3(32'hbc996e44),
	.w4(32'hbc2f2470),
	.w5(32'h3c62862a),
	.w6(32'hbd0e8fe2),
	.w7(32'hbca85bae),
	.w8(32'h3c80c745),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e72b7),
	.w1(32'hbc3474c0),
	.w2(32'h3ad91955),
	.w3(32'hbabf3fb3),
	.w4(32'hbbbdb555),
	.w5(32'h3cb310ee),
	.w6(32'h3b83b959),
	.w7(32'hbbac3c16),
	.w8(32'h3c91afd3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb625d8),
	.w1(32'h3b63f1e3),
	.w2(32'hbc33d06a),
	.w3(32'h3cbbe093),
	.w4(32'h3ceac463),
	.w5(32'hbb6d54bd),
	.w6(32'h3ceeb037),
	.w7(32'h3ccdef8a),
	.w8(32'h3c4a93ec),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc847b7a),
	.w1(32'hbc2da3fc),
	.w2(32'h3a4b06fd),
	.w3(32'hbbf4cd8f),
	.w4(32'hba20c69d),
	.w5(32'h3c1026a3),
	.w6(32'h3ca8ec2c),
	.w7(32'h3c50917e),
	.w8(32'hbab20ac5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaf7d1),
	.w1(32'hbbbf04b7),
	.w2(32'h3ad7157c),
	.w3(32'h3b5c1d0c),
	.w4(32'hba9dc0ad),
	.w5(32'hbad26ac7),
	.w6(32'hbb207e0c),
	.w7(32'hbbd23539),
	.w8(32'hbb544970),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba922426),
	.w1(32'h3bbb6e87),
	.w2(32'h3c020ec8),
	.w3(32'hbbbc4f54),
	.w4(32'h3bc689fc),
	.w5(32'h3b988ff7),
	.w6(32'h3b8f9a14),
	.w7(32'h3c914316),
	.w8(32'hbc0c6e51),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf6db4),
	.w1(32'hbc1e408e),
	.w2(32'h39a94c09),
	.w3(32'hbb176948),
	.w4(32'hbc6aee69),
	.w5(32'hbbbe18c5),
	.w6(32'hb8541734),
	.w7(32'hbc4d19b8),
	.w8(32'hbbe2cb1b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c56b0),
	.w1(32'h3b57baea),
	.w2(32'hbb84b755),
	.w3(32'hbb9a317b),
	.w4(32'h3b536e38),
	.w5(32'hbbd48548),
	.w6(32'hbc4af5a9),
	.w7(32'hbb337b59),
	.w8(32'h3afcd996),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04b07c),
	.w1(32'hbbb58ec2),
	.w2(32'hbb77fa3f),
	.w3(32'hbc1dc5df),
	.w4(32'hbbc0cb3e),
	.w5(32'hbc01238c),
	.w6(32'h3ba5b89c),
	.w7(32'h3ba0cb13),
	.w8(32'hbc003f4f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc94a42),
	.w1(32'h39af29d8),
	.w2(32'h3c9d1609),
	.w3(32'hbc1dc29a),
	.w4(32'hb9b91038),
	.w5(32'h3c87eafb),
	.w6(32'hbbde4bb3),
	.w7(32'hbb68b168),
	.w8(32'h3c45b920),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e8818),
	.w1(32'h3c9699db),
	.w2(32'h3c476ece),
	.w3(32'h3c42972d),
	.w4(32'h3c4bd5d8),
	.w5(32'h3c2125a8),
	.w6(32'h3ba447a2),
	.w7(32'h3bb2d2d5),
	.w8(32'h3ba16822),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad6bf7),
	.w1(32'h3c0ad32c),
	.w2(32'hbb2bbb0b),
	.w3(32'h3bcefb56),
	.w4(32'h3c29047f),
	.w5(32'h3bac343d),
	.w6(32'h3bbdf386),
	.w7(32'h3bdf8ac5),
	.w8(32'hbadf015c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b964263),
	.w1(32'h3b86afe0),
	.w2(32'hbb0f7ea5),
	.w3(32'h3ab73c37),
	.w4(32'hbb98b5a9),
	.w5(32'hbb6ac57d),
	.w6(32'h3acb33d7),
	.w7(32'hbb68848a),
	.w8(32'hbb7e9bbd),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6c878),
	.w1(32'hbbbf4b64),
	.w2(32'hba91d962),
	.w3(32'hbc000860),
	.w4(32'hbc1622b2),
	.w5(32'hbbd2e0a4),
	.w6(32'hbbba6f01),
	.w7(32'hbc14876e),
	.w8(32'hbba9f544),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30c097),
	.w1(32'h39cdcbe3),
	.w2(32'hbc09ae0b),
	.w3(32'hbbe05746),
	.w4(32'hbbe79c01),
	.w5(32'hbba1cd3f),
	.w6(32'hbc02c103),
	.w7(32'hbbe2c6c2),
	.w8(32'h3c884dee),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc295462),
	.w1(32'hbbc55a78),
	.w2(32'h3ae0474c),
	.w3(32'hbc147c28),
	.w4(32'hbc10bdf3),
	.w5(32'h3b10450d),
	.w6(32'h3c8b13f0),
	.w7(32'h3c8e14a9),
	.w8(32'h3b746ac9),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b663320),
	.w1(32'h3b3f995d),
	.w2(32'h3a8cffa2),
	.w3(32'hba09a14a),
	.w4(32'hbb45938d),
	.w5(32'hb9546143),
	.w6(32'h3aee9307),
	.w7(32'hb9d18bcd),
	.w8(32'hba8a38bf),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05373c),
	.w1(32'h3b79d77b),
	.w2(32'h3b2c89c2),
	.w3(32'h3b33a1ae),
	.w4(32'h3be155be),
	.w5(32'h3b7d6e08),
	.w6(32'h3b2fa590),
	.w7(32'h3bd23539),
	.w8(32'h3c27553f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4eae2),
	.w1(32'hba18b975),
	.w2(32'hbbb2815b),
	.w3(32'h3b904fda),
	.w4(32'h3af745b7),
	.w5(32'hbb093387),
	.w6(32'h3c4f2a9f),
	.w7(32'h3c0ca7d0),
	.w8(32'hbbc1176a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0219d3),
	.w1(32'hbc1693ad),
	.w2(32'h3c048d93),
	.w3(32'hbbe05320),
	.w4(32'hbbe06c8f),
	.w5(32'h3b85f400),
	.w6(32'hbbefbd1d),
	.w7(32'hbc05140d),
	.w8(32'h3c271e53),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabdc19),
	.w1(32'h3b9bdc6c),
	.w2(32'hbbb9b19e),
	.w3(32'hbb94b392),
	.w4(32'hbb6c970d),
	.w5(32'hbb52b7e7),
	.w6(32'hbc5e3350),
	.w7(32'hbc5fb789),
	.w8(32'hbbb1636b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18ef96),
	.w1(32'hbb0c89a3),
	.w2(32'hb9bccede),
	.w3(32'hba75a925),
	.w4(32'hbbd62223),
	.w5(32'h3bb2011d),
	.w6(32'hbb70cb4a),
	.w7(32'hbbadb86f),
	.w8(32'h3b5aa313),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a051e),
	.w1(32'hbbc0ea62),
	.w2(32'h3ae1eb42),
	.w3(32'hb96cf4ee),
	.w4(32'hbac4c387),
	.w5(32'hbb9a57e3),
	.w6(32'hbc254208),
	.w7(32'hbc6b1bae),
	.w8(32'hbc295600),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde3887),
	.w1(32'hbc0f92ca),
	.w2(32'h3b087c49),
	.w3(32'hbbddd137),
	.w4(32'hbc201bef),
	.w5(32'hb9c7705c),
	.w6(32'hbc41161e),
	.w7(32'hbc1e5659),
	.w8(32'hbab0ee14),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb801777),
	.w1(32'hbb187c56),
	.w2(32'hbad77578),
	.w3(32'hbc147bf1),
	.w4(32'hbbd90108),
	.w5(32'hbbdf8eba),
	.w6(32'hbba3e244),
	.w7(32'hbb9432dd),
	.w8(32'hbbb7a076),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0273b5),
	.w1(32'hbb94a0cc),
	.w2(32'h3ad2d4ee),
	.w3(32'hbbca88c0),
	.w4(32'hbb9eda0a),
	.w5(32'h3bac61d8),
	.w6(32'hbbbf09f2),
	.w7(32'hbb9523a8),
	.w8(32'h3c0fa00a),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb10b3e),
	.w1(32'h3c1c5f57),
	.w2(32'hbc10d691),
	.w3(32'h3c20c27c),
	.w4(32'h3c0ab300),
	.w5(32'h3a91fa31),
	.w6(32'h3c67a6fc),
	.w7(32'h3bcfe655),
	.w8(32'hbc09289d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8296fb),
	.w1(32'h3a2a748d),
	.w2(32'hb7a2d953),
	.w3(32'hbbca2a33),
	.w4(32'hbab27fc6),
	.w5(32'h3a450b54),
	.w6(32'hbbfe0ca3),
	.w7(32'h3a91c0e8),
	.w8(32'h3aaae19c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf87787),
	.w1(32'hbaa77207),
	.w2(32'hbb0d821c),
	.w3(32'h39052e4a),
	.w4(32'hba1ca9dc),
	.w5(32'hbb0bdc5a),
	.w6(32'h3a83d3c1),
	.w7(32'h394ec3d2),
	.w8(32'h3aab2e44),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb346e8),
	.w1(32'hbb1162b7),
	.w2(32'hbb13f7f7),
	.w3(32'h3b15c4c3),
	.w4(32'hbb7fe00a),
	.w5(32'h3c056c54),
	.w6(32'h3badab8b),
	.w7(32'h3bc4e7bb),
	.w8(32'hbb0fdb70),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93a786),
	.w1(32'hbc80b7fe),
	.w2(32'hbac64b04),
	.w3(32'hbc4da353),
	.w4(32'hbc36681b),
	.w5(32'hbab5ce93),
	.w6(32'hbc3e9af8),
	.w7(32'hbc345b22),
	.w8(32'hbb5bdb2b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b407e),
	.w1(32'h3b35b16b),
	.w2(32'h3c1d0062),
	.w3(32'h39835260),
	.w4(32'hba1f98c4),
	.w5(32'h3bf5bcb0),
	.w6(32'hbb93886e),
	.w7(32'hbaad2881),
	.w8(32'h3b04da89),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6e241),
	.w1(32'h39edcffa),
	.w2(32'h3c1d8f8b),
	.w3(32'h3bd29cae),
	.w4(32'h3b8bec80),
	.w5(32'h3c2a2f95),
	.w6(32'h3baa9c26),
	.w7(32'hbbbf6145),
	.w8(32'h38e69cab),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dfac7),
	.w1(32'h3b5582ab),
	.w2(32'h3b85f2a1),
	.w3(32'h3b870b2b),
	.w4(32'h3b88b2e6),
	.w5(32'h3b9ac23d),
	.w6(32'h3ba65490),
	.w7(32'h3aafccae),
	.w8(32'h3b1b192e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6088b6),
	.w1(32'h3b05576e),
	.w2(32'hb9f63dac),
	.w3(32'h3acf90df),
	.w4(32'h3aec0d7e),
	.w5(32'h3b58d75b),
	.w6(32'h3ab2eaa9),
	.w7(32'hba39e6dd),
	.w8(32'hbbcbd22d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a1a73),
	.w1(32'h3c0cf8f3),
	.w2(32'h3a5e5afe),
	.w3(32'hbb46b582),
	.w4(32'hbaf00fc3),
	.w5(32'h396ac5a1),
	.w6(32'hbc562537),
	.w7(32'hbc36eaac),
	.w8(32'hba1519b4),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d14d0),
	.w1(32'hba61b442),
	.w2(32'hbbc9fd8f),
	.w3(32'h3afa461e),
	.w4(32'h3a8bedaf),
	.w5(32'hbb65318a),
	.w6(32'h3a58718e),
	.w7(32'hba9e8a7d),
	.w8(32'h3b8ec690),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94f35c),
	.w1(32'hbada6c26),
	.w2(32'h3b7bf6be),
	.w3(32'hbc550de3),
	.w4(32'h3b24a700),
	.w5(32'h39bae562),
	.w6(32'hbc494a5a),
	.w7(32'h3a07b497),
	.w8(32'hbb942b0c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b5a7b),
	.w1(32'hbb4c13b0),
	.w2(32'h3c5a513e),
	.w3(32'hbbe97df9),
	.w4(32'hbbc9b40b),
	.w5(32'h39d4271c),
	.w6(32'hbc25a337),
	.w7(32'hbbfdf4c0),
	.w8(32'hbbf8e09d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c641a23),
	.w1(32'h3b7fe135),
	.w2(32'h3b2ffd85),
	.w3(32'h3bf0a289),
	.w4(32'h3bc81229),
	.w5(32'h3b674641),
	.w6(32'hbbba6192),
	.w7(32'h3b3e1524),
	.w8(32'h3a97d0f6),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306716),
	.w1(32'h3c21aac5),
	.w2(32'hbbcf4ff6),
	.w3(32'hbc41474f),
	.w4(32'hbafc438c),
	.w5(32'hbb1fe0f7),
	.w6(32'hbc102fc5),
	.w7(32'hbb8c1974),
	.w8(32'hbbd6c30b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64fae2),
	.w1(32'hbb138f21),
	.w2(32'h3aa78d11),
	.w3(32'hba8b4cc3),
	.w4(32'hbb7b47c4),
	.w5(32'hbb058791),
	.w6(32'hbc13573d),
	.w7(32'hbbe58751),
	.w8(32'hbc30431a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f9186),
	.w1(32'h3a987fc1),
	.w2(32'h3c4ec7d4),
	.w3(32'h3bb3f7b1),
	.w4(32'h3bf8841a),
	.w5(32'h3c5d00b6),
	.w6(32'h3afbff4d),
	.w7(32'h3c207f50),
	.w8(32'h3c7a3938),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf71abf),
	.w1(32'hbc93b15c),
	.w2(32'hbb41bba6),
	.w3(32'hbb09626e),
	.w4(32'hbcc5dcda),
	.w5(32'hbbacd5b1),
	.w6(32'h3a2e033b),
	.w7(32'hbc7eea45),
	.w8(32'hbb5f5968),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a1666),
	.w1(32'hbbf326e3),
	.w2(32'h3be0e025),
	.w3(32'hbb2c7f2e),
	.w4(32'hba3a9a9d),
	.w5(32'hbbb44242),
	.w6(32'hbaa31820),
	.w7(32'hb91d8fe6),
	.w8(32'hbc2faf8a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45b4de),
	.w1(32'hbb96ae13),
	.w2(32'h3a75294a),
	.w3(32'hbc239686),
	.w4(32'hbb94b00f),
	.w5(32'hbb8dd9b7),
	.w6(32'hbc023553),
	.w7(32'h3b894d3f),
	.w8(32'hbc41505e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dc0d0),
	.w1(32'h3cfd09f1),
	.w2(32'hbb56b86e),
	.w3(32'h3b0dd5d3),
	.w4(32'h3c56ca53),
	.w5(32'h391d469f),
	.w6(32'hbaaabefe),
	.w7(32'h3a2d0f32),
	.w8(32'h3c31410f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c177eb),
	.w1(32'hbc1f67b8),
	.w2(32'h3c299d1f),
	.w3(32'h3c5fdd52),
	.w4(32'h3c0a0982),
	.w5(32'h3b11a11e),
	.w6(32'h3c93fdd7),
	.w7(32'h3c8a891d),
	.w8(32'h3aea5edf),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c146ade),
	.w1(32'hbadfffa4),
	.w2(32'hb8914d75),
	.w3(32'h3c0c115b),
	.w4(32'h3bc570ec),
	.w5(32'hbb0afd11),
	.w6(32'h3bf06d77),
	.w7(32'h3b93aada),
	.w8(32'hba99121f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38c56e),
	.w1(32'hbb980758),
	.w2(32'h392fdde7),
	.w3(32'hb93beff8),
	.w4(32'hb8a3f48b),
	.w5(32'h3ab1474b),
	.w6(32'hba159fa7),
	.w7(32'hbaf3081c),
	.w8(32'h3b86d1cd),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc5d88),
	.w1(32'h3bbfbde3),
	.w2(32'h3bd302ad),
	.w3(32'h3bf953a6),
	.w4(32'hbbd5a6cd),
	.w5(32'h3c0b95d0),
	.w6(32'h3c021d02),
	.w7(32'hbaff326c),
	.w8(32'hbbaf8461),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e23a5),
	.w1(32'h3c8d1f79),
	.w2(32'h3ba4d62a),
	.w3(32'hbbab70f2),
	.w4(32'h3aa0b496),
	.w5(32'hbbad6d8e),
	.w6(32'hbc98e8fd),
	.w7(32'hbbab3ef7),
	.w8(32'hbc4a7958),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5a688),
	.w1(32'h3ca1468d),
	.w2(32'h395784c8),
	.w3(32'h3ab35d69),
	.w4(32'h3adf4a78),
	.w5(32'h3ac57bc8),
	.w6(32'hbaa69266),
	.w7(32'h3b7c210d),
	.w8(32'hbba93ad7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c260d9d),
	.w1(32'h3c898653),
	.w2(32'hbb04453b),
	.w3(32'hbb7b64cf),
	.w4(32'h3c2912a2),
	.w5(32'hbbf3dfdb),
	.w6(32'hbc835588),
	.w7(32'h3b65b9fa),
	.w8(32'hbad2d291),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8e0cc),
	.w1(32'h3c0a0ff7),
	.w2(32'h3c283841),
	.w3(32'h3c183b57),
	.w4(32'h3c1c6bc5),
	.w5(32'h3b75c459),
	.w6(32'h399736bd),
	.w7(32'h3b8ccdbd),
	.w8(32'hbbe0809c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc021433),
	.w1(32'hbb60d480),
	.w2(32'hb9bd6c53),
	.w3(32'hbb8c3dc3),
	.w4(32'h3b3fd8ed),
	.w5(32'h39cb1802),
	.w6(32'hbbd9b314),
	.w7(32'hbb323c85),
	.w8(32'hbbe81a08),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c8321),
	.w1(32'h3ac1c770),
	.w2(32'hba236f13),
	.w3(32'h3b6c29fb),
	.w4(32'h3c235a32),
	.w5(32'hbb961178),
	.w6(32'h3b0acec2),
	.w7(32'h3c1689be),
	.w8(32'hbb8d5a29),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb894565e),
	.w1(32'hba354725),
	.w2(32'h3c2a05da),
	.w3(32'hbac2f0c3),
	.w4(32'hbb2bffae),
	.w5(32'h3c33737f),
	.w6(32'hbbd50293),
	.w7(32'hbb0b6981),
	.w8(32'h3bd05000),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44655c),
	.w1(32'h3a13dfe9),
	.w2(32'h3b2eb6c1),
	.w3(32'h3a6d669d),
	.w4(32'hbbd02746),
	.w5(32'h3b5f6b19),
	.w6(32'hbba9d434),
	.w7(32'hbc062aa8),
	.w8(32'hbb0b259d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb867b7c),
	.w1(32'hb9eb5d28),
	.w2(32'h3aaa98eb),
	.w3(32'hbb40294f),
	.w4(32'h3b0264af),
	.w5(32'hba137b6d),
	.w6(32'hbbcd4997),
	.w7(32'hbb250835),
	.w8(32'hbb689db6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb97348),
	.w1(32'h39ba08e2),
	.w2(32'h3b154f6d),
	.w3(32'hbb8b348c),
	.w4(32'hbb3f2443),
	.w5(32'h3c413172),
	.w6(32'hbbe7b8f7),
	.w7(32'hbbacae09),
	.w8(32'h3c5ca984),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b226133),
	.w1(32'hbb1b14ca),
	.w2(32'hbb0bee05),
	.w3(32'h3b76c52b),
	.w4(32'hbc42c238),
	.w5(32'hbc1a605a),
	.w6(32'h3c5fefb5),
	.w7(32'h3c33210a),
	.w8(32'hbb95346c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6a5df),
	.w1(32'h3ad40599),
	.w2(32'h3beeec20),
	.w3(32'h3b845ca4),
	.w4(32'h3b14b5c2),
	.w5(32'h3ba87865),
	.w6(32'h3b067a27),
	.w7(32'hbb8a646a),
	.w8(32'h3c50b574),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad37c23),
	.w1(32'hbc0b0ca6),
	.w2(32'hba889df1),
	.w3(32'hb9e4c525),
	.w4(32'hbc347bda),
	.w5(32'hbb6f3113),
	.w6(32'hbb96dba9),
	.w7(32'hbbdb92fd),
	.w8(32'hbb5db5b1),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8778ff),
	.w1(32'hbb1a9301),
	.w2(32'h36807044),
	.w3(32'hbb0bfaa4),
	.w4(32'hbb2acdd4),
	.w5(32'hbc4f1745),
	.w6(32'hbbab3296),
	.w7(32'hbb8e16bd),
	.w8(32'hba3b2435),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb3502),
	.w1(32'hbb899cfd),
	.w2(32'hbb2cf2e7),
	.w3(32'hbc348856),
	.w4(32'h3bc4d0a9),
	.w5(32'hbb9aba62),
	.w6(32'h3bbdf534),
	.w7(32'h3c45cb54),
	.w8(32'hbbd6a458),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a885cf6),
	.w1(32'h3bf350f7),
	.w2(32'h3b3550d5),
	.w3(32'hbb3191da),
	.w4(32'h3bc7bdb4),
	.w5(32'h3ad30b14),
	.w6(32'hbc0331ae),
	.w7(32'hba62a039),
	.w8(32'h3aed92da),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb852916),
	.w1(32'hbb8de195),
	.w2(32'h3b7d3f8e),
	.w3(32'hbb3f017e),
	.w4(32'hbaa02f06),
	.w5(32'h3a2c522e),
	.w6(32'hbb19d2a1),
	.w7(32'hbac2348c),
	.w8(32'hb9a63991),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3435e0),
	.w1(32'hb9e54119),
	.w2(32'hbbc39506),
	.w3(32'hbae0dd04),
	.w4(32'hbc1712c8),
	.w5(32'hbc01f7f6),
	.w6(32'hbbf1b9aa),
	.w7(32'hbc22b9a3),
	.w8(32'hbc25eeb4),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be18450),
	.w1(32'h3c61cc30),
	.w2(32'hbb1e1a8d),
	.w3(32'hbb64b980),
	.w4(32'h3c8fcf70),
	.w5(32'hbabb23fa),
	.w6(32'hbc108f5f),
	.w7(32'h3baecfb2),
	.w8(32'hba97f5a4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb994c23),
	.w1(32'hbb68cc79),
	.w2(32'hbac664aa),
	.w3(32'hbb7563f2),
	.w4(32'hbb012247),
	.w5(32'hbb281085),
	.w6(32'hbb7e5c22),
	.w7(32'hbb362af6),
	.w8(32'hbbe9596e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba77012),
	.w1(32'hbab1bab3),
	.w2(32'h3bc809f0),
	.w3(32'hbb17c5fa),
	.w4(32'hbb86cd7e),
	.w5(32'h3bcf5c20),
	.w6(32'hbad236f6),
	.w7(32'h3aecd064),
	.w8(32'h3ba1f1d8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07722),
	.w1(32'h3be81533),
	.w2(32'hba02160c),
	.w3(32'h3ba8ece6),
	.w4(32'h3b36bf75),
	.w5(32'hb844e3e5),
	.w6(32'h3bbfb68c),
	.w7(32'h3b333310),
	.w8(32'h3bbe89c4),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95312c),
	.w1(32'hbc37ff43),
	.w2(32'hbc44059f),
	.w3(32'h3c3e6e56),
	.w4(32'hbaa97b2b),
	.w5(32'hbc82acd8),
	.w6(32'h3c5d4083),
	.w7(32'h3c3c3bf3),
	.w8(32'hbbfc04f5),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7974b),
	.w1(32'h3c74db53),
	.w2(32'h3b546877),
	.w3(32'hbbd6e277),
	.w4(32'h3c7a405b),
	.w5(32'h3b4105b3),
	.w6(32'hbc4073e2),
	.w7(32'hba507809),
	.w8(32'h3b3eae08),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54a2b9),
	.w1(32'hb939aafd),
	.w2(32'h3b7a2f61),
	.w3(32'h3b51bc92),
	.w4(32'h3b726309),
	.w5(32'h3b23ea77),
	.w6(32'h39f24922),
	.w7(32'h3b05b53a),
	.w8(32'h3babe674),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb8917),
	.w1(32'hba30da7d),
	.w2(32'hbc018754),
	.w3(32'h3bd705fa),
	.w4(32'hb971fce5),
	.w5(32'hbc401c07),
	.w6(32'h3c2260f9),
	.w7(32'h3bcd1ca3),
	.w8(32'hbc607adb),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f444c),
	.w1(32'h3c8f41e8),
	.w2(32'hbc275434),
	.w3(32'hbbbc3c60),
	.w4(32'h3d0071f4),
	.w5(32'hbc448639),
	.w6(32'hbb126bf4),
	.w7(32'h3ca894dc),
	.w8(32'hbc8f4e87),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbfd69),
	.w1(32'h3c8492a2),
	.w2(32'h3ad5ce84),
	.w3(32'hbbc9d2ed),
	.w4(32'h3cf398e5),
	.w5(32'h3b971526),
	.w6(32'h3be47c87),
	.w7(32'h3ce51045),
	.w8(32'h3b97693c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a867e73),
	.w1(32'hbbfe4fd3),
	.w2(32'hbb89e9ec),
	.w3(32'h3c16a977),
	.w4(32'hba14efe6),
	.w5(32'hba918e34),
	.w6(32'h3b4acdfe),
	.w7(32'h3c343081),
	.w8(32'hbab78b83),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05fd3e),
	.w1(32'hb81c7e11),
	.w2(32'hbb6b2e1c),
	.w3(32'h3b7918f4),
	.w4(32'h3b1f76e1),
	.w5(32'hbb84c748),
	.w6(32'h3b11ceb0),
	.w7(32'hb96a3977),
	.w8(32'hbb99bd3e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6595c),
	.w1(32'hbb287ed8),
	.w2(32'hba727710),
	.w3(32'hbbf91f62),
	.w4(32'hbb845c7d),
	.w5(32'h3a18c9a1),
	.w6(32'hbc20f3c9),
	.w7(32'hbbdbefda),
	.w8(32'hb8177f29),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39078691),
	.w1(32'h39c973cd),
	.w2(32'hbc2cad43),
	.w3(32'h3a327a0a),
	.w4(32'h3acc87ff),
	.w5(32'hb7dec77c),
	.w6(32'h3afd028f),
	.w7(32'h3b7a3689),
	.w8(32'h3c0e6729),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc538ffa),
	.w1(32'hbb774d5c),
	.w2(32'hbaeb055f),
	.w3(32'hbb9b49eb),
	.w4(32'hbc82d07b),
	.w5(32'hbb1471b3),
	.w6(32'hbb98ecc3),
	.w7(32'hbc5bc839),
	.w8(32'h3b556373),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c040756),
	.w1(32'h3bce8bb8),
	.w2(32'hbaee98e8),
	.w3(32'h3bdde59a),
	.w4(32'h3c5c6ebe),
	.w5(32'hbc04ff99),
	.w6(32'hbb677793),
	.w7(32'h3c03cbe7),
	.w8(32'hbba129a1),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00d504),
	.w1(32'hbc85338f),
	.w2(32'h3baf1291),
	.w3(32'h3bfc5f57),
	.w4(32'hbb92693a),
	.w5(32'h3b66bf46),
	.w6(32'h3af24fca),
	.w7(32'h3b99cbcf),
	.w8(32'hbb75ed85),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef6da8),
	.w1(32'h3c048918),
	.w2(32'hbbd3bdae),
	.w3(32'h3bfde584),
	.w4(32'h3badc1f6),
	.w5(32'hbc05b1fe),
	.w6(32'h3ad151e9),
	.w7(32'h3a7a4b80),
	.w8(32'hbbe625d4),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba801f90),
	.w1(32'h3b175769),
	.w2(32'h3b3041fa),
	.w3(32'hbb748b43),
	.w4(32'h3b4cf679),
	.w5(32'h3b9f7577),
	.w6(32'hbc18bd1a),
	.w7(32'h3b99154d),
	.w8(32'h3b7609ef),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86f7f0),
	.w1(32'h3b5a1b47),
	.w2(32'hbae5ec7c),
	.w3(32'h3b9e2e47),
	.w4(32'h3b58de13),
	.w5(32'h3ad169a8),
	.w6(32'h3a23c133),
	.w7(32'h3b01a6ab),
	.w8(32'hbc1597b7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5ba1b),
	.w1(32'h3cb62c5b),
	.w2(32'h3c3d8360),
	.w3(32'h3a879a28),
	.w4(32'h3c47b4f8),
	.w5(32'h3a02a89e),
	.w6(32'hbc5f0a39),
	.w7(32'hbc0d5d77),
	.w8(32'hbc216b98),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbc864),
	.w1(32'h3c5d71b8),
	.w2(32'h3c1691b7),
	.w3(32'h3bb76d41),
	.w4(32'h3c1f857d),
	.w5(32'h3c39cde0),
	.w6(32'hbc4e8914),
	.w7(32'h38b4c003),
	.w8(32'h3c0b900a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9561d),
	.w1(32'hbac61736),
	.w2(32'h3b8c617f),
	.w3(32'hbb9fc29e),
	.w4(32'h3b33980a),
	.w5(32'h3c59b40b),
	.w6(32'hbbe9f541),
	.w7(32'hbb7ff481),
	.w8(32'h3c413514),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb911d),
	.w1(32'h3b04cd1b),
	.w2(32'h3af7fd06),
	.w3(32'hbb2525b4),
	.w4(32'hbb81601c),
	.w5(32'h3b43e006),
	.w6(32'h3b2b34ec),
	.w7(32'hba9cb9ab),
	.w8(32'hbb8207e1),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7f47c),
	.w1(32'hbb894e94),
	.w2(32'hbb0cd5b8),
	.w3(32'h3b292ceb),
	.w4(32'hba844efb),
	.w5(32'hbaba157d),
	.w6(32'hb5f80c59),
	.w7(32'hbb1c864d),
	.w8(32'h3af9ea02),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb571d2f),
	.w1(32'hbb32f498),
	.w2(32'hbbb01a92),
	.w3(32'hba2c09d9),
	.w4(32'hbacc67ff),
	.w5(32'hbbe640ea),
	.w6(32'h3acc04ed),
	.w7(32'h3adbfb88),
	.w8(32'hbc33b980),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b162fed),
	.w1(32'h3cac2986),
	.w2(32'hbc45742a),
	.w3(32'h3aa8177c),
	.w4(32'h3c868f51),
	.w5(32'hbc64e9a4),
	.w6(32'hbc0f3e22),
	.w7(32'h3b972084),
	.w8(32'hba97d052),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8637f6),
	.w1(32'h3bba3406),
	.w2(32'h3a9b1d78),
	.w3(32'hb9b3bc82),
	.w4(32'hbba58590),
	.w5(32'h3b1170d7),
	.w6(32'hbb7ecb9a),
	.w7(32'hba656de7),
	.w8(32'h3b3bafb2),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bfa8d),
	.w1(32'hb9d324b5),
	.w2(32'h3b9137fe),
	.w3(32'h3adf4b2b),
	.w4(32'hba9312db),
	.w5(32'h3afa44f7),
	.w6(32'hb9919661),
	.w7(32'hba4c6b8b),
	.w8(32'h3c0bf203),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb695ab0),
	.w1(32'hbc979646),
	.w2(32'h3af48361),
	.w3(32'hb94cafd9),
	.w4(32'hbc4b90e5),
	.w5(32'h3a8e0024),
	.w6(32'hbbad8b5f),
	.w7(32'hbc0a1776),
	.w8(32'hbbffc27e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3dd2e),
	.w1(32'h3c3e99db),
	.w2(32'h3bba4468),
	.w3(32'h3b8d203d),
	.w4(32'h3c61c6fc),
	.w5(32'h3b7a4aef),
	.w6(32'hbc6240fd),
	.w7(32'h3bae4b9e),
	.w8(32'h3c097df7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd134),
	.w1(32'hbb9dade5),
	.w2(32'h3c290ed8),
	.w3(32'hbb7ff7d4),
	.w4(32'hbbaab71e),
	.w5(32'h3c46055f),
	.w6(32'h3a463f1c),
	.w7(32'hbb1025da),
	.w8(32'h3b5465e6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a3886),
	.w1(32'hbc36efba),
	.w2(32'h3aab1746),
	.w3(32'h3b1a68ae),
	.w4(32'hbbf6d921),
	.w5(32'hbbf09dcc),
	.w6(32'h3c95363b),
	.w7(32'hb88f875e),
	.w8(32'hba34e458),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc056b5),
	.w1(32'hbb640446),
	.w2(32'h3be88905),
	.w3(32'h3bd2d575),
	.w4(32'h3bf18ac3),
	.w5(32'h3a8ce7a3),
	.w6(32'h3c86f94b),
	.w7(32'h3c8b7584),
	.w8(32'hbc03d270),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca570a),
	.w1(32'h3c0e6a1c),
	.w2(32'h3bcc5ef7),
	.w3(32'h3b1d27b3),
	.w4(32'h3bca898e),
	.w5(32'h3bf839f6),
	.w6(32'hbc046959),
	.w7(32'hbb37c877),
	.w8(32'h39e54c99),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba813289),
	.w1(32'h3b270410),
	.w2(32'h3c02941c),
	.w3(32'h3bb614a9),
	.w4(32'h3bf17e85),
	.w5(32'h3c2444b7),
	.w6(32'hba885702),
	.w7(32'h3b7455c3),
	.w8(32'h3c0dea1d),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b746b),
	.w1(32'h3bad7e77),
	.w2(32'hbaf8093d),
	.w3(32'h3be47d23),
	.w4(32'h3bddd1e6),
	.w5(32'hbb1cb087),
	.w6(32'h3bab7865),
	.w7(32'h3c1d1012),
	.w8(32'hbb6584ec),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a1f0e),
	.w1(32'h3b87569b),
	.w2(32'h3a108cbb),
	.w3(32'h3b22d648),
	.w4(32'h3b61a5ab),
	.w5(32'h39d65af2),
	.w6(32'hbb33fc2b),
	.w7(32'hb92d8092),
	.w8(32'hbbaef21f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b294f4f),
	.w1(32'h3ae21341),
	.w2(32'hb66a1bdb),
	.w3(32'h3b3fd0fc),
	.w4(32'h3b0274a3),
	.w5(32'hbb216875),
	.w6(32'hbb2fbced),
	.w7(32'h3a62f297),
	.w8(32'h3b01a5f3),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4c022),
	.w1(32'hbb981f0f),
	.w2(32'hbbd61b55),
	.w3(32'hbbbb22a5),
	.w4(32'hbc21027d),
	.w5(32'hb85d9d1c),
	.w6(32'hbb9593d8),
	.w7(32'h3ad2a4c9),
	.w8(32'hbb2037a4),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96d7f1),
	.w1(32'hbbb5b7b2),
	.w2(32'h3c228771),
	.w3(32'h3b9c7085),
	.w4(32'hbc2f642e),
	.w5(32'hbb7e93e2),
	.w6(32'h3bea78ca),
	.w7(32'h3be81dc2),
	.w8(32'h3bbaae8b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b454012),
	.w1(32'hbc1728ff),
	.w2(32'h3c37c0c9),
	.w3(32'h3b7ee1a9),
	.w4(32'h3af5e349),
	.w5(32'h3c255967),
	.w6(32'h3b3aeabb),
	.w7(32'hbabcab22),
	.w8(32'h3c28ea31),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb989c3b),
	.w1(32'hbc20bcca),
	.w2(32'hba864337),
	.w3(32'hbaa21576),
	.w4(32'hbc8506f8),
	.w5(32'h3b3e7ead),
	.w6(32'hbc2db220),
	.w7(32'hbcb01914),
	.w8(32'h3bb277ae),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b496b),
	.w1(32'hbaeb297f),
	.w2(32'h3b96325a),
	.w3(32'h3ae3292c),
	.w4(32'h3a0813bb),
	.w5(32'h3bda0541),
	.w6(32'h3bce1f84),
	.w7(32'h3b8de958),
	.w8(32'h3b12e79c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6e082),
	.w1(32'hbba509b2),
	.w2(32'h3c1ba859),
	.w3(32'hbb2b90ee),
	.w4(32'hbbc6ccd0),
	.w5(32'h3c6380f3),
	.w6(32'hbc572fe1),
	.w7(32'hbca68bee),
	.w8(32'h3bf4243e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad72b8a),
	.w1(32'hbb75f4ba),
	.w2(32'h3b94136d),
	.w3(32'h3b72ae0c),
	.w4(32'hbc5b3642),
	.w5(32'h3bd0d817),
	.w6(32'hbb8171e4),
	.w7(32'hbc59b3ac),
	.w8(32'hbb75efc8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b446402),
	.w1(32'h3b0bfcb3),
	.w2(32'hba6ac519),
	.w3(32'h3b9d87f4),
	.w4(32'h3c074375),
	.w5(32'hba97de20),
	.w6(32'hba7b9cee),
	.w7(32'h3baea06f),
	.w8(32'hba4b7bc4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10af7a),
	.w1(32'h3b4d77b2),
	.w2(32'hbba7e3e6),
	.w3(32'hbb74cbe2),
	.w4(32'hbb9e7e2d),
	.w5(32'hbb9abdc8),
	.w6(32'hbadd6d9f),
	.w7(32'hbac3aa6d),
	.w8(32'h3ae72206),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d9c3c),
	.w1(32'h39301185),
	.w2(32'hbb1e7288),
	.w3(32'hbc4639ac),
	.w4(32'hbb952b6f),
	.w5(32'hba2ac427),
	.w6(32'hbc19913b),
	.w7(32'hbbd77ff3),
	.w8(32'hbb9577c1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcaf34),
	.w1(32'h3ac89508),
	.w2(32'hbab9463f),
	.w3(32'hb726240e),
	.w4(32'hbb3ebd17),
	.w5(32'hbc38ebcf),
	.w6(32'hbb099cf7),
	.w7(32'hbb32f9ea),
	.w8(32'hbb12cab0),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a3b3b),
	.w1(32'h3bdc3c1d),
	.w2(32'h3bb6f267),
	.w3(32'hbb67346d),
	.w4(32'h3c8012b0),
	.w5(32'h3adb02f9),
	.w6(32'h3bb5eb87),
	.w7(32'h3c1dbe91),
	.w8(32'h3bc066b3),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22430d),
	.w1(32'hbbb2b980),
	.w2(32'h3bef05fe),
	.w3(32'h3ba341a7),
	.w4(32'hbb8692d2),
	.w5(32'h3c3ac4f8),
	.w6(32'h3c7bba6a),
	.w7(32'h3c2e14c3),
	.w8(32'h3bb128d0),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b9038),
	.w1(32'hbac5e4d9),
	.w2(32'hb92ad4e3),
	.w3(32'h3bb00867),
	.w4(32'hbc20ec1e),
	.w5(32'hbb1d8992),
	.w6(32'h3a4746dc),
	.w7(32'hbc31d8bf),
	.w8(32'hbb8c35e6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ac494),
	.w1(32'h3b15b7f0),
	.w2(32'h3b05ec01),
	.w3(32'h38accd3b),
	.w4(32'hba99701a),
	.w5(32'hba29109c),
	.w6(32'hbb825c11),
	.w7(32'hbbac11f9),
	.w8(32'hbad407c5),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fc355),
	.w1(32'h3bc0a389),
	.w2(32'h3a81999c),
	.w3(32'h372bf344),
	.w4(32'hb9302bbc),
	.w5(32'hb99934b7),
	.w6(32'hbb79b365),
	.w7(32'hba7f6fe8),
	.w8(32'hbbb73c27),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa6887),
	.w1(32'hbb1904a4),
	.w2(32'h3b10ac0e),
	.w3(32'h3a2a7d54),
	.w4(32'h3a0fe979),
	.w5(32'h3b14e57d),
	.w6(32'hbc1932b3),
	.w7(32'h37b049e9),
	.w8(32'h3b185514),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9151b05),
	.w1(32'hbb6547da),
	.w2(32'h38f54f33),
	.w3(32'h393dcf2d),
	.w4(32'hbb9f21bb),
	.w5(32'h3ba3ef81),
	.w6(32'hba29c022),
	.w7(32'hb92fb2b9),
	.w8(32'h3b9a4702),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae577e9),
	.w1(32'h3bfdfcb3),
	.w2(32'h3b3e1399),
	.w3(32'h3b83f56f),
	.w4(32'hba253e5a),
	.w5(32'h3b441ba2),
	.w6(32'h3c0110f0),
	.w7(32'hbb9a2f70),
	.w8(32'hba84c8b8),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0390bd),
	.w1(32'hbaf93b54),
	.w2(32'hbadf46d5),
	.w3(32'h3bd8062a),
	.w4(32'hbbdef4c5),
	.w5(32'hba0419dd),
	.w6(32'h3bb6bddc),
	.w7(32'h3b21ca11),
	.w8(32'h3b18f305),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba27aa7),
	.w1(32'hbb8f812c),
	.w2(32'h3bd3f4a5),
	.w3(32'hba5e73ed),
	.w4(32'hbb1832a0),
	.w5(32'h3b614986),
	.w6(32'h3a07695b),
	.w7(32'h3b0ff40a),
	.w8(32'hbb3daabf),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule