module layer_10_featuremap_280(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a492f),
	.w1(32'h3a723366),
	.w2(32'h39933ca4),
	.w3(32'h3a94b258),
	.w4(32'h3a6ed1ce),
	.w5(32'h39295267),
	.w6(32'h3a8826ba),
	.w7(32'h39d7b9a0),
	.w8(32'h39f7979b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a467269),
	.w1(32'h3a32e13d),
	.w2(32'h39b6c103),
	.w3(32'hb9942980),
	.w4(32'h38ddea08),
	.w5(32'hba49400a),
	.w6(32'h395ee9d1),
	.w7(32'h394bc765),
	.w8(32'hba93ab4a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83c13e),
	.w1(32'h3a328b55),
	.w2(32'h3a914c0b),
	.w3(32'hb82023f3),
	.w4(32'h3985a317),
	.w5(32'h397884e4),
	.w6(32'h3aa13057),
	.w7(32'h3a6c5482),
	.w8(32'h39161724),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e64523),
	.w1(32'hba03f9ba),
	.w2(32'hb8daea7d),
	.w3(32'hb9993ccd),
	.w4(32'hb921d4ae),
	.w5(32'hb972a6d7),
	.w6(32'hb9d8b691),
	.w7(32'hb95fa31b),
	.w8(32'hba04c244),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab8679),
	.w1(32'hba624adb),
	.w2(32'hbacdd4e4),
	.w3(32'hb99f5607),
	.w4(32'hba19dbd7),
	.w5(32'h38689a00),
	.w6(32'hba2c7152),
	.w7(32'hbb106d89),
	.w8(32'h384c6591),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a25037),
	.w1(32'hb8297d4f),
	.w2(32'hba07e358),
	.w3(32'h39c9fba7),
	.w4(32'h38711cda),
	.w5(32'h39c8d918),
	.w6(32'h393b5de7),
	.w7(32'hb9c65098),
	.w8(32'h39b4cb70),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995ecbc),
	.w1(32'hb973a046),
	.w2(32'hb8e75a49),
	.w3(32'hb92073cc),
	.w4(32'h398831f3),
	.w5(32'h3a16af72),
	.w6(32'hb9c855eb),
	.w7(32'hb85d8071),
	.w8(32'hb9337bf6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91385b1),
	.w1(32'h38375cfe),
	.w2(32'h39172574),
	.w3(32'hb80bc238),
	.w4(32'h3979ab81),
	.w5(32'h3a524e0b),
	.w6(32'hb9b4d4e7),
	.w7(32'h3810b213),
	.w8(32'h39fe1f86),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8d219),
	.w1(32'hb8566d70),
	.w2(32'h39086b6a),
	.w3(32'h39ab3e5e),
	.w4(32'h39e001ed),
	.w5(32'hb8864e9d),
	.w6(32'hb90fcfad),
	.w7(32'hb904a433),
	.w8(32'h387d8b9d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a381fc),
	.w1(32'hba3176c7),
	.w2(32'hba6775ca),
	.w3(32'h36ed334b),
	.w4(32'hb9d3543e),
	.w5(32'h39d05828),
	.w6(32'h38da1a1f),
	.w7(32'hba074fe5),
	.w8(32'h3a7f5863),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01bc0a),
	.w1(32'hb88ee93e),
	.w2(32'hba4fcc12),
	.w3(32'h3a77f336),
	.w4(32'h391f855b),
	.w5(32'h3a50873d),
	.w6(32'h3a0c8309),
	.w7(32'hba4857fa),
	.w8(32'h3a0045fd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a111544),
	.w1(32'h3a251dba),
	.w2(32'h39aa30a2),
	.w3(32'h3a1d7c6c),
	.w4(32'h3a5c8166),
	.w5(32'hb9a0ee70),
	.w6(32'h3985ac7e),
	.w7(32'h39ba36df),
	.w8(32'hba360084),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a60af2),
	.w1(32'hb9c9e239),
	.w2(32'hb995d8f6),
	.w3(32'h3a32f575),
	.w4(32'h3a4f916e),
	.w5(32'hbaebedb6),
	.w6(32'hb7021f98),
	.w7(32'hb9a151e9),
	.w8(32'hba6400a6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3ac69),
	.w1(32'hbb8663dc),
	.w2(32'h3b00ed3a),
	.w3(32'hbb964d90),
	.w4(32'h3ae2c799),
	.w5(32'h39ae2734),
	.w6(32'hbb37a1e0),
	.w7(32'h3a87b9cb),
	.w8(32'h3978783f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388c7f95),
	.w1(32'hb9d9bb5e),
	.w2(32'hb85e3a0a),
	.w3(32'hb9b1a7d1),
	.w4(32'hb9a8bf5a),
	.w5(32'hb8ea5db5),
	.w6(32'hba2eb7e7),
	.w7(32'hb9ef8fae),
	.w8(32'hb968c2f5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d98518),
	.w1(32'h39040185),
	.w2(32'h3a06012c),
	.w3(32'hb84d0ff6),
	.w4(32'h39d7bd34),
	.w5(32'hb908027e),
	.w6(32'h39cb6ad6),
	.w7(32'h391256b5),
	.w8(32'hb8ae0b78),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39873fc8),
	.w1(32'h3a08a837),
	.w2(32'h388db534),
	.w3(32'h39758b00),
	.w4(32'h3a0afcdb),
	.w5(32'h38e8a8be),
	.w6(32'h38eb8768),
	.w7(32'hb8fbaf13),
	.w8(32'h38f2fd03),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92500be),
	.w1(32'hb95ad20a),
	.w2(32'hb9a8be5b),
	.w3(32'h39c33433),
	.w4(32'h3916b5c5),
	.w5(32'hba20f976),
	.w6(32'h382ed9b2),
	.w7(32'h395155e8),
	.w8(32'hba44d146),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80d9ac),
	.w1(32'hba598a09),
	.w2(32'hba9c0496),
	.w3(32'h37cbbaa1),
	.w4(32'hb9e154a9),
	.w5(32'hb9c13e6c),
	.w6(32'hba1789e0),
	.w7(32'hba40f1d4),
	.w8(32'hba2a82a4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba569095),
	.w1(32'hba7d3efd),
	.w2(32'h393c028d),
	.w3(32'hba90d1f4),
	.w4(32'hb8da3f75),
	.w5(32'hba018b0e),
	.w6(32'hb903448c),
	.w7(32'hb95b9bbb),
	.w8(32'hba62b53f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f3584),
	.w1(32'h38bbb7dd),
	.w2(32'h396a64d9),
	.w3(32'h3a16ec61),
	.w4(32'h39e245ab),
	.w5(32'h39ebd83d),
	.w6(32'h3992b642),
	.w7(32'h37446333),
	.w8(32'h39a57c24),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b8ebe),
	.w1(32'h39e8bc74),
	.w2(32'h3a700aaa),
	.w3(32'h3973e946),
	.w4(32'h39b5b602),
	.w5(32'hbadf71ea),
	.w6(32'h380b2114),
	.w7(32'h39ab796c),
	.w8(32'hbaa0a8f2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae82daa),
	.w1(32'h3b3bb7a5),
	.w2(32'h3b9d4cf5),
	.w3(32'h3946808e),
	.w4(32'h3abf73fa),
	.w5(32'hb986c503),
	.w6(32'hb999977a),
	.w7(32'h3b8005ca),
	.w8(32'hb9b0d83f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a2fcc),
	.w1(32'hba08ac8b),
	.w2(32'hb923ae4f),
	.w3(32'h38cd09c4),
	.w4(32'h3967049d),
	.w5(32'h3a3482b2),
	.w6(32'h36ad3f16),
	.w7(32'hb8e099ee),
	.w8(32'h3a0fd94a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37802d5d),
	.w1(32'h388889a3),
	.w2(32'hba18352a),
	.w3(32'hb986f1d0),
	.w4(32'h38f4f369),
	.w5(32'h3a5ed998),
	.w6(32'hb7d89974),
	.w7(32'hba1867f2),
	.w8(32'h38e7e062),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a013a8b),
	.w1(32'hb7e72d4e),
	.w2(32'hb9b7cbd4),
	.w3(32'h395dd3cf),
	.w4(32'hb93fd25a),
	.w5(32'hb8f12470),
	.w6(32'h390797d7),
	.w7(32'hb70b38f8),
	.w8(32'h37ac3ec3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dbb464),
	.w1(32'h390af419),
	.w2(32'h3a11d4f5),
	.w3(32'h39113068),
	.w4(32'h39e94b54),
	.w5(32'h3966a948),
	.w6(32'hb7a6956f),
	.w7(32'h3a346bae),
	.w8(32'hb803d9a1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0b1d1),
	.w1(32'h3a388f14),
	.w2(32'h39e9b5f6),
	.w3(32'h3a919aff),
	.w4(32'h3ab5161f),
	.w5(32'h39a38cbf),
	.w6(32'h3a342f96),
	.w7(32'h3a090110),
	.w8(32'hb9a111c7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac356ac),
	.w1(32'hbb9845cc),
	.w2(32'hbb8efc60),
	.w3(32'hbb4bfbe3),
	.w4(32'hbb3cbdf2),
	.w5(32'hb8b95d1e),
	.w6(32'hbb4c3aa6),
	.w7(32'hbb94ab02),
	.w8(32'h3995a6cd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e05c71),
	.w1(32'hba538a84),
	.w2(32'hb9ccb73a),
	.w3(32'hb993ed3c),
	.w4(32'hb9a01864),
	.w5(32'h3a82e97c),
	.w6(32'hb7c9ff1e),
	.w7(32'h38c83225),
	.w8(32'h3a594330),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ec5c7),
	.w1(32'h3a99c0ed),
	.w2(32'h3ab78471),
	.w3(32'h3ac1f698),
	.w4(32'h3983615f),
	.w5(32'hb9570d04),
	.w6(32'h39f02430),
	.w7(32'h3a0ca453),
	.w8(32'h39a89368),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d9c0d),
	.w1(32'hb9c6feb5),
	.w2(32'hba797446),
	.w3(32'h39e2adb1),
	.w4(32'h39c9bd76),
	.w5(32'h3aade3a6),
	.w6(32'h38d36688),
	.w7(32'hb9ec84eb),
	.w8(32'h3abf3c0f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a898397),
	.w1(32'hba0bae4a),
	.w2(32'hba232ec5),
	.w3(32'h38c6e21b),
	.w4(32'hb41c22ce),
	.w5(32'h3a0bb873),
	.w6(32'hb996e0f0),
	.w7(32'hba0d4d2d),
	.w8(32'h39e3f0a9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bedaea),
	.w1(32'h38f5efcf),
	.w2(32'hb9bc2168),
	.w3(32'h3a00022b),
	.w4(32'hb87af0ec),
	.w5(32'hba9452e2),
	.w6(32'h398e822c),
	.w7(32'hb9924908),
	.w8(32'hb980ae4c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9763576),
	.w1(32'hb9bd5cc3),
	.w2(32'hba115105),
	.w3(32'h3ab84dfa),
	.w4(32'h3ab08003),
	.w5(32'hb99c2b93),
	.w6(32'hb8e040a3),
	.w7(32'h3a2eb29c),
	.w8(32'hba1ff9f3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26675f),
	.w1(32'hba071ebb),
	.w2(32'hb9991205),
	.w3(32'h36924b68),
	.w4(32'hba25d826),
	.w5(32'hb9af216d),
	.w6(32'hb9b1c172),
	.w7(32'hb9b932f8),
	.w8(32'hb9a6e5d1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7723d3),
	.w1(32'h39b1f2ec),
	.w2(32'hb8f848fd),
	.w3(32'h3a43d6e9),
	.w4(32'h3a5326df),
	.w5(32'hb989098d),
	.w6(32'h39ce9e8b),
	.w7(32'h3a58cb73),
	.w8(32'h38a17769),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b44a3f),
	.w1(32'h3942eb60),
	.w2(32'hbaa63aa7),
	.w3(32'h39ad8360),
	.w4(32'hba1f3f02),
	.w5(32'hba78db3b),
	.w6(32'h38fb6ac0),
	.w7(32'hba07f9e8),
	.w8(32'hb9f49cc1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd5fe1),
	.w1(32'hb908ac57),
	.w2(32'hb99b981f),
	.w3(32'h38214fbc),
	.w4(32'h38e0b457),
	.w5(32'hba3c7a96),
	.w6(32'hb951b48f),
	.w7(32'h38c8a314),
	.w8(32'hb9a79519),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b5f3b),
	.w1(32'h39f94215),
	.w2(32'h3a2a7749),
	.w3(32'h39d62523),
	.w4(32'h3a485da3),
	.w5(32'h3ab9e3e8),
	.w6(32'h39c92da8),
	.w7(32'h39ba891d),
	.w8(32'h3adfe960),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe3f97),
	.w1(32'h3a8a9c0a),
	.w2(32'h3a1f0029),
	.w3(32'h3a7f5a74),
	.w4(32'h39f97941),
	.w5(32'hb7c07f59),
	.w6(32'h3ad6ea2c),
	.w7(32'h39f14976),
	.w8(32'hba067887),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4636f),
	.w1(32'hba681bca),
	.w2(32'hba7cd760),
	.w3(32'hba1c46dd),
	.w4(32'hba127ad2),
	.w5(32'hba1ded2d),
	.w6(32'hba3797ae),
	.w7(32'hba0e2d82),
	.w8(32'hb90b9575),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ae138),
	.w1(32'hba124566),
	.w2(32'hbabeba15),
	.w3(32'hb9e2d54c),
	.w4(32'hba863120),
	.w5(32'h39848104),
	.w6(32'h3894bed2),
	.w7(32'hba74e3a6),
	.w8(32'h3a60c64f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c1731),
	.w1(32'h3955f1c7),
	.w2(32'h39975b09),
	.w3(32'h3aaa638d),
	.w4(32'h3a8b4fbc),
	.w5(32'h3a77df45),
	.w6(32'h3ac4c865),
	.w7(32'h39ad352c),
	.w8(32'h380373d0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3861fe0b),
	.w1(32'hba80aadd),
	.w2(32'hba44d13b),
	.w3(32'hb987c55f),
	.w4(32'hb9e4f383),
	.w5(32'h3852d99b),
	.w6(32'hba966ab7),
	.w7(32'hb9de76f2),
	.w8(32'h38733a8e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e500c1),
	.w1(32'h39897e30),
	.w2(32'h3a8a8cd0),
	.w3(32'h3a6690ad),
	.w4(32'h3a8c64c0),
	.w5(32'hb9143cb5),
	.w6(32'h3a775f22),
	.w7(32'h3a18a3d9),
	.w8(32'hba0a1d9e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e802d7),
	.w1(32'hb9d398fd),
	.w2(32'hb9e52ba4),
	.w3(32'h38e37760),
	.w4(32'h37e70f7d),
	.w5(32'h3a93bcdf),
	.w6(32'h396f42d5),
	.w7(32'hb936f108),
	.w8(32'h3a8ceffc),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c4c19),
	.w1(32'h3995d83c),
	.w2(32'h3a01abcb),
	.w3(32'h39ec8715),
	.w4(32'h3a11c550),
	.w5(32'h395aae91),
	.w6(32'h39181ebe),
	.w7(32'h39244c19),
	.w8(32'hb99b7ce8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f53376),
	.w1(32'hb99f715e),
	.w2(32'hb9004154),
	.w3(32'h3a26a6d4),
	.w4(32'h39c9e6d1),
	.w5(32'h3a344b78),
	.w6(32'hb9ea8d28),
	.w7(32'hb97362df),
	.w8(32'h39f35771),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7fc57),
	.w1(32'h3a457bc2),
	.w2(32'h3a6ef2d0),
	.w3(32'h3a376184),
	.w4(32'h3a717b7f),
	.w5(32'hbb48c9a9),
	.w6(32'h3987da88),
	.w7(32'h3a3eedff),
	.w8(32'hbb860d60),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb096cae),
	.w1(32'hba216155),
	.w2(32'h3a6cffff),
	.w3(32'hbaf58455),
	.w4(32'h3a24f350),
	.w5(32'hba73a910),
	.w6(32'hb802d0e5),
	.w7(32'h3a5183ca),
	.w8(32'hba32fa01),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba927b93),
	.w1(32'hb9d53970),
	.w2(32'hba27c27d),
	.w3(32'hba7cac95),
	.w4(32'hba5624f4),
	.w5(32'h3a45873a),
	.w6(32'hb9cc2ff2),
	.w7(32'hb9ffe031),
	.w8(32'hba8165d5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2509f),
	.w1(32'hbb895349),
	.w2(32'hbb83534a),
	.w3(32'hbb661a1b),
	.w4(32'hbb579bfa),
	.w5(32'h3a8c3c13),
	.w6(32'hbb4a1847),
	.w7(32'hbba4031a),
	.w8(32'h3a7e2823),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a814b29),
	.w1(32'h3a404473),
	.w2(32'h3a7c854e),
	.w3(32'h39eecc6b),
	.w4(32'h3a640fcc),
	.w5(32'h39eb6bc3),
	.w6(32'h39648600),
	.w7(32'h3a9cc734),
	.w8(32'h3a2c2806),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79a309),
	.w1(32'h3a6e668c),
	.w2(32'hba40043d),
	.w3(32'h3a75bc70),
	.w4(32'hb92e543b),
	.w5(32'h3750b159),
	.w6(32'h3a91aaf0),
	.w7(32'hb9898f79),
	.w8(32'h3a18be8e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8ca62),
	.w1(32'h3aa1a6a5),
	.w2(32'h389951a9),
	.w3(32'h3a918f5a),
	.w4(32'h396445a2),
	.w5(32'h396de4ff),
	.w6(32'h3aa081b2),
	.w7(32'hb7cbd49e),
	.w8(32'h396955be),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa25dc),
	.w1(32'h3a4c9908),
	.w2(32'h399e976d),
	.w3(32'h3a406bbc),
	.w4(32'hb824f25e),
	.w5(32'hb95617c5),
	.w6(32'h3a0e3d8e),
	.w7(32'h399d43eb),
	.w8(32'h39a26754),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3955208b),
	.w1(32'hb9ff8340),
	.w2(32'hba1f381e),
	.w3(32'hba026bca),
	.w4(32'h39860ab2),
	.w5(32'h3a302ccc),
	.w6(32'h39912687),
	.w7(32'hb9f34937),
	.w8(32'h39d67134),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b93346),
	.w1(32'h38d47054),
	.w2(32'h392000d0),
	.w3(32'h39bbad80),
	.w4(32'h39be0396),
	.w5(32'hbaaeae38),
	.w6(32'hb98b1753),
	.w7(32'h37ffc296),
	.w8(32'hbada9302),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa3165),
	.w1(32'hba362f34),
	.w2(32'hb9117d5a),
	.w3(32'hba76e11b),
	.w4(32'hba33eda2),
	.w5(32'hb8f220ed),
	.w6(32'hb8bc1c13),
	.w7(32'hba072b00),
	.w8(32'h3752d7e3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3863cfe9),
	.w1(32'hb7e5bf48),
	.w2(32'hb7061198),
	.w3(32'h39149a36),
	.w4(32'h39cabc5b),
	.w5(32'h3a413376),
	.w6(32'h37bca029),
	.w7(32'h39d58995),
	.w8(32'h3a06754c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11ac02),
	.w1(32'h3a2e9cfc),
	.w2(32'h3a04d8f6),
	.w3(32'h39c10916),
	.w4(32'h3a05597f),
	.w5(32'hbb2f5cc7),
	.w6(32'h3a27d62c),
	.w7(32'h3a38c464),
	.w8(32'hbb4408de),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc45c3),
	.w1(32'hbaa0cc5e),
	.w2(32'hbaf87dba),
	.w3(32'hb9c74ebb),
	.w4(32'h3a3d3aa9),
	.w5(32'hb9b2c82b),
	.w6(32'hbab4a2cd),
	.w7(32'hba9f7c20),
	.w8(32'hb8a0de19),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f4f16c),
	.w1(32'hb9af0dd0),
	.w2(32'hb9f5c2d0),
	.w3(32'h38a43998),
	.w4(32'hba40e67e),
	.w5(32'h3b28a9cb),
	.w6(32'hba518f0a),
	.w7(32'h38a4c6c8),
	.w8(32'h3b3d7e54),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b236305),
	.w1(32'h3b503131),
	.w2(32'hba8152d9),
	.w3(32'h3bb01200),
	.w4(32'h3a163256),
	.w5(32'hb8cbd43d),
	.w6(32'h3b760681),
	.w7(32'h39ac9c67),
	.w8(32'h382c576e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39feface),
	.w1(32'hba9f443c),
	.w2(32'hbb15e5dd),
	.w3(32'h397bc52a),
	.w4(32'hb9b254f3),
	.w5(32'h391d933d),
	.w6(32'hb9e45807),
	.w7(32'hbace53a2),
	.w8(32'hb9fa75a9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4c3e9),
	.w1(32'hb99ded2b),
	.w2(32'h3923e9f2),
	.w3(32'hb888e04f),
	.w4(32'h39cd5616),
	.w5(32'hba04163d),
	.w6(32'hb9901042),
	.w7(32'hb81a122a),
	.w8(32'hba7451eb),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba835ef0),
	.w1(32'hbac3f94c),
	.w2(32'hb9b7a2b7),
	.w3(32'hbaf6393a),
	.w4(32'hbb0c6bec),
	.w5(32'h3b85f584),
	.w6(32'hbb27be02),
	.w7(32'hbb0735fa),
	.w8(32'h3ba39206),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c78a6),
	.w1(32'h3b8416d0),
	.w2(32'hbb0b5dd1),
	.w3(32'h3baaa6b5),
	.w4(32'hb9975be6),
	.w5(32'h3a320f59),
	.w6(32'h3b9bf316),
	.w7(32'hba97419c),
	.w8(32'h3983e537),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eada51),
	.w1(32'h3a5f9658),
	.w2(32'h3903e822),
	.w3(32'h3a9274ef),
	.w4(32'h39e32420),
	.w5(32'h39e51436),
	.w6(32'h39d45754),
	.w7(32'h38e3e9fc),
	.w8(32'h3a3c56c4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ce588),
	.w1(32'h39b6c833),
	.w2(32'hb8e7d29b),
	.w3(32'h39aa87f3),
	.w4(32'hb90c64bf),
	.w5(32'hb90f6459),
	.w6(32'hb909cc02),
	.w7(32'hb97bc27d),
	.w8(32'hba2f3aaf),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0242fd),
	.w1(32'h38e33b12),
	.w2(32'h3a07fed1),
	.w3(32'h372668fa),
	.w4(32'h395b7cda),
	.w5(32'h3953ea7e),
	.w6(32'hb84abd19),
	.w7(32'h38f874fd),
	.w8(32'h379cf5a9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9048f7f),
	.w1(32'h392a3301),
	.w2(32'h39f7d08c),
	.w3(32'h388425ce),
	.w4(32'hb9dcfdc9),
	.w5(32'hba835d85),
	.w6(32'h39cc151a),
	.w7(32'h39ca69da),
	.w8(32'hb9a59377),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d262e),
	.w1(32'h397e7a84),
	.w2(32'hb589cb7c),
	.w3(32'hb9aff348),
	.w4(32'hb8281bf8),
	.w5(32'hb91ce71a),
	.w6(32'hb964a5c4),
	.w7(32'h38f7b2b8),
	.w8(32'hb98e2a38),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98abba3),
	.w1(32'hb9a69656),
	.w2(32'hb949f696),
	.w3(32'h3913d36e),
	.w4(32'h38f3bf52),
	.w5(32'h39919388),
	.w6(32'hb958ac4e),
	.w7(32'hb9cb241e),
	.w8(32'h39a7c55e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d6278),
	.w1(32'h38ebd9ee),
	.w2(32'hb98ddd70),
	.w3(32'h3a49e28d),
	.w4(32'hb75eb0d1),
	.w5(32'h39384ef7),
	.w6(32'h39d6fe86),
	.w7(32'hba26c184),
	.w8(32'h39fe7db8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f3873b),
	.w1(32'h3a910c29),
	.w2(32'h38fc0bd1),
	.w3(32'h3a51c43f),
	.w4(32'hba2cbfe7),
	.w5(32'h38eb6a66),
	.w6(32'h39fd74cb),
	.w7(32'h39898e09),
	.w8(32'h39890bd8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c314f6),
	.w1(32'h3996d61a),
	.w2(32'h39f3000a),
	.w3(32'h39b10fe1),
	.w4(32'h3913f6a4),
	.w5(32'h3938fd72),
	.w6(32'h39c7314a),
	.w7(32'h39b1c582),
	.w8(32'h38d0e771),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3042f1),
	.w1(32'h38fe2b67),
	.w2(32'hb978b9b2),
	.w3(32'h39a20b6a),
	.w4(32'h3916e9bf),
	.w5(32'h3874c55d),
	.w6(32'h388aa56a),
	.w7(32'hb9d8dcf1),
	.w8(32'hb9b8a0a6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9555030),
	.w1(32'hb761a6e3),
	.w2(32'h398029f8),
	.w3(32'h39c64cb9),
	.w4(32'h3a0c2550),
	.w5(32'h3a8f8891),
	.w6(32'hb9c04efe),
	.w7(32'hb99511e4),
	.w8(32'h3ad2f00a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fb316),
	.w1(32'h3a9106ce),
	.w2(32'h3a948337),
	.w3(32'h3a8b82cd),
	.w4(32'h39b67f15),
	.w5(32'h3a5fb0ab),
	.w6(32'h3a947deb),
	.w7(32'h3a36530c),
	.w8(32'hb7ab7bb5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4a5a3),
	.w1(32'h39c25553),
	.w2(32'h392641fd),
	.w3(32'h3a58503d),
	.w4(32'hb91a94d1),
	.w5(32'h3b4cfb00),
	.w6(32'h3847d8be),
	.w7(32'hb989cb3b),
	.w8(32'h3ba842ea),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90558b),
	.w1(32'h3bc99a01),
	.w2(32'h3a80b142),
	.w3(32'h3bce6434),
	.w4(32'h3b0a792a),
	.w5(32'h391b7bc1),
	.w6(32'h3bcc9b1e),
	.w7(32'h3b1d7a5f),
	.w8(32'h3a04997b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ecae1),
	.w1(32'hba5837ee),
	.w2(32'h38375347),
	.w3(32'hba81ac2b),
	.w4(32'hba9b9179),
	.w5(32'hb9bae0a7),
	.w6(32'hba530bbc),
	.w7(32'hba1cdbbc),
	.w8(32'h39b1b874),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecc97f),
	.w1(32'h3b2dd4bb),
	.w2(32'h3b374fb6),
	.w3(32'h39e3ef67),
	.w4(32'h374d6388),
	.w5(32'h3a81ffc1),
	.w6(32'h39f167c4),
	.w7(32'h3ade545d),
	.w8(32'h3a850981),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d8e19),
	.w1(32'h3a88dd70),
	.w2(32'hb9264b36),
	.w3(32'h3adfa248),
	.w4(32'h3a5d6834),
	.w5(32'h391503a0),
	.w6(32'h3abfbec0),
	.w7(32'h39ce063f),
	.w8(32'hb9b7fbb8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d3d81),
	.w1(32'h3a191d3f),
	.w2(32'h388bfd02),
	.w3(32'h379f615a),
	.w4(32'h3a6f9351),
	.w5(32'h3a5fa7e3),
	.w6(32'h3a3d898e),
	.w7(32'h3a80cbdf),
	.w8(32'hb9ca2678),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76ea21),
	.w1(32'hb9c79273),
	.w2(32'h38f6ac4a),
	.w3(32'hb8f0631b),
	.w4(32'hba77a3dd),
	.w5(32'h39f103b0),
	.w6(32'h3908f0b5),
	.w7(32'hb8260856),
	.w8(32'h39875578),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd1c25),
	.w1(32'hb9193a27),
	.w2(32'h39888eab),
	.w3(32'hb90ddcba),
	.w4(32'h3a03589b),
	.w5(32'h3a82354d),
	.w6(32'hb9f971b7),
	.w7(32'hb86fb631),
	.w8(32'h3a663c97),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f5092),
	.w1(32'hba2aa2f5),
	.w2(32'h39ff5bc4),
	.w3(32'hb8d91716),
	.w4(32'h398f0791),
	.w5(32'h39c80715),
	.w6(32'hb9af226c),
	.w7(32'h39fd97d3),
	.w8(32'h39ad9756),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b71989),
	.w1(32'hb95b80c4),
	.w2(32'hb994915b),
	.w3(32'h38ef41da),
	.w4(32'h3827812f),
	.w5(32'h3a1a6d22),
	.w6(32'hb93431dc),
	.w7(32'hb7c827f3),
	.w8(32'h3a831def),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fcfa0),
	.w1(32'hbad95186),
	.w2(32'hb8ca3429),
	.w3(32'hba87e42c),
	.w4(32'hba072318),
	.w5(32'h392d693b),
	.w6(32'hbab2fd50),
	.w7(32'hb9686717),
	.w8(32'h3a28692e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d358aa),
	.w1(32'hba57f925),
	.w2(32'hba0580f3),
	.w3(32'hb9b7aef0),
	.w4(32'h3a764cae),
	.w5(32'hbaecec0d),
	.w6(32'hba0499af),
	.w7(32'h3a022ef8),
	.w8(32'hbabb46e8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b7940),
	.w1(32'hba3cc67f),
	.w2(32'hb92ebe55),
	.w3(32'hba976ca9),
	.w4(32'hba4b59f5),
	.w5(32'h3943aa23),
	.w6(32'hb9a5e511),
	.w7(32'hba3c0cd3),
	.w8(32'h393975c4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86ac5d0),
	.w1(32'h37f7ec37),
	.w2(32'hb957ab68),
	.w3(32'h3999762c),
	.w4(32'h39341321),
	.w5(32'hb9a8a808),
	.w6(32'h393f004e),
	.w7(32'hb75224c1),
	.w8(32'hba1fb7fe),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8669fd),
	.w1(32'h37d0c65b),
	.w2(32'hb93ad305),
	.w3(32'h38547441),
	.w4(32'hb99a3568),
	.w5(32'hb9ef6e94),
	.w6(32'h398232ff),
	.w7(32'h393d574b),
	.w8(32'hb9926a98),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d00e6),
	.w1(32'hb7bed2ae),
	.w2(32'h3962a816),
	.w3(32'h383d668d),
	.w4(32'h39098de5),
	.w5(32'h38387473),
	.w6(32'h39a7c80b),
	.w7(32'h38bd8f82),
	.w8(32'h3a86c5f6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cd427),
	.w1(32'h3a9ad305),
	.w2(32'h3b0550e5),
	.w3(32'h3a5959a6),
	.w4(32'h3a1f689d),
	.w5(32'hbb912f07),
	.w6(32'h399c3faa),
	.w7(32'h3a7abd3d),
	.w8(32'hbb9c3385),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4693b9),
	.w1(32'hbbb51393),
	.w2(32'hbb51da36),
	.w3(32'hbba36698),
	.w4(32'hbbb5053e),
	.w5(32'hbc305276),
	.w6(32'hbba6ca83),
	.w7(32'hbb2fb98e),
	.w8(32'hbc3a4d95),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41bb59),
	.w1(32'hbc8888e9),
	.w2(32'hbc1152d3),
	.w3(32'hbbccfe4c),
	.w4(32'hbc7bec6e),
	.w5(32'h3b45085e),
	.w6(32'hba91c1cb),
	.w7(32'hbc864ad3),
	.w8(32'hbc0b5f99),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf9b77),
	.w1(32'hbbfe0750),
	.w2(32'hbb9492df),
	.w3(32'h3a7eb1d5),
	.w4(32'h3bbefb59),
	.w5(32'h3b521b41),
	.w6(32'hbb633104),
	.w7(32'h3b459ef1),
	.w8(32'hb95a83a2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0f08b),
	.w1(32'h3ba52686),
	.w2(32'h3a65f4a3),
	.w3(32'hba860c4f),
	.w4(32'h3b39551e),
	.w5(32'h3b003d9b),
	.w6(32'hbbcbbce7),
	.w7(32'hbbb05274),
	.w8(32'h3941a87d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe4bbb),
	.w1(32'hbb27e142),
	.w2(32'h3b440e85),
	.w3(32'hba83ecbe),
	.w4(32'h3b131cc3),
	.w5(32'hbb9e7464),
	.w6(32'hbc1285a4),
	.w7(32'hba8c0547),
	.w8(32'h3b2d07ff),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97e053),
	.w1(32'h3bbf80cc),
	.w2(32'h3b8460a2),
	.w3(32'hbaaf70f1),
	.w4(32'hbbb81a60),
	.w5(32'hbbd2b035),
	.w6(32'h3c106a99),
	.w7(32'h3bac9129),
	.w8(32'hbb67cf3f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0865a),
	.w1(32'h3b3e0549),
	.w2(32'hbb4c9349),
	.w3(32'hbb8fdfe1),
	.w4(32'h3bceb22b),
	.w5(32'hb73e2116),
	.w6(32'hbb50dc6c),
	.w7(32'hba5d1fa0),
	.w8(32'hbb5d3359),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9565e6),
	.w1(32'hbb921129),
	.w2(32'hba79d373),
	.w3(32'h3bb37089),
	.w4(32'h3b8825ee),
	.w5(32'hbc85aeb0),
	.w6(32'h3baa9b20),
	.w7(32'hbaf7823b),
	.w8(32'hbc7744e9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08ce3a),
	.w1(32'hbbfe1d6b),
	.w2(32'hbb01860b),
	.w3(32'hbbe4288f),
	.w4(32'hbc259039),
	.w5(32'h3b56d73b),
	.w6(32'hbc1c2ceb),
	.w7(32'hbc3a47d7),
	.w8(32'hbb00dfea),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7dd02a),
	.w1(32'h3baf4942),
	.w2(32'h3bb13499),
	.w3(32'h3a5003df),
	.w4(32'h3b8148f0),
	.w5(32'hbb81a652),
	.w6(32'h392ac3c5),
	.w7(32'hb9e18889),
	.w8(32'hbb85a584),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb734973),
	.w1(32'hbbf91f7a),
	.w2(32'hbbdc03cc),
	.w3(32'hbba938b2),
	.w4(32'hbbe91a7b),
	.w5(32'h3c555d79),
	.w6(32'hbb856816),
	.w7(32'hbbc85007),
	.w8(32'h3b5e1820),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53be02),
	.w1(32'h3adccb5c),
	.w2(32'h3ba19f9b),
	.w3(32'h3b7662f8),
	.w4(32'h3bf03caa),
	.w5(32'h3b581ea1),
	.w6(32'hbc5ca714),
	.w7(32'h39bdd3bb),
	.w8(32'hbbfaac93),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac3c00),
	.w1(32'hbb9e8b20),
	.w2(32'h3b2e0029),
	.w3(32'hbb28dc3e),
	.w4(32'hbc2ea495),
	.w5(32'hbaded99b),
	.w6(32'hbc1e840d),
	.w7(32'hbc427a81),
	.w8(32'hbae29a3e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8ac53),
	.w1(32'h3bd4dac6),
	.w2(32'h3b50e6aa),
	.w3(32'hb8c7053c),
	.w4(32'hbae16df2),
	.w5(32'h3c1563a6),
	.w6(32'hbbc82c63),
	.w7(32'h3b26e1f6),
	.w8(32'h3b7ff03f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6283e),
	.w1(32'hbbf1b487),
	.w2(32'hbb92b41b),
	.w3(32'h3b024186),
	.w4(32'hb999e8b3),
	.w5(32'h3ba7c9f7),
	.w6(32'hbbf22270),
	.w7(32'hbc0ca8e4),
	.w8(32'h3bb81e69),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be77a40),
	.w1(32'h3b2938dd),
	.w2(32'hba21c85a),
	.w3(32'h3b1ed1a7),
	.w4(32'h3950d7e9),
	.w5(32'hbbc3686d),
	.w6(32'h3a1d3737),
	.w7(32'hbadcef57),
	.w8(32'hbc2c944d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27ba59),
	.w1(32'hbbc65ccd),
	.w2(32'hbc1219dc),
	.w3(32'h3be020b6),
	.w4(32'h3b7ec32a),
	.w5(32'h3bf49463),
	.w6(32'h3bb3f3c5),
	.w7(32'h3bd3e600),
	.w8(32'h3b4b2518),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac945f3),
	.w1(32'h39824838),
	.w2(32'hbb4a0c26),
	.w3(32'h3b5e2db2),
	.w4(32'h3ae659b0),
	.w5(32'h3aa9b0e1),
	.w6(32'hbc14da0f),
	.w7(32'hbb5ae272),
	.w8(32'h3aabb101),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a8081),
	.w1(32'h3ab9e254),
	.w2(32'h3b2d869a),
	.w3(32'h3b7e2b15),
	.w4(32'h3b99429a),
	.w5(32'hbc2be4b9),
	.w6(32'h3c41b413),
	.w7(32'h3c1990ab),
	.w8(32'h3b16b8f6),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b227127),
	.w1(32'h3a81425a),
	.w2(32'hbbb199d6),
	.w3(32'hbbde9116),
	.w4(32'hbbc1748d),
	.w5(32'hbb19e13b),
	.w6(32'h3b63566e),
	.w7(32'hbbd0dbd5),
	.w8(32'hbbc282c7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b5b88),
	.w1(32'hbbe0162b),
	.w2(32'hbab45a97),
	.w3(32'hbbd291c7),
	.w4(32'hbbb70e70),
	.w5(32'hbbd06a4c),
	.w6(32'hbba7a259),
	.w7(32'hbb6309ab),
	.w8(32'hbb95d5f0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba705117),
	.w1(32'hbc44dfcf),
	.w2(32'hb9dcca66),
	.w3(32'hbc3ad90a),
	.w4(32'hbc16169b),
	.w5(32'h3adf02ba),
	.w6(32'hbcb8d38a),
	.w7(32'hbb8afcd8),
	.w8(32'h3b28f2af),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b939bbe),
	.w1(32'hbb8c94cd),
	.w2(32'hbb601c74),
	.w3(32'hb9f8044c),
	.w4(32'hbbd0ca79),
	.w5(32'h3999a1ce),
	.w6(32'hbc1b409d),
	.w7(32'hbbe2867e),
	.w8(32'hb97b96c7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b8690c),
	.w1(32'h3ba236d4),
	.w2(32'hbb87579b),
	.w3(32'h3b3269cd),
	.w4(32'hb9e8c5ee),
	.w5(32'h3bc5dbc6),
	.w6(32'hbaf6d8f5),
	.w7(32'hbbd788ef),
	.w8(32'h3b8b012b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0093d5),
	.w1(32'h3b833843),
	.w2(32'h3bd606aa),
	.w3(32'h3ace3e31),
	.w4(32'h3b65af9e),
	.w5(32'h3c2b5b14),
	.w6(32'hbbe0a110),
	.w7(32'hbbb39830),
	.w8(32'h3c1e0160),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b390a38),
	.w1(32'h3c382fb6),
	.w2(32'h3b883a0f),
	.w3(32'h3c21f629),
	.w4(32'hbb2e2b5c),
	.w5(32'hbabf227e),
	.w6(32'h3c34e50f),
	.w7(32'h3b9f2492),
	.w8(32'h3be4a50e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6adfc),
	.w1(32'h3b130f69),
	.w2(32'h3b8e8e2e),
	.w3(32'hbaf9299b),
	.w4(32'h398f9efc),
	.w5(32'hbbdbead4),
	.w6(32'hbb15e6ff),
	.w7(32'hb849af30),
	.w8(32'h3b366431),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7fed6),
	.w1(32'h3bfbb86b),
	.w2(32'h3b293858),
	.w3(32'h3ba38497),
	.w4(32'h3b8713b1),
	.w5(32'hbb074ac8),
	.w6(32'h3c329c62),
	.w7(32'h3a5ccbb7),
	.w8(32'hbbdd2afc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb804806),
	.w1(32'h3b28dd19),
	.w2(32'hba77782b),
	.w3(32'hbb2f458f),
	.w4(32'h3a89f7e9),
	.w5(32'h3aeeede5),
	.w6(32'hba1a87ec),
	.w7(32'hbba17b00),
	.w8(32'h3b1709ff),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae66fb1),
	.w1(32'hbb193c69),
	.w2(32'hbaac9fbd),
	.w3(32'h3a321502),
	.w4(32'h3babf4b4),
	.w5(32'h3c741b02),
	.w6(32'hbb57be78),
	.w7(32'h3b09c1e3),
	.w8(32'h3af42613),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3eb867),
	.w1(32'hbc30b546),
	.w2(32'hbaba9b82),
	.w3(32'hba7bb25b),
	.w4(32'h3bdc4e77),
	.w5(32'h3b2bdfe9),
	.w6(32'hbd207863),
	.w7(32'hbc529bf7),
	.w8(32'hbbbc8f53),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8383b8),
	.w1(32'hb9fe9424),
	.w2(32'h3bdc8a7d),
	.w3(32'hbb40e8d4),
	.w4(32'h3b7af371),
	.w5(32'h3b898063),
	.w6(32'hbc378bed),
	.w7(32'h3aaae164),
	.w8(32'hbb92d17d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6ea48),
	.w1(32'hbc5226ee),
	.w2(32'hbb59ad5a),
	.w3(32'h3ba2bdfd),
	.w4(32'h3a807837),
	.w5(32'hbbdc90d0),
	.w6(32'hbc405a89),
	.w7(32'hbbcd5a20),
	.w8(32'hbbcc6873),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e8cc5),
	.w1(32'hbb1316ed),
	.w2(32'hbb9791db),
	.w3(32'hba9b9894),
	.w4(32'hbb91ff2f),
	.w5(32'hbb3d074e),
	.w6(32'h3b453f7b),
	.w7(32'hba59307a),
	.w8(32'hbb90f335),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6db462),
	.w1(32'h3b8a972c),
	.w2(32'h3b3567af),
	.w3(32'h3b58d9a9),
	.w4(32'hbb13b89a),
	.w5(32'h3afed1df),
	.w6(32'hbc15194c),
	.w7(32'hbaaa2619),
	.w8(32'hbb46ffac),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b445bf9),
	.w1(32'hba8a4e13),
	.w2(32'hba945e53),
	.w3(32'hbaa9a34b),
	.w4(32'hbae26813),
	.w5(32'hbc262ccd),
	.w6(32'hbbf33ef8),
	.w7(32'hbbb407c0),
	.w8(32'hbc710eeb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33eaf1),
	.w1(32'hbc3c3708),
	.w2(32'hbc46a196),
	.w3(32'hbc19f6a0),
	.w4(32'hbba0c9e9),
	.w5(32'hbbcd9839),
	.w6(32'hbc3fa749),
	.w7(32'hbc348347),
	.w8(32'hbc72d1d0),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ad55e),
	.w1(32'hbc86bdb9),
	.w2(32'hbc8d8444),
	.w3(32'hbc5fee31),
	.w4(32'hbc633204),
	.w5(32'h3ba48682),
	.w6(32'hbcb4513c),
	.w7(32'hbcd7ac2a),
	.w8(32'hba8d407f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8326ea),
	.w1(32'hbbcdde9f),
	.w2(32'hbb81ba84),
	.w3(32'hbb379f1b),
	.w4(32'hbb387131),
	.w5(32'h3b5ae6e8),
	.w6(32'hbc32314f),
	.w7(32'hbbf780a5),
	.w8(32'hba9c6695),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16e671),
	.w1(32'h398292ff),
	.w2(32'h3a92be92),
	.w3(32'h3a86dca6),
	.w4(32'hbad87ad9),
	.w5(32'hbbae7ee7),
	.w6(32'hbb387f67),
	.w7(32'h38c3af4b),
	.w8(32'hbaee2c81),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2efdc5),
	.w1(32'hbbca61aa),
	.w2(32'hbb8e7122),
	.w3(32'hba931c84),
	.w4(32'hbb7fdce9),
	.w5(32'h3b2cf7e1),
	.w6(32'hbb5daca0),
	.w7(32'hbb82e6e0),
	.w8(32'hbb91d6b5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39088cae),
	.w1(32'hbbd90b17),
	.w2(32'hbb7780e9),
	.w3(32'h3bd5cd03),
	.w4(32'h3a6eff46),
	.w5(32'h3bc5681f),
	.w6(32'hbc2210d7),
	.w7(32'hbc93ca5e),
	.w8(32'h3c18dfc8),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd9b17),
	.w1(32'h3b44fa29),
	.w2(32'h3bca9337),
	.w3(32'h3bc118ec),
	.w4(32'h3bc3e217),
	.w5(32'hbb9bd3de),
	.w6(32'h3be9e689),
	.w7(32'h3b82aaa8),
	.w8(32'hbb14aecb),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccef00),
	.w1(32'h3b1660ba),
	.w2(32'hb6da08a6),
	.w3(32'h3acbac82),
	.w4(32'h3b1edfe7),
	.w5(32'hbb3157ee),
	.w6(32'hbbb24261),
	.w7(32'h3b87596d),
	.w8(32'hbc7637e3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a5a77),
	.w1(32'hbc46c420),
	.w2(32'hbc1bd5fb),
	.w3(32'hbc2900f0),
	.w4(32'hbc5519e5),
	.w5(32'h3ae41e42),
	.w6(32'hbc5d1ae5),
	.w7(32'hbc8fd272),
	.w8(32'hbab25731),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08e694),
	.w1(32'hb9bee1e4),
	.w2(32'h3a6e6306),
	.w3(32'hbb6d6407),
	.w4(32'h3a47bdba),
	.w5(32'h3c05eaa6),
	.w6(32'hbc57fdef),
	.w7(32'hbbc1b6f2),
	.w8(32'h3aa370ee),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf8d08),
	.w1(32'h3a807e22),
	.w2(32'h3bcbbcaf),
	.w3(32'hbb114847),
	.w4(32'h3c4b90a9),
	.w5(32'hbb7d754e),
	.w6(32'hbbe497f6),
	.w7(32'hbbac6413),
	.w8(32'hbb682bba),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d22c0),
	.w1(32'hbb906024),
	.w2(32'hbb9b7a9c),
	.w3(32'hb843d93a),
	.w4(32'hbb52ebcc),
	.w5(32'hbc2f13b8),
	.w6(32'hbbade1b4),
	.w7(32'hbb87a2f2),
	.w8(32'hbc4ca73d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8728dd),
	.w1(32'hbb9365a7),
	.w2(32'hba3a7072),
	.w3(32'hbc445e11),
	.w4(32'hbc2c0c69),
	.w5(32'hbabd3b2b),
	.w6(32'hbc832e8c),
	.w7(32'hbc2fca63),
	.w8(32'hbab89589),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb31449),
	.w1(32'h3b2a2963),
	.w2(32'hbbe3f89c),
	.w3(32'h3c263582),
	.w4(32'h3b9d38b9),
	.w5(32'h3bee500f),
	.w6(32'h3bb07c6a),
	.w7(32'h3bb68868),
	.w8(32'h3944985c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9593a8f),
	.w1(32'h3c23d93c),
	.w2(32'h3c464011),
	.w3(32'h3be3168d),
	.w4(32'h3b35fc5a),
	.w5(32'h3abea775),
	.w6(32'hbb28e92f),
	.w7(32'h3b87f55c),
	.w8(32'h3b5a4a15),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88e1a8),
	.w1(32'h3b2d6870),
	.w2(32'h3a8e9398),
	.w3(32'h3ba68fe3),
	.w4(32'h3bdd42a7),
	.w5(32'h3b161581),
	.w6(32'h3c5094cf),
	.w7(32'h3ba7b166),
	.w8(32'hb90c3371),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3c05d),
	.w1(32'hbae02fe3),
	.w2(32'h3afec889),
	.w3(32'hbb3f3f03),
	.w4(32'hbb2b4b85),
	.w5(32'hbaebc105),
	.w6(32'hbc281021),
	.w7(32'hbba11884),
	.w8(32'hbba7f139),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d1b5f),
	.w1(32'h3ba7c469),
	.w2(32'hb9ac45dd),
	.w3(32'h3a0fa8aa),
	.w4(32'hbc1a8b79),
	.w5(32'h3bd76e27),
	.w6(32'hbcbcb33b),
	.w7(32'hbbb8b48a),
	.w8(32'h3b554301),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba140e52),
	.w1(32'h3b2d11fa),
	.w2(32'hbb42dcd4),
	.w3(32'h398bb9d0),
	.w4(32'h3a80ce6d),
	.w5(32'hbacd1e74),
	.w6(32'h3a8cda25),
	.w7(32'h3b1149a7),
	.w8(32'hbc1545e1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0441bf),
	.w1(32'hbba86aa0),
	.w2(32'hbb8a96a0),
	.w3(32'hbc503122),
	.w4(32'hba2c6b51),
	.w5(32'hba4e6a34),
	.w6(32'hbc1357d9),
	.w7(32'hbc228b18),
	.w8(32'hbb0d9d59),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb03aed),
	.w1(32'hbbb211f0),
	.w2(32'h3a896f6e),
	.w3(32'hbb0e8d21),
	.w4(32'h3bbc7179),
	.w5(32'h3c86efda),
	.w6(32'hbb8e1969),
	.w7(32'hb9c7856c),
	.w8(32'h3b9320d6),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7491ca),
	.w1(32'h3a959cb8),
	.w2(32'h3c25e6b6),
	.w3(32'h3b907354),
	.w4(32'h3c04e207),
	.w5(32'hbb20f456),
	.w6(32'hbc8aec94),
	.w7(32'h3b9d3958),
	.w8(32'h3a80ba02),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1176db),
	.w1(32'hb9fe7926),
	.w2(32'h3a0b82ef),
	.w3(32'h3b122b01),
	.w4(32'hba7cac8a),
	.w5(32'h3baea2de),
	.w6(32'h3bb45977),
	.w7(32'h3ba1f6bc),
	.w8(32'h3b0415ab),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba528312),
	.w1(32'h3c439094),
	.w2(32'h3b5db163),
	.w3(32'h3bc32ae2),
	.w4(32'h3abe63bb),
	.w5(32'hb9583e52),
	.w6(32'h3b050734),
	.w7(32'h3a29efec),
	.w8(32'hbbba90d2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01c8eb),
	.w1(32'h3b1743aa),
	.w2(32'hbc20a24b),
	.w3(32'hbba227cf),
	.w4(32'hbbbc575e),
	.w5(32'h3b53b395),
	.w6(32'hbb2e9eb8),
	.w7(32'hbb333c39),
	.w8(32'h3bbdb13d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3a74e),
	.w1(32'h3b35ca6c),
	.w2(32'hb99636d5),
	.w3(32'h3c14074e),
	.w4(32'h3a853fd1),
	.w5(32'hbb764d9b),
	.w6(32'h3c69ccc4),
	.w7(32'h3b52aec6),
	.w8(32'hb9ed5b24),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd756c),
	.w1(32'hb921a1e7),
	.w2(32'h3b1c7549),
	.w3(32'hbc84fc79),
	.w4(32'hbae5e6ff),
	.w5(32'hbb942937),
	.w6(32'hbcb6b625),
	.w7(32'h3b7bd308),
	.w8(32'hbbfc60c5),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a5f0c),
	.w1(32'h3a32e3a4),
	.w2(32'h3ab0247d),
	.w3(32'h3b849e9d),
	.w4(32'hbb41e5bc),
	.w5(32'h3a892fd3),
	.w6(32'h3a182908),
	.w7(32'hbbd7d9e1),
	.w8(32'h3ad66f5d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ef58e),
	.w1(32'hbb5d967c),
	.w2(32'hbba5c99e),
	.w3(32'h39ecbcaf),
	.w4(32'h3b6b84bc),
	.w5(32'h3be5dcaf),
	.w6(32'h3c2d1282),
	.w7(32'h3bd1d085),
	.w8(32'h3acf3507),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea0287),
	.w1(32'hbafcd3ae),
	.w2(32'h3b8f9218),
	.w3(32'h3c2d8f00),
	.w4(32'hbaa3aafc),
	.w5(32'h3a888f85),
	.w6(32'hbba48859),
	.w7(32'hbbd6e863),
	.w8(32'h3b6a8173),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7149a3),
	.w1(32'h3c2b1ead),
	.w2(32'h3b818bb2),
	.w3(32'h3a85aebf),
	.w4(32'h3b112812),
	.w5(32'hbbc21a46),
	.w6(32'h3b89dce3),
	.w7(32'h3ade7c59),
	.w8(32'hbbb43134),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd8493),
	.w1(32'hbbfad6d7),
	.w2(32'hbadd9478),
	.w3(32'hbc23ffe9),
	.w4(32'h3b97fc58),
	.w5(32'h3ba4bfb7),
	.w6(32'hbc642401),
	.w7(32'h3a47505d),
	.w8(32'h3a81a57b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa84e7e),
	.w1(32'h3ba42fb7),
	.w2(32'h3bd00917),
	.w3(32'h3bd09db9),
	.w4(32'h3ac314c3),
	.w5(32'hbb82a230),
	.w6(32'h3b197974),
	.w7(32'h3b813fbb),
	.w8(32'hbb9ee7f1),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c68f9),
	.w1(32'h3a9bf2f6),
	.w2(32'hbc036553),
	.w3(32'hbc0cbd01),
	.w4(32'hbc21ee3a),
	.w5(32'hb94b6d38),
	.w6(32'h3bbf1cfd),
	.w7(32'hbba5561a),
	.w8(32'hbaee5a83),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba325216),
	.w1(32'hbbbfdde9),
	.w2(32'h38ff84ff),
	.w3(32'h3b891bf0),
	.w4(32'hb986a74b),
	.w5(32'hba9c656f),
	.w6(32'hbb956839),
	.w7(32'hbb1902e6),
	.w8(32'hbc22fe67),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb868946),
	.w1(32'h39b0d86e),
	.w2(32'hbad1bd20),
	.w3(32'hbb3229f1),
	.w4(32'h3b9b2511),
	.w5(32'hbc5a7f9a),
	.w6(32'hba88db37),
	.w7(32'hbba49ec7),
	.w8(32'hbbf0a4d8),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a742f),
	.w1(32'hbc177d6d),
	.w2(32'hbb0114f4),
	.w3(32'hbb2d0047),
	.w4(32'hbb9208f4),
	.w5(32'hbb5e6082),
	.w6(32'hbc38206d),
	.w7(32'hbaa67ad5),
	.w8(32'hbb8beb73),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fba17),
	.w1(32'h3b834485),
	.w2(32'h3b30430f),
	.w3(32'h3b6dce16),
	.w4(32'hba9ce018),
	.w5(32'hbb8b75e3),
	.w6(32'h3aa61ad6),
	.w7(32'hbae9b333),
	.w8(32'hbb299a39),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb985c22),
	.w1(32'hbab794b8),
	.w2(32'hbb840c0e),
	.w3(32'hbb3eed69),
	.w4(32'hbb5d3e7e),
	.w5(32'hbb0e253a),
	.w6(32'hbb0530ba),
	.w7(32'h3af002fb),
	.w8(32'hbbe50b2a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5c0f3),
	.w1(32'hbb3de59d),
	.w2(32'h399d0d7e),
	.w3(32'hba7a7658),
	.w4(32'hbae98b02),
	.w5(32'hbc0393da),
	.w6(32'h3b6fd965),
	.w7(32'hbbec62b8),
	.w8(32'hbc36f444),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21f9c9),
	.w1(32'hbc6c1c62),
	.w2(32'hbc177bc8),
	.w3(32'hbc49c212),
	.w4(32'hbc145dc7),
	.w5(32'h3c7517a6),
	.w6(32'hbc1d77d4),
	.w7(32'hbc379943),
	.w8(32'h3c370c1e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c333291),
	.w1(32'h3bb7157a),
	.w2(32'h3bb026e6),
	.w3(32'h3be38b94),
	.w4(32'h3c11f510),
	.w5(32'h3c134775),
	.w6(32'h3bdf23dc),
	.w7(32'h3c042800),
	.w8(32'h3b97495e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba81457),
	.w1(32'h3b70641d),
	.w2(32'h3c13e739),
	.w3(32'h3bcaf0ea),
	.w4(32'h3aa9eb0c),
	.w5(32'h3b9364af),
	.w6(32'hbb97c1e5),
	.w7(32'h3bccc0f7),
	.w8(32'h3ac6a6a0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6bea5),
	.w1(32'hba6b49b2),
	.w2(32'h3a5807a5),
	.w3(32'h3b29bfb7),
	.w4(32'h3c055dce),
	.w5(32'h3bc06578),
	.w6(32'h3be57888),
	.w7(32'h3b3fe9f6),
	.w8(32'h3a6f2ca0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6d070),
	.w1(32'h3a74d84c),
	.w2(32'hbbb8c735),
	.w3(32'h3b500325),
	.w4(32'hbb5c48a3),
	.w5(32'hbc519662),
	.w6(32'h39efb526),
	.w7(32'hbc13d578),
	.w8(32'hbc4011df),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc088e4f),
	.w1(32'hbbea9e84),
	.w2(32'hbc2f521b),
	.w3(32'hbb11ae92),
	.w4(32'hbb0f9716),
	.w5(32'hbb0b44cc),
	.w6(32'hbb87b3fa),
	.w7(32'hbb860fcd),
	.w8(32'hba0ed693),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bb4b4),
	.w1(32'hbbb1bcab),
	.w2(32'h39f95b92),
	.w3(32'h3b8b279c),
	.w4(32'hbba5259e),
	.w5(32'hba820a7c),
	.w6(32'hbc037443),
	.w7(32'hbb8e1d28),
	.w8(32'hbb38b85e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b694c52),
	.w1(32'h3ac5a783),
	.w2(32'hbbfa93ba),
	.w3(32'h3b1bc905),
	.w4(32'hbb7adc32),
	.w5(32'hbb9e7437),
	.w6(32'h3b0bee5f),
	.w7(32'hbbe07d98),
	.w8(32'h3b5b70a1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ae5026),
	.w1(32'h3bb320f2),
	.w2(32'hbb5f0fb9),
	.w3(32'h3bcd7484),
	.w4(32'h3b879b9b),
	.w5(32'h3a558ede),
	.w6(32'h3c1b8fbd),
	.w7(32'h3be80f2d),
	.w8(32'h3ac2d5a0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb01273),
	.w1(32'hba1310eb),
	.w2(32'h3b1f6085),
	.w3(32'hbb82342a),
	.w4(32'hba8d11ec),
	.w5(32'h3bf7336e),
	.w6(32'h3bb3924b),
	.w7(32'h3b978592),
	.w8(32'h3b857a10),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e36b0a),
	.w1(32'h3b62df1d),
	.w2(32'h3b8dcb51),
	.w3(32'h3b57ac6f),
	.w4(32'h3b45d503),
	.w5(32'hbaa3a2f8),
	.w6(32'h3c2e5f74),
	.w7(32'h3c2ca825),
	.w8(32'h3ab41762),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bd4d3),
	.w1(32'h3b660ec7),
	.w2(32'h3b86aa10),
	.w3(32'h3b523b70),
	.w4(32'hb9f78999),
	.w5(32'h3a5beccc),
	.w6(32'h3be217c4),
	.w7(32'h3ba218ba),
	.w8(32'hbba52761),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb113697),
	.w1(32'hbbfd2f73),
	.w2(32'hbbcee4ab),
	.w3(32'hbb9421ef),
	.w4(32'h3a9cfd59),
	.w5(32'h3b7f9e86),
	.w6(32'hba95c250),
	.w7(32'hbb14ef47),
	.w8(32'h3c8445fe),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c010b87),
	.w1(32'h3c902b4a),
	.w2(32'h3c54c6d4),
	.w3(32'h3b9ba13c),
	.w4(32'h3c98855d),
	.w5(32'h3a3cb6f6),
	.w6(32'h3d2403fc),
	.w7(32'h3d05e3bc),
	.w8(32'hba6c1fb2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf00c1d),
	.w1(32'hba93ccfc),
	.w2(32'hbb22b461),
	.w3(32'h3b1bfcd5),
	.w4(32'hbb44a863),
	.w5(32'hbba39242),
	.w6(32'h3b15cd6a),
	.w7(32'hbb3040ba),
	.w8(32'hbbd9fb5a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed029b),
	.w1(32'hbbb497d7),
	.w2(32'hbc05d588),
	.w3(32'hbc0e2589),
	.w4(32'hbc13670f),
	.w5(32'h3b05a61a),
	.w6(32'hbb9edec3),
	.w7(32'hbc3f584e),
	.w8(32'h3b9194dc),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b292ec),
	.w1(32'h3ae003b2),
	.w2(32'h3942aad7),
	.w3(32'hba0b1e86),
	.w4(32'h3b0da385),
	.w5(32'h3b16415f),
	.w6(32'h39f354e7),
	.w7(32'h39ae33f6),
	.w8(32'hbaccecf1),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b05be),
	.w1(32'hbb225ad8),
	.w2(32'h3b017d2d),
	.w3(32'h39a9ae4f),
	.w4(32'h3b045a8d),
	.w5(32'hbbe125c8),
	.w6(32'hbb973a3e),
	.w7(32'h3bb0525c),
	.w8(32'h3b81ae14),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad24f62),
	.w1(32'hbb802544),
	.w2(32'hbc0e243d),
	.w3(32'hbbac93a4),
	.w4(32'hbb8489ee),
	.w5(32'h3b502a67),
	.w6(32'h37171b4b),
	.w7(32'h3a7be179),
	.w8(32'h3c2d7443),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c2ee8),
	.w1(32'h3b23b6b5),
	.w2(32'h3bad4383),
	.w3(32'h3bb961b7),
	.w4(32'h3b982aae),
	.w5(32'hbc1e64a9),
	.w6(32'h3aca698c),
	.w7(32'h3b518017),
	.w8(32'hbb82ec08),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf360a9),
	.w1(32'hbc42b295),
	.w2(32'hbc82e601),
	.w3(32'hbbaf44b2),
	.w4(32'hbc1ebabc),
	.w5(32'hb9a91a55),
	.w6(32'hbc01c1ab),
	.w7(32'hbcc1a679),
	.w8(32'hbad138b8),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e438e),
	.w1(32'hbc031934),
	.w2(32'hbbbd1ee9),
	.w3(32'hbaa03773),
	.w4(32'hbab1e5b9),
	.w5(32'hbb469950),
	.w6(32'hbb9b7417),
	.w7(32'hbb8f925d),
	.w8(32'hbb6efdf6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91dba4),
	.w1(32'hbb07ce97),
	.w2(32'h3a4d0603),
	.w3(32'hbb2bfe46),
	.w4(32'h3b280490),
	.w5(32'hbabecbb9),
	.w6(32'hbc059459),
	.w7(32'h3ba0158f),
	.w8(32'hba949796),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb962e07b),
	.w1(32'h3b2bb425),
	.w2(32'hbb303c6a),
	.w3(32'h3b039c87),
	.w4(32'hbb290a66),
	.w5(32'hbb9c58cc),
	.w6(32'h3c83e6b8),
	.w7(32'hbbd23b68),
	.w8(32'hbbc5e67b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24bd04),
	.w1(32'hbbae9cf4),
	.w2(32'h39bad539),
	.w3(32'hbbabb866),
	.w4(32'hba2bb17a),
	.w5(32'hbb731961),
	.w6(32'hbc55a170),
	.w7(32'hbb2bb643),
	.w8(32'hbc47b88e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e907f),
	.w1(32'h3b135c48),
	.w2(32'hbbe079d6),
	.w3(32'hbbb8799f),
	.w4(32'hbae0f3a6),
	.w5(32'h3a667e0d),
	.w6(32'hbc672cc0),
	.w7(32'hbc9b063a),
	.w8(32'hbb6e82b7),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13ed66),
	.w1(32'hbb25dc54),
	.w2(32'h3c39dfd9),
	.w3(32'h3a93d1af),
	.w4(32'hbaf190dc),
	.w5(32'h39664b1a),
	.w6(32'hbb8378bf),
	.w7(32'h3bfca4e4),
	.w8(32'h3b0e8b2e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fc506),
	.w1(32'h3bfeabe3),
	.w2(32'h3bef0552),
	.w3(32'h3b96acfe),
	.w4(32'hbb65d356),
	.w5(32'hb9cfca29),
	.w6(32'h3c948fb7),
	.w7(32'h3b996168),
	.w8(32'h3bb1fe7a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf6dd7),
	.w1(32'hbbfa66a9),
	.w2(32'hbabc3d4c),
	.w3(32'h3bc24a4d),
	.w4(32'h3b28efcd),
	.w5(32'h3b52e669),
	.w6(32'hbbd596fa),
	.w7(32'hbc1bb87e),
	.w8(32'h3b9bb6f0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae033ae),
	.w1(32'h3bd5b461),
	.w2(32'h3bfa5fcc),
	.w3(32'h3c027cb2),
	.w4(32'h386bcb38),
	.w5(32'hbb0e47e2),
	.w6(32'h3b51bed7),
	.w7(32'h3b3e927c),
	.w8(32'hbb045131),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbaee2),
	.w1(32'hbb03382b),
	.w2(32'h3b769e8b),
	.w3(32'h3a0eda69),
	.w4(32'h3b2b0d25),
	.w5(32'hbc8e6f36),
	.w6(32'hbc2ccfdc),
	.w7(32'hbb3d41a2),
	.w8(32'hbc83272e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc316852),
	.w1(32'hbc22f606),
	.w2(32'hbc294859),
	.w3(32'hbc10d281),
	.w4(32'hbc1edf25),
	.w5(32'hbc2a792f),
	.w6(32'hbc0f6d22),
	.w7(32'hbc29beaa),
	.w8(32'hbc1620af),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98daea),
	.w1(32'hbc7ebcff),
	.w2(32'hbc50204a),
	.w3(32'hbbf437a0),
	.w4(32'hbc6a32e8),
	.w5(32'h3bf2b3e5),
	.w6(32'hbbb64908),
	.w7(32'hbc462d4b),
	.w8(32'hba9d0faf),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44ff0e),
	.w1(32'hbbc203f6),
	.w2(32'hbbeb7e19),
	.w3(32'hbb4c8cf6),
	.w4(32'hbb317d86),
	.w5(32'hbb3f617d),
	.w6(32'hbc78367f),
	.w7(32'hbc5525cb),
	.w8(32'hbb388f25),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ea920),
	.w1(32'hbb392765),
	.w2(32'h3b3cede9),
	.w3(32'h3a8cec48),
	.w4(32'hbab194e4),
	.w5(32'hbb4a2aaa),
	.w6(32'hbbb669b1),
	.w7(32'h3abbd06d),
	.w8(32'hbb4089e7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab12c61),
	.w1(32'h3ad8d4b9),
	.w2(32'h3b6946b0),
	.w3(32'h3996b2ef),
	.w4(32'hbb10c98d),
	.w5(32'hbb8544f5),
	.w6(32'h3a5f340f),
	.w7(32'h3a75fe27),
	.w8(32'hb9d1dcf0),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d8fdc),
	.w1(32'hbbba123c),
	.w2(32'hbb372209),
	.w3(32'hbb5ee993),
	.w4(32'hbbeb024b),
	.w5(32'h3bcc0c85),
	.w6(32'hbc60b81e),
	.w7(32'hbc351111),
	.w8(32'h3c099421),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1dd94),
	.w1(32'h3c909ac1),
	.w2(32'h3c90fa1d),
	.w3(32'h3bc470de),
	.w4(32'h3c0d59dd),
	.w5(32'h3b2cbc14),
	.w6(32'h3c821ba8),
	.w7(32'h3c82b8ac),
	.w8(32'h3bd06817),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfae012),
	.w1(32'hbaf17200),
	.w2(32'h3a0cfe60),
	.w3(32'h3b365092),
	.w4(32'h3afa8dfe),
	.w5(32'h3b3ad9a0),
	.w6(32'hbadfd00e),
	.w7(32'h39b16b64),
	.w8(32'h3a2b6ee8),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c67aa),
	.w1(32'h39fc8d1d),
	.w2(32'h3b04d1c9),
	.w3(32'h3b9c3223),
	.w4(32'hbb8f5276),
	.w5(32'hbb405256),
	.w6(32'hbb55fa54),
	.w7(32'hbaf8c2a4),
	.w8(32'hbc514ad9),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7fd01),
	.w1(32'hbbefb384),
	.w2(32'hbadb18f4),
	.w3(32'hbbf39750),
	.w4(32'hbbd52078),
	.w5(32'hbaa82824),
	.w6(32'hbc33be54),
	.w7(32'hbc6c6118),
	.w8(32'h3a9374c6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b089f),
	.w1(32'h3c70cce2),
	.w2(32'h3c095721),
	.w3(32'h3b1bc22e),
	.w4(32'h3b65a661),
	.w5(32'h398eeb78),
	.w6(32'h39d46e11),
	.w7(32'h3baed66d),
	.w8(32'hbb840c1c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ae6ba),
	.w1(32'hbc29c1a5),
	.w2(32'hbc429600),
	.w3(32'hbbe67702),
	.w4(32'hbb2c43dd),
	.w5(32'h3c13d38a),
	.w6(32'hbc254992),
	.w7(32'hbc250321),
	.w8(32'h3ac99a23),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef10f1),
	.w1(32'hba2a23cd),
	.w2(32'hbc470592),
	.w3(32'hbb07f279),
	.w4(32'h3a7a24cc),
	.w5(32'h3bb37b1c),
	.w6(32'hbc753ebd),
	.w7(32'hbc440d7e),
	.w8(32'hbb35448e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58e806),
	.w1(32'h3af019c5),
	.w2(32'h3b74b538),
	.w3(32'h3b3722d0),
	.w4(32'hbbd147f9),
	.w5(32'hbc0f5724),
	.w6(32'hbb18141d),
	.w7(32'hbb10c4cd),
	.w8(32'hbc0c4ddd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf499b7),
	.w1(32'hbb9690b3),
	.w2(32'hbbff1a05),
	.w3(32'hbbd0298d),
	.w4(32'hba7d9763),
	.w5(32'hbb547c27),
	.w6(32'hbbe9ac81),
	.w7(32'hbb308aff),
	.w8(32'hbc40f8f5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39462211),
	.w1(32'hbba7d218),
	.w2(32'hbc0296b1),
	.w3(32'hbb386747),
	.w4(32'h3b7adacb),
	.w5(32'h3a9decc9),
	.w6(32'hbc3d141e),
	.w7(32'h3bb62558),
	.w8(32'hbabca03e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a679c5),
	.w1(32'h3b5804db),
	.w2(32'h3bf8fd16),
	.w3(32'h3abe40ab),
	.w4(32'h3b36a4e4),
	.w5(32'hbac683b5),
	.w6(32'h3a3614c7),
	.w7(32'h3bdd649a),
	.w8(32'hbba2a64b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b152e19),
	.w1(32'hbb9f0058),
	.w2(32'hbb86e5fb),
	.w3(32'hbbe8408b),
	.w4(32'h3b6d84cf),
	.w5(32'hbc13e0cd),
	.w6(32'hbc9d6e16),
	.w7(32'hbb9447a3),
	.w8(32'hbc6ffad3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb876dc5),
	.w1(32'hbc8dd031),
	.w2(32'hbbe4403f),
	.w3(32'hb9d83435),
	.w4(32'h3b81e2d5),
	.w5(32'h3aa0c4c2),
	.w6(32'hbca3910b),
	.w7(32'hbc4e34e8),
	.w8(32'h3be0a193),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcf92e),
	.w1(32'h3bc88290),
	.w2(32'h3a933de3),
	.w3(32'h3c031beb),
	.w4(32'hba67252b),
	.w5(32'h3b7bc8b6),
	.w6(32'h3cb8e40f),
	.w7(32'h3be45f34),
	.w8(32'h3ac06693),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf0294),
	.w1(32'h3bc663c7),
	.w2(32'h3a8b790b),
	.w3(32'hbc255a32),
	.w4(32'h39736cb9),
	.w5(32'hb68c5815),
	.w6(32'hbc9658fd),
	.w7(32'h3af594be),
	.w8(32'hb78bff01),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb53744e6),
	.w1(32'hb549d3a7),
	.w2(32'h36be926b),
	.w3(32'hb7e0e431),
	.w4(32'hb66d8610),
	.w5(32'h3780104e),
	.w6(32'hb8560437),
	.w7(32'hb7a97b58),
	.w8(32'hb753d261),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b65cfe),
	.w1(32'hb9b08a59),
	.w2(32'hb99d22fe),
	.w3(32'hb989cf97),
	.w4(32'hb8fef2fb),
	.w5(32'hb98b4415),
	.w6(32'hb90df0d9),
	.w7(32'hb8f603d1),
	.w8(32'hb93cdd89),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d64b12),
	.w1(32'hb8d3501c),
	.w2(32'hb8a9f7a4),
	.w3(32'hb868f1fd),
	.w4(32'hb8cbb793),
	.w5(32'hb90ee16d),
	.w6(32'hb86dd0ba),
	.w7(32'hb88f18da),
	.w8(32'hb8af4d07),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369611b0),
	.w1(32'hb6e0e496),
	.w2(32'h37254333),
	.w3(32'hb6d10249),
	.w4(32'hb66c1487),
	.w5(32'hb62c42cb),
	.w6(32'hb8330097),
	.w7(32'hb7480aab),
	.w8(32'hb717de03),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8413f65),
	.w1(32'hb8a0acda),
	.w2(32'hb7c93823),
	.w3(32'h37ce0fb7),
	.w4(32'h3640b8b0),
	.w5(32'hb8380956),
	.w6(32'h3810b077),
	.w7(32'hb81c8a42),
	.w8(32'hb8e8afee),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb864905a),
	.w1(32'hb7684114),
	.w2(32'hb7c38bcb),
	.w3(32'h3867709d),
	.w4(32'h382f1745),
	.w5(32'h37a7281f),
	.w6(32'hb7dce841),
	.w7(32'hb74c3b58),
	.w8(32'hb729745b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36df6905),
	.w1(32'hb7a34b11),
	.w2(32'hb81f7fa1),
	.w3(32'h37898185),
	.w4(32'h378ee67b),
	.w5(32'h37d06826),
	.w6(32'hb7bdcd62),
	.w7(32'hb7d189c3),
	.w8(32'h371fe7ba),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d46410),
	.w1(32'h37d520dd),
	.w2(32'h384b85b1),
	.w3(32'h3806bf55),
	.w4(32'h3893388b),
	.w5(32'h38b0dd0a),
	.w6(32'h3826261b),
	.w7(32'h37ce3c04),
	.w8(32'h38b66416),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a346c1),
	.w1(32'hb5400824),
	.w2(32'h374e7066),
	.w3(32'hb7225c92),
	.w4(32'hb5a86eeb),
	.w5(32'h369e086f),
	.w6(32'hb722219d),
	.w7(32'h3765570c),
	.w8(32'h3761ac69),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c092c3),
	.w1(32'hb8931cb5),
	.w2(32'h38719630),
	.w3(32'hb8c0bd8d),
	.w4(32'hb736f43c),
	.w5(32'h3828dacc),
	.w6(32'hb88e9962),
	.w7(32'h37d3fe55),
	.w8(32'h3804f03f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b89c92),
	.w1(32'hb721f219),
	.w2(32'h34c258b0),
	.w3(32'hb688b2ca),
	.w4(32'h33ff4434),
	.w5(32'hb7107f02),
	.w6(32'hb6ca521d),
	.w7(32'hb73ab433),
	.w8(32'hb72fff0c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7360d6b),
	.w1(32'hb7c15950),
	.w2(32'hb7ce93fb),
	.w3(32'hb8362fe5),
	.w4(32'hb7beda21),
	.w5(32'h366c590d),
	.w6(32'hb84ae5da),
	.w7(32'hb7e66b1b),
	.w8(32'h37c3ba8d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37891eec),
	.w1(32'hb6ce1889),
	.w2(32'h3712b046),
	.w3(32'hb7bd599b),
	.w4(32'h35a30467),
	.w5(32'h3866f8be),
	.w6(32'h37d67062),
	.w7(32'hb7480225),
	.w8(32'h3502afc5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982580a),
	.w1(32'hb9836db2),
	.w2(32'hb8d6df0d),
	.w3(32'hb8ea9b66),
	.w4(32'hb8fff70e),
	.w5(32'hb8b5be68),
	.w6(32'hb84de74e),
	.w7(32'hb892d7bf),
	.w8(32'hb89a37ab),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c29933),
	.w1(32'h38558103),
	.w2(32'h393c1cdc),
	.w3(32'h3944d593),
	.w4(32'h390e9c4a),
	.w5(32'h3962e3d0),
	.w6(32'h38fc8b28),
	.w7(32'h372dca32),
	.w8(32'h39279684),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f5357),
	.w1(32'hb945b1aa),
	.w2(32'hb9406840),
	.w3(32'hb8bcf195),
	.w4(32'hb9069566),
	.w5(32'hb900fbce),
	.w6(32'hb878988e),
	.w7(32'hb8cdc48b),
	.w8(32'hb81af9e8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80386ad),
	.w1(32'hb764e1da),
	.w2(32'h36e47be5),
	.w3(32'h3709f6ed),
	.w4(32'hb7183fda),
	.w5(32'h37a08cf0),
	.w6(32'hb70ed8d3),
	.w7(32'hb76f6651),
	.w8(32'h379f7446),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fd54dd),
	.w1(32'hb731293b),
	.w2(32'h36979ba4),
	.w3(32'hb6f9e474),
	.w4(32'hb71efbf0),
	.w5(32'hb73cdcc4),
	.w6(32'hb74aa9c9),
	.w7(32'hb78ab242),
	.w8(32'hb747990d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7076146),
	.w1(32'h3802b183),
	.w2(32'h37697f87),
	.w3(32'h373e3946),
	.w4(32'h3766c41c),
	.w5(32'h3729d4cc),
	.w6(32'h37289b09),
	.w7(32'h3826e434),
	.w8(32'h37c05dfb),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37864330),
	.w1(32'hb773f269),
	.w2(32'h360d2e83),
	.w3(32'h3761463a),
	.w4(32'h36785f61),
	.w5(32'h3706ebbd),
	.w6(32'hb7ebb87b),
	.w7(32'h358c03bf),
	.w8(32'hb77c81fc),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb847b137),
	.w1(32'hb8294769),
	.w2(32'h384b541c),
	.w3(32'hb877cb51),
	.w4(32'h3831532d),
	.w5(32'h385d1faa),
	.w6(32'hb879cc0e),
	.w7(32'h37c6cd6c),
	.w8(32'h363049dc),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86d7744),
	.w1(32'hb91395c6),
	.w2(32'hb88b6c9f),
	.w3(32'hb8592ff3),
	.w4(32'hb8f80a1d),
	.w5(32'hb8093169),
	.w6(32'hb8e2521d),
	.w7(32'hb8e89523),
	.w8(32'hb8b60530),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b8e5a5),
	.w1(32'h390629ac),
	.w2(32'h38908ad9),
	.w3(32'h384e26b2),
	.w4(32'h38b49b5f),
	.w5(32'h381f479c),
	.w6(32'h37755e5f),
	.w7(32'h385d29ed),
	.w8(32'h384deafb),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385c4160),
	.w1(32'h38a42691),
	.w2(32'h37ceb7b0),
	.w3(32'h383feef8),
	.w4(32'h37a015b8),
	.w5(32'h3832140f),
	.w6(32'h38529ced),
	.w7(32'h379016a7),
	.w8(32'h377c5580),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63b9add),
	.w1(32'hb82f70b3),
	.w2(32'h380ec3e1),
	.w3(32'hb86420c3),
	.w4(32'hb7e3d64f),
	.w5(32'h381ddb29),
	.w6(32'hb8c704f5),
	.w7(32'hb7522519),
	.w8(32'h38554148),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386dcd93),
	.w1(32'h38306880),
	.w2(32'h3826734f),
	.w3(32'h37977fc2),
	.w4(32'h37802b09),
	.w5(32'h37913f4c),
	.w6(32'h37eb9a52),
	.w7(32'h3798112e),
	.w8(32'h3721e186),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68a83a3),
	.w1(32'hb7a1847a),
	.w2(32'h364cface),
	.w3(32'hb7526e45),
	.w4(32'hb6cc6233),
	.w5(32'h3731c360),
	.w6(32'hb7f17c1a),
	.w7(32'hb66c1aec),
	.w8(32'hb77b9fc4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ee6c56),
	.w1(32'h37373ebd),
	.w2(32'h388466da),
	.w3(32'h37f40165),
	.w4(32'h3803d267),
	.w5(32'h37ca3231),
	.w6(32'h3837204d),
	.w7(32'h384b40c9),
	.w8(32'h38a2782c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cee50a),
	.w1(32'hb8132d18),
	.w2(32'hb67fa50f),
	.w3(32'hb7b9247b),
	.w4(32'hb829b64a),
	.w5(32'h34953fd5),
	.w6(32'hb7e061f8),
	.w7(32'hb753e05b),
	.w8(32'hb6a29c3e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b08e70),
	.w1(32'hb73a334b),
	.w2(32'h380a426d),
	.w3(32'h372d18fc),
	.w4(32'hb81c7ad6),
	.w5(32'h37b7ce83),
	.w6(32'hb7807014),
	.w7(32'hb7b72063),
	.w8(32'h3777b2b5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule