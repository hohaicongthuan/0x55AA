module layer_10_featuremap_389(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31e715),
	.w1(32'h3a143c69),
	.w2(32'hba382dc4),
	.w3(32'hbbacd15e),
	.w4(32'h3a9eda6a),
	.w5(32'hba78107c),
	.w6(32'h3b0cc7d7),
	.w7(32'h3b8359b3),
	.w8(32'h3acab2d5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fbe9e),
	.w1(32'hbb78d628),
	.w2(32'hbaeabfb8),
	.w3(32'hbaca821a),
	.w4(32'hbbaae4ae),
	.w5(32'hbb29072a),
	.w6(32'hb9fe71ca),
	.w7(32'hbb272ba0),
	.w8(32'h3b4113a6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa97c9),
	.w1(32'hbaf63c11),
	.w2(32'h3a8754b5),
	.w3(32'hbb49c487),
	.w4(32'hbaeab603),
	.w5(32'hbb92a644),
	.w6(32'hbb25f084),
	.w7(32'h3a868ef2),
	.w8(32'h3a8416f4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dad08),
	.w1(32'h3a99862d),
	.w2(32'hbb9da9e0),
	.w3(32'hbabe0df5),
	.w4(32'hbb7ef87b),
	.w5(32'hbb04405c),
	.w6(32'h3ba529cd),
	.w7(32'hbb08c1f2),
	.w8(32'hbade341f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9bf8e),
	.w1(32'h3b75a011),
	.w2(32'h3a1f0cda),
	.w3(32'h3b7a0cf4),
	.w4(32'h3b1ccde6),
	.w5(32'hbb989a1d),
	.w6(32'hbb660cdb),
	.w7(32'hb90d8d65),
	.w8(32'hbb4b6124),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3eb760),
	.w1(32'hbab5b464),
	.w2(32'hbad7f316),
	.w3(32'hb9b84e31),
	.w4(32'hbb2cf8c5),
	.w5(32'hb9955090),
	.w6(32'h3a73c91c),
	.w7(32'hbb213a82),
	.w8(32'h3b3e7d01),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f7c8d),
	.w1(32'h3bcb5a11),
	.w2(32'h3c34dcda),
	.w3(32'hbb2f86ca),
	.w4(32'h3bc77173),
	.w5(32'h3b253b1f),
	.w6(32'hba93ab14),
	.w7(32'h3c0278d5),
	.w8(32'h39b906f4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b417de3),
	.w1(32'h3c14ed3b),
	.w2(32'hbaea76ac),
	.w3(32'h3b679d22),
	.w4(32'h3c4b4d80),
	.w5(32'h3a01ed97),
	.w6(32'h3aa01597),
	.w7(32'h3c0e7f35),
	.w8(32'hbb34353c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe98410),
	.w1(32'h38c26f19),
	.w2(32'h3a071b92),
	.w3(32'h39b8dae5),
	.w4(32'h3b68b93b),
	.w5(32'hbbbab021),
	.w6(32'h39bfb1ff),
	.w7(32'h3b8ea36e),
	.w8(32'hbbbb1fb7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb632f2e),
	.w1(32'h3ae3e966),
	.w2(32'h3ac7c4b3),
	.w3(32'h3a09bfbe),
	.w4(32'hbb49be9e),
	.w5(32'h3b195173),
	.w6(32'h3ac8b9ed),
	.w7(32'h3a0925d1),
	.w8(32'h3c00e770),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00b7d4),
	.w1(32'hb87e755f),
	.w2(32'hba0d2bbd),
	.w3(32'hb981f420),
	.w4(32'h3a8c908b),
	.w5(32'h3b65ac97),
	.w6(32'h3b058ed2),
	.w7(32'hbb82b893),
	.w8(32'hbb24dda6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba760d17),
	.w1(32'hbb882791),
	.w2(32'h3b6ff39f),
	.w3(32'h39af632a),
	.w4(32'hbb8140e7),
	.w5(32'h3ac370bb),
	.w6(32'h3a4a8b0a),
	.w7(32'h3a7714c3),
	.w8(32'hbb1927be),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8987ea),
	.w1(32'hbbf99681),
	.w2(32'h39a2fff0),
	.w3(32'hbbca1622),
	.w4(32'hbc0a3e39),
	.w5(32'h3c02b453),
	.w6(32'hbba9826e),
	.w7(32'hbb858d15),
	.w8(32'h3c75a198),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c284783),
	.w1(32'h3bee0f63),
	.w2(32'h3b130d78),
	.w3(32'hba5792b8),
	.w4(32'hbafac5d5),
	.w5(32'hbb71b8b3),
	.w6(32'hbb2fbc09),
	.w7(32'hbb28cbbf),
	.w8(32'hbb296a94),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2571fd),
	.w1(32'h3bd859f7),
	.w2(32'h3b4f4410),
	.w3(32'hba16728c),
	.w4(32'h39178a9f),
	.w5(32'hbb118925),
	.w6(32'h3b3cb82c),
	.w7(32'hbb07e618),
	.w8(32'h3a815617),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba414e88),
	.w1(32'h3a307449),
	.w2(32'h3bf0b114),
	.w3(32'hbab076ed),
	.w4(32'h39a78ad3),
	.w5(32'h3c19f74e),
	.w6(32'h3b829f72),
	.w7(32'h3b0e2d41),
	.w8(32'h3bc8eb93),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00d314),
	.w1(32'h384010fb),
	.w2(32'h3b146e24),
	.w3(32'hbb893056),
	.w4(32'hbb0c6800),
	.w5(32'h3a39fdb7),
	.w6(32'hba73d598),
	.w7(32'hbb1624e0),
	.w8(32'hbaa33ac6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb5729),
	.w1(32'hbabc428f),
	.w2(32'hbb4b9788),
	.w3(32'hbab054b9),
	.w4(32'hbb68da19),
	.w5(32'h3ac7f672),
	.w6(32'hb9d437a1),
	.w7(32'h3b6aa96a),
	.w8(32'h3b4a3400),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5228e),
	.w1(32'h3bf4ca95),
	.w2(32'h3ba0aee8),
	.w3(32'h3afe1cdc),
	.w4(32'h3b89d3de),
	.w5(32'h3aaaf88c),
	.w6(32'h3875d888),
	.w7(32'h3b5a5697),
	.w8(32'hbb9c910d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a215f),
	.w1(32'hb5cd63d8),
	.w2(32'hbbc591fe),
	.w3(32'hba9ff20e),
	.w4(32'hba14e464),
	.w5(32'hbc0bdc5a),
	.w6(32'h3a0a6194),
	.w7(32'hbba6f7fc),
	.w8(32'hbc0f18ac),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab33bb3),
	.w1(32'h3a9f47e1),
	.w2(32'h3a25a741),
	.w3(32'hbb97051d),
	.w4(32'h3b214fbc),
	.w5(32'hb921e608),
	.w6(32'hbb8fa464),
	.w7(32'h3a7fc4e4),
	.w8(32'hbb417354),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b4d8c),
	.w1(32'hbb9d3a6c),
	.w2(32'hbaf727f8),
	.w3(32'hbbc460ab),
	.w4(32'hbb5e36ed),
	.w5(32'hbb6745bd),
	.w6(32'hbba33f3a),
	.w7(32'hbb99d790),
	.w8(32'hbabc7eaa),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4651ee),
	.w1(32'hba0dff44),
	.w2(32'hbb52e71e),
	.w3(32'hba5ff8d8),
	.w4(32'hbc003800),
	.w5(32'hbb0cb7bf),
	.w6(32'h3bc168b5),
	.w7(32'h3bbab764),
	.w8(32'h3c739fe8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1182a),
	.w1(32'hba85a9ef),
	.w2(32'hbb6677c5),
	.w3(32'hbb656cca),
	.w4(32'hbb3c5f2c),
	.w5(32'hbbbc6e39),
	.w6(32'h3b058ab6),
	.w7(32'h39f60639),
	.w8(32'hb9cf119b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c5958),
	.w1(32'hbbbf7bd9),
	.w2(32'hbba0da32),
	.w3(32'hbba9f85f),
	.w4(32'hbb873967),
	.w5(32'hbadc3e21),
	.w6(32'h3b42e3bf),
	.w7(32'h3b85e7fd),
	.w8(32'hb9c51055),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33639e),
	.w1(32'h3b265c9c),
	.w2(32'hbb0f3d70),
	.w3(32'hbaca1a4c),
	.w4(32'h3ac7d47b),
	.w5(32'hbbb67700),
	.w6(32'hbb545563),
	.w7(32'h3a1517be),
	.w8(32'h39073392),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb393107),
	.w1(32'hbab90f22),
	.w2(32'h3c11398c),
	.w3(32'h3a8f56e4),
	.w4(32'h3b7e4867),
	.w5(32'h39f9b305),
	.w6(32'h3b9515d8),
	.w7(32'h3b57e839),
	.w8(32'hbb0202e9),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc173fea),
	.w1(32'h3b3460b4),
	.w2(32'h3a819f96),
	.w3(32'hbaea23a6),
	.w4(32'h3b43a56a),
	.w5(32'h3a9488f2),
	.w6(32'hbbb4686d),
	.w7(32'h3b299e7d),
	.w8(32'h3afa5b36),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398966ef),
	.w1(32'hbbb26b39),
	.w2(32'hbbaf964a),
	.w3(32'hbac1d569),
	.w4(32'hbbce962b),
	.w5(32'hb99495ef),
	.w6(32'h3ae6027a),
	.w7(32'hba95754e),
	.w8(32'hb96d6085),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44d9a0),
	.w1(32'hbb44a095),
	.w2(32'hbb167b9e),
	.w3(32'hbb9b9c5f),
	.w4(32'h3a2cff62),
	.w5(32'h39b8acb2),
	.w6(32'hbc0ab40d),
	.w7(32'h3b4ccc57),
	.w8(32'h3ac2a99d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a405a6d),
	.w1(32'h3bf2182e),
	.w2(32'h3bea9103),
	.w3(32'hbaea726a),
	.w4(32'h3af2c3b4),
	.w5(32'h3b9da1c6),
	.w6(32'hbac6499e),
	.w7(32'h3b21aa4d),
	.w8(32'h3b08de16),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0e1f2),
	.w1(32'hbb444c23),
	.w2(32'hbb7ae1c6),
	.w3(32'h3b05e426),
	.w4(32'hbb5956fe),
	.w5(32'hba9339b9),
	.w6(32'hbab1a456),
	.w7(32'hbb782bff),
	.w8(32'h3bd3c16f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c70cd4),
	.w1(32'hbb727e51),
	.w2(32'hbba3c1c5),
	.w3(32'h392bc474),
	.w4(32'hba675213),
	.w5(32'hbbaee595),
	.w6(32'h3b65933f),
	.w7(32'hbb45beed),
	.w8(32'hbb042783),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e78c7),
	.w1(32'hb95f4c8e),
	.w2(32'hbac53e4f),
	.w3(32'hba806e34),
	.w4(32'h3b32bf48),
	.w5(32'h39cae70a),
	.w6(32'h3b7f6c92),
	.w7(32'h3b090617),
	.w8(32'h39f3260e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb944208),
	.w1(32'h3ba644e8),
	.w2(32'h3baccd86),
	.w3(32'hbb3ff8be),
	.w4(32'hbb1295b0),
	.w5(32'h3b877660),
	.w6(32'h3b729236),
	.w7(32'hba35f601),
	.w8(32'h3b9dac8f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dc909),
	.w1(32'hbbac2a3f),
	.w2(32'hb9fc8949),
	.w3(32'h3b88a6bb),
	.w4(32'hbbfd9789),
	.w5(32'h3b929501),
	.w6(32'h3a5f0dad),
	.w7(32'h3a75d896),
	.w8(32'h3bc0f67f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef584b),
	.w1(32'h3aac9ebd),
	.w2(32'h3b3961c2),
	.w3(32'h3bc56280),
	.w4(32'h3b86638c),
	.w5(32'hbb1584ac),
	.w6(32'h3b0ac775),
	.w7(32'hbba201fe),
	.w8(32'hbb99bce0),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd39466),
	.w1(32'hbb8f42f6),
	.w2(32'h3ab050dc),
	.w3(32'hbb39f7f8),
	.w4(32'hbbb75a5d),
	.w5(32'h3bae2766),
	.w6(32'hbb65dc2f),
	.w7(32'hb938cfe8),
	.w8(32'h3c78bf86),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bf851),
	.w1(32'hbb574732),
	.w2(32'h3ad0c462),
	.w3(32'h39db6317),
	.w4(32'h3ad61566),
	.w5(32'hb98e23f5),
	.w6(32'hba3ef0f9),
	.w7(32'h3af131c5),
	.w8(32'hba964f3b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbb270),
	.w1(32'h38874035),
	.w2(32'hbb9a58cb),
	.w3(32'h39a74ff1),
	.w4(32'hbb806b3b),
	.w5(32'hb9d60e7c),
	.w6(32'hbb12c26b),
	.w7(32'hbb0b306b),
	.w8(32'h3b9bf3df),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dd449),
	.w1(32'h3bbaee33),
	.w2(32'hbb7f4109),
	.w3(32'hbaef6afb),
	.w4(32'hbaafe080),
	.w5(32'hbba6e8e1),
	.w6(32'hbac521ea),
	.w7(32'hbbd6c6fa),
	.w8(32'h3a7ba562),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c520308),
	.w1(32'h3b2ace91),
	.w2(32'h3b96917c),
	.w3(32'h3c129ef4),
	.w4(32'h3bac74b0),
	.w5(32'h3ac30cc2),
	.w6(32'h3b37e8df),
	.w7(32'hba3a47c4),
	.w8(32'hbb682aff),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3493a0),
	.w1(32'h39fbffb6),
	.w2(32'h3abffa91),
	.w3(32'h3b017c47),
	.w4(32'hbb9c3bce),
	.w5(32'h3bbb5074),
	.w6(32'h3a6d5bba),
	.w7(32'hbb14b712),
	.w8(32'h3bcf79b4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28ab01),
	.w1(32'hba641ca2),
	.w2(32'hba9ba7e7),
	.w3(32'hbac33f41),
	.w4(32'h3b0e86de),
	.w5(32'hbb18d77c),
	.w6(32'h3b4b2d95),
	.w7(32'h3b284112),
	.w8(32'hba2b4bdf),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebefa0),
	.w1(32'hbabb8c57),
	.w2(32'hbafe3558),
	.w3(32'hbb82a130),
	.w4(32'h3b0d186a),
	.w5(32'h3b62b610),
	.w6(32'hbbfb116e),
	.w7(32'h3b202a69),
	.w8(32'h3ad4b44a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf314fd),
	.w1(32'hbb85147b),
	.w2(32'h3c1fb630),
	.w3(32'h3adb927c),
	.w4(32'hbbc97143),
	.w5(32'h3bff116b),
	.w6(32'h3beefb98),
	.w7(32'h3b3afdb2),
	.w8(32'h3c122b35),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b80bd),
	.w1(32'hba991a7b),
	.w2(32'hba9ea1c0),
	.w3(32'hbaeeb98a),
	.w4(32'hbbef558a),
	.w5(32'hbabc9dff),
	.w6(32'h3b506ca9),
	.w7(32'hbbcf50b7),
	.w8(32'h3b2828fe),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b272a45),
	.w1(32'h3aa2bdcb),
	.w2(32'hb9cf966c),
	.w3(32'h3a94c887),
	.w4(32'hb93e50c8),
	.w5(32'hbb4f8d92),
	.w6(32'h3b570311),
	.w7(32'h3b70a450),
	.w8(32'h3a9a9f73),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c32e5),
	.w1(32'h3bcc634e),
	.w2(32'h3bacf617),
	.w3(32'hba89f3fb),
	.w4(32'h3c2b4d16),
	.w5(32'h39f5eef0),
	.w6(32'hbb477195),
	.w7(32'h3bc7f6ea),
	.w8(32'hbb8ecf0d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb1e1e),
	.w1(32'hbb4873a8),
	.w2(32'hba44ad63),
	.w3(32'hbb3eae88),
	.w4(32'hbb114c24),
	.w5(32'h3bd4c0a9),
	.w6(32'hba9af8e5),
	.w7(32'h3a898487),
	.w8(32'h3c381324),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becabe6),
	.w1(32'h3aabbf34),
	.w2(32'h3ac5bf0a),
	.w3(32'h3b50ecac),
	.w4(32'hbb8cb3ee),
	.w5(32'h3b812a98),
	.w6(32'h3a2ba70c),
	.w7(32'hbaa3a3cd),
	.w8(32'h3b0befc8),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ae506),
	.w1(32'hba94ce81),
	.w2(32'h3b953003),
	.w3(32'h3b84a9be),
	.w4(32'hbaa9f61f),
	.w5(32'hbb54bcaf),
	.w6(32'h3b5bb11d),
	.w7(32'h3ad8b901),
	.w8(32'hbacd6df5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d11c1),
	.w1(32'h3b45ef13),
	.w2(32'hba2f5cac),
	.w3(32'h39895895),
	.w4(32'h3b45a8f4),
	.w5(32'h3a77c00a),
	.w6(32'hba99344d),
	.w7(32'h3bd2175f),
	.w8(32'hbb2ee15d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9a6b8),
	.w1(32'hbac0889b),
	.w2(32'hb9a7115e),
	.w3(32'h3a91afb8),
	.w4(32'h3ad9fef1),
	.w5(32'hbb3297c0),
	.w6(32'hba95c3ba),
	.w7(32'h3b83e8d3),
	.w8(32'hba341c07),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81a3b8),
	.w1(32'hbaa6bbdc),
	.w2(32'hb938ba70),
	.w3(32'h39db0fd2),
	.w4(32'hbb06ee82),
	.w5(32'h3ba35d0e),
	.w6(32'h3ba6c884),
	.w7(32'hb850701f),
	.w8(32'h3c48e198),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2248e),
	.w1(32'hbbc13a8d),
	.w2(32'h395c752f),
	.w3(32'hbb4062c0),
	.w4(32'hbba9e0d6),
	.w5(32'hbb0ec2cc),
	.w6(32'hbb242a27),
	.w7(32'hba8db5a2),
	.w8(32'h3bd26696),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa14582),
	.w1(32'h3b45a549),
	.w2(32'h3ad13111),
	.w3(32'hbaee64d1),
	.w4(32'h3b32cc9e),
	.w5(32'h3a8e43a2),
	.w6(32'h3b934189),
	.w7(32'h39ea139b),
	.w8(32'h38ef47cd),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba950f37),
	.w1(32'hbac71173),
	.w2(32'hba85720d),
	.w3(32'h39638d0e),
	.w4(32'h3a872d97),
	.w5(32'hbbdca24d),
	.w6(32'h3b8a8404),
	.w7(32'hbb2d048e),
	.w8(32'hbbed2f3f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59fb7d),
	.w1(32'h3b11baa8),
	.w2(32'h3a10a620),
	.w3(32'h38f51cdc),
	.w4(32'hbb089a16),
	.w5(32'h3b858653),
	.w6(32'h3a6f29bd),
	.w7(32'h393fc4e4),
	.w8(32'h3ab91e72),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf708a5),
	.w1(32'hbbd12f66),
	.w2(32'hbb66eed3),
	.w3(32'hbba97332),
	.w4(32'hbb64e580),
	.w5(32'hbbfd9e70),
	.w6(32'hb9b38fa5),
	.w7(32'h3ade46b7),
	.w8(32'h3b816991),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb968f66),
	.w1(32'h3a24f620),
	.w2(32'h3b921c8f),
	.w3(32'hbc04a8ea),
	.w4(32'hbb033411),
	.w5(32'hbbb880fe),
	.w6(32'h3a763f05),
	.w7(32'hbb5ddb4f),
	.w8(32'hbb11b1c2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadc217),
	.w1(32'h3987f60d),
	.w2(32'hbac5c02f),
	.w3(32'hbb577af8),
	.w4(32'hb8db5643),
	.w5(32'hbbd45172),
	.w6(32'h3979dc3d),
	.w7(32'hbb89165f),
	.w8(32'hbad31494),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb174b12),
	.w1(32'hb9d6e241),
	.w2(32'hbae6dc01),
	.w3(32'hbb6c9771),
	.w4(32'hbbab0948),
	.w5(32'h3b449a94),
	.w6(32'h39f3304c),
	.w7(32'h39bee40e),
	.w8(32'h3bb0fa7e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99f972),
	.w1(32'hb961c22e),
	.w2(32'h39c22f28),
	.w3(32'h3b4c1132),
	.w4(32'h3a26fa0e),
	.w5(32'hba169b3a),
	.w6(32'hbb122059),
	.w7(32'h3b841f02),
	.w8(32'hbab98625),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafba572),
	.w1(32'h3a9abd4d),
	.w2(32'hba4f98d1),
	.w3(32'hba6d2cc5),
	.w4(32'hbab8dfed),
	.w5(32'h3a90b253),
	.w6(32'h3b1356dc),
	.w7(32'hba46a6b7),
	.w8(32'h3b8aa12b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9433ec),
	.w1(32'h3b8f1230),
	.w2(32'h3b9cb819),
	.w3(32'h3b35c12f),
	.w4(32'h3c106cb8),
	.w5(32'hbb51dafc),
	.w6(32'h3b0489e1),
	.w7(32'h3b15f0a8),
	.w8(32'hbc0917be),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08a296),
	.w1(32'hbc0b9776),
	.w2(32'hbb99c5e2),
	.w3(32'h3ac64739),
	.w4(32'hbb1b2a78),
	.w5(32'hbaf3a051),
	.w6(32'hbb88694a),
	.w7(32'hbb0e6502),
	.w8(32'hb9830858),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3e492),
	.w1(32'h3a920af7),
	.w2(32'h3be8b5d2),
	.w3(32'hbbb376dc),
	.w4(32'hbacd71c8),
	.w5(32'h39a1d6e4),
	.w6(32'h3bc1eb09),
	.w7(32'h3ba19769),
	.w8(32'h3bccaeec),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba843372),
	.w1(32'hba13b4df),
	.w2(32'hbba52dfd),
	.w3(32'h3b2a24c5),
	.w4(32'hbb8a5333),
	.w5(32'hbc13f78f),
	.w6(32'h3c0ac722),
	.w7(32'hbb5dae04),
	.w8(32'hbb8ed37b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24f927),
	.w1(32'h3bed3e79),
	.w2(32'hba3ce239),
	.w3(32'hbb6e0c02),
	.w4(32'hbc1bd0ac),
	.w5(32'hb90e9c1f),
	.w6(32'hba61e40f),
	.w7(32'h3b8ed65a),
	.w8(32'h3bc84057),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f181c),
	.w1(32'h3b0fa356),
	.w2(32'h3a90916f),
	.w3(32'h3a784aa7),
	.w4(32'hb9a7e95d),
	.w5(32'hbaf7b8ae),
	.w6(32'h3bb8187f),
	.w7(32'hba3fae9f),
	.w8(32'h3b0b51af),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cbf68),
	.w1(32'h3b17033f),
	.w2(32'h3c0346cd),
	.w3(32'hbb67d3a8),
	.w4(32'hbb0db9e3),
	.w5(32'hbb157595),
	.w6(32'h3a34a8cd),
	.w7(32'hbb27c2fb),
	.w8(32'h3a6e290d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9e262),
	.w1(32'h3b7270c7),
	.w2(32'hbc06ed61),
	.w3(32'hba4e109c),
	.w4(32'hbb839c81),
	.w5(32'hbaa165fc),
	.w6(32'hbbaecd33),
	.w7(32'h3c285763),
	.w8(32'h3bebb13f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d8d2f),
	.w1(32'h37a29808),
	.w2(32'hbb397a36),
	.w3(32'hbb79d36b),
	.w4(32'hbba5b589),
	.w5(32'h3afd7781),
	.w6(32'hbb898900),
	.w7(32'hbacbd892),
	.w8(32'hbb130820),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2f254),
	.w1(32'hbbfef119),
	.w2(32'h3a02eb0a),
	.w3(32'h398b593d),
	.w4(32'hbc7eca20),
	.w5(32'hbc7282ea),
	.w6(32'h3afe2360),
	.w7(32'hbae7b310),
	.w8(32'hb9840e02),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba839977),
	.w1(32'hbae05b23),
	.w2(32'h3b3c7ffb),
	.w3(32'hbc981446),
	.w4(32'hbb9698f3),
	.w5(32'h3babebad),
	.w6(32'hba65c6f4),
	.w7(32'hbab4aa64),
	.w8(32'hbb1ca08c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84bf94),
	.w1(32'hbabc33d1),
	.w2(32'hb9de9a4c),
	.w3(32'h3ada8bf5),
	.w4(32'h3af7601d),
	.w5(32'hbbd0c399),
	.w6(32'hba0b926b),
	.w7(32'h3c0a09d9),
	.w8(32'h3c3b17bb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b890d74),
	.w1(32'h3bcf0ed3),
	.w2(32'h3bdf94ee),
	.w3(32'hbadadc0a),
	.w4(32'hba6638d8),
	.w5(32'h3bb5b1c8),
	.w6(32'h3b430e5a),
	.w7(32'h3bcd1964),
	.w8(32'h3b83a224),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7f77f),
	.w1(32'hba48387b),
	.w2(32'h3bd940e7),
	.w3(32'h3b0b8f6a),
	.w4(32'hbafbf61b),
	.w5(32'hb97bd6a4),
	.w6(32'h3a380e07),
	.w7(32'h3b15f047),
	.w8(32'h3bd5f72b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8573cf),
	.w1(32'hbc6ef4c8),
	.w2(32'hbc04e3fd),
	.w3(32'h3b2cf0ba),
	.w4(32'h3b699934),
	.w5(32'hbbbb4639),
	.w6(32'h3a857202),
	.w7(32'hbc10cf35),
	.w8(32'h3bb9f6aa),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae50b35),
	.w1(32'h3bfaa173),
	.w2(32'h3c301481),
	.w3(32'hbc1832ac),
	.w4(32'hbb0d4a6b),
	.w5(32'hbbd3c970),
	.w6(32'h38b60194),
	.w7(32'hbaef110d),
	.w8(32'h39f2f046),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3fcf8),
	.w1(32'h39a9d591),
	.w2(32'h3be3cdb7),
	.w3(32'h3bbe4565),
	.w4(32'h3b3785d9),
	.w5(32'h3ab2f6eb),
	.w6(32'h3b5da045),
	.w7(32'h3aad4fc4),
	.w8(32'h3ae6fc14),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41207c),
	.w1(32'hbaa941c0),
	.w2(32'h39d8750e),
	.w3(32'h3b4a9110),
	.w4(32'h3a985557),
	.w5(32'h3b41857b),
	.w6(32'hb6ba88fa),
	.w7(32'h3b33030b),
	.w8(32'h3a6e1435),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96dbab),
	.w1(32'h3b15996e),
	.w2(32'h3a84a437),
	.w3(32'h3a6eb9c8),
	.w4(32'hbad4a7cc),
	.w5(32'hbb401117),
	.w6(32'h3ace70b6),
	.w7(32'hbc0ccde7),
	.w8(32'hbb33906c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ee8d5),
	.w1(32'h3b251b72),
	.w2(32'h3bce27af),
	.w3(32'h3c12104a),
	.w4(32'h38d797ca),
	.w5(32'h3aa22a9e),
	.w6(32'hbbd97ef5),
	.w7(32'hbae4fa05),
	.w8(32'hb9d71cd7),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cea60),
	.w1(32'hbb9143be),
	.w2(32'hbc4d1cba),
	.w3(32'hbb9d6966),
	.w4(32'h3b918710),
	.w5(32'hbb1f0578),
	.w6(32'hbabbfcb0),
	.w7(32'hbb20d5d7),
	.w8(32'hbc54b271),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ebc3a),
	.w1(32'h3ac1e2af),
	.w2(32'hbc496ab6),
	.w3(32'hbb86a4c3),
	.w4(32'h3a2385b2),
	.w5(32'h3c05ad0b),
	.w6(32'hbbf45b79),
	.w7(32'h3bd0849c),
	.w8(32'h3c19a809),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95f699),
	.w1(32'hbabc95d8),
	.w2(32'hbc1fd8c0),
	.w3(32'hbba4c577),
	.w4(32'h3af9e9c4),
	.w5(32'h3cbc71d0),
	.w6(32'h3afc286e),
	.w7(32'hba84ac7e),
	.w8(32'hbb13b8bb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9b16a),
	.w1(32'h3abf0621),
	.w2(32'hb91ee5b6),
	.w3(32'hbadf9531),
	.w4(32'hbb24bf7f),
	.w5(32'hbbf2f242),
	.w6(32'hbb9a26fe),
	.w7(32'h3be959ed),
	.w8(32'h3c8d7662),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba273dcb),
	.w1(32'hbb91c8f1),
	.w2(32'h39c4c1d1),
	.w3(32'hbbde902c),
	.w4(32'hba809b11),
	.w5(32'hb99378bd),
	.w6(32'h3a6633a1),
	.w7(32'h3c11390f),
	.w8(32'h3b74f8e3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f7c43),
	.w1(32'hbc41136e),
	.w2(32'hbab80862),
	.w3(32'h3b213733),
	.w4(32'hbbbf7f6c),
	.w5(32'hbb9385ba),
	.w6(32'hbbcc5cb1),
	.w7(32'hbbed7e15),
	.w8(32'hbb0e5b9e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd38ed5),
	.w1(32'h3a8750f8),
	.w2(32'hbc1fd650),
	.w3(32'h372550e1),
	.w4(32'h3c907b86),
	.w5(32'h3d613e51),
	.w6(32'hbbc5607a),
	.w7(32'h3b9d9316),
	.w8(32'h3b654062),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbde86),
	.w1(32'h3a8322cd),
	.w2(32'h3b2454bd),
	.w3(32'h3cc56e12),
	.w4(32'hb9bcb398),
	.w5(32'h3b1b2836),
	.w6(32'h3bb27095),
	.w7(32'hbb575a35),
	.w8(32'hba846fdd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf0fa5),
	.w1(32'h3a4869de),
	.w2(32'h3b781b15),
	.w3(32'hbb053671),
	.w4(32'h3b3eaaa9),
	.w5(32'h3a248174),
	.w6(32'hbb09d2a6),
	.w7(32'h3ba57523),
	.w8(32'hba985a6b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb800594),
	.w1(32'hbb6d15d9),
	.w2(32'hbb5c80fb),
	.w3(32'h3b970579),
	.w4(32'h3c0620b5),
	.w5(32'h3c886c22),
	.w6(32'hbb9a4a38),
	.w7(32'h3b70c426),
	.w8(32'h3c410e5d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5ae72),
	.w1(32'hbb127ee2),
	.w2(32'hbbdf703d),
	.w3(32'hbbc33b4a),
	.w4(32'h39a13ca4),
	.w5(32'hbbd47c94),
	.w6(32'h3b90a098),
	.w7(32'hba3fb95c),
	.w8(32'hbb9f0cb9),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ff2de),
	.w1(32'hbad19053),
	.w2(32'hbc2163ee),
	.w3(32'hbb60c72b),
	.w4(32'h3b94efc2),
	.w5(32'h3af66347),
	.w6(32'hba0ce0c0),
	.w7(32'h3b27cf1a),
	.w8(32'h3ae480ce),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb3c3a),
	.w1(32'h3b59719e),
	.w2(32'h3b850e81),
	.w3(32'h3ad227d5),
	.w4(32'hbb93a7a1),
	.w5(32'hbbba452f),
	.w6(32'h3b921d42),
	.w7(32'h3bf00d9f),
	.w8(32'h39df1119),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38267558),
	.w1(32'hbb201050),
	.w2(32'h3b69e493),
	.w3(32'hbb393c05),
	.w4(32'hbba984ec),
	.w5(32'hbbf5db7e),
	.w6(32'hbb22fda9),
	.w7(32'h3bf1115b),
	.w8(32'h3be62a3e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e0f44),
	.w1(32'h3b03970a),
	.w2(32'h3c400bd4),
	.w3(32'h3b6e2b70),
	.w4(32'hbbac18b2),
	.w5(32'hbc03d68e),
	.w6(32'h3ba1742c),
	.w7(32'hb88e7582),
	.w8(32'h3a7373c8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde453c),
	.w1(32'h39e7ed49),
	.w2(32'hbb0df8d5),
	.w3(32'hba8e4d18),
	.w4(32'h3b57aa97),
	.w5(32'h3b295ec5),
	.w6(32'hbc1ce20a),
	.w7(32'h3be06ae1),
	.w8(32'h3c2d1b7d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ddc95),
	.w1(32'hbbc4293a),
	.w2(32'hbba9ef64),
	.w3(32'hbbf90cd4),
	.w4(32'hbb49c389),
	.w5(32'hbb0d5c7c),
	.w6(32'h3ba050ea),
	.w7(32'hbafa6379),
	.w8(32'h3b1182f9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1c102),
	.w1(32'h3aff888a),
	.w2(32'h3b1c41f7),
	.w3(32'h3b710e99),
	.w4(32'h3b10109f),
	.w5(32'h3bf85a1b),
	.w6(32'hbb0e4da3),
	.w7(32'h3b56a91d),
	.w8(32'h3b9d2941),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af08152),
	.w1(32'h3b1a0e6e),
	.w2(32'h3b0cef91),
	.w3(32'hba139860),
	.w4(32'h3b3a643e),
	.w5(32'h3b976a6e),
	.w6(32'h3b1fcd3c),
	.w7(32'hbb097dc2),
	.w8(32'h3bbca50d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb40d99),
	.w1(32'hba383322),
	.w2(32'hbb2bea73),
	.w3(32'h3ba6daff),
	.w4(32'h3aae28aa),
	.w5(32'hba885b24),
	.w6(32'h3ba78f41),
	.w7(32'hbb9f50e5),
	.w8(32'h3bc61081),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a6f11),
	.w1(32'hbadb4eb0),
	.w2(32'h388da96c),
	.w3(32'hbb83f0df),
	.w4(32'h3ac5af19),
	.w5(32'h3bb5b62a),
	.w6(32'h3bb2664e),
	.w7(32'h3bf4eb36),
	.w8(32'h3c3012b2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4446dd),
	.w1(32'h3b34e781),
	.w2(32'h3b9ca0f7),
	.w3(32'h3b992e4a),
	.w4(32'h3bbc99b4),
	.w5(32'h3b115c74),
	.w6(32'h3a917acb),
	.w7(32'hba1874ae),
	.w8(32'hbb3e1b7e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04f627),
	.w1(32'h3c6277b4),
	.w2(32'hba47c605),
	.w3(32'h3bd8d7e3),
	.w4(32'h38d7bda6),
	.w5(32'hbb093298),
	.w6(32'h3af92903),
	.w7(32'hbbe08f1d),
	.w8(32'hbbe40744),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fd2ff),
	.w1(32'hbb3548a8),
	.w2(32'h3bb4bd4f),
	.w3(32'h3bcc09e9),
	.w4(32'hbb44beb2),
	.w5(32'hbbc77179),
	.w6(32'h3b92e8ba),
	.w7(32'h3ae174e6),
	.w8(32'h3b5d878f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e32c6),
	.w1(32'hbc0c13d6),
	.w2(32'hbc1d0c3c),
	.w3(32'hbb3d6ad1),
	.w4(32'h3b1d6aef),
	.w5(32'h3cc7e884),
	.w6(32'h3957203a),
	.w7(32'h3ba20d25),
	.w8(32'h3c20575c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f2944),
	.w1(32'hbbb14013),
	.w2(32'h3a2b2906),
	.w3(32'h399c4e0b),
	.w4(32'h3c167789),
	.w5(32'h3c105281),
	.w6(32'h3b6168bc),
	.w7(32'h3b41a4a5),
	.w8(32'hbb1ff73f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4deb18),
	.w1(32'hbb68f6bc),
	.w2(32'hbbf24cef),
	.w3(32'h3c363296),
	.w4(32'hbc030586),
	.w5(32'hbbe6ec66),
	.w6(32'hbb42641c),
	.w7(32'hba0c2147),
	.w8(32'hbbe05672),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b280a),
	.w1(32'hbb59d885),
	.w2(32'hbbcc5180),
	.w3(32'hbb816329),
	.w4(32'hbbc26761),
	.w5(32'hb99a6e1c),
	.w6(32'h3b3e98a6),
	.w7(32'h3ae7978a),
	.w8(32'hbaead0c2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80aa31),
	.w1(32'hba993be6),
	.w2(32'hbb33c9ec),
	.w3(32'h3b816d45),
	.w4(32'h3b58a043),
	.w5(32'h3c07e7c8),
	.w6(32'h3bb61a9e),
	.w7(32'h3b043a4c),
	.w8(32'h3b31ce7b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf59291),
	.w1(32'h3bed6701),
	.w2(32'h3b5aabf9),
	.w3(32'h3c0ba22d),
	.w4(32'h3b932e0f),
	.w5(32'h3c1cca26),
	.w6(32'h3b64d9f6),
	.w7(32'h3a68ca43),
	.w8(32'h3b4e0caf),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9ba3f),
	.w1(32'h3c0e3e51),
	.w2(32'h3ba05317),
	.w3(32'h3aa44748),
	.w4(32'hb9ffb9bb),
	.w5(32'hb9926987),
	.w6(32'h3c04d5f4),
	.w7(32'h3abd36cf),
	.w8(32'h3c129606),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae17bdd),
	.w1(32'h3b763660),
	.w2(32'hba804a0b),
	.w3(32'h3aac4a84),
	.w4(32'h3ba29255),
	.w5(32'h3c0f04b9),
	.w6(32'h3b43c7e2),
	.w7(32'h3ad0f37a),
	.w8(32'h3b6d964d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f176b),
	.w1(32'h3b4d65f8),
	.w2(32'h3b9db132),
	.w3(32'h3b1a426b),
	.w4(32'hba17d4be),
	.w5(32'hbc474d8c),
	.w6(32'h3ad858d0),
	.w7(32'h3bbd1f60),
	.w8(32'hbb0d461b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c23cd),
	.w1(32'h3bb3e355),
	.w2(32'hbb53ba9f),
	.w3(32'h3a78593d),
	.w4(32'h3b2a2da9),
	.w5(32'h3c4d3a85),
	.w6(32'h3b1479d0),
	.w7(32'hbb29e248),
	.w8(32'h3adbbf98),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe549e1),
	.w1(32'h3aab87d7),
	.w2(32'hbb80fd34),
	.w3(32'h3b211b56),
	.w4(32'hbbf711e6),
	.w5(32'hba953fdd),
	.w6(32'h3b508270),
	.w7(32'hbb52bf9e),
	.w8(32'hbbb2d024),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae06c96),
	.w1(32'hbb003b7b),
	.w2(32'h3af6db13),
	.w3(32'hbb91aa93),
	.w4(32'h39dafc8f),
	.w5(32'hbb9ceef6),
	.w6(32'h3a027be7),
	.w7(32'h3aea1000),
	.w8(32'h3b438a06),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e26b2),
	.w1(32'hbc10e6da),
	.w2(32'h3bbba0c3),
	.w3(32'hbb529dd8),
	.w4(32'hbb6b2bce),
	.w5(32'hbbff2ced),
	.w6(32'hbb323418),
	.w7(32'hbaaecdd8),
	.w8(32'h3b44649d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb67e5),
	.w1(32'hba41ff71),
	.w2(32'hbb596674),
	.w3(32'h3af68929),
	.w4(32'h3bfe2f31),
	.w5(32'h3c238e94),
	.w6(32'h3b0e1b6b),
	.w7(32'h3c02b9cd),
	.w8(32'h3be01006),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc378c1c),
	.w1(32'hbad9ff98),
	.w2(32'hb938444c),
	.w3(32'h3abe9c75),
	.w4(32'hbb7ea059),
	.w5(32'hbbb953f2),
	.w6(32'h3b819536),
	.w7(32'hbb20505a),
	.w8(32'h3ad03ff9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb981bfb),
	.w1(32'h3ac8f300),
	.w2(32'h3c7311d6),
	.w3(32'h3b9d3ab6),
	.w4(32'hbbdb0c97),
	.w5(32'h3b8916b5),
	.w6(32'h3a357250),
	.w7(32'h3a8dece5),
	.w8(32'h3b5149cd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19c1d6),
	.w1(32'h39c99522),
	.w2(32'h3b6b4568),
	.w3(32'h3b0d8642),
	.w4(32'h3bb69a8f),
	.w5(32'h3b3e997b),
	.w6(32'hbb6860ba),
	.w7(32'hb9d9fc50),
	.w8(32'hbb2f1315),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93e4cb),
	.w1(32'hbc0aba14),
	.w2(32'hbb8e1c90),
	.w3(32'h3a4f6e93),
	.w4(32'hbb0b0ca3),
	.w5(32'h3b7be8d2),
	.w6(32'h3b0756f4),
	.w7(32'hbb9d322f),
	.w8(32'hbb3d48e5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f2afa),
	.w1(32'hbabd6217),
	.w2(32'hbb3ae748),
	.w3(32'h39209c56),
	.w4(32'hbb6e7721),
	.w5(32'hb9bb69b5),
	.w6(32'h3aeb327d),
	.w7(32'h3b9567a5),
	.w8(32'h3b71af8f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe61a5b),
	.w1(32'h3aad3cf7),
	.w2(32'h3ba55a49),
	.w3(32'hbbc4777c),
	.w4(32'hba8b0d93),
	.w5(32'hbbc5a010),
	.w6(32'hbb435eca),
	.w7(32'h3bfbc14d),
	.w8(32'h3bfebf9c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cff2e),
	.w1(32'hbb31146e),
	.w2(32'hbbae5ce3),
	.w3(32'h3a8b5e06),
	.w4(32'hba86bf6e),
	.w5(32'hbb8c1874),
	.w6(32'h3795a780),
	.w7(32'hbabafe96),
	.w8(32'hbbeaf508),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f2f92),
	.w1(32'h3a3af9c2),
	.w2(32'hbb73db82),
	.w3(32'hbb3c4bc8),
	.w4(32'h3bf06a45),
	.w5(32'h3c9c53c7),
	.w6(32'h38292ce8),
	.w7(32'h3b643cee),
	.w8(32'h3c286426),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3b65a),
	.w1(32'hbc033b02),
	.w2(32'h3a6a173c),
	.w3(32'h3c2bb366),
	.w4(32'h3b239eb6),
	.w5(32'hbb990d26),
	.w6(32'h3b5aea7d),
	.w7(32'h3baf6914),
	.w8(32'h3b9b1b76),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76a5ad),
	.w1(32'hba1986c0),
	.w2(32'h3a9e2751),
	.w3(32'hbb910d92),
	.w4(32'hbae93c31),
	.w5(32'hbb8eb3d0),
	.w6(32'hba624bff),
	.w7(32'h3a172189),
	.w8(32'h3a52a1cd),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c84df),
	.w1(32'h3a970af7),
	.w2(32'h3bedf0fe),
	.w3(32'h3ab1c295),
	.w4(32'hbb6a9e63),
	.w5(32'hbbec4bd4),
	.w6(32'h3a2f2290),
	.w7(32'h3b5ef9be),
	.w8(32'hbb8e339e),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5353af),
	.w1(32'h3bcdf2ae),
	.w2(32'h3bbc0848),
	.w3(32'h3a380136),
	.w4(32'hbb3e4b08),
	.w5(32'h3af435b0),
	.w6(32'h3bb1216d),
	.w7(32'hbba8e690),
	.w8(32'hbbc5b284),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c4694),
	.w1(32'h3bcbbfad),
	.w2(32'h3ba5479c),
	.w3(32'hbb5af886),
	.w4(32'h3c36ea5e),
	.w5(32'hbab05d63),
	.w6(32'hbb9d478c),
	.w7(32'h3b3e8225),
	.w8(32'hbb501fad),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba585aa9),
	.w1(32'hbb7d0523),
	.w2(32'hbb85bfa9),
	.w3(32'h3c2439c1),
	.w4(32'hbb42b5df),
	.w5(32'hbc0c4efb),
	.w6(32'hb86f8b9c),
	.w7(32'hbbc3bb39),
	.w8(32'hb91dfb00),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6102d),
	.w1(32'hbb00be4f),
	.w2(32'h3b270925),
	.w3(32'hbbbee59d),
	.w4(32'h3a53f096),
	.w5(32'hb9b4ffb4),
	.w6(32'h3adc98fc),
	.w7(32'h3b76f803),
	.w8(32'h3b905e5c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1738c),
	.w1(32'hbba0881a),
	.w2(32'hbb623bd5),
	.w3(32'hbb60e0f8),
	.w4(32'hbb201232),
	.w5(32'hbb79802d),
	.w6(32'h3be6848d),
	.w7(32'h3b8593b6),
	.w8(32'h376d3ff4),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4de5d9),
	.w1(32'hbbee54b8),
	.w2(32'hbb95483d),
	.w3(32'hbc15960b),
	.w4(32'hbb124263),
	.w5(32'hbb6363a4),
	.w6(32'hbb3c18ef),
	.w7(32'hbb7267d6),
	.w8(32'h3a9ff2f7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ac4b6),
	.w1(32'hbaa5897c),
	.w2(32'hbab56b5c),
	.w3(32'hbbd92ec1),
	.w4(32'h3ad290df),
	.w5(32'hbb99ac57),
	.w6(32'hbab119d2),
	.w7(32'hb9bdd5ad),
	.w8(32'h3b42d917),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73ce34),
	.w1(32'hba36f0ec),
	.w2(32'hbc2a62a6),
	.w3(32'hbb5efd35),
	.w4(32'h3bbc76db),
	.w5(32'h3c4ae398),
	.w6(32'hbb56d9e4),
	.w7(32'h3ae00083),
	.w8(32'h3c097406),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ad360),
	.w1(32'h3b7f60a5),
	.w2(32'h3c1d97e4),
	.w3(32'hba595e40),
	.w4(32'h3a5165aa),
	.w5(32'h3ba0bba1),
	.w6(32'h3b9dd0af),
	.w7(32'h3bcfe00b),
	.w8(32'h3a2577d7),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c7985),
	.w1(32'hbafc047a),
	.w2(32'hba3fa245),
	.w3(32'h3b8c8d5e),
	.w4(32'hbaac63ba),
	.w5(32'hbb8cb0d4),
	.w6(32'hba61c026),
	.w7(32'hbb70411d),
	.w8(32'h3a27fac9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0c974),
	.w1(32'h3b9be68a),
	.w2(32'h3c35357e),
	.w3(32'hbbd8f6b5),
	.w4(32'hbb9d5601),
	.w5(32'h3a9402d4),
	.w6(32'hbbc17e3a),
	.w7(32'hbbd538e0),
	.w8(32'hbb8cb925),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf99620),
	.w1(32'hbb9f8974),
	.w2(32'hbb15af56),
	.w3(32'h3b46948c),
	.w4(32'h3b9967e2),
	.w5(32'hbba40925),
	.w6(32'hbbbefafa),
	.w7(32'h3ae43668),
	.w8(32'h3aa52bde),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb834ada),
	.w1(32'h3ad815e5),
	.w2(32'hba36d1c4),
	.w3(32'hbbdf605c),
	.w4(32'h3a999941),
	.w5(32'hbbcb94bc),
	.w6(32'hbb8a8100),
	.w7(32'hbb37d525),
	.w8(32'hba3a4468),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb882f83),
	.w1(32'hbbd58d8c),
	.w2(32'h3c038769),
	.w3(32'hbb267286),
	.w4(32'h3a3784e7),
	.w5(32'hbc16c7e3),
	.w6(32'hba0765a2),
	.w7(32'h3b9c3004),
	.w8(32'h3b7fc746),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81cc23),
	.w1(32'h3b9c4091),
	.w2(32'h3b49be8a),
	.w3(32'hbbfed9bf),
	.w4(32'h3b9f2f3a),
	.w5(32'h3b716345),
	.w6(32'hbbf83d01),
	.w7(32'hbb05acf5),
	.w8(32'hbc251d44),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3575c2),
	.w1(32'h3b986e03),
	.w2(32'h3c079047),
	.w3(32'hb96ed5a9),
	.w4(32'h3bce5ece),
	.w5(32'hbb4dee52),
	.w6(32'hbb9515b7),
	.w7(32'h3ba20a77),
	.w8(32'h3bd525dd),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53c838),
	.w1(32'h3afc0bc2),
	.w2(32'h3c7a96a0),
	.w3(32'hbad57867),
	.w4(32'hbb8a415f),
	.w5(32'hbc34233a),
	.w6(32'h3b334f87),
	.w7(32'hb8fa09ce),
	.w8(32'h3c24de2c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5a2a2),
	.w1(32'hbab79012),
	.w2(32'hbaad6339),
	.w3(32'hbaf8ca7a),
	.w4(32'hbbca86fe),
	.w5(32'hbc1a2c08),
	.w6(32'h3b90f1fa),
	.w7(32'hbb25dd30),
	.w8(32'hbb9e9c94),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc634e8f),
	.w1(32'hbbb8136c),
	.w2(32'hbc0f8955),
	.w3(32'hbc981e27),
	.w4(32'hbb38cc79),
	.w5(32'h3bceebdd),
	.w6(32'hbc7be4a6),
	.w7(32'hbb4616f0),
	.w8(32'h3ab41482),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb69d2f),
	.w1(32'h3bdfc20e),
	.w2(32'h3c549e85),
	.w3(32'hbbd30556),
	.w4(32'hbb0b08c5),
	.w5(32'hbb8d1694),
	.w6(32'hbbf8405c),
	.w7(32'h3b42cc2e),
	.w8(32'hbbb4bd54),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e8400),
	.w1(32'h3a070591),
	.w2(32'hbba7caad),
	.w3(32'h3c5786e6),
	.w4(32'h3a7ebc39),
	.w5(32'hbb7de8b6),
	.w6(32'h3b58a6e0),
	.w7(32'hbacd5ff6),
	.w8(32'hb9054d3c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3d112),
	.w1(32'h3ab46a1f),
	.w2(32'hbb10e134),
	.w3(32'hbc0c49b9),
	.w4(32'hba507a02),
	.w5(32'hbbacd04b),
	.w6(32'hba5f0351),
	.w7(32'h39937e3f),
	.w8(32'hbb28b1b7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a321c),
	.w1(32'h3beb063a),
	.w2(32'h3c6bcd46),
	.w3(32'hbaa9c78b),
	.w4(32'hbb385192),
	.w5(32'hbbf9efa9),
	.w6(32'hbb20446f),
	.w7(32'hbb1893ec),
	.w8(32'hbb168a9d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0afe3),
	.w1(32'hbb9d7ede),
	.w2(32'hbafd304e),
	.w3(32'hbbb4052e),
	.w4(32'hbb46e7d3),
	.w5(32'hbba73dc0),
	.w6(32'h3b10e90a),
	.w7(32'hbb975c53),
	.w8(32'hbba10582),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7861c5),
	.w1(32'h3c22d3e5),
	.w2(32'h3c72ed37),
	.w3(32'hb983f01f),
	.w4(32'hba98e2be),
	.w5(32'hbbdeef74),
	.w6(32'hbb896bf3),
	.w7(32'h3b94044c),
	.w8(32'h3b1bcfcd),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1faa20),
	.w1(32'hbb181765),
	.w2(32'hbb511df1),
	.w3(32'hbbb19eed),
	.w4(32'hb9ea0bd1),
	.w5(32'hba22c726),
	.w6(32'h3a80613e),
	.w7(32'h3b7a9269),
	.w8(32'h392565b3),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b225e),
	.w1(32'hbb20f16a),
	.w2(32'hbb715283),
	.w3(32'hbb475c9d),
	.w4(32'hbc2b9901),
	.w5(32'hbc01a8b9),
	.w6(32'hbb356c34),
	.w7(32'h3c0317e3),
	.w8(32'h3acb48c0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8728b9),
	.w1(32'h3bc8ef2e),
	.w2(32'h3c53df37),
	.w3(32'hbc1a409d),
	.w4(32'hbb6f5877),
	.w5(32'hbb1fe165),
	.w6(32'hbb5b6803),
	.w7(32'h3bdadfd3),
	.w8(32'h3c2a3365),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd76ba0),
	.w1(32'h3bacd267),
	.w2(32'h3b051d5d),
	.w3(32'h3b50bba2),
	.w4(32'h3bbc4204),
	.w5(32'hbb4e427d),
	.w6(32'h3b98689f),
	.w7(32'h3bebafd7),
	.w8(32'h3b0125a2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bea14),
	.w1(32'hb988434c),
	.w2(32'h3a7fdefd),
	.w3(32'h3c1f7ae1),
	.w4(32'h3b11a3c9),
	.w5(32'h3b02860a),
	.w6(32'hbbcac2c1),
	.w7(32'hba27f888),
	.w8(32'h3b25ca63),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f4abb),
	.w1(32'hbaca8ada),
	.w2(32'hba402594),
	.w3(32'h3a6d5f0b),
	.w4(32'h3bd7077c),
	.w5(32'h3afa4652),
	.w6(32'h3b3ac1a2),
	.w7(32'h3c234888),
	.w8(32'hb6ae58d8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8f9b1),
	.w1(32'hbbdfd44d),
	.w2(32'hbabf2c12),
	.w3(32'hbb465db7),
	.w4(32'hbb9c944c),
	.w5(32'h3ad87f5c),
	.w6(32'hba9061c9),
	.w7(32'h39cd914a),
	.w8(32'h3b58ef87),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a505e04),
	.w1(32'h3b0b4eff),
	.w2(32'hbb95332d),
	.w3(32'hbaec6561),
	.w4(32'h3c2a3a5b),
	.w5(32'h3c1d5951),
	.w6(32'h3b285715),
	.w7(32'h3b597ba6),
	.w8(32'h3b4f7dbd),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2efa69),
	.w1(32'h3a470bd6),
	.w2(32'h3b66faed),
	.w3(32'h3c304756),
	.w4(32'hbacce92e),
	.w5(32'h3b2eeff2),
	.w6(32'h3bdf93c7),
	.w7(32'hbaccc5ff),
	.w8(32'h3b326871),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb873f76),
	.w1(32'h39f6c0a4),
	.w2(32'h3ae76e89),
	.w3(32'hb9ee227a),
	.w4(32'hbb8fe855),
	.w5(32'hbbc4943f),
	.w6(32'h3bc5ae39),
	.w7(32'h3b8c1251),
	.w8(32'h3c14d7f0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a2859),
	.w1(32'hbbcb2fca),
	.w2(32'hbbbcb5bc),
	.w3(32'hbb30d804),
	.w4(32'h3b28c8ec),
	.w5(32'hb9ba37b9),
	.w6(32'h3b3ca689),
	.w7(32'h3b57bb73),
	.w8(32'hbb4bb05a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be2d9),
	.w1(32'h39be584f),
	.w2(32'h3b4c20ac),
	.w3(32'hb6f6251c),
	.w4(32'h3bcfd5d1),
	.w5(32'hbb2f3e2f),
	.w6(32'hbaf59840),
	.w7(32'h3bc3c680),
	.w8(32'h3ab5d98c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390460e6),
	.w1(32'h3a9171a3),
	.w2(32'h3b355ee7),
	.w3(32'hbb310b60),
	.w4(32'hba0f1d71),
	.w5(32'hbbf426e3),
	.w6(32'hba498b51),
	.w7(32'h3b624c85),
	.w8(32'hbb8b82a0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e03ad),
	.w1(32'h3ba23307),
	.w2(32'h3b573595),
	.w3(32'h39f00196),
	.w4(32'hb9160d4a),
	.w5(32'hbbf3b893),
	.w6(32'hbbc43926),
	.w7(32'h3b9ad4b5),
	.w8(32'h3b797ab8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8980ed3),
	.w1(32'hba403ee2),
	.w2(32'hb94764ed),
	.w3(32'hbb4cf784),
	.w4(32'h3b33dcb4),
	.w5(32'h3bc668bd),
	.w6(32'hbadb2cce),
	.w7(32'hb8d01a34),
	.w8(32'h3b00da71),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6de561),
	.w1(32'h3b8731de),
	.w2(32'hbbb7d8aa),
	.w3(32'h3a799fae),
	.w4(32'h3bded55a),
	.w5(32'h3ccba046),
	.w6(32'h3b08a501),
	.w7(32'h3a9ae871),
	.w8(32'h3aa680d6),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc117354),
	.w1(32'h3a32b11b),
	.w2(32'hbbfa4dee),
	.w3(32'h3c028bcf),
	.w4(32'h37d62942),
	.w5(32'hbb9ea9ae),
	.w6(32'h3b4b03d5),
	.w7(32'hba06a44e),
	.w8(32'hba2f57a6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f09520),
	.w1(32'h3b55b337),
	.w2(32'h3ad82ea2),
	.w3(32'h3b8e085f),
	.w4(32'h3a1dfd54),
	.w5(32'h39ae511f),
	.w6(32'h3ba8c5b5),
	.w7(32'hba6f83b5),
	.w8(32'h3ba1a7b7),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74adcb),
	.w1(32'h3bafcd87),
	.w2(32'hbb0b3f08),
	.w3(32'h3b861fbe),
	.w4(32'hbac6d10d),
	.w5(32'hba4bda1c),
	.w6(32'h3abaa599),
	.w7(32'hbb095b37),
	.w8(32'hbb4d6edb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1d52a),
	.w1(32'h3b33d47b),
	.w2(32'h3ae4a1bb),
	.w3(32'h3bc0864c),
	.w4(32'hbabdec93),
	.w5(32'hbbcfdfbb),
	.w6(32'hba3db142),
	.w7(32'h3aee1dc7),
	.w8(32'hbbd1cd23),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade6eed),
	.w1(32'hbb5cd7cd),
	.w2(32'hbb95d086),
	.w3(32'hbb3b72ed),
	.w4(32'hb9f2fb7c),
	.w5(32'h3b88f9a8),
	.w6(32'h3be48a3e),
	.w7(32'hbaa1fc78),
	.w8(32'hba122856),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb774b29e),
	.w1(32'h3b946fe0),
	.w2(32'h3bc504e6),
	.w3(32'hbbb5d8b7),
	.w4(32'hbb5a810a),
	.w5(32'h3af31645),
	.w6(32'h3b81af1d),
	.w7(32'h3b89df14),
	.w8(32'h3b8ea8a6),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18ae3e),
	.w1(32'h3bb5a1b8),
	.w2(32'h3a32614a),
	.w3(32'h3ba396b4),
	.w4(32'h3bdaba34),
	.w5(32'h3c3fb101),
	.w6(32'h3ba4395d),
	.w7(32'h3a729bc4),
	.w8(32'hba8fbe3a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f34ff),
	.w1(32'hba9c9005),
	.w2(32'h3a716eec),
	.w3(32'h3bc532a6),
	.w4(32'h3b03c6d5),
	.w5(32'h3b7d554b),
	.w6(32'hbc36594f),
	.w7(32'h3b9407b1),
	.w8(32'h3c2d2b74),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2680b4),
	.w1(32'hbb62fad2),
	.w2(32'h39bf451d),
	.w3(32'h3977a03c),
	.w4(32'hbb25d8ec),
	.w5(32'hba757e98),
	.w6(32'h3b605d34),
	.w7(32'h3b3daf67),
	.w8(32'h3c213727),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b902215),
	.w1(32'h39d84c2f),
	.w2(32'h3b40174d),
	.w3(32'hbb06f8d3),
	.w4(32'h3b19a420),
	.w5(32'h3b5b0a49),
	.w6(32'h3a30b810),
	.w7(32'h3bc059f7),
	.w8(32'h3bd1bcc0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac49d4f),
	.w1(32'h3b2d6859),
	.w2(32'h3b753556),
	.w3(32'h3b9cea68),
	.w4(32'hba8dbdc9),
	.w5(32'hbbd29d7d),
	.w6(32'h3b0003ac),
	.w7(32'h3c032a15),
	.w8(32'hbb21afb9),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11b0e6),
	.w1(32'hbbeb4cb8),
	.w2(32'hbbb5e2b0),
	.w3(32'hbbb62782),
	.w4(32'hbb8869e7),
	.w5(32'hbc25ed73),
	.w6(32'h3accbad5),
	.w7(32'hba69a6a0),
	.w8(32'hbae05f6d),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaf91a),
	.w1(32'h3c06462d),
	.w2(32'hbc477705),
	.w3(32'hbb85ccd9),
	.w4(32'h3a77ffa6),
	.w5(32'h3d3541bd),
	.w6(32'h39a648e2),
	.w7(32'hba012acb),
	.w8(32'hb9b3f268),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc543bcc),
	.w1(32'h3b951a5d),
	.w2(32'hbc0cc64d),
	.w3(32'h3c23f2ad),
	.w4(32'h3c07bb07),
	.w5(32'h3cabe242),
	.w6(32'h3c656a2f),
	.w7(32'h3bed26fb),
	.w8(32'hbb966821),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cda4a),
	.w1(32'hbae3d339),
	.w2(32'h3b7c161b),
	.w3(32'h3c8082e4),
	.w4(32'hbbe16081),
	.w5(32'hbbd6c021),
	.w6(32'h3b8f3363),
	.w7(32'h3acfc16b),
	.w8(32'hbb66a478),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39cbba),
	.w1(32'hbbe8941b),
	.w2(32'hbb9dee29),
	.w3(32'hba68cc78),
	.w4(32'h3bce7464),
	.w5(32'hbb48eeec),
	.w6(32'hbb8aa68c),
	.w7(32'h3b8b9532),
	.w8(32'hbac0cbbe),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf62c89),
	.w1(32'h3b694238),
	.w2(32'h3b628c61),
	.w3(32'hbbaa9895),
	.w4(32'hba3ec255),
	.w5(32'hbb9bb63b),
	.w6(32'hbbb82201),
	.w7(32'h3c43be33),
	.w8(32'h3c8af0c2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d345c),
	.w1(32'h3ad91600),
	.w2(32'h3b8a457b),
	.w3(32'hbab84041),
	.w4(32'h3ab760c5),
	.w5(32'h3b043eab),
	.w6(32'h3c62018d),
	.w7(32'hb931bc5c),
	.w8(32'h3b74b5c1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd01f76),
	.w1(32'h3b43f089),
	.w2(32'h3a7ee4ec),
	.w3(32'h3bc2d136),
	.w4(32'h3bb29bfb),
	.w5(32'h3ba2a4a8),
	.w6(32'h3be3dfb6),
	.w7(32'hbaa444b1),
	.w8(32'h3b9f275e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1875e3),
	.w1(32'h3b17b80d),
	.w2(32'h3b1e03b0),
	.w3(32'h3baa5110),
	.w4(32'h3ac94bfc),
	.w5(32'h3b1c338e),
	.w6(32'h3a975697),
	.w7(32'hba9f639f),
	.w8(32'h3b3be2ea),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ea901),
	.w1(32'hbb6eae8b),
	.w2(32'h3b8eb7cb),
	.w3(32'h3bc9bc4a),
	.w4(32'h39bffcc0),
	.w5(32'hbc1d7442),
	.w6(32'h3bc1c25b),
	.w7(32'h3bad2f6f),
	.w8(32'h3a91a646),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb949187),
	.w1(32'h3b3577f7),
	.w2(32'hbc0e3207),
	.w3(32'hbb36d3dc),
	.w4(32'hb9afc3b7),
	.w5(32'hbc44c3a4),
	.w6(32'hbb756468),
	.w7(32'hbbaa88ad),
	.w8(32'hbc1ba5c4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b201e5),
	.w1(32'h3c333462),
	.w2(32'hbb42199b),
	.w3(32'hbb9283e6),
	.w4(32'h3b05cbdf),
	.w5(32'h3ab58ff9),
	.w6(32'hbb97f273),
	.w7(32'h3b8ebb37),
	.w8(32'h3c18b68a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcac87),
	.w1(32'hbc30473e),
	.w2(32'hbb6f4602),
	.w3(32'hbc2ed609),
	.w4(32'hbbc58c18),
	.w5(32'hbb39bd61),
	.w6(32'hbc262cee),
	.w7(32'hbbe08f53),
	.w8(32'hbc0235a9),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12ffeb),
	.w1(32'h39caad76),
	.w2(32'hbb5baf18),
	.w3(32'hbb6b35ff),
	.w4(32'hbc2d661c),
	.w5(32'h3c2bd6cf),
	.w6(32'h3b2f69fc),
	.w7(32'hb9894416),
	.w8(32'h3b5ca735),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3523b6),
	.w1(32'h3c2fe5a3),
	.w2(32'h3bd5abe0),
	.w3(32'h3b1664ae),
	.w4(32'h3ab6f081),
	.w5(32'hbb2f0c63),
	.w6(32'h3a5d20ca),
	.w7(32'hbb1a2712),
	.w8(32'hbbfcaa09),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dc797),
	.w1(32'hbbbedf4a),
	.w2(32'hbadb77ac),
	.w3(32'h3a9be200),
	.w4(32'hbbd75a2d),
	.w5(32'hba93cd54),
	.w6(32'h3ac83758),
	.w7(32'hbb79db40),
	.w8(32'h3ad9ca24),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0b998),
	.w1(32'h3ac5bef2),
	.w2(32'hbb885e7b),
	.w3(32'hbbb8716b),
	.w4(32'hbc693eb2),
	.w5(32'hbbccc4dc),
	.w6(32'h3b6fb6bc),
	.w7(32'hbc12bfc6),
	.w8(32'hbc366535),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9408c1b),
	.w1(32'hbbb2b422),
	.w2(32'hbb52560f),
	.w3(32'hbbcf8dc0),
	.w4(32'hbb93a86a),
	.w5(32'h3bbb3a46),
	.w6(32'hbb31105f),
	.w7(32'hbae71100),
	.w8(32'h39e5fbf2),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16239b),
	.w1(32'h3bf08117),
	.w2(32'hbc003fa8),
	.w3(32'hbb68f2dd),
	.w4(32'h3b83ed7a),
	.w5(32'hbb95cfc1),
	.w6(32'h39970bb0),
	.w7(32'h3c196b23),
	.w8(32'h3c3bdf1f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8060af),
	.w1(32'hbb52649e),
	.w2(32'h3bd27568),
	.w3(32'hbaca4cfb),
	.w4(32'hbc3b0b15),
	.w5(32'h3c401872),
	.w6(32'hbb385cd8),
	.w7(32'hbc094bc9),
	.w8(32'hbc884d6c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08c755),
	.w1(32'h3b3cf2dd),
	.w2(32'h3bb98e33),
	.w3(32'h3bd82ee4),
	.w4(32'h3a5c2bce),
	.w5(32'hbc053fbb),
	.w6(32'hbb96eec5),
	.w7(32'h3afb2f59),
	.w8(32'hbb2b97fd),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7beae2e),
	.w1(32'hba31ec9a),
	.w2(32'hbb771106),
	.w3(32'hbbd77534),
	.w4(32'hbc12074b),
	.w5(32'h3b9da380),
	.w6(32'hbbecb3f5),
	.w7(32'hbc59b9bf),
	.w8(32'hbb223e8f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babf8b6),
	.w1(32'h3c1c8a45),
	.w2(32'h3c4c2531),
	.w3(32'h3bb28753),
	.w4(32'h3c4c6c88),
	.w5(32'hba18779e),
	.w6(32'hbb554d67),
	.w7(32'h3cb11ff3),
	.w8(32'h3ca7cca6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e5d45),
	.w1(32'h3c7b5d4e),
	.w2(32'h3ccd2905),
	.w3(32'hbbea392f),
	.w4(32'h3ba95510),
	.w5(32'h3b9366a4),
	.w6(32'hb6296cc2),
	.w7(32'hbc0fdea0),
	.w8(32'hbc9bf291),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76bba4),
	.w1(32'h3b31d960),
	.w2(32'hbaf48037),
	.w3(32'hbb47c17c),
	.w4(32'hbb40fc88),
	.w5(32'hbc136d4e),
	.w6(32'hbc2de124),
	.w7(32'hbba463cc),
	.w8(32'hbbe9b11d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a7820),
	.w1(32'hbb377a30),
	.w2(32'hba33954e),
	.w3(32'hbc41bad0),
	.w4(32'hbc00e8e2),
	.w5(32'hbc08897e),
	.w6(32'hbbafdd99),
	.w7(32'h3b78d1f3),
	.w8(32'hbc1b62c3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398701f2),
	.w1(32'hba81f70b),
	.w2(32'h3c33a6c5),
	.w3(32'hbb36474a),
	.w4(32'hbb59ed31),
	.w5(32'h3bdaf9b8),
	.w6(32'h3bd14f7f),
	.w7(32'h3b8834ae),
	.w8(32'hbb8ea162),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1b2aa),
	.w1(32'hbc384741),
	.w2(32'hbbce72ed),
	.w3(32'hba26d548),
	.w4(32'hbc156692),
	.w5(32'h3bcbf2e7),
	.w6(32'hba7789df),
	.w7(32'hbbb759d9),
	.w8(32'hbba8f2c7),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5eb4c3),
	.w1(32'hbc1c9c18),
	.w2(32'hbc759eee),
	.w3(32'h3c994adc),
	.w4(32'hbbaaa9b9),
	.w5(32'h3a5b1b8e),
	.w6(32'h3c4fb98c),
	.w7(32'h3a33aff3),
	.w8(32'h3c4a29dc),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc913515),
	.w1(32'h3b4f5131),
	.w2(32'hbbc5d1e0),
	.w3(32'hbb7ce4c8),
	.w4(32'hba687a72),
	.w5(32'h3bc22392),
	.w6(32'h3acba81d),
	.w7(32'h3b54b7fc),
	.w8(32'h3b3cbea8),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf6988),
	.w1(32'h3b0d25ef),
	.w2(32'h38a135b2),
	.w3(32'hbb1b9feb),
	.w4(32'hba76909e),
	.w5(32'hbc04db6e),
	.w6(32'hbb5c243f),
	.w7(32'hbba0d6fc),
	.w8(32'h3b62dd2c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b5fde),
	.w1(32'hb9f5554c),
	.w2(32'h3c22b39b),
	.w3(32'hbb3dd912),
	.w4(32'h3b2a9e0e),
	.w5(32'h3b43893e),
	.w6(32'h3a858339),
	.w7(32'hbb9335e9),
	.w8(32'hbbd3eb70),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8954e4),
	.w1(32'h3c01aef1),
	.w2(32'h3b37be5e),
	.w3(32'h3c5a6733),
	.w4(32'h3a1960a5),
	.w5(32'h3bd4af87),
	.w6(32'h3c1709dd),
	.w7(32'h3c114f6d),
	.w8(32'h3c00eebb),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb572257),
	.w1(32'hbb400206),
	.w2(32'hbc214bf1),
	.w3(32'h3aa7608f),
	.w4(32'h3c511b92),
	.w5(32'h3c1c207e),
	.w6(32'h3bff4b27),
	.w7(32'h3bca48cd),
	.w8(32'h3c067c7c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4111ec),
	.w1(32'h3c0c5590),
	.w2(32'h3bb27de5),
	.w3(32'hbbdf2cb3),
	.w4(32'h3b277f9d),
	.w5(32'h3afde24c),
	.w6(32'h3bc21bbd),
	.w7(32'h3c176a0d),
	.w8(32'h3b9da6c8),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd9c86),
	.w1(32'h3bc751b6),
	.w2(32'hb926fe73),
	.w3(32'hbb74d76e),
	.w4(32'h3b46960d),
	.w5(32'hbc45b70f),
	.w6(32'hba149d6c),
	.w7(32'h3c11e041),
	.w8(32'hbacceb15),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5caf4d),
	.w1(32'h3b87386a),
	.w2(32'h3a2c8b36),
	.w3(32'hbbf39019),
	.w4(32'h3c8275f2),
	.w5(32'h3b9156ef),
	.w6(32'hbba1ee00),
	.w7(32'h3b30b53c),
	.w8(32'h3b6e5097),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b8fe9),
	.w1(32'hbc46d757),
	.w2(32'hbcb5f53f),
	.w3(32'hbc22bdfc),
	.w4(32'hbc451fd5),
	.w5(32'h3bfef079),
	.w6(32'h3ae6250e),
	.w7(32'h3b125796),
	.w8(32'h3c18acf8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e428a),
	.w1(32'hba2aadf1),
	.w2(32'h3beedb93),
	.w3(32'hba502bba),
	.w4(32'hbbe680e2),
	.w5(32'hbbc694e8),
	.w6(32'h3c277ff2),
	.w7(32'hbb9e7359),
	.w8(32'hbc737659),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb771db),
	.w1(32'hbb48ce99),
	.w2(32'hbbdb05b2),
	.w3(32'hbbc13509),
	.w4(32'h398bdece),
	.w5(32'hbc0e5d0b),
	.w6(32'hbc17160d),
	.w7(32'hbb7ed74d),
	.w8(32'hbbe521c5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0627c0),
	.w1(32'h3b3853f5),
	.w2(32'h3a7c70d4),
	.w3(32'h3b71270d),
	.w4(32'hb9d9ade7),
	.w5(32'h3b1b0eee),
	.w6(32'hbadae5f0),
	.w7(32'hbb735fe7),
	.w8(32'h3adb73ad),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39baf285),
	.w1(32'hbc156e51),
	.w2(32'hbc5d7e21),
	.w3(32'h3c59aeca),
	.w4(32'hbc4e2b2f),
	.w5(32'h3bff78db),
	.w6(32'h3c80889f),
	.w7(32'h3b002c36),
	.w8(32'h3c4acc0d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f7716),
	.w1(32'hbb23e82a),
	.w2(32'hbbacb8d6),
	.w3(32'h3caea45a),
	.w4(32'h3b064810),
	.w5(32'hba089c3f),
	.w6(32'h3c6a9781),
	.w7(32'h3b2855f4),
	.w8(32'h3bc0996a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeebc84),
	.w1(32'hbb20c9cf),
	.w2(32'h3a365743),
	.w3(32'hbbcc19b7),
	.w4(32'hb902c64f),
	.w5(32'h3ae66d1f),
	.w6(32'hbacdbe87),
	.w7(32'h3b240252),
	.w8(32'hbc0bb71f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6ac15),
	.w1(32'h3850ec21),
	.w2(32'hbc17e40f),
	.w3(32'h3b40b526),
	.w4(32'hbb51ff95),
	.w5(32'h3af44ddf),
	.w6(32'hba313078),
	.w7(32'h3b4e14b1),
	.w8(32'h3a8a4e9f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f99b6),
	.w1(32'hbb337837),
	.w2(32'h3c591db7),
	.w3(32'hbbedf48a),
	.w4(32'h3a029163),
	.w5(32'hbb96e634),
	.w6(32'h3b84e14c),
	.w7(32'hbbb06be2),
	.w8(32'hbc7bad8d),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f6155),
	.w1(32'h3b374d5c),
	.w2(32'hbc088015),
	.w3(32'hba94998c),
	.w4(32'hbb81c3b2),
	.w5(32'hb9b23463),
	.w6(32'hbb43b4d8),
	.w7(32'hb9443f36),
	.w8(32'hb9857d75),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09a1fd),
	.w1(32'h3c3be75d),
	.w2(32'h3c332742),
	.w3(32'h38e16598),
	.w4(32'h3bcd7d70),
	.w5(32'hbbcbdfb6),
	.w6(32'hbad85db3),
	.w7(32'hbaf6ada5),
	.w8(32'hbc01e327),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be931ce),
	.w1(32'h3b92abb8),
	.w2(32'h3c4d6fe1),
	.w3(32'hbb70510b),
	.w4(32'h3b8ce443),
	.w5(32'hbbb564a2),
	.w6(32'hbc2e13fc),
	.w7(32'hbbe86d2c),
	.w8(32'hbca0a106),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1600d),
	.w1(32'hbbdca4a8),
	.w2(32'hba822c1a),
	.w3(32'hbbd9e75b),
	.w4(32'hbbb66299),
	.w5(32'h3b165e56),
	.w6(32'hbbdaa103),
	.w7(32'hba2b068c),
	.w8(32'h3a44569c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd4c41),
	.w1(32'hbb9095c4),
	.w2(32'h3bc8b9ac),
	.w3(32'hbbda594a),
	.w4(32'hbaa474e7),
	.w5(32'h3b95c7b0),
	.w6(32'hbb8b60cc),
	.w7(32'h3979db0d),
	.w8(32'h3b1c46d3),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba874c2),
	.w1(32'hb9a01b88),
	.w2(32'hbc57f923),
	.w3(32'hbb70ba59),
	.w4(32'hbbb68b50),
	.w5(32'hbaa73e39),
	.w6(32'hbbf20ee2),
	.w7(32'hbb382cf0),
	.w8(32'h3a8ac78c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ecc6a),
	.w1(32'hbc1fd6b8),
	.w2(32'h3b610126),
	.w3(32'hb8dd3cee),
	.w4(32'h3bff7235),
	.w5(32'hbc3c8354),
	.w6(32'h39ad677c),
	.w7(32'hbaa6fa39),
	.w8(32'h3c75bf39),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb864cb7),
	.w1(32'hb98e4582),
	.w2(32'h3c2d7b24),
	.w3(32'h3bcbe322),
	.w4(32'h3add1b67),
	.w5(32'h3c0e85e1),
	.w6(32'h3c25b0b7),
	.w7(32'hbc0e88af),
	.w8(32'hbc958c26),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ff235),
	.w1(32'hb9b62ec7),
	.w2(32'h3b9e3125),
	.w3(32'h3c0a825f),
	.w4(32'hbb545df0),
	.w5(32'h3c187f54),
	.w6(32'hb990cad0),
	.w7(32'h3a95174c),
	.w8(32'h3bba040c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5ee4b),
	.w1(32'hbb87162f),
	.w2(32'hbb06e1f8),
	.w3(32'hbba51d57),
	.w4(32'hbb8579c5),
	.w5(32'h3b4f9e9d),
	.w6(32'h39c373ae),
	.w7(32'hbb12734d),
	.w8(32'h3b8ed46f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b416890),
	.w1(32'hb7a2a807),
	.w2(32'hbbe42d77),
	.w3(32'hbb807958),
	.w4(32'h3b8b8aaa),
	.w5(32'h3bedd12f),
	.w6(32'hbc1e923f),
	.w7(32'h3be8b3e4),
	.w8(32'h3ca934ec),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87abdf),
	.w1(32'hba265584),
	.w2(32'h3bfc8265),
	.w3(32'hbb65e47e),
	.w4(32'hb5d169bb),
	.w5(32'h3943cdeb),
	.w6(32'h3b165eaa),
	.w7(32'hbb108d6f),
	.w8(32'hbba7de19),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc93081),
	.w1(32'h3b4adf48),
	.w2(32'h3b1f0ac4),
	.w3(32'h3b62b8b2),
	.w4(32'h3a0dd501),
	.w5(32'h3ba1f4ea),
	.w6(32'hb91c2f7b),
	.w7(32'hbc1cfb47),
	.w8(32'hbbdb9eff),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5795ab),
	.w1(32'h3b3c0725),
	.w2(32'h3b1bbd80),
	.w3(32'h3b7b6dbc),
	.w4(32'h3aee227e),
	.w5(32'hba77cd67),
	.w6(32'hbba77af0),
	.w7(32'hba7587ef),
	.w8(32'hba1c2b9c),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cb290),
	.w1(32'h3b5387f6),
	.w2(32'hbb4d64b9),
	.w3(32'h3b9fedb6),
	.w4(32'hbbe415bb),
	.w5(32'h3c0dc9fc),
	.w6(32'h3acf9af1),
	.w7(32'h3b7fa3c1),
	.w8(32'h3bb39031),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a43e4),
	.w1(32'hbc2cff75),
	.w2(32'hbc199d41),
	.w3(32'hbb40c3b4),
	.w4(32'hbba681dc),
	.w5(32'h3a4b7d72),
	.w6(32'h3bc482ac),
	.w7(32'hbb20daad),
	.w8(32'h3aec1caf),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbeefc1),
	.w1(32'h3b58b49a),
	.w2(32'hbbb5896c),
	.w3(32'hbb83b9e2),
	.w4(32'h38d89417),
	.w5(32'hbc01e0eb),
	.w6(32'h3a533857),
	.w7(32'h3b5d000a),
	.w8(32'h3aeb8737),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0141af),
	.w1(32'h3b6224a1),
	.w2(32'h3bdf87a4),
	.w3(32'hbb405d7c),
	.w4(32'h3b295d42),
	.w5(32'h3c007e62),
	.w6(32'h3a06dc14),
	.w7(32'hbb740de6),
	.w8(32'hbb2ec254),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b202b),
	.w1(32'hbbc27133),
	.w2(32'hbbb72e58),
	.w3(32'h3c131028),
	.w4(32'hbb842771),
	.w5(32'hbb22e631),
	.w6(32'hbc391628),
	.w7(32'hbb59f493),
	.w8(32'hbc1d3b1b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18a6a7),
	.w1(32'h3b5410ee),
	.w2(32'h3c3d96ae),
	.w3(32'hbc1065cf),
	.w4(32'hb934dd4a),
	.w5(32'h3b131023),
	.w6(32'hbb5fee25),
	.w7(32'hbb9b49e1),
	.w8(32'hbc323f50),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63906b),
	.w1(32'hbbb4075a),
	.w2(32'hbb74ea77),
	.w3(32'h3b0f26af),
	.w4(32'hbbed2e13),
	.w5(32'h3be32241),
	.w6(32'hbc2ff8b5),
	.w7(32'hbb53052e),
	.w8(32'hbbde5750),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d0c5d),
	.w1(32'hb9d30c0d),
	.w2(32'hbb5aa0a5),
	.w3(32'h3bdcaabf),
	.w4(32'hbad58645),
	.w5(32'h3a951828),
	.w6(32'hbc0a4982),
	.w7(32'hbbdadaba),
	.w8(32'hbbdf689c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d19e12),
	.w1(32'hbb495690),
	.w2(32'hbc3b6b7d),
	.w3(32'hbb80aa8b),
	.w4(32'hbb9aafdd),
	.w5(32'hbbbe2fec),
	.w6(32'h3b6184db),
	.w7(32'hbc654064),
	.w8(32'hbc3770e4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72bd1f),
	.w1(32'hbc138695),
	.w2(32'hbc8267a0),
	.w3(32'hbb9bbf93),
	.w4(32'hbc98ccfd),
	.w5(32'hbc3a0777),
	.w6(32'hbb6ba669),
	.w7(32'hbaed34a6),
	.w8(32'hbb38caf4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule