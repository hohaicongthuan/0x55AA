module layer_10_featuremap_394(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac62c2),
	.w1(32'h3b0f25b4),
	.w2(32'h3b52527e),
	.w3(32'h3c15f690),
	.w4(32'hbaa188b2),
	.w5(32'hbb3de653),
	.w6(32'h3b418b03),
	.w7(32'h39cae787),
	.w8(32'h3b75176b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcedaa0),
	.w1(32'hba9ade29),
	.w2(32'hbac98860),
	.w3(32'hb8609d94),
	.w4(32'hbb377f38),
	.w5(32'h3a1ae3dc),
	.w6(32'h3b97ec3e),
	.w7(32'h3a0e3aa8),
	.w8(32'h3a61ce5e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e8a3e),
	.w1(32'hb9d7c27f),
	.w2(32'hbb802b8a),
	.w3(32'hbb8f440f),
	.w4(32'h3aca3a71),
	.w5(32'h3c034392),
	.w6(32'hbbfa2c9f),
	.w7(32'hbb8fd9e0),
	.w8(32'hbbf5f8a6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcb936),
	.w1(32'hbbbd0e86),
	.w2(32'h3c199632),
	.w3(32'hbb654761),
	.w4(32'h3b5342d3),
	.w5(32'h3a52c03e),
	.w6(32'hb9fc98d9),
	.w7(32'h3af20c74),
	.w8(32'hbb426c5c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7338b3),
	.w1(32'hb92830e5),
	.w2(32'hbb35c3af),
	.w3(32'hbb6370a2),
	.w4(32'hbb21fc52),
	.w5(32'hbb0886bb),
	.w6(32'hba3e380f),
	.w7(32'h3a51fa6c),
	.w8(32'hbbed5a69),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b823c8),
	.w1(32'h3adbef76),
	.w2(32'hbbc6b54c),
	.w3(32'hba9647b7),
	.w4(32'hbb925ae8),
	.w5(32'h3b396d51),
	.w6(32'hbb83a61d),
	.w7(32'h3b2b39fa),
	.w8(32'h3c7a9263),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8842c2),
	.w1(32'h39cdd78b),
	.w2(32'h3bb5c0f8),
	.w3(32'hbba8eee8),
	.w4(32'h3b80bb82),
	.w5(32'hbad17cdb),
	.w6(32'hb94d720b),
	.w7(32'hb9602422),
	.w8(32'hbb3585de),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fca04),
	.w1(32'h3a93db74),
	.w2(32'h3b96e7ad),
	.w3(32'hbc02aca7),
	.w4(32'h3977d13b),
	.w5(32'hbbde59ae),
	.w6(32'h3aa61786),
	.w7(32'h3c2df903),
	.w8(32'h3bb836fa),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c5a81),
	.w1(32'h3b5a2425),
	.w2(32'h3bb1fd5d),
	.w3(32'h3b8063d1),
	.w4(32'h39cad6e3),
	.w5(32'hbbb1944d),
	.w6(32'h3bf663d2),
	.w7(32'hbb536272),
	.w8(32'hbb181b31),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b348f73),
	.w1(32'hb8ac4680),
	.w2(32'hba6a8cb2),
	.w3(32'hbbad1e71),
	.w4(32'hba9e56b1),
	.w5(32'hbbc0cbae),
	.w6(32'hbb0b241a),
	.w7(32'hbbb51337),
	.w8(32'hbbd08a7e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1eec0f),
	.w1(32'h3b1a0506),
	.w2(32'h3a6b81f8),
	.w3(32'hbb2d3297),
	.w4(32'hbb2bc2e0),
	.w5(32'hbbc07dec),
	.w6(32'hba93091d),
	.w7(32'h3b105e84),
	.w8(32'hbb4a378b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fbe36),
	.w1(32'h3bbbb8d1),
	.w2(32'h3bcda833),
	.w3(32'hbb4977ce),
	.w4(32'hbbaacf60),
	.w5(32'h3a620e4b),
	.w6(32'hbb220994),
	.w7(32'hbb49c0bb),
	.w8(32'hbbcd90c8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7d749),
	.w1(32'h3b62b560),
	.w2(32'hbbe5ecb3),
	.w3(32'hbbcb29e2),
	.w4(32'h3a46041a),
	.w5(32'hb9a62274),
	.w6(32'hbbd0226a),
	.w7(32'hbbbcc8f7),
	.w8(32'hbc13e8bd),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b8413),
	.w1(32'hba812f52),
	.w2(32'h3a190e6e),
	.w3(32'hba378efa),
	.w4(32'h3b31059f),
	.w5(32'h3bded1e6),
	.w6(32'hbb6bf4a1),
	.w7(32'h3b49acd1),
	.w8(32'hbc21706e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47b3ca),
	.w1(32'hbb8d6cdd),
	.w2(32'hbb8c1084),
	.w3(32'h3ba6a5b0),
	.w4(32'hbb1421b7),
	.w5(32'hba547a7d),
	.w6(32'hbb220b75),
	.w7(32'hbb4d66f9),
	.w8(32'hbb8b584d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc1251),
	.w1(32'hbb6dfb0b),
	.w2(32'hbc07a0d0),
	.w3(32'hb88448f3),
	.w4(32'hbb99d96e),
	.w5(32'hbba036bf),
	.w6(32'h3b10214d),
	.w7(32'hbbcc224d),
	.w8(32'hbb915f68),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab2b4b),
	.w1(32'hbb0ec65f),
	.w2(32'h3a3a65cc),
	.w3(32'h3ac00f31),
	.w4(32'hbaa2e431),
	.w5(32'hba193bfc),
	.w6(32'h3b6edf43),
	.w7(32'hbb861132),
	.w8(32'hbc0a506a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb98b77),
	.w1(32'h3b12b489),
	.w2(32'hbb3c98d3),
	.w3(32'hbb937a23),
	.w4(32'hba422177),
	.w5(32'hbb2acfd7),
	.w6(32'h3b371bd0),
	.w7(32'h3b885990),
	.w8(32'h3bb0246d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccb3ad),
	.w1(32'h3ad291a8),
	.w2(32'hbb3ac216),
	.w3(32'hbbb2bacc),
	.w4(32'hbb8fd1eb),
	.w5(32'hbb116275),
	.w6(32'h3b9e9554),
	.w7(32'hbb920f25),
	.w8(32'h3ad4cb40),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74e9ef),
	.w1(32'hbab00ec3),
	.w2(32'hba32683e),
	.w3(32'hbb13e460),
	.w4(32'hbabd54b9),
	.w5(32'hbb87bbe4),
	.w6(32'hbb229dcf),
	.w7(32'h3bac81dc),
	.w8(32'hbafcc6bd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb412a5),
	.w1(32'hb9be7723),
	.w2(32'hbb7f111e),
	.w3(32'h3ab08734),
	.w4(32'hbba58d9d),
	.w5(32'h3af4b2cc),
	.w6(32'h3bfb8a2a),
	.w7(32'hbb10f140),
	.w8(32'h3afd150c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb013001),
	.w1(32'h3bdc2184),
	.w2(32'hbbb02ebb),
	.w3(32'hbbafd334),
	.w4(32'hbb7141b5),
	.w5(32'h3befbfe6),
	.w6(32'hbb85c79a),
	.w7(32'h3b391793),
	.w8(32'h3c4d5f30),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20b184),
	.w1(32'hbb1d85e8),
	.w2(32'h3938d3b2),
	.w3(32'h3a9c5e38),
	.w4(32'h3bb8efe3),
	.w5(32'hbb2851ba),
	.w6(32'h3c3085c6),
	.w7(32'hbab6d055),
	.w8(32'h3c0adf34),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb47de6),
	.w1(32'hbb0346b9),
	.w2(32'hbc01c557),
	.w3(32'h3bda0af4),
	.w4(32'h39eb1c50),
	.w5(32'hbbe3c6de),
	.w6(32'hb93802bf),
	.w7(32'hbad4d9c8),
	.w8(32'hbb3e93b5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1c748),
	.w1(32'hbab9c3f2),
	.w2(32'hbc252243),
	.w3(32'hbb8a22b3),
	.w4(32'h3b0c42cf),
	.w5(32'hbbe6f438),
	.w6(32'h3aee7ac2),
	.w7(32'h3bc0b045),
	.w8(32'h3baa9b92),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f704b),
	.w1(32'hbbbff148),
	.w2(32'hb92c9ad1),
	.w3(32'hbbbd46ed),
	.w4(32'hbb63caa8),
	.w5(32'h3ce7847d),
	.w6(32'h3c47c6f3),
	.w7(32'h3b18459e),
	.w8(32'h3cc6be2b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba687cb8),
	.w1(32'hb8e811fc),
	.w2(32'hbb46624d),
	.w3(32'h3c47083c),
	.w4(32'hbb3da183),
	.w5(32'h3bfba38c),
	.w6(32'h3cbbc3df),
	.w7(32'h3b79db39),
	.w8(32'h3c344686),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75b045),
	.w1(32'h3bdfbfd9),
	.w2(32'h39164468),
	.w3(32'h3c37e372),
	.w4(32'h3c10c82a),
	.w5(32'hbb401653),
	.w6(32'hbbe134f4),
	.w7(32'h3ab223db),
	.w8(32'hbc015d7a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bdf96),
	.w1(32'h3a65e482),
	.w2(32'h3a549ba6),
	.w3(32'hbb2c453e),
	.w4(32'hbb39bd4d),
	.w5(32'hbc017d24),
	.w6(32'hbb0d01a9),
	.w7(32'hbc249d63),
	.w8(32'hbb24436f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94fadb),
	.w1(32'h3bcdc9f1),
	.w2(32'h3b90d796),
	.w3(32'hbbf8331b),
	.w4(32'h3b48667b),
	.w5(32'h398a9127),
	.w6(32'h38883168),
	.w7(32'hbabe5a2e),
	.w8(32'hbba3e0f0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac83d1),
	.w1(32'hbb0b83bd),
	.w2(32'h3b807f7d),
	.w3(32'h398804c7),
	.w4(32'hbb5eeab3),
	.w5(32'hbb3dc560),
	.w6(32'hbbd4db53),
	.w7(32'h3b3ee402),
	.w8(32'hbafacbef),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfade8),
	.w1(32'h3b8c4490),
	.w2(32'h3b5f730d),
	.w3(32'hbbbf5d5e),
	.w4(32'hbaa5240a),
	.w5(32'h3b304877),
	.w6(32'h38af0840),
	.w7(32'h3ac8ba0b),
	.w8(32'h3aa8f6ce),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06e8e3),
	.w1(32'h36ba608a),
	.w2(32'h399fb79d),
	.w3(32'hb956b31c),
	.w4(32'h3b1e3d05),
	.w5(32'h3afa3be6),
	.w6(32'hbb7d4c9e),
	.w7(32'hbab9a797),
	.w8(32'hbba0be67),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b5aa9),
	.w1(32'h3b794d48),
	.w2(32'h3c11ee96),
	.w3(32'hbaf40234),
	.w4(32'h3bf95dfc),
	.w5(32'hbc0ebc7c),
	.w6(32'h3aa09b85),
	.w7(32'h3b421c86),
	.w8(32'h3a901aaf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a55e9),
	.w1(32'h3a5d0d5e),
	.w2(32'h3abd2760),
	.w3(32'hba0b19c5),
	.w4(32'h3aef6d6e),
	.w5(32'h3ad281a3),
	.w6(32'h3c076a43),
	.w7(32'h3bdca2cb),
	.w8(32'h3b419a17),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7be84e),
	.w1(32'hb9ab3f36),
	.w2(32'h3b6007f6),
	.w3(32'h3a9d5284),
	.w4(32'hba8b49b9),
	.w5(32'hba4da6c4),
	.w6(32'h3c255b56),
	.w7(32'hbae487d1),
	.w8(32'hba395051),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98e8e9),
	.w1(32'h3b4a762c),
	.w2(32'hbb129d48),
	.w3(32'hbb0184b3),
	.w4(32'hba4c5c80),
	.w5(32'h3ba35b8b),
	.w6(32'hbb706999),
	.w7(32'h3b649cfa),
	.w8(32'hbbabd5a5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a54741),
	.w1(32'hbbcce0a8),
	.w2(32'hbad6d6aa),
	.w3(32'h3baf8512),
	.w4(32'h3afd77b7),
	.w5(32'h39f0354d),
	.w6(32'hbbc694b6),
	.w7(32'hbb90bdc7),
	.w8(32'hbbb58f75),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81ac2c),
	.w1(32'h3a921ec9),
	.w2(32'hb960ecb7),
	.w3(32'hbac1ad00),
	.w4(32'h3b8d3cd8),
	.w5(32'hbaf25d25),
	.w6(32'hbc2afd91),
	.w7(32'hb9ff31ae),
	.w8(32'hbb9cea63),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1500c0),
	.w1(32'hbb0c22d1),
	.w2(32'h3afd5c53),
	.w3(32'h3ac07a73),
	.w4(32'h3bba2398),
	.w5(32'h3ae273a9),
	.w6(32'hb83b0b21),
	.w7(32'h3b7335b7),
	.w8(32'hba30a573),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d2849),
	.w1(32'h395afa27),
	.w2(32'h3b8dd72b),
	.w3(32'h3aff8e28),
	.w4(32'h3bbb3df9),
	.w5(32'h3c682765),
	.w6(32'h3b00f355),
	.w7(32'hbacc7ce3),
	.w8(32'hbbe58dee),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47f64f),
	.w1(32'hbaff1cac),
	.w2(32'hbb709f2a),
	.w3(32'h3b45119b),
	.w4(32'hbb0db012),
	.w5(32'h3b12269b),
	.w6(32'hbb27f797),
	.w7(32'hbb96c58b),
	.w8(32'hbbed3973),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d19d9),
	.w1(32'h3baf1225),
	.w2(32'h3b3ede4f),
	.w3(32'hbbb1dee0),
	.w4(32'h3b86cf76),
	.w5(32'h3b1a509b),
	.w6(32'hbc07be80),
	.w7(32'hb9e99f06),
	.w8(32'h3a816201),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba948331),
	.w1(32'hbc060cf4),
	.w2(32'hbb68145f),
	.w3(32'hbb7525cd),
	.w4(32'hbb8080a2),
	.w5(32'hbb7a3524),
	.w6(32'h3b53a294),
	.w7(32'h3ad8a5dc),
	.w8(32'hbb06027d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab21f8b),
	.w1(32'hbabcb901),
	.w2(32'hbba6b8fb),
	.w3(32'hbbebca27),
	.w4(32'hbab6587e),
	.w5(32'hbb54d4a9),
	.w6(32'hbaec7e97),
	.w7(32'hbb4b05de),
	.w8(32'hba3efea0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a58862),
	.w1(32'hbba15b89),
	.w2(32'hb9b18df1),
	.w3(32'h3ad8a0dc),
	.w4(32'hbb969583),
	.w5(32'hbbe39bd3),
	.w6(32'h3afbfb89),
	.w7(32'hb978a847),
	.w8(32'h398ea3d4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0293c0),
	.w1(32'hba81364f),
	.w2(32'hbc0a7b15),
	.w3(32'h3aef1b53),
	.w4(32'h3b671f69),
	.w5(32'h3c00f96c),
	.w6(32'h3b572a0d),
	.w7(32'h3be9d959),
	.w8(32'h3c1aa29a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dd7a6),
	.w1(32'hbac02d54),
	.w2(32'h3bc3cc75),
	.w3(32'h39ff5f21),
	.w4(32'hba9d3244),
	.w5(32'hba748e43),
	.w6(32'h3c741a96),
	.w7(32'h3c101f94),
	.w8(32'h3bbc71f6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadea8a4),
	.w1(32'h3b9efa1d),
	.w2(32'h3b759cbc),
	.w3(32'hbbd1f1a4),
	.w4(32'h3b2261e8),
	.w5(32'h39b5db31),
	.w6(32'hbb606a6d),
	.w7(32'hb9fea664),
	.w8(32'hbba04b60),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b936908),
	.w1(32'h3b9140ce),
	.w2(32'h3c0e6825),
	.w3(32'h3c2afb29),
	.w4(32'hba8e417e),
	.w5(32'h3b8eb6fc),
	.w6(32'h3bbfe7be),
	.w7(32'h3b89d281),
	.w8(32'h3c445e19),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef6a15),
	.w1(32'h398331c1),
	.w2(32'hba2e6c54),
	.w3(32'h3c0cd67e),
	.w4(32'hbaf28ff8),
	.w5(32'h3add6618),
	.w6(32'h3a4ddcd5),
	.w7(32'hbbbf893e),
	.w8(32'h39ca9cc4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91fe1f),
	.w1(32'hbaa6a929),
	.w2(32'h3b8b610a),
	.w3(32'hbb5b0261),
	.w4(32'hbb203c0b),
	.w5(32'hbbd5216b),
	.w6(32'hba11218c),
	.w7(32'h3b7c0f3c),
	.w8(32'h3bbdbbea),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c72ea),
	.w1(32'h3b99a140),
	.w2(32'h394bad3e),
	.w3(32'hbb952343),
	.w4(32'h39070ae6),
	.w5(32'hbbc4de41),
	.w6(32'h3abe6ed4),
	.w7(32'h3a58b5b6),
	.w8(32'h3bd8e984),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb583f5e),
	.w1(32'h3bb697a9),
	.w2(32'h39a4acde),
	.w3(32'hbb2a6d6e),
	.w4(32'h3ada7d87),
	.w5(32'hbb95277d),
	.w6(32'h3c23a8d7),
	.w7(32'h3bc68a33),
	.w8(32'h3c4fa384),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88a612),
	.w1(32'hbb149336),
	.w2(32'hbb53daa2),
	.w3(32'h3b366b89),
	.w4(32'h3bbeddf2),
	.w5(32'hbbf397b3),
	.w6(32'h3bdb36ab),
	.w7(32'h3b7449e4),
	.w8(32'hbb68e35d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6cce6),
	.w1(32'h3b7a2361),
	.w2(32'h3b89c026),
	.w3(32'hba133a71),
	.w4(32'h3ac4ca0f),
	.w5(32'h39b73250),
	.w6(32'h3b6f63aa),
	.w7(32'h3a0c721b),
	.w8(32'h3be14138),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4330f7),
	.w1(32'h3b123a0f),
	.w2(32'h3bb8ad66),
	.w3(32'hba2d2285),
	.w4(32'h3ba01b78),
	.w5(32'h3c31c489),
	.w6(32'h3ba2c8f7),
	.w7(32'h3b56ed3d),
	.w8(32'h39b41f65),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b75de),
	.w1(32'hba706686),
	.w2(32'hbb838a13),
	.w3(32'h3bc4763e),
	.w4(32'hbba9e6fa),
	.w5(32'hbb56698f),
	.w6(32'hbae70d07),
	.w7(32'hbb791735),
	.w8(32'h3b9398d7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8deb56),
	.w1(32'h3bd143ea),
	.w2(32'hbad47923),
	.w3(32'hbafa3648),
	.w4(32'h3c122a5f),
	.w5(32'hbb438f3f),
	.w6(32'hbbbf8410),
	.w7(32'h3b0f1f51),
	.w8(32'hbb31633f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0edc85),
	.w1(32'hbabb2159),
	.w2(32'hbc012a19),
	.w3(32'h3b529910),
	.w4(32'h3a41c5e5),
	.w5(32'h3bbb54be),
	.w6(32'h3b79bf5a),
	.w7(32'h3ac6c219),
	.w8(32'h3a5a0a6e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6a641),
	.w1(32'h3a303acd),
	.w2(32'hbb0be425),
	.w3(32'h3bbb261d),
	.w4(32'h3ba61d83),
	.w5(32'h3cb51048),
	.w6(32'h3c658f04),
	.w7(32'h3c1b752f),
	.w8(32'h3b915746),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb06964),
	.w1(32'h3b917f72),
	.w2(32'h3bd729d7),
	.w3(32'h3beeda85),
	.w4(32'h3b76514b),
	.w5(32'h3bae9e0f),
	.w6(32'hb9af4852),
	.w7(32'h3bb511ba),
	.w8(32'hb9b7c1e8),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b445912),
	.w1(32'hbb351808),
	.w2(32'hbbacdb64),
	.w3(32'h3b2a52ef),
	.w4(32'h3ab32999),
	.w5(32'hbb551cb9),
	.w6(32'h3ba63b6f),
	.w7(32'hbc0a9bd7),
	.w8(32'h3a64e3a2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9814cf),
	.w1(32'h3bd8f91c),
	.w2(32'h3bc139e7),
	.w3(32'hbb797ef5),
	.w4(32'h3b0c29ea),
	.w5(32'h3b1b3ca7),
	.w6(32'h3b75db00),
	.w7(32'hbb269dc0),
	.w8(32'hba09f821),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd4a5f),
	.w1(32'h3b943c50),
	.w2(32'h3c2b2135),
	.w3(32'h3b2ea7b1),
	.w4(32'h3b6ebcea),
	.w5(32'h3aeb67ae),
	.w6(32'h3aef08f1),
	.w7(32'hba0f7315),
	.w8(32'hb8ad8e83),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c298d4c),
	.w1(32'h3ad9181e),
	.w2(32'h3b907bf4),
	.w3(32'h3bd2c76b),
	.w4(32'h396d21f2),
	.w5(32'h3b0ee21b),
	.w6(32'h3b105025),
	.w7(32'hba935be1),
	.w8(32'h3b7a252f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b7de5),
	.w1(32'h398cb5b0),
	.w2(32'hbb2b9954),
	.w3(32'h3badbd47),
	.w4(32'hbb733505),
	.w5(32'hbb897357),
	.w6(32'h3b6ff260),
	.w7(32'hbc0ed4a5),
	.w8(32'h3afa2cfe),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a99ed),
	.w1(32'h3b439c03),
	.w2(32'h3bc04e4f),
	.w3(32'h3abb8184),
	.w4(32'h3b712cbe),
	.w5(32'hba55ae5e),
	.w6(32'h3ae1cc1e),
	.w7(32'h3afbb759),
	.w8(32'hba16ff15),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03a17a),
	.w1(32'h38e31d12),
	.w2(32'hbba4f756),
	.w3(32'h3ac830a7),
	.w4(32'h3ac13a24),
	.w5(32'hbbbea8b6),
	.w6(32'h3bdf89c7),
	.w7(32'hb883aa6c),
	.w8(32'hbb6844a4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05ea3d),
	.w1(32'hbbc13151),
	.w2(32'hbbc02e4a),
	.w3(32'hbc174f3b),
	.w4(32'hbb21060a),
	.w5(32'hbbe16f8b),
	.w6(32'hba8759be),
	.w7(32'hbb9b0806),
	.w8(32'hbc1be1c9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9b2ae),
	.w1(32'hbb8c4e0c),
	.w2(32'hbb88717c),
	.w3(32'h3b347b37),
	.w4(32'hbaa7b260),
	.w5(32'h3b61deaa),
	.w6(32'h3b46b2c6),
	.w7(32'hba9f64e6),
	.w8(32'hbbb672d9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b045dc4),
	.w1(32'h3b13fdf4),
	.w2(32'hbae59d3e),
	.w3(32'h3b156571),
	.w4(32'h3ab5287e),
	.w5(32'h3c7475e5),
	.w6(32'h3a87d764),
	.w7(32'h3a0a7fff),
	.w8(32'hba704a27),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b015b),
	.w1(32'hba6b0571),
	.w2(32'hbb3e53a8),
	.w3(32'h3b6e1e46),
	.w4(32'hbb885e7b),
	.w5(32'hbbc7314e),
	.w6(32'h384b0a4c),
	.w7(32'h3aebd91d),
	.w8(32'h3a8b96d5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85efbd),
	.w1(32'hbad1b5ea),
	.w2(32'h3b3a03a2),
	.w3(32'hbb0138c8),
	.w4(32'hbbd70805),
	.w5(32'hbc579b60),
	.w6(32'h3c272870),
	.w7(32'hbc07d6cc),
	.w8(32'hbc3e32b4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d75d8),
	.w1(32'hbc2817d0),
	.w2(32'hbc43bf19),
	.w3(32'hbbec3a53),
	.w4(32'hbcd4da26),
	.w5(32'hbd34fd29),
	.w6(32'hbb4891b1),
	.w7(32'hbbfbd953),
	.w8(32'hbc4c9715),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadba96),
	.w1(32'hbbbc7467),
	.w2(32'hbb551669),
	.w3(32'hbd00b0cb),
	.w4(32'hbc060a68),
	.w5(32'hbb816222),
	.w6(32'hbc2aef9f),
	.w7(32'hbc3537c1),
	.w8(32'hbbdc72ac),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e4f56),
	.w1(32'h3b46660d),
	.w2(32'h3a9fe1e5),
	.w3(32'hbc1220a8),
	.w4(32'h3aa00a50),
	.w5(32'hbb67a77f),
	.w6(32'hbbaff3b0),
	.w7(32'h3bd086af),
	.w8(32'h3b310c39),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99fe3a),
	.w1(32'hbbcc985d),
	.w2(32'h3ac0a057),
	.w3(32'h3ba13433),
	.w4(32'h3be189a8),
	.w5(32'h3d371d26),
	.w6(32'h3b38639e),
	.w7(32'h3ba97bb6),
	.w8(32'h3c4c4845),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4433c8),
	.w1(32'hbb1517c4),
	.w2(32'hbad89cf5),
	.w3(32'h3b751e96),
	.w4(32'hb94c9864),
	.w5(32'h3bd1b6d4),
	.w6(32'h3bf407f2),
	.w7(32'h3b2b6bdc),
	.w8(32'h3b86e2b1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf2ccf),
	.w1(32'h3b2d9e4a),
	.w2(32'hbbced5db),
	.w3(32'hba3da53b),
	.w4(32'hbb8c74d3),
	.w5(32'hbba683c1),
	.w6(32'h3c2ab671),
	.w7(32'hbab13673),
	.w8(32'hba1de79c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985b3ca),
	.w1(32'h3c0ddb53),
	.w2(32'h3c4de2ee),
	.w3(32'hbba3fc28),
	.w4(32'hba23a099),
	.w5(32'hbaf58a31),
	.w6(32'hbb2c1673),
	.w7(32'h3c75844b),
	.w8(32'h3bdd63b0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4066b9),
	.w1(32'hbc15c1c3),
	.w2(32'hbbc9f6a5),
	.w3(32'h3b01ba2f),
	.w4(32'hbbb0a7cb),
	.w5(32'h3b4737b5),
	.w6(32'h3c7e3832),
	.w7(32'hbb9d4932),
	.w8(32'h3b48a846),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ff306),
	.w1(32'h3c82fb18),
	.w2(32'h3c7c98be),
	.w3(32'h3a7bee59),
	.w4(32'h3c8688ad),
	.w5(32'h3cdfb428),
	.w6(32'h3ae8868a),
	.w7(32'h3c7d3bf4),
	.w8(32'h3c808aa5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c974980),
	.w1(32'h3ba9efc4),
	.w2(32'hbbdb02d8),
	.w3(32'h3c4ed624),
	.w4(32'hbc106533),
	.w5(32'hbbb49d9a),
	.w6(32'h3c2ffd74),
	.w7(32'h3bc77df6),
	.w8(32'h3b4bd4ed),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b531e8a),
	.w1(32'hbbde2c23),
	.w2(32'hbc386176),
	.w3(32'hb8ccad98),
	.w4(32'h39bf33c6),
	.w5(32'h3c426960),
	.w6(32'hb97e9fc4),
	.w7(32'h3b8be9ab),
	.w8(32'h3c63b60d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c5e24),
	.w1(32'h3c2bf649),
	.w2(32'h3abb4823),
	.w3(32'hbba4ade2),
	.w4(32'hbb333309),
	.w5(32'h3b2aabee),
	.w6(32'h3b84d980),
	.w7(32'hbbdb798d),
	.w8(32'hbbf487d9),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8c265),
	.w1(32'hbb7e67ac),
	.w2(32'hbb81a88d),
	.w3(32'h3bb1bb35),
	.w4(32'h3b903906),
	.w5(32'h3cd7efc9),
	.w6(32'h3b8114fa),
	.w7(32'h3c0b2960),
	.w8(32'h3c260792),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba88687),
	.w1(32'h3af0ad38),
	.w2(32'h3b00aa39),
	.w3(32'h3acccc67),
	.w4(32'h3bfe3d89),
	.w5(32'h3d2a4b3d),
	.w6(32'hb9c496fd),
	.w7(32'h3bf72277),
	.w8(32'h3ce316c9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed4f13),
	.w1(32'hbad44ba2),
	.w2(32'h38a29cce),
	.w3(32'h3b040d1e),
	.w4(32'hbb65f4a7),
	.w5(32'h3b8250b2),
	.w6(32'h3c95a0ed),
	.w7(32'h3b8ff0f7),
	.w8(32'h3c298455),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82ee50),
	.w1(32'hbb2d8b5d),
	.w2(32'hbbf3a37a),
	.w3(32'h3b48b74c),
	.w4(32'hbb970c4c),
	.w5(32'h3bd7f494),
	.w6(32'h3ab23057),
	.w7(32'h3b074ce6),
	.w8(32'h3c100044),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f02b8),
	.w1(32'hba6dff59),
	.w2(32'hbc025f1f),
	.w3(32'h3b65aa1d),
	.w4(32'h3acb9eb5),
	.w5(32'hba266dab),
	.w6(32'hbb295272),
	.w7(32'h39d01521),
	.w8(32'hbb5ebc5f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1c124),
	.w1(32'h3aaa5af1),
	.w2(32'hbb88cd81),
	.w3(32'h3bac7f86),
	.w4(32'h3b342db9),
	.w5(32'h3ae8e0ed),
	.w6(32'hba9611b1),
	.w7(32'hbb74de25),
	.w8(32'hbba3ab3d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3f331),
	.w1(32'hbbb29507),
	.w2(32'hbc847f57),
	.w3(32'h3b9099fb),
	.w4(32'hbc1f7c6b),
	.w5(32'hbbdf9734),
	.w6(32'hbb952dce),
	.w7(32'h3acdd6cd),
	.w8(32'hba5bf876),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf50ce),
	.w1(32'hbcdb5992),
	.w2(32'hbd262219),
	.w3(32'hbc1380c0),
	.w4(32'hbd1bc1f5),
	.w5(32'hbd71e65f),
	.w6(32'h3bd4559c),
	.w7(32'hbc0eff75),
	.w8(32'hbcfb9f0d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7eaa5),
	.w1(32'h3a50fc29),
	.w2(32'hbc143e61),
	.w3(32'hbd21e0f4),
	.w4(32'h3c20cc6b),
	.w5(32'h3c90179a),
	.w6(32'hbcbbc99b),
	.w7(32'h3a546d14),
	.w8(32'h3a9a03a2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8c967),
	.w1(32'h3b018346),
	.w2(32'hbac792bd),
	.w3(32'h3bbe7003),
	.w4(32'h373d7a55),
	.w5(32'hba8eba7f),
	.w6(32'hbb0f7c57),
	.w7(32'hbbcb2317),
	.w8(32'hbb85c7c8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4b8a3),
	.w1(32'hbb474741),
	.w2(32'hbbd949d5),
	.w3(32'h3bf1cb33),
	.w4(32'hbb3f4359),
	.w5(32'h3b385816),
	.w6(32'hbb5cc512),
	.w7(32'hbbafd51e),
	.w8(32'h3bc01c60),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc435416),
	.w1(32'hbbf28715),
	.w2(32'hbc464b6f),
	.w3(32'hbb7a65f5),
	.w4(32'hb9d47b4f),
	.w5(32'h3b355038),
	.w6(32'h3c3b9cca),
	.w7(32'h3c54e8b7),
	.w8(32'h3c07e7ce),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24dc4d),
	.w1(32'hbb1e8c18),
	.w2(32'hbbcaa427),
	.w3(32'hba8cf73e),
	.w4(32'hbb690051),
	.w5(32'h3b97b085),
	.w6(32'h3b77bcde),
	.w7(32'hbb1be6ab),
	.w8(32'hb932f5e0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a892e),
	.w1(32'hbb7012aa),
	.w2(32'hbb7db7dd),
	.w3(32'hbb1d0abe),
	.w4(32'hbb16e7cc),
	.w5(32'h3ae5a78f),
	.w6(32'h3c19174c),
	.w7(32'h3c115646),
	.w8(32'h3c159263),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b869b8c),
	.w1(32'hbc062bb3),
	.w2(32'hbbc5a2fe),
	.w3(32'h3bc09910),
	.w4(32'h3a9f258a),
	.w5(32'h3a874d0b),
	.w6(32'h3bd948b9),
	.w7(32'h3b0914f7),
	.w8(32'h3c19451a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc192308),
	.w1(32'hbb78a753),
	.w2(32'hbc1bfba7),
	.w3(32'h3b7abd86),
	.w4(32'h3bd024a9),
	.w5(32'hbab5147c),
	.w6(32'h3c1fe4d8),
	.w7(32'h3c51f2ad),
	.w8(32'h3bae9d09),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399cba7b),
	.w1(32'hbcba8daf),
	.w2(32'hbc905cbc),
	.w3(32'h3b7e266b),
	.w4(32'hbc5bd736),
	.w5(32'h3d3f7e6a),
	.w6(32'h3b9a2ecb),
	.w7(32'hbc682e62),
	.w8(32'h3cf81531),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc549e19),
	.w1(32'h3b138cf5),
	.w2(32'hbc8a9206),
	.w3(32'h3b4925ac),
	.w4(32'h3ba3d0b2),
	.w5(32'h3d252978),
	.w6(32'hbc21cb63),
	.w7(32'hbc9083f4),
	.w8(32'h3b54e877),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0bd0d2),
	.w1(32'h3a65798d),
	.w2(32'hb9a50de3),
	.w3(32'hbb095025),
	.w4(32'hbc619cd4),
	.w5(32'hbc91babe),
	.w6(32'h3bef2afc),
	.w7(32'h3b7494b0),
	.w8(32'hbc65030a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb888994),
	.w1(32'hbb92b15b),
	.w2(32'hb9977c9d),
	.w3(32'hbc89e62b),
	.w4(32'hbc40fb22),
	.w5(32'hbbdbc471),
	.w6(32'hbb9d7a79),
	.w7(32'hbbec533e),
	.w8(32'hbbe1a931),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95487f8),
	.w1(32'h3b8d62c6),
	.w2(32'h3baa1476),
	.w3(32'hbb81659b),
	.w4(32'h3983567c),
	.w5(32'hbc059876),
	.w6(32'hbb351696),
	.w7(32'hbb6ada12),
	.w8(32'hbbd385b4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83d40a),
	.w1(32'h3b8752d6),
	.w2(32'hbbb1c538),
	.w3(32'h3b3f14fa),
	.w4(32'h3b3d9561),
	.w5(32'h39b12d05),
	.w6(32'hba1f7850),
	.w7(32'h3b2a0f8b),
	.w8(32'h3bd10f9b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb59e2c),
	.w1(32'h3a3264f7),
	.w2(32'hbc325cca),
	.w3(32'h3ae915dd),
	.w4(32'hbb904719),
	.w5(32'hbb4e782e),
	.w6(32'h3b8d3726),
	.w7(32'h3b844651),
	.w8(32'hbba585e2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99002d),
	.w1(32'hbc3c39b1),
	.w2(32'hbc2209ac),
	.w3(32'hbb9a977b),
	.w4(32'hbbf29726),
	.w5(32'hbb4dbcd1),
	.w6(32'hbbb28858),
	.w7(32'h3c4b11e0),
	.w8(32'hbacac0db),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b555173),
	.w1(32'h3c3546a4),
	.w2(32'hbac2472e),
	.w3(32'hbb972229),
	.w4(32'h3ba2b19d),
	.w5(32'h3982063b),
	.w6(32'hbbd1769f),
	.w7(32'hbafa174d),
	.w8(32'h3bcf4ec8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f392b),
	.w1(32'hbb1c694e),
	.w2(32'hbbc44cf5),
	.w3(32'h3b5da362),
	.w4(32'hb9d48c39),
	.w5(32'h3b8d1dd0),
	.w6(32'hba8314c5),
	.w7(32'h3aa07d51),
	.w8(32'h3b085902),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a775e63),
	.w1(32'h3b6369a2),
	.w2(32'h3b8aabf6),
	.w3(32'hba66f491),
	.w4(32'h3c580c2a),
	.w5(32'h3c4a508a),
	.w6(32'h3bf30722),
	.w7(32'h3c93ad1e),
	.w8(32'h3bf92d87),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44c2e7),
	.w1(32'h3a067f23),
	.w2(32'h3d6a34a8),
	.w3(32'h3bc2084f),
	.w4(32'hbcae1a00),
	.w5(32'hbc8403f7),
	.w6(32'hbb9aa594),
	.w7(32'hbcc87f82),
	.w8(32'hbd386141),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75d1c3),
	.w1(32'hbb71beba),
	.w2(32'hba0e6013),
	.w3(32'h3b8bc719),
	.w4(32'hbbb38736),
	.w5(32'hbc02cf91),
	.w6(32'hbc11a987),
	.w7(32'hbbc3ba9c),
	.w8(32'hbc6932cd),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b594cdb),
	.w1(32'h3a9881eb),
	.w2(32'hbab7d183),
	.w3(32'h39f173a7),
	.w4(32'h3b82380d),
	.w5(32'h3b49d115),
	.w6(32'h39837371),
	.w7(32'h3b817ca4),
	.w8(32'hb999b3d3),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad2125),
	.w1(32'hbc37b527),
	.w2(32'hbc4aa2bd),
	.w3(32'hba1b39cd),
	.w4(32'h3a338094),
	.w5(32'hbc913905),
	.w6(32'h3b64c4d7),
	.w7(32'h3c10c885),
	.w8(32'hbc570cc6),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20e2de),
	.w1(32'hbc6cd239),
	.w2(32'hbd0fe4fd),
	.w3(32'hbb8140f7),
	.w4(32'hbca3dbe4),
	.w5(32'hbd1bb711),
	.w6(32'hbbc4cbaa),
	.w7(32'hbbe50796),
	.w8(32'hbcc4710a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae34d3),
	.w1(32'hbae303f3),
	.w2(32'h3b8ba7a8),
	.w3(32'hbd0a2163),
	.w4(32'h3b561001),
	.w5(32'h3c95c048),
	.w6(32'hbc497620),
	.w7(32'h3ba91886),
	.w8(32'h3c2edc40),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25c005),
	.w1(32'hbca18073),
	.w2(32'hbc4888ca),
	.w3(32'h3bc111ce),
	.w4(32'h3b4a829d),
	.w5(32'hbc0fddbc),
	.w6(32'h3c071b26),
	.w7(32'h3c591d13),
	.w8(32'hbbba454f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6363d8),
	.w1(32'h3a25c88c),
	.w2(32'h3bc2f2e1),
	.w3(32'h3b77a7b9),
	.w4(32'h3b376fef),
	.w5(32'hbbd1716a),
	.w6(32'hbc43725e),
	.w7(32'h3bfecf8b),
	.w8(32'h3ab71440),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24ed55),
	.w1(32'h3b92e660),
	.w2(32'h3b030a53),
	.w3(32'hbb8f509b),
	.w4(32'hb9b49d70),
	.w5(32'h3c046379),
	.w6(32'hbb3b4401),
	.w7(32'hb9c39451),
	.w8(32'h3c19b19b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe54cf),
	.w1(32'h399568cc),
	.w2(32'h3b36856f),
	.w3(32'h3bc1ca8f),
	.w4(32'h3b270182),
	.w5(32'h3c82f7a9),
	.w6(32'h3afb9e80),
	.w7(32'h3ac6d0ad),
	.w8(32'hbb2dc6fa),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51b337),
	.w1(32'h3b0899ed),
	.w2(32'h3b6d0328),
	.w3(32'h3c25ca51),
	.w4(32'hbb0c06c2),
	.w5(32'hbc0c3a2a),
	.w6(32'hbbb5050d),
	.w7(32'h3aa96970),
	.w8(32'hbb169c25),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b04ea),
	.w1(32'hbc1b2a7d),
	.w2(32'hbb0a386c),
	.w3(32'h3ae9e157),
	.w4(32'hbc032757),
	.w5(32'h3bb5d28e),
	.w6(32'h3a683d26),
	.w7(32'h3ae4d7b0),
	.w8(32'hbb748a80),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ba0fa),
	.w1(32'hbb087dd3),
	.w2(32'h3a2a6b44),
	.w3(32'hbbc35ac3),
	.w4(32'hbaf3ccc1),
	.w5(32'hbbe12948),
	.w6(32'hbb8474a2),
	.w7(32'hbc42fd10),
	.w8(32'hbc884960),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b5d01),
	.w1(32'hbb4ec3f6),
	.w2(32'hb99788dd),
	.w3(32'h3c15c22e),
	.w4(32'hbb692030),
	.w5(32'h3bc7f8a5),
	.w6(32'h3c058ba2),
	.w7(32'hbc80be7e),
	.w8(32'hbb686b9f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba833c4d),
	.w1(32'h3b815bf3),
	.w2(32'hbb988bbe),
	.w3(32'h3b3cec20),
	.w4(32'hbc1c6d0f),
	.w5(32'hbbdc73b0),
	.w6(32'h3c243e89),
	.w7(32'hbadebfa6),
	.w8(32'hbb13f6fb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3d08f),
	.w1(32'hb8910144),
	.w2(32'hbaec1e55),
	.w3(32'hbc44ce4f),
	.w4(32'hbbd125ef),
	.w5(32'hbbb01c47),
	.w6(32'hbc159ae8),
	.w7(32'h3b18bbf9),
	.w8(32'hbb840c4a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b65a7),
	.w1(32'hba6acee6),
	.w2(32'hbc2e8297),
	.w3(32'hbaac0d77),
	.w4(32'hbad06d7a),
	.w5(32'hbba48e35),
	.w6(32'hbc0d6070),
	.w7(32'hbba03e5b),
	.w8(32'hbb4ec54d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13dc3f),
	.w1(32'hbcfa28b8),
	.w2(32'hbc75ad99),
	.w3(32'hba6a05af),
	.w4(32'hbc039c95),
	.w5(32'h3bbcd5e6),
	.w6(32'hb9a0cded),
	.w7(32'hbbb6d0b2),
	.w8(32'h3ba780e4),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a471a),
	.w1(32'hbbca5231),
	.w2(32'hbb19b639),
	.w3(32'h3ba6e15f),
	.w4(32'hbb81c251),
	.w5(32'hbbbbe245),
	.w6(32'hba937398),
	.w7(32'h39872d2a),
	.w8(32'hbc2b6d7f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c09a2),
	.w1(32'h391c5322),
	.w2(32'hbb6aac4d),
	.w3(32'h3947f00d),
	.w4(32'h3b0c0775),
	.w5(32'h3ac9699d),
	.w6(32'h3c1b99f3),
	.w7(32'h3bb210d3),
	.w8(32'h3ba77b67),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91ee08),
	.w1(32'hbb266701),
	.w2(32'h3b4edb43),
	.w3(32'h3b9ec371),
	.w4(32'h3c24ea55),
	.w5(32'h3aae19e1),
	.w6(32'h3bef0215),
	.w7(32'hbb15f5d2),
	.w8(32'hbb849064),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7065c),
	.w1(32'h3bd3cb87),
	.w2(32'h3b8c29d6),
	.w3(32'hbba7a6d3),
	.w4(32'hbbc91473),
	.w5(32'h3c77a0c3),
	.w6(32'h3b8166ce),
	.w7(32'h38b6c259),
	.w8(32'h3bb17007),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c54a9),
	.w1(32'hbc6649be),
	.w2(32'hbc4dc125),
	.w3(32'h3b324cb5),
	.w4(32'hbcbee295),
	.w5(32'hbd322ae3),
	.w6(32'hbb276dcd),
	.w7(32'hbc1bcd70),
	.w8(32'hbcae9d86),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab3474),
	.w1(32'hbad40f55),
	.w2(32'hbc3e3488),
	.w3(32'hbcb7a645),
	.w4(32'h3babe850),
	.w5(32'h3abd3ab1),
	.w6(32'hbc94fa71),
	.w7(32'hbbe259df),
	.w8(32'hbb1ba200),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6e741),
	.w1(32'hba110a78),
	.w2(32'hbbada2ac),
	.w3(32'h3b9fe55c),
	.w4(32'hbbac43b9),
	.w5(32'h3b40209a),
	.w6(32'h3ce2181f),
	.w7(32'h3c30b2c7),
	.w8(32'h3b8dc6d6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0b7af),
	.w1(32'hbbb8e973),
	.w2(32'h3ada5353),
	.w3(32'hbb1ae635),
	.w4(32'hbc314826),
	.w5(32'h39c51f45),
	.w6(32'h3bf37815),
	.w7(32'hbc770100),
	.w8(32'hbc8bc516),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7348b4),
	.w1(32'hbb8c582f),
	.w2(32'h3bd609c3),
	.w3(32'hbb845c0f),
	.w4(32'h3ac63931),
	.w5(32'h3b3155b3),
	.w6(32'hbc3ac3e3),
	.w7(32'hbb8dfad0),
	.w8(32'hbb5cfa74),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade0a0b),
	.w1(32'h3b65d207),
	.w2(32'h3ac3577e),
	.w3(32'h3b2a6590),
	.w4(32'hba0b5522),
	.w5(32'hbb7a05ab),
	.w6(32'hbb4e65f2),
	.w7(32'hbc355de2),
	.w8(32'hbbeaa2ff),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb935d3f),
	.w1(32'h3bc8bbf9),
	.w2(32'hbbb6afd5),
	.w3(32'hb9db7f0b),
	.w4(32'h3c80cb9e),
	.w5(32'h3d29c81c),
	.w6(32'h3bd6ff29),
	.w7(32'hbbed27e0),
	.w8(32'h3b610626),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed8aa8),
	.w1(32'hbc06af69),
	.w2(32'hbbef3dd8),
	.w3(32'h3c19f4f0),
	.w4(32'hbab8ddb3),
	.w5(32'hbb987dc2),
	.w6(32'hb999966d),
	.w7(32'h3a1a4511),
	.w8(32'hbc020682),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27a20a),
	.w1(32'hba66aba3),
	.w2(32'h3ba507d9),
	.w3(32'h3b08d451),
	.w4(32'hb9fe3811),
	.w5(32'hbc09bb6d),
	.w6(32'hbbfca8bf),
	.w7(32'h37532605),
	.w8(32'hbbe2a8e2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a9a82),
	.w1(32'h391d8506),
	.w2(32'hbbc1c19e),
	.w3(32'h394b6063),
	.w4(32'hbaafaf66),
	.w5(32'hbc47c6e2),
	.w6(32'hbbcd222a),
	.w7(32'h3c0996d7),
	.w8(32'h3aa283ab),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b516e85),
	.w1(32'hbb772953),
	.w2(32'h39d9a2bd),
	.w3(32'hbac76bf2),
	.w4(32'hbb4017d0),
	.w5(32'h3b8c6235),
	.w6(32'hbb8372e0),
	.w7(32'hbb9cb943),
	.w8(32'hbbc61f6c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9151985),
	.w1(32'hbbb38a1a),
	.w2(32'h3ba2ae7a),
	.w3(32'h3c106830),
	.w4(32'hbbb1b8f2),
	.w5(32'hbaa477df),
	.w6(32'hbb25bca6),
	.w7(32'hbad37a89),
	.w8(32'h3a66d206),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bb081),
	.w1(32'h3bd547bb),
	.w2(32'hb9c75cd4),
	.w3(32'h3b44419d),
	.w4(32'h3b14fd7a),
	.w5(32'h3b88572c),
	.w6(32'h3bd5149f),
	.w7(32'hba9bca60),
	.w8(32'h399c18f6),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b463853),
	.w1(32'h3bdee1b6),
	.w2(32'h3c365057),
	.w3(32'hbb0fe8d3),
	.w4(32'h3a63c643),
	.w5(32'hbb451f32),
	.w6(32'h39a143fc),
	.w7(32'hbb4a8871),
	.w8(32'hbad22636),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3a199),
	.w1(32'hba82545e),
	.w2(32'hbb19b082),
	.w3(32'hbb0a28d6),
	.w4(32'hba147889),
	.w5(32'hbaa21f7a),
	.w6(32'h3b982351),
	.w7(32'h3b5a95b2),
	.w8(32'h3ac8693e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c195894),
	.w1(32'hbb834081),
	.w2(32'hbbacf948),
	.w3(32'h3b9e0951),
	.w4(32'hbb10af90),
	.w5(32'hbaef2e03),
	.w6(32'h3c01fce5),
	.w7(32'h3b3ad701),
	.w8(32'h3bc65844),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8631c),
	.w1(32'h3c29f0a8),
	.w2(32'h3bedfe12),
	.w3(32'h3b105b46),
	.w4(32'hba84bd97),
	.w5(32'hbb8be458),
	.w6(32'h3b9c69b9),
	.w7(32'h38d646e7),
	.w8(32'h3a98eca0),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05cc41),
	.w1(32'hbb63fa2e),
	.w2(32'h3a15802c),
	.w3(32'hbb28ee16),
	.w4(32'h3c10d52c),
	.w5(32'h3c161df0),
	.w6(32'hb976b15b),
	.w7(32'hbb6f3106),
	.w8(32'hbc1e1baa),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7837c),
	.w1(32'hbaa69792),
	.w2(32'hbb8e1209),
	.w3(32'h3b8b986d),
	.w4(32'h3bcb2bbd),
	.w5(32'hbc11694b),
	.w6(32'hbb332980),
	.w7(32'h3b8eda9b),
	.w8(32'h3a358588),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c2588),
	.w1(32'h3be9acc8),
	.w2(32'hbb25090b),
	.w3(32'hbb672e33),
	.w4(32'h3bd1f74b),
	.w5(32'h3956e82e),
	.w6(32'h3b7fddea),
	.w7(32'h3c5f4bec),
	.w8(32'h3b9b68af),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10af0f),
	.w1(32'hbb8c1cb8),
	.w2(32'hbb469c87),
	.w3(32'h3bbc4765),
	.w4(32'hb95bb976),
	.w5(32'h3b2fc373),
	.w6(32'h3c1c086b),
	.w7(32'hbc10eee1),
	.w8(32'hbbd2cfba),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa0c9f),
	.w1(32'h3a1c7efa),
	.w2(32'hba9b6c44),
	.w3(32'hbb478c92),
	.w4(32'hb96a0fca),
	.w5(32'hbb1a258f),
	.w6(32'hbbe0f9e8),
	.w7(32'hbaa482da),
	.w8(32'hbb806ef6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd701a),
	.w1(32'hbb5951a6),
	.w2(32'hbb2a258d),
	.w3(32'h3c01940b),
	.w4(32'h3bf7263b),
	.w5(32'h3c105238),
	.w6(32'h3b71e3fd),
	.w7(32'hbbb0779d),
	.w8(32'h3b9efc3d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7fa87),
	.w1(32'h3a3d1c17),
	.w2(32'hbb536ca5),
	.w3(32'h3c07c7e7),
	.w4(32'h3acb0002),
	.w5(32'h3a776d0d),
	.w6(32'h3aa03246),
	.w7(32'h3aa45056),
	.w8(32'h3c0da116),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb925c3b),
	.w1(32'hbc5e72ab),
	.w2(32'hbb242801),
	.w3(32'hbb595942),
	.w4(32'h3ba5011c),
	.w5(32'hbc0dc8d7),
	.w6(32'h3b314b54),
	.w7(32'h3c92b695),
	.w8(32'hbb1e2bbf),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48980f),
	.w1(32'h3b81357e),
	.w2(32'hbbff8163),
	.w3(32'hb9fdddc3),
	.w4(32'h3b5018bb),
	.w5(32'h3ce5818f),
	.w6(32'hbb99d291),
	.w7(32'h3abec8b3),
	.w8(32'h3ba7b1aa),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81e634),
	.w1(32'h3bcb7ff9),
	.w2(32'hbb4d5450),
	.w3(32'h3bc70af9),
	.w4(32'h398f3cc1),
	.w5(32'h3c62d89b),
	.w6(32'hbb3c2938),
	.w7(32'h3b644cd1),
	.w8(32'h3b4364ab),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a3afc),
	.w1(32'h3c95460c),
	.w2(32'h3d22825b),
	.w3(32'h3ac63407),
	.w4(32'h3cb6a96a),
	.w5(32'h3d85ca6d),
	.w6(32'h3b834baa),
	.w7(32'h3c86fc25),
	.w8(32'h3d1c0536),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab9c3b),
	.w1(32'h3a80e6ba),
	.w2(32'h3b820af3),
	.w3(32'h3cd7f1ca),
	.w4(32'hbbdd17eb),
	.w5(32'hba901440),
	.w6(32'h3c6f2a7f),
	.w7(32'hbb82f762),
	.w8(32'hbc1df67c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3f5a6),
	.w1(32'hbb2c9814),
	.w2(32'hbc719a36),
	.w3(32'hb9e9f2a6),
	.w4(32'hbc850ba2),
	.w5(32'hbc857932),
	.w6(32'hb7955f33),
	.w7(32'hbc675d03),
	.w8(32'hbcb97a26),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9111b),
	.w1(32'hb57a16c9),
	.w2(32'hbb456f44),
	.w3(32'h3b0eaac6),
	.w4(32'h3ba573fc),
	.w5(32'h3bc4bb4d),
	.w6(32'hbbddfc3b),
	.w7(32'hba1c38f3),
	.w8(32'h3a390a02),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb3901),
	.w1(32'hbc03dc3f),
	.w2(32'hbc7233a2),
	.w3(32'hbad0b6c1),
	.w4(32'hbc34d633),
	.w5(32'hbc447050),
	.w6(32'hbc0701aa),
	.w7(32'hbaeb23f1),
	.w8(32'hbc015180),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba649c3),
	.w1(32'hba4ad8a2),
	.w2(32'hbb9b1523),
	.w3(32'hbae1c8ae),
	.w4(32'h3bad23a0),
	.w5(32'h3c1a89a1),
	.w6(32'hbc1210b7),
	.w7(32'h3ba6b148),
	.w8(32'h3ba6a74d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9b1a4),
	.w1(32'hbc942e59),
	.w2(32'hbd3d5236),
	.w3(32'hbb40bc3c),
	.w4(32'h3b980c27),
	.w5(32'hbc1e4af3),
	.w6(32'h3c09856a),
	.w7(32'h3c410f9c),
	.w8(32'h3d0aa484),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8af5c5),
	.w1(32'hbbeeb67e),
	.w2(32'hbc65f5ea),
	.w3(32'hbb50aa6c),
	.w4(32'hbbf115d4),
	.w5(32'hbc5c279f),
	.w6(32'h3b90e720),
	.w7(32'h399173e4),
	.w8(32'hbbddc9f2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2413f),
	.w1(32'h3bb040e9),
	.w2(32'h3b594c5f),
	.w3(32'hba97eb00),
	.w4(32'h3b41871b),
	.w5(32'hbbcb0ebd),
	.w6(32'hbaea7ad6),
	.w7(32'h3b89fdfd),
	.w8(32'hbbd627a0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13dbe3),
	.w1(32'hba007c18),
	.w2(32'hbb3f2f35),
	.w3(32'h3c0f60b6),
	.w4(32'h3ab266f5),
	.w5(32'hbc298d05),
	.w6(32'h3c029d7e),
	.w7(32'h3acd91d9),
	.w8(32'h3b9e18ee),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eced2f),
	.w1(32'hbbb7790d),
	.w2(32'hbc082744),
	.w3(32'hb98c505a),
	.w4(32'hbb0e89a0),
	.w5(32'hbadded74),
	.w6(32'hbabdcca5),
	.w7(32'h38fb0302),
	.w8(32'hba16f223),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93ca7e),
	.w1(32'hbb8b21c5),
	.w2(32'h398f671b),
	.w3(32'h3b581ee1),
	.w4(32'hbb59291a),
	.w5(32'hba6bc220),
	.w6(32'h3b801094),
	.w7(32'hbb69e5a8),
	.w8(32'hbbe4b947),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f9efb),
	.w1(32'hbc33cafa),
	.w2(32'hbbd4e49e),
	.w3(32'hbb07ad48),
	.w4(32'hbc7eef31),
	.w5(32'hbc0feb05),
	.w6(32'h3b45d210),
	.w7(32'hbba1bf96),
	.w8(32'hbbf2f1c4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07161f),
	.w1(32'hb9f3ed34),
	.w2(32'h3aacaeb3),
	.w3(32'hbc4b2925),
	.w4(32'h3a7e3cec),
	.w5(32'h3c3fbb49),
	.w6(32'hba94e451),
	.w7(32'h3bc69745),
	.w8(32'h3bc3fe95),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c56e85),
	.w1(32'h3c227ccd),
	.w2(32'h3b83bdfe),
	.w3(32'h3b9d016b),
	.w4(32'h3b9bdf87),
	.w5(32'h3c0648f5),
	.w6(32'h3af9de6a),
	.w7(32'hbc247fa0),
	.w8(32'h3b99eeb2),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0493a7),
	.w1(32'hbc98414a),
	.w2(32'hbbe92d8b),
	.w3(32'hbbf79916),
	.w4(32'hbbbe7548),
	.w5(32'hbcaadd0a),
	.w6(32'h3b616734),
	.w7(32'h3abe9fe0),
	.w8(32'hbb10d740),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b17bb),
	.w1(32'hbb9cba8b),
	.w2(32'hbb8644f1),
	.w3(32'hbbb47345),
	.w4(32'hbb263f0c),
	.w5(32'hbb06f698),
	.w6(32'hbc40b01b),
	.w7(32'hbac7ef39),
	.w8(32'hb89eba59),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5cc11),
	.w1(32'h3ba9ab12),
	.w2(32'h3be6ef67),
	.w3(32'hbbc90519),
	.w4(32'hbaf98b92),
	.w5(32'h3c21f685),
	.w6(32'hbb0e1d12),
	.w7(32'hb905d325),
	.w8(32'hba466cad),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f7aae),
	.w1(32'h3b4b2a7a),
	.w2(32'h3c4de138),
	.w3(32'hbb49295f),
	.w4(32'h3c77373f),
	.w5(32'h3ca672c7),
	.w6(32'h3b1dfe19),
	.w7(32'h3c225137),
	.w8(32'h3ca45581),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f2009),
	.w1(32'h3c76ddd9),
	.w2(32'h3cfa4260),
	.w3(32'h3c5f7e61),
	.w4(32'h3c5847e1),
	.w5(32'h3d371a22),
	.w6(32'h3c89b6f1),
	.w7(32'h3a93ffa3),
	.w8(32'h3c925f0a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62ad63),
	.w1(32'hbb9d8734),
	.w2(32'hbbb2c6f3),
	.w3(32'h3cc4f471),
	.w4(32'h3b81f5e3),
	.w5(32'h3bb136e3),
	.w6(32'h3c82d940),
	.w7(32'h3b8e7427),
	.w8(32'h3c195900),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb4856),
	.w1(32'h3c145eb2),
	.w2(32'hbb00d67f),
	.w3(32'h3a1b1cc9),
	.w4(32'hbb94471e),
	.w5(32'h3d01b4b6),
	.w6(32'h3c0deb01),
	.w7(32'hbca2da29),
	.w8(32'hbc31d154),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc816994),
	.w1(32'hbc2508f1),
	.w2(32'hbb883ab3),
	.w3(32'h3ba472e5),
	.w4(32'hbbc37741),
	.w5(32'hba40e1c0),
	.w6(32'h3c31e2f3),
	.w7(32'hbb8a7216),
	.w8(32'hbb37314c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85ae42),
	.w1(32'h3b4f6801),
	.w2(32'h3b0181fc),
	.w3(32'h3b9e84a9),
	.w4(32'h3c1eeccc),
	.w5(32'h3ae9b4c5),
	.w6(32'h3ad9220b),
	.w7(32'h39a56a43),
	.w8(32'h3bbdf2e8),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb238473),
	.w1(32'hba83b9b1),
	.w2(32'hbb37cc0f),
	.w3(32'hbb9dbdc1),
	.w4(32'h3c1a2eac),
	.w5(32'h3a70cdf0),
	.w6(32'h3ae5d6fa),
	.w7(32'h3c15780e),
	.w8(32'h3c4bf7fb),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b588b),
	.w1(32'hba5f64ec),
	.w2(32'hbc0a1dd7),
	.w3(32'hbb4393ed),
	.w4(32'h3b0276cb),
	.w5(32'h3b315ef7),
	.w6(32'h3bda88a7),
	.w7(32'h3b967d6e),
	.w8(32'hbad2389a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a814cc7),
	.w1(32'hb9ab44e7),
	.w2(32'hbb9b93c3),
	.w3(32'hba8d86a0),
	.w4(32'h3be94f8c),
	.w5(32'h3bc00709),
	.w6(32'hbb61b95e),
	.w7(32'hb9cf694b),
	.w8(32'hbb64235a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4a66e),
	.w1(32'hbbea6629),
	.w2(32'hbc4a7a41),
	.w3(32'h3c1b3662),
	.w4(32'hbb98604e),
	.w5(32'hbc99137d),
	.w6(32'h3abb1193),
	.w7(32'h3beae3da),
	.w8(32'hbc84ba5a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c386676),
	.w1(32'hbb05fa30),
	.w2(32'h3c0eed3d),
	.w3(32'hbab3cf3e),
	.w4(32'hbaf271a4),
	.w5(32'h3b447c0a),
	.w6(32'hbc5e2311),
	.w7(32'h3bf9aed6),
	.w8(32'h3c7d518d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf39791),
	.w1(32'hbb6b8356),
	.w2(32'h3a98df72),
	.w3(32'hbb6b2e56),
	.w4(32'hbb002d06),
	.w5(32'hbad81112),
	.w6(32'hba53c571),
	.w7(32'h3ba33f2d),
	.w8(32'h3b24fd36),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba185d0a),
	.w1(32'h3bbf4a00),
	.w2(32'h3bcb73cd),
	.w3(32'hbb75135c),
	.w4(32'hbb399a7d),
	.w5(32'h3ab7e4de),
	.w6(32'h3acc31cd),
	.w7(32'h3b9a8292),
	.w8(32'h3bc9e97d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59dac0),
	.w1(32'hba17029d),
	.w2(32'hbb8c5ad2),
	.w3(32'hbb6c7ef8),
	.w4(32'hbb1f5992),
	.w5(32'hbc089972),
	.w6(32'h3c004819),
	.w7(32'h3abf4a8c),
	.w8(32'h3ba8ca13),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc9e59),
	.w1(32'h3b7e3c77),
	.w2(32'hbaceedfd),
	.w3(32'hb8063326),
	.w4(32'h3b6e76b3),
	.w5(32'h3c23a3fb),
	.w6(32'hbb1866ed),
	.w7(32'hbc252b3e),
	.w8(32'hbbbf84bc),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba06412),
	.w1(32'h38fcd5dd),
	.w2(32'hbbae1358),
	.w3(32'hb911c8ad),
	.w4(32'hbc364451),
	.w5(32'h3baf1af7),
	.w6(32'hbb98c66a),
	.w7(32'hbc145176),
	.w8(32'hbc7978a2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9caf89),
	.w1(32'hbaac315f),
	.w2(32'hba207026),
	.w3(32'hbb3b3762),
	.w4(32'h391e1fc6),
	.w5(32'h3a0ac58a),
	.w6(32'hbc1a7e67),
	.w7(32'h3852524f),
	.w8(32'h3b77bef4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b24afe),
	.w1(32'h3b13cf38),
	.w2(32'h3ae2b5f5),
	.w3(32'hbb61de82),
	.w4(32'hbb63714e),
	.w5(32'hbb80aace),
	.w6(32'hb9ad9d71),
	.w7(32'h3ab4c964),
	.w8(32'h3bd28f79),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f5845),
	.w1(32'hba4fd880),
	.w2(32'hbaa3b910),
	.w3(32'h3b0306c0),
	.w4(32'h39ad19fb),
	.w5(32'hb9eca8ec),
	.w6(32'h3bff7991),
	.w7(32'hbb01a08f),
	.w8(32'hbba64410),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c255e),
	.w1(32'h3b19940d),
	.w2(32'h3ba34b99),
	.w3(32'hb9510fda),
	.w4(32'h3b6847f0),
	.w5(32'hbb68deae),
	.w6(32'hbaf564eb),
	.w7(32'hb8d848f1),
	.w8(32'h3b915a14),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd56ae),
	.w1(32'hbb5aaa3b),
	.w2(32'h3affa577),
	.w3(32'hbbb7b4c6),
	.w4(32'hbb444838),
	.w5(32'hbabcfdab),
	.w6(32'h3c0f0f1b),
	.w7(32'hbb28a112),
	.w8(32'hbb3a491b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1530ab),
	.w1(32'hba423113),
	.w2(32'hbb9027f0),
	.w3(32'h3ae4a47d),
	.w4(32'h3a184d0e),
	.w5(32'h3c001122),
	.w6(32'hbb9fbaa9),
	.w7(32'h3bea0724),
	.w8(32'h3a399a72),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a8fda),
	.w1(32'hbbd72c76),
	.w2(32'hbb1d84ec),
	.w3(32'h3c1c8f95),
	.w4(32'h3ab65937),
	.w5(32'h3ab25b1e),
	.w6(32'hb912d2cc),
	.w7(32'h3c41da01),
	.w8(32'hba902469),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39003da7),
	.w1(32'h3b975de4),
	.w2(32'h3b5c5e71),
	.w3(32'h3c0eec46),
	.w4(32'h3b9b9d2f),
	.w5(32'h3b3de459),
	.w6(32'hbaa158f5),
	.w7(32'h3b6a5490),
	.w8(32'h3b822a22),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5557d),
	.w1(32'h3b1d6352),
	.w2(32'h3a86464b),
	.w3(32'h3b76f537),
	.w4(32'hbaf26d85),
	.w5(32'hbb4ff483),
	.w6(32'h3bb42447),
	.w7(32'hbbb54255),
	.w8(32'hbb077548),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b093408),
	.w1(32'hbbd0957f),
	.w2(32'hbc093d9d),
	.w3(32'h39ee8305),
	.w4(32'hbb19c933),
	.w5(32'h3bee72b4),
	.w6(32'hbaad2d34),
	.w7(32'h3bbf88c5),
	.w8(32'hbaf7bacb),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9917fc3),
	.w1(32'hbc09ae5a),
	.w2(32'hbbfbf0af),
	.w3(32'h3a77a927),
	.w4(32'hba816a16),
	.w5(32'hbbc64504),
	.w6(32'hbba154cf),
	.w7(32'hba214e77),
	.w8(32'hbaffe5bb),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec13c2),
	.w1(32'h3b043670),
	.w2(32'h3b87a039),
	.w3(32'hbc13440b),
	.w4(32'hbb07a5d8),
	.w5(32'h3b5886d9),
	.w6(32'h3b609a76),
	.w7(32'h3b85137b),
	.w8(32'h3ba1401d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a316f6b),
	.w1(32'h3b0a860b),
	.w2(32'hbaa89be1),
	.w3(32'h3b9ef6c8),
	.w4(32'h3b2c0d08),
	.w5(32'h3b1fa074),
	.w6(32'h3b647451),
	.w7(32'hb9a1963e),
	.w8(32'h3915633e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b799e0d),
	.w1(32'hbb2e8654),
	.w2(32'hbaf29007),
	.w3(32'h3adacce3),
	.w4(32'hba8e71b1),
	.w5(32'h3a7182ca),
	.w6(32'h3b0f7762),
	.w7(32'hbb369907),
	.w8(32'hbb5e0a0a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc692a),
	.w1(32'hb9f1e792),
	.w2(32'h3a0648ce),
	.w3(32'hbb7ed11f),
	.w4(32'h3a4787c0),
	.w5(32'hba06ee18),
	.w6(32'hbb6ad97a),
	.w7(32'h38a6e176),
	.w8(32'h3bb913d1),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd56873),
	.w1(32'hbbb23bc8),
	.w2(32'h3b40eff2),
	.w3(32'hbb0aa709),
	.w4(32'hbb3429fb),
	.w5(32'hbb01f946),
	.w6(32'h3bef1a02),
	.w7(32'h3a9b7b95),
	.w8(32'hbbe30b69),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e9b37),
	.w1(32'hbbd69cd2),
	.w2(32'hbbb86585),
	.w3(32'hba50cd35),
	.w4(32'hbb898941),
	.w5(32'hbbb053d7),
	.w6(32'h3aea7c9f),
	.w7(32'h3b000431),
	.w8(32'h3aa3906d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7edd70),
	.w1(32'hbb36ff99),
	.w2(32'hbac5b76d),
	.w3(32'hbb620c6a),
	.w4(32'hbb74a406),
	.w5(32'hbacdf4e0),
	.w6(32'hbb06144c),
	.w7(32'h39ae6899),
	.w8(32'hbb1ffdc3),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb766ca2),
	.w1(32'hbb8dc2fd),
	.w2(32'h3aa72898),
	.w3(32'h3a8a9d67),
	.w4(32'h3b09fb2a),
	.w5(32'h3bb07ba5),
	.w6(32'hbb1f68a5),
	.w7(32'hb927dc0a),
	.w8(32'hbb7ddb20),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a932fb0),
	.w1(32'hbb3b889c),
	.w2(32'hbbbf65c4),
	.w3(32'h382ba593),
	.w4(32'hbad08ee6),
	.w5(32'h3c74379b),
	.w6(32'h3a182c9b),
	.w7(32'h3c6e0ce2),
	.w8(32'h3c03f5cb),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21f511),
	.w1(32'h3a883bfd),
	.w2(32'hb953284d),
	.w3(32'h3cb2748f),
	.w4(32'h39bb9c90),
	.w5(32'h3a05be76),
	.w6(32'hbaeb29d6),
	.w7(32'h3ab094ae),
	.w8(32'h3af63320),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc2ed5),
	.w1(32'hbb63d5c9),
	.w2(32'hbb33b950),
	.w3(32'hb9edb03f),
	.w4(32'hbbc234e8),
	.w5(32'hbbb4a212),
	.w6(32'h3bb097e8),
	.w7(32'hba48e53d),
	.w8(32'hba639869),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa324b),
	.w1(32'hba925f2c),
	.w2(32'hba25a0c3),
	.w3(32'hbbc4e98f),
	.w4(32'hbb8a9123),
	.w5(32'hba3bb001),
	.w6(32'h3b85e9f4),
	.w7(32'h3bba41eb),
	.w8(32'h3b76b715),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d5559),
	.w1(32'hbb2e6395),
	.w2(32'hbac5b42b),
	.w3(32'hbb599fdc),
	.w4(32'hbb18dd22),
	.w5(32'hbbdd5349),
	.w6(32'hbb394c38),
	.w7(32'h3acec247),
	.w8(32'hbb82ebb9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaca12),
	.w1(32'h3ad7d58d),
	.w2(32'h3b53fe84),
	.w3(32'h3a4bdc70),
	.w4(32'hb9a6332f),
	.w5(32'hbbc9ab3c),
	.w6(32'h3aee594c),
	.w7(32'hbbd87a00),
	.w8(32'hbbaaf112),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a55cf9),
	.w1(32'h3b9004ea),
	.w2(32'hbacc3209),
	.w3(32'hbbb265c5),
	.w4(32'h3b1b96cd),
	.w5(32'h39888cff),
	.w6(32'hba1c4708),
	.w7(32'hba4b7d6c),
	.w8(32'hb9367e64),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb9c4a),
	.w1(32'hbb48f1a7),
	.w2(32'h3b487dcb),
	.w3(32'hb8990bad),
	.w4(32'hbb822c1a),
	.w5(32'h3b0c7c2b),
	.w6(32'h3b285208),
	.w7(32'hbb562fa2),
	.w8(32'hbc1fa0e5),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf74ec6),
	.w1(32'hbaf53ddf),
	.w2(32'hbbdcca73),
	.w3(32'h3b4730c5),
	.w4(32'hbb0cf0a2),
	.w5(32'h3c0ad7dd),
	.w6(32'hbb2a7267),
	.w7(32'h3ba59a2d),
	.w8(32'hb99282b6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ab497),
	.w1(32'h3a3b8038),
	.w2(32'hbbee7ccb),
	.w3(32'h3c74bea8),
	.w4(32'hbbf5c252),
	.w5(32'h3a6cfc98),
	.w6(32'hbb658642),
	.w7(32'h3c1b2c91),
	.w8(32'h3b6e3941),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24d2b6),
	.w1(32'hbad9f1f1),
	.w2(32'hbb2a8ddb),
	.w3(32'h3c386a80),
	.w4(32'hbbb166b8),
	.w5(32'hbb987129),
	.w6(32'hbba637ff),
	.w7(32'hbbbf8dc1),
	.w8(32'hbad1ca23),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60ab8d),
	.w1(32'h3b398738),
	.w2(32'hba229005),
	.w3(32'hbb3b8081),
	.w4(32'hbbafae91),
	.w5(32'hbb5feffd),
	.w6(32'hbacbfa27),
	.w7(32'h3ad91f78),
	.w8(32'h3b4fc01b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b7645),
	.w1(32'hbb95c901),
	.w2(32'hbbc071ad),
	.w3(32'h39e68017),
	.w4(32'hbb683152),
	.w5(32'hbb145d99),
	.w6(32'h3b09f0cd),
	.w7(32'hba4c445e),
	.w8(32'hbc389e21),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59c312),
	.w1(32'hba45b096),
	.w2(32'hbb46332e),
	.w3(32'hb9e8b679),
	.w4(32'hbbfcb8ae),
	.w5(32'hba759f1f),
	.w6(32'hbadf03c1),
	.w7(32'h3bf4c72c),
	.w8(32'h3bdfe2eb),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb418b08),
	.w1(32'hbae366f7),
	.w2(32'hbbbc6545),
	.w3(32'h3c079b97),
	.w4(32'hbb4c4fc2),
	.w5(32'hba71c57f),
	.w6(32'h3af9a8e6),
	.w7(32'hbc01f991),
	.w8(32'hbc0a57d5),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54e6fb),
	.w1(32'hbb00fb06),
	.w2(32'hbb763bb9),
	.w3(32'hba23e50e),
	.w4(32'hbc3edbf7),
	.w5(32'hb9a69dd2),
	.w6(32'h3b3a86d0),
	.w7(32'h3c9b1e21),
	.w8(32'h3c8ba65a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1de63),
	.w1(32'hbb579301),
	.w2(32'hbabe24b0),
	.w3(32'h3c67281c),
	.w4(32'hbb8f11ed),
	.w5(32'hbac9d64f),
	.w6(32'h3ba10f4f),
	.w7(32'h39b10d69),
	.w8(32'hbb808bd3),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c55d7),
	.w1(32'hba51ef2e),
	.w2(32'h3ba43697),
	.w3(32'h3ae32e85),
	.w4(32'h3aeb37cd),
	.w5(32'hbb8e486f),
	.w6(32'hbbb9e48f),
	.w7(32'hbba0f254),
	.w8(32'h3b584f1b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a614b02),
	.w1(32'h3a37ea7c),
	.w2(32'hba588e38),
	.w3(32'hbbf05d95),
	.w4(32'hbb348f51),
	.w5(32'hba05ddff),
	.w6(32'h3bbe6d40),
	.w7(32'h3ad11010),
	.w8(32'h3b6fc90c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35160d),
	.w1(32'h3a1e5eb9),
	.w2(32'h3b524876),
	.w3(32'hbb06793a),
	.w4(32'h3b0706f8),
	.w5(32'h394af02a),
	.w6(32'h3aa0383a),
	.w7(32'hbb10a8a1),
	.w8(32'hbacc11b5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0e506),
	.w1(32'h38d4b74d),
	.w2(32'hb94bd2ff),
	.w3(32'hbbf42ad8),
	.w4(32'h38a18029),
	.w5(32'hbb2acee7),
	.w6(32'h39ed7803),
	.w7(32'hbb8ea042),
	.w8(32'h3ae6a920),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7ae52),
	.w1(32'h3b1b8c5d),
	.w2(32'h3ad86b71),
	.w3(32'hba6638a9),
	.w4(32'h38c2b11f),
	.w5(32'hbb744ff6),
	.w6(32'h3b33011f),
	.w7(32'hbad68b29),
	.w8(32'h3a8737c2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a878bc5),
	.w1(32'hba279621),
	.w2(32'h3ac5f97a),
	.w3(32'hb95d047a),
	.w4(32'hbb3b596e),
	.w5(32'hbba241ed),
	.w6(32'h3a388d64),
	.w7(32'hbb7eef72),
	.w8(32'h3ac63608),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d9e4b),
	.w1(32'h3b6d329d),
	.w2(32'h39dc9baf),
	.w3(32'hb8d21d44),
	.w4(32'h3996325b),
	.w5(32'h3982e821),
	.w6(32'hba8e6e9f),
	.w7(32'hbb9a3dc8),
	.w8(32'hbb65e717),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35e3b8),
	.w1(32'h3bd19e71),
	.w2(32'hbaa857ff),
	.w3(32'hbbabe1a6),
	.w4(32'hbb2f63e8),
	.w5(32'hbbcf7bba),
	.w6(32'hbb5a8d4f),
	.w7(32'hbbb4bbeb),
	.w8(32'hbb4aa404),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd9e99),
	.w1(32'hbb2ba82d),
	.w2(32'hbb93289e),
	.w3(32'hbb4f35f4),
	.w4(32'hbb92a27e),
	.w5(32'h3c2666dc),
	.w6(32'h3ada7545),
	.w7(32'h3c063d67),
	.w8(32'h3b5798ab),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07a7e0),
	.w1(32'hbbce6cf0),
	.w2(32'h39294d9c),
	.w3(32'h3c7dcfe7),
	.w4(32'h3c4b6fc3),
	.w5(32'hbb2d9abb),
	.w6(32'hbb3a7002),
	.w7(32'hbbbd08dd),
	.w8(32'h3b8bdfd5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ecf74),
	.w1(32'hb93abc57),
	.w2(32'h3aae177d),
	.w3(32'hbb97ef61),
	.w4(32'hbb333390),
	.w5(32'hbba07522),
	.w6(32'hba74d91c),
	.w7(32'hbae6969a),
	.w8(32'h39e7402a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e38fba),
	.w1(32'hbb0c23fc),
	.w2(32'hbb4ad8e7),
	.w3(32'hbbb3528d),
	.w4(32'hb9d530fd),
	.w5(32'h3b4b6eb0),
	.w6(32'h3b2de564),
	.w7(32'hbb80ee89),
	.w8(32'h3ae2829e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03d4a4),
	.w1(32'h3a0635b4),
	.w2(32'h3b1f7343),
	.w3(32'h3b57a4ab),
	.w4(32'hbb5e7fe9),
	.w5(32'hbb1ebd9f),
	.w6(32'h3ae1d371),
	.w7(32'hba9ff3d4),
	.w8(32'hbb39e4d4),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94b704),
	.w1(32'h3bb654d1),
	.w2(32'h3b017dcf),
	.w3(32'hbb136755),
	.w4(32'hbab8cc76),
	.w5(32'hbc065ef3),
	.w6(32'hba611f79),
	.w7(32'hbbbe6705),
	.w8(32'h38bc7af3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31c272),
	.w1(32'hbbfc77c0),
	.w2(32'hbc48c19f),
	.w3(32'hbc4d57bd),
	.w4(32'hbb3f93a0),
	.w5(32'h3c82dcbf),
	.w6(32'h3b20aba0),
	.w7(32'h3c2f7255),
	.w8(32'h3b4a1ff5),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e71da),
	.w1(32'hbbbb72f7),
	.w2(32'hba0054c0),
	.w3(32'h3c6ca296),
	.w4(32'h3a427f57),
	.w5(32'hba50b1dc),
	.w6(32'hbb1c9a5f),
	.w7(32'hbb29f9ac),
	.w8(32'hbb2c6dc4),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1324e),
	.w1(32'h3ac1efbc),
	.w2(32'h3be88667),
	.w3(32'h3aec4505),
	.w4(32'h3b9bfc7a),
	.w5(32'h3b0f8f74),
	.w6(32'hbb0a12dc),
	.w7(32'h397ce5b6),
	.w8(32'h3aba5614),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f439a),
	.w1(32'hbb2f08c4),
	.w2(32'hbbb63eb7),
	.w3(32'h3a14eee3),
	.w4(32'hbbcee64e),
	.w5(32'hbabe8746),
	.w6(32'h3b273096),
	.w7(32'h3b33ed2e),
	.w8(32'hba546b6b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba504250),
	.w1(32'h3ad69ffd),
	.w2(32'hb9ce390c),
	.w3(32'h3b8bd62b),
	.w4(32'hba9bba5d),
	.w5(32'h3c578ea6),
	.w6(32'h3a3b95a6),
	.w7(32'h3bc9dc66),
	.w8(32'h3b4585d1),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd951f8),
	.w1(32'h3b56d384),
	.w2(32'hbb80a605),
	.w3(32'h3c7ee870),
	.w4(32'hba5598da),
	.w5(32'h3b4d87f6),
	.w6(32'h3a93be44),
	.w7(32'h3ac877da),
	.w8(32'hbb63e89b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba92228),
	.w1(32'h3b200cbb),
	.w2(32'h3b934083),
	.w3(32'h3bdacdcd),
	.w4(32'hbb71a67e),
	.w5(32'hbbe9e2a2),
	.w6(32'hbb5321ad),
	.w7(32'hbb96565e),
	.w8(32'h37b3e690),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1519c5),
	.w1(32'hb9a1ba77),
	.w2(32'h3b2e683c),
	.w3(32'hbbc017b7),
	.w4(32'h3c030238),
	.w5(32'hb9e5e9fb),
	.w6(32'h3b6bf60b),
	.w7(32'hbb922ea7),
	.w8(32'h3bcc54c2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ee59b0),
	.w1(32'h3b6b21ec),
	.w2(32'h3b0d67ce),
	.w3(32'hba233234),
	.w4(32'hba92f3be),
	.w5(32'hbbbba108),
	.w6(32'h3b6bab3f),
	.w7(32'h3b4046bc),
	.w8(32'hba659a76),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cbbd7),
	.w1(32'hbb94aaa9),
	.w2(32'hbbe11321),
	.w3(32'hbaf0034c),
	.w4(32'hbacb25db),
	.w5(32'hbb34dea0),
	.w6(32'h3b8dbd4d),
	.w7(32'h3bdfc31b),
	.w8(32'h3ab0cec5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule