module layer_10_featuremap_270(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9df81b),
	.w1(32'hbbe14e5b),
	.w2(32'hba992a29),
	.w3(32'hbc28ffa3),
	.w4(32'hbb6f0d91),
	.w5(32'hbbc17e22),
	.w6(32'hbad45257),
	.w7(32'h3983b9a1),
	.w8(32'h3b598d8d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bfc4b),
	.w1(32'hbba4ea92),
	.w2(32'hbc3ffe42),
	.w3(32'hbac63603),
	.w4(32'hbb0f5760),
	.w5(32'hba0fc688),
	.w6(32'h3b4ce151),
	.w7(32'hbc3005ce),
	.w8(32'hbae176ea),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70aa2a),
	.w1(32'hbc40f5da),
	.w2(32'h3b94eb7c),
	.w3(32'hbbcfa84e),
	.w4(32'h3a05d515),
	.w5(32'hbb53cf35),
	.w6(32'hbc4b5b7e),
	.w7(32'hbb7b6151),
	.w8(32'hbb9b8196),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab90fa2),
	.w1(32'hbafad56e),
	.w2(32'hb8c83e5a),
	.w3(32'hbb2ee150),
	.w4(32'hba1d5bed),
	.w5(32'h3bc72a7a),
	.w6(32'hbbc54eea),
	.w7(32'hbb3b732a),
	.w8(32'h3aea993e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aafc99),
	.w1(32'h3a8d0a29),
	.w2(32'h3c36e37a),
	.w3(32'h3c403bc4),
	.w4(32'h3c24c9ae),
	.w5(32'hbb8f2edb),
	.w6(32'h3c2498c7),
	.w7(32'h3c511ec2),
	.w8(32'hbb759f0d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4afc04),
	.w1(32'hbb5125b4),
	.w2(32'h39ab9ef0),
	.w3(32'hbba3b8fd),
	.w4(32'hbab4646d),
	.w5(32'hba81ea87),
	.w6(32'hbb442c31),
	.w7(32'hbb1b820f),
	.w8(32'hbb1489fc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4406de),
	.w1(32'hbb9808dc),
	.w2(32'hba742ec9),
	.w3(32'hbb96f07f),
	.w4(32'hba96b226),
	.w5(32'hbb79fe56),
	.w6(32'hbbd3aa2b),
	.w7(32'hbbba7bdf),
	.w8(32'hbbf72705),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5f98e),
	.w1(32'hbc463837),
	.w2(32'hbc2008b7),
	.w3(32'hbc4c06f1),
	.w4(32'hbbd789cf),
	.w5(32'hbc23a71d),
	.w6(32'hbc672cc1),
	.w7(32'hbc66eb22),
	.w8(32'hbc686e41),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f1e93),
	.w1(32'hbc89038b),
	.w2(32'hbc430310),
	.w3(32'hbc62f2b9),
	.w4(32'hbc482a7e),
	.w5(32'hbbc8a258),
	.w6(32'hbc4301b0),
	.w7(32'hbc70add6),
	.w8(32'hbbaec878),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30352a),
	.w1(32'hbb311780),
	.w2(32'hb985e717),
	.w3(32'hbb802301),
	.w4(32'hba9d3c2a),
	.w5(32'hbb085504),
	.w6(32'hbb11d3d1),
	.w7(32'hb9a4d13d),
	.w8(32'hbb0c78b6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5194ba),
	.w1(32'h39b4f695),
	.w2(32'h39ad32b6),
	.w3(32'hbb8ec11a),
	.w4(32'hb92840be),
	.w5(32'h3ba184e6),
	.w6(32'hbb5ddf13),
	.w7(32'hb9063d16),
	.w8(32'hbb88865c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcefabd),
	.w1(32'hbb30074a),
	.w2(32'h3bdf81e2),
	.w3(32'h3bbfd34f),
	.w4(32'h3bd763f0),
	.w5(32'h3b919bd5),
	.w6(32'hbc3912fc),
	.w7(32'h38fbf506),
	.w8(32'h3ba4d110),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d6856a),
	.w1(32'hbab9e265),
	.w2(32'h3aa96fc4),
	.w3(32'h3c4841a3),
	.w4(32'h3bf4559b),
	.w5(32'h3b45d26d),
	.w6(32'h3c2b834a),
	.w7(32'h3bf75c8a),
	.w8(32'h3bcb4ec7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0105aa),
	.w1(32'h3b928b53),
	.w2(32'h3b9ce71b),
	.w3(32'h3b5b8be8),
	.w4(32'hbb861018),
	.w5(32'h3b62634f),
	.w6(32'h3bc7e137),
	.w7(32'h3b53f786),
	.w8(32'hba66e898),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1163c8),
	.w1(32'hbba14e5c),
	.w2(32'h3b5a1b06),
	.w3(32'hbaa2ab37),
	.w4(32'h39a40e3e),
	.w5(32'hbb970c55),
	.w6(32'hbb9298f1),
	.w7(32'hbb375f72),
	.w8(32'h3a9b2dfe),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb942273),
	.w1(32'hbba887d3),
	.w2(32'h38b3de00),
	.w3(32'hbb7a2e99),
	.w4(32'h3abae9ce),
	.w5(32'hbbfefadd),
	.w6(32'h3bda4fc5),
	.w7(32'h3a54fd7d),
	.w8(32'hbb947bee),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa94d65),
	.w1(32'hbb44c7e5),
	.w2(32'hbb4cad34),
	.w3(32'hbc06a975),
	.w4(32'hbb9e705b),
	.w5(32'h3bafb265),
	.w6(32'hba9c8edd),
	.w7(32'hbc2b5daa),
	.w8(32'h3aa24511),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb027e67),
	.w1(32'h3b1366d0),
	.w2(32'h3c03fa6f),
	.w3(32'h3c09b1ce),
	.w4(32'h3bd1d51b),
	.w5(32'hba7d183f),
	.w6(32'hbc17f316),
	.w7(32'h3c0b2463),
	.w8(32'hbc165da9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b824cd7),
	.w1(32'h3c689de4),
	.w2(32'h3c61dda7),
	.w3(32'hba4ee3b7),
	.w4(32'hbb1d6dd0),
	.w5(32'h3a827f29),
	.w6(32'hbc7ec7e1),
	.w7(32'h3c465427),
	.w8(32'h39f4c19e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2faa8f),
	.w1(32'hbb1daa1d),
	.w2(32'hbb3556a4),
	.w3(32'hbb22d28c),
	.w4(32'hbafb57e1),
	.w5(32'hbb12f652),
	.w6(32'hbb36fc2b),
	.w7(32'hbb0c7e64),
	.w8(32'hba0b4913),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb101056),
	.w1(32'hbb8bd1cf),
	.w2(32'hbba6de3d),
	.w3(32'hba2ec747),
	.w4(32'hbb9f1510),
	.w5(32'hbb392d29),
	.w6(32'h3b5a9d23),
	.w7(32'hbb05f7b9),
	.w8(32'hbbf1c6fc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813037),
	.w1(32'hbb21fa48),
	.w2(32'hbb6b4e67),
	.w3(32'hba3573b8),
	.w4(32'hbb1568eb),
	.w5(32'hbbc3234f),
	.w6(32'hba5bd5ef),
	.w7(32'hbb65c8ac),
	.w8(32'hbbc33fcd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d9a84),
	.w1(32'hba948e71),
	.w2(32'hbbb1f366),
	.w3(32'hbc0702b4),
	.w4(32'hbbcc9eda),
	.w5(32'hbbe41468),
	.w6(32'hbc57b8b0),
	.w7(32'h3af391f4),
	.w8(32'hbc0a71a1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b7e47),
	.w1(32'hbbf5f0a8),
	.w2(32'hbc561333),
	.w3(32'hb8f33a7a),
	.w4(32'hbbde9191),
	.w5(32'h3b0bd20c),
	.w6(32'h3b4a151b),
	.w7(32'hbbd69919),
	.w8(32'h3aaf3b81),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16bf4b),
	.w1(32'hbc2266cd),
	.w2(32'hbb84d38f),
	.w3(32'h3baaf94b),
	.w4(32'hbb7481e1),
	.w5(32'hba85ed5d),
	.w6(32'h3b72adb7),
	.w7(32'hbaf7d316),
	.w8(32'hbb46dd28),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0760f),
	.w1(32'hbb501582),
	.w2(32'h3ba83c05),
	.w3(32'hbb9cc82f),
	.w4(32'h3a5c1bf9),
	.w5(32'h3b1000b4),
	.w6(32'hbbc5a0c9),
	.w7(32'hbb749076),
	.w8(32'hb8afee38),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41826d),
	.w1(32'hbba93a97),
	.w2(32'h3b455948),
	.w3(32'hbbc80c8e),
	.w4(32'h3b090464),
	.w5(32'hbb81df07),
	.w6(32'hbbd51a7e),
	.w7(32'hbb836ea9),
	.w8(32'hbb4e3c18),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6698f5),
	.w1(32'hbbe1b539),
	.w2(32'hbb48b9e5),
	.w3(32'hbbcb13a8),
	.w4(32'hbb97071c),
	.w5(32'hbc1a85a1),
	.w6(32'hba1fa32e),
	.w7(32'hbbb0ceae),
	.w8(32'hbaca6b56),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc189bc1),
	.w1(32'hbb931685),
	.w2(32'hb98df44d),
	.w3(32'hbba40b6f),
	.w4(32'hbac8e79c),
	.w5(32'h3b0d54bc),
	.w6(32'hbae96134),
	.w7(32'h3af999a7),
	.w8(32'hbaa7eda5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ea46d),
	.w1(32'hbb6b82b0),
	.w2(32'hbb991923),
	.w3(32'h3a3a3134),
	.w4(32'hb8dc437f),
	.w5(32'h3c1e3ffe),
	.w6(32'h3be1d6e6),
	.w7(32'hbb0b83dc),
	.w8(32'h3b7e5f44),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c78f6f),
	.w1(32'h3bf5c4db),
	.w2(32'h3bc77c03),
	.w3(32'h3b58a22e),
	.w4(32'h3ba47b41),
	.w5(32'hbc07138b),
	.w6(32'hbb68c64b),
	.w7(32'h3c248b99),
	.w8(32'hbbcf0c02),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd55d1d),
	.w1(32'hbb08c354),
	.w2(32'hbb2bd5dc),
	.w3(32'h3a1618f5),
	.w4(32'h3b24852a),
	.w5(32'h3c507670),
	.w6(32'hbc1f858a),
	.w7(32'hbb9f7d8e),
	.w8(32'h39990a03),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c0600),
	.w1(32'hba86f28d),
	.w2(32'h3c0e302b),
	.w3(32'hba268235),
	.w4(32'hbb8f1ae5),
	.w5(32'h3b7880cc),
	.w6(32'hbce8d5ce),
	.w7(32'h3b3537b5),
	.w8(32'h3b6d9d31),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e77ddb),
	.w1(32'h3b98bfad),
	.w2(32'h39459742),
	.w3(32'h3b980d29),
	.w4(32'h3ae4bddd),
	.w5(32'h3ab62813),
	.w6(32'hbc161f58),
	.w7(32'h3a2e7daa),
	.w8(32'hbbb59096),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24378d),
	.w1(32'hb9a26c57),
	.w2(32'h3b2bc82e),
	.w3(32'h3b7f8e58),
	.w4(32'h3b389859),
	.w5(32'h3c2b3f62),
	.w6(32'h3a202ca9),
	.w7(32'h3b8d4420),
	.w8(32'h3c2a3ccc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c131f7f),
	.w1(32'h3bcaf1eb),
	.w2(32'h3c391dcd),
	.w3(32'h3c1ab9b3),
	.w4(32'h3b3073e2),
	.w5(32'h3a276c51),
	.w6(32'hbc0ae8f7),
	.w7(32'h3c1febc2),
	.w8(32'hbbde779b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a1bae),
	.w1(32'h3c041fd3),
	.w2(32'h3b0b1682),
	.w3(32'hbc239f6b),
	.w4(32'h3ab003bc),
	.w5(32'hbbde13de),
	.w6(32'hbcc77770),
	.w7(32'hbbb805b5),
	.w8(32'hbbafd421),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14d8cf),
	.w1(32'hbb6ca6fb),
	.w2(32'h3a800ea9),
	.w3(32'hbc454a14),
	.w4(32'hbac6c95c),
	.w5(32'h3a9eb5a6),
	.w6(32'hbba9bd05),
	.w7(32'hbacad5b7),
	.w8(32'h3c37b040),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a820d97),
	.w1(32'hbb5eaf25),
	.w2(32'hbc529baa),
	.w3(32'h3b93ba3d),
	.w4(32'hbbe6401c),
	.w5(32'hbc419d38),
	.w6(32'h3c9dbbdb),
	.w7(32'hbac081b0),
	.w8(32'hbc171661),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22f711),
	.w1(32'h3c6681ca),
	.w2(32'h3c7752ce),
	.w3(32'hbb3a8e57),
	.w4(32'h3b457bad),
	.w5(32'hbae35913),
	.w6(32'h3b70f10e),
	.w7(32'h3c82e8f9),
	.w8(32'hbafebac2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaff72),
	.w1(32'hbb665025),
	.w2(32'h3a0e6a04),
	.w3(32'h3b7fa2e7),
	.w4(32'h3af5f387),
	.w5(32'h3b03db5f),
	.w6(32'hba88c812),
	.w7(32'h3bef4804),
	.w8(32'hbb8aa858),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d6b48),
	.w1(32'h393f2d7a),
	.w2(32'h3c11c95c),
	.w3(32'hbb92c347),
	.w4(32'h3b09c1b5),
	.w5(32'h3b3c4c55),
	.w6(32'hbc1e1bea),
	.w7(32'hbb5ddf7f),
	.w8(32'hb9a5728d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63e50a),
	.w1(32'h3c503e8e),
	.w2(32'h3c050549),
	.w3(32'h3b5647a0),
	.w4(32'hba024d49),
	.w5(32'hbbaf6fb1),
	.w6(32'hbbc786c5),
	.w7(32'h3b66173e),
	.w8(32'hbb5d6cc1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f5c12),
	.w1(32'hbc683f52),
	.w2(32'hbc4b4824),
	.w3(32'hbc485529),
	.w4(32'hbaffd2f7),
	.w5(32'hbbd0d3ca),
	.w6(32'hbc9396c2),
	.w7(32'hbc498fb3),
	.w8(32'hbc64bb38),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3016d1),
	.w1(32'hbc1921f9),
	.w2(32'h3b13bd33),
	.w3(32'hbc953157),
	.w4(32'hbb929e75),
	.w5(32'h3a776d91),
	.w6(32'hbd15eeee),
	.w7(32'hbc15a592),
	.w8(32'hba7437a1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92e14e),
	.w1(32'hbab92e66),
	.w2(32'hbb3f11b9),
	.w3(32'h39acb3e8),
	.w4(32'h3b5ba247),
	.w5(32'hbadad28d),
	.w6(32'h3b69392e),
	.w7(32'h3a9d3fc8),
	.w8(32'hbb83874f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9828570),
	.w1(32'hbc233b85),
	.w2(32'h3b96ea35),
	.w3(32'hbbc54774),
	.w4(32'h3bb8525b),
	.w5(32'hbbd277a8),
	.w6(32'hbc6f002d),
	.w7(32'h3b260f65),
	.w8(32'hbbcf25d9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cf1eb),
	.w1(32'hbc78672c),
	.w2(32'hbc76204b),
	.w3(32'hbc0a91dc),
	.w4(32'hbc59e51a),
	.w5(32'hbb3f2736),
	.w6(32'h3a946f59),
	.w7(32'hbc85a2bf),
	.w8(32'hbc4b5a0a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e9040),
	.w1(32'hbc2097b3),
	.w2(32'hbbc88a54),
	.w3(32'hba48a3eb),
	.w4(32'hbb44a033),
	.w5(32'hbae8062b),
	.w6(32'hbbef38cb),
	.w7(32'hbbf6e2d7),
	.w8(32'hbbe1bca0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4fe90),
	.w1(32'hbc124f57),
	.w2(32'hbb91f935),
	.w3(32'hbc008c3b),
	.w4(32'hbb8cf131),
	.w5(32'h3c126f58),
	.w6(32'hbbc0ddd4),
	.w7(32'hbc05699a),
	.w8(32'h3bbdd771),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace5bdd),
	.w1(32'h3aa42578),
	.w2(32'hbb9143cb),
	.w3(32'h3c9c84b9),
	.w4(32'hbb3e043f),
	.w5(32'hbad147f3),
	.w6(32'h3badb18a),
	.w7(32'hbc3a4e05),
	.w8(32'h3b9f8d04),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bb9bb),
	.w1(32'h3c06c962),
	.w2(32'hb98a6a6f),
	.w3(32'h3be85d0a),
	.w4(32'h3c41e7fc),
	.w5(32'hbbf97670),
	.w6(32'hbc6226dd),
	.w7(32'h3c20e537),
	.w8(32'hbc01a68b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1792dd),
	.w1(32'h3b98e244),
	.w2(32'h3bb4766e),
	.w3(32'hbbdb0e28),
	.w4(32'hbb8502b7),
	.w5(32'h3c17a705),
	.w6(32'hbbcd8d7a),
	.w7(32'h3ba9e633),
	.w8(32'hba151183),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb877aac),
	.w1(32'hbc48a17d),
	.w2(32'h3c4b10f8),
	.w3(32'hbc106946),
	.w4(32'h3c3a61f7),
	.w5(32'hbb388d71),
	.w6(32'hbc6958f0),
	.w7(32'h3b6c4204),
	.w8(32'h3b813da5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea166e),
	.w1(32'h3b898ce7),
	.w2(32'h3b30538c),
	.w3(32'hb988280a),
	.w4(32'h3b0979b6),
	.w5(32'h3bb40cfa),
	.w6(32'h39f9b8c8),
	.w7(32'h3ab5e206),
	.w8(32'h3b47a6ca),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b495d5b),
	.w1(32'hba8cfce1),
	.w2(32'h3a9dfe43),
	.w3(32'h3b294c2e),
	.w4(32'h399275f8),
	.w5(32'h3b235e82),
	.w6(32'h39fa24d6),
	.w7(32'h3ab9b91b),
	.w8(32'hb8cfa3e0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb052c5a),
	.w1(32'hbbd35393),
	.w2(32'hbba5c11c),
	.w3(32'h3b0d7f4f),
	.w4(32'h3b3a372d),
	.w5(32'hbad269f8),
	.w6(32'hb97ce183),
	.w7(32'h3b4224f7),
	.w8(32'hbb90657f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ecd04),
	.w1(32'h3a991e01),
	.w2(32'h3b88e10b),
	.w3(32'hbbabd26d),
	.w4(32'h3afdfac1),
	.w5(32'h3a6dac79),
	.w6(32'hbbbd2af2),
	.w7(32'h3ba3236b),
	.w8(32'hbb8aa0cb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e705),
	.w1(32'hbbeeeb99),
	.w2(32'hb9a52100),
	.w3(32'hbb985cf4),
	.w4(32'hba8ead9b),
	.w5(32'h3b866caf),
	.w6(32'hbb8bc525),
	.w7(32'hbbcd3578),
	.w8(32'hbbea0f59),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4266d),
	.w1(32'h3a790947),
	.w2(32'h3ba111b0),
	.w3(32'hba752baf),
	.w4(32'hbb64602a),
	.w5(32'hbb005d04),
	.w6(32'hbc57c9cb),
	.w7(32'hbb9de357),
	.w8(32'h3716a3b3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2a9f4),
	.w1(32'hbc096531),
	.w2(32'hbbcb3271),
	.w3(32'hbb51cad1),
	.w4(32'hbb763ae1),
	.w5(32'h3931e7a2),
	.w6(32'hb94929a1),
	.w7(32'hbb662150),
	.w8(32'hbb6e155e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82cf33),
	.w1(32'hbb8ce36a),
	.w2(32'hba94660f),
	.w3(32'hbbd8ddbe),
	.w4(32'hbb25c36b),
	.w5(32'h3b6e3ac4),
	.w6(32'hbbb6869f),
	.w7(32'hbc1a8841),
	.w8(32'hbbd2abde),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd5db7),
	.w1(32'hb9e9e4c7),
	.w2(32'hbb39e87a),
	.w3(32'h3c6c1d5f),
	.w4(32'h3b78cb32),
	.w5(32'h3b4f0ffe),
	.w6(32'h3a444c98),
	.w7(32'h395df710),
	.w8(32'h39b1eff0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e53ae),
	.w1(32'hb963e9f2),
	.w2(32'hba98dc1e),
	.w3(32'h3bd74be9),
	.w4(32'h3b702594),
	.w5(32'hbb054d0b),
	.w6(32'h3b9f2ed1),
	.w7(32'h3bda02a5),
	.w8(32'hbb1a721d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01b9fc),
	.w1(32'h3b832460),
	.w2(32'h389eb9f1),
	.w3(32'h3b58851f),
	.w4(32'h3ad3a49d),
	.w5(32'hbb9b622e),
	.w6(32'hbb823780),
	.w7(32'h3b4644d1),
	.w8(32'hbb14400a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77f2e0),
	.w1(32'h3bbb5c15),
	.w2(32'hbaa2e626),
	.w3(32'hbab7704d),
	.w4(32'hbb841cb0),
	.w5(32'hbc0e12ec),
	.w6(32'hbaa2bc3e),
	.w7(32'h3af922de),
	.w8(32'hbc12aa0d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03caaf),
	.w1(32'hbbe31fbf),
	.w2(32'hbbb5ffdb),
	.w3(32'hbc7ec42d),
	.w4(32'hbbd3496d),
	.w5(32'hbad2b9e5),
	.w6(32'hbbb4b90a),
	.w7(32'hbbb32af5),
	.w8(32'hbb42aa9c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a380e),
	.w1(32'hbc90315d),
	.w2(32'hbc5985cc),
	.w3(32'hbc214d7c),
	.w4(32'hbc53c2b0),
	.w5(32'h3c06080d),
	.w6(32'hbbe005c2),
	.w7(32'hbcb0313b),
	.w8(32'h3bb8ccde),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b508233),
	.w1(32'hbb6d670e),
	.w2(32'hbbf1ae82),
	.w3(32'hb97029c1),
	.w4(32'hbba413a4),
	.w5(32'h3c258b71),
	.w6(32'hbc1712eb),
	.w7(32'hbc0f8e19),
	.w8(32'h3b6c7f7a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5fe28f),
	.w1(32'h3c26f2fc),
	.w2(32'h3c3dee8e),
	.w3(32'h3bae3afc),
	.w4(32'h3bb4e31d),
	.w5(32'h3aae0b07),
	.w6(32'hbc4a4bbd),
	.w7(32'hbaa72e34),
	.w8(32'hbbb2b0f3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39903530),
	.w1(32'h3ae3d0e8),
	.w2(32'h3b6266fe),
	.w3(32'hbb6a1588),
	.w4(32'h3b25eb02),
	.w5(32'hba94f130),
	.w6(32'hbc777136),
	.w7(32'hbb29ede1),
	.w8(32'h3b2e35fe),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85c006),
	.w1(32'hbb666c73),
	.w2(32'hbb5f462d),
	.w3(32'h3c2b0365),
	.w4(32'h3aa66301),
	.w5(32'hbb0de2cf),
	.w6(32'h3c1f20f5),
	.w7(32'h37e03cda),
	.w8(32'h3bce5f8c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14c905),
	.w1(32'h38f35e77),
	.w2(32'hb9357fc0),
	.w3(32'h3a840387),
	.w4(32'hbaed3915),
	.w5(32'h3b32907d),
	.w6(32'h3bd65e15),
	.w7(32'hbb7daf89),
	.w8(32'h3bd5b2c4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dfff9),
	.w1(32'h3bbe5fef),
	.w2(32'h3ad38cd6),
	.w3(32'h3b4b396a),
	.w4(32'h3b7b7a18),
	.w5(32'hbc18bbf2),
	.w6(32'hbc5bf615),
	.w7(32'hbc067919),
	.w8(32'hbc08ad82),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1e79a),
	.w1(32'hbb98d7d1),
	.w2(32'hbb2ae17e),
	.w3(32'hbc401b9a),
	.w4(32'hbba0c5e6),
	.w5(32'h3bc24bbf),
	.w6(32'hbab245c8),
	.w7(32'hbb5681da),
	.w8(32'h3bb1dd81),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a80c4e),
	.w1(32'hba008770),
	.w2(32'hbba99c58),
	.w3(32'h3c59f74c),
	.w4(32'h3a194e9e),
	.w5(32'hba9a5632),
	.w6(32'hb741c01c),
	.w7(32'h3baacc61),
	.w8(32'hbb56f601),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e344f),
	.w1(32'h3a9a273d),
	.w2(32'hbb8543e3),
	.w3(32'hbab3fa9c),
	.w4(32'hbb8e5ec6),
	.w5(32'hbbce6648),
	.w6(32'hbb2c2060),
	.w7(32'h3ac700d8),
	.w8(32'hbc15c0d5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0502e6),
	.w1(32'h3be621f3),
	.w2(32'h3be3078d),
	.w3(32'h3b93acd8),
	.w4(32'h3c09f999),
	.w5(32'hb93ab99d),
	.w6(32'hbbda4493),
	.w7(32'h3c633a3a),
	.w8(32'h3b811024),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c300ce8),
	.w1(32'h3c729c7d),
	.w2(32'h3c696c2c),
	.w3(32'h3ba6dcac),
	.w4(32'h3bf1d284),
	.w5(32'hbc0e142a),
	.w6(32'h3b9d3379),
	.w7(32'h3c80b791),
	.w8(32'hbc1c5419),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52887d),
	.w1(32'hbc86b231),
	.w2(32'hbc3487a9),
	.w3(32'hbc4b1613),
	.w4(32'hbbe3e0cc),
	.w5(32'h3b491d22),
	.w6(32'hbc00ff9d),
	.w7(32'hbc670a79),
	.w8(32'hbb9af4ae),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e3921),
	.w1(32'hba91d74c),
	.w2(32'hbbfbde92),
	.w3(32'hbbedf204),
	.w4(32'hbc009165),
	.w5(32'h3c319661),
	.w6(32'hbc64ee2c),
	.w7(32'hbc3557f8),
	.w8(32'h3bf2005b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80055f),
	.w1(32'h3c9c67f3),
	.w2(32'h3cb2877f),
	.w3(32'h3b640ff1),
	.w4(32'h3bcaab50),
	.w5(32'h3bb4b0bc),
	.w6(32'hbc1794ca),
	.w7(32'h3c365b8b),
	.w8(32'h3b0e3330),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c079d9a),
	.w1(32'h3b7bac06),
	.w2(32'h3bb4f18b),
	.w3(32'h3b856803),
	.w4(32'hba64c698),
	.w5(32'hba2a7dd8),
	.w6(32'hbb0137c7),
	.w7(32'h3bbbf190),
	.w8(32'hbb8b7baa),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a290843),
	.w1(32'h3c2e436f),
	.w2(32'h3c5b967c),
	.w3(32'h3bf3f7bd),
	.w4(32'h3bdb779e),
	.w5(32'hbbeca3a1),
	.w6(32'h3c86e067),
	.w7(32'h3c54acbc),
	.w8(32'hbb61fd4a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b295805),
	.w1(32'h3b9ec4fb),
	.w2(32'h3c0a361d),
	.w3(32'hbb91c79c),
	.w4(32'hbaf1e1f5),
	.w5(32'h3ba26070),
	.w6(32'h3963bb47),
	.w7(32'h3b497407),
	.w8(32'h3b4fc1e4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9095dc6),
	.w1(32'hbba60ae8),
	.w2(32'hbc35dced),
	.w3(32'hbbb21d4b),
	.w4(32'hbc14b4c7),
	.w5(32'h3ad2353a),
	.w6(32'h3ab3c73e),
	.w7(32'hbbdb561d),
	.w8(32'hba72dabc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae46682),
	.w1(32'hbc20ac9e),
	.w2(32'h3c45f359),
	.w3(32'hbb786c68),
	.w4(32'h3c394094),
	.w5(32'h3bd393ae),
	.w6(32'hbc243294),
	.w7(32'h3bb7b157),
	.w8(32'h3a4bb2ee),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2e62e),
	.w1(32'h3b2e3c5c),
	.w2(32'hbbcc0bc1),
	.w3(32'h3b700f93),
	.w4(32'hbb534cdb),
	.w5(32'hbb1ae145),
	.w6(32'h3a81b425),
	.w7(32'hbb8abc72),
	.w8(32'hbb60655b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae80a9),
	.w1(32'hbc252a35),
	.w2(32'hbb9aa79f),
	.w3(32'hbc094045),
	.w4(32'hbb60d7a5),
	.w5(32'hbbd785c0),
	.w6(32'hbc0b0131),
	.w7(32'hbbfec246),
	.w8(32'hbbef9280),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee0cfc),
	.w1(32'hbbc0d3b9),
	.w2(32'hbba7d5be),
	.w3(32'h3af04993),
	.w4(32'hba83aa4e),
	.w5(32'hbc02ad32),
	.w6(32'h3b91df92),
	.w7(32'hb8f63106),
	.w8(32'hbc42fc69),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc8e9c),
	.w1(32'hbb0818d3),
	.w2(32'hba8518a2),
	.w3(32'hbb6080fe),
	.w4(32'hba7ff3ef),
	.w5(32'h3b213a74),
	.w6(32'h3ab353e5),
	.w7(32'h3b9518ec),
	.w8(32'h3b0e3809),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ec3df),
	.w1(32'h3b181b97),
	.w2(32'h3a39d882),
	.w3(32'hbb37d350),
	.w4(32'h3aaf9155),
	.w5(32'hba5989e8),
	.w6(32'hbb78c996),
	.w7(32'h3ae08768),
	.w8(32'h3bca4fe8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2af564),
	.w1(32'hbbf9eb72),
	.w2(32'hb9c086e9),
	.w3(32'hbc12c5ac),
	.w4(32'h3b25f24b),
	.w5(32'hbb4d64ff),
	.w6(32'hbc21bb7f),
	.w7(32'hbb5d4afb),
	.w8(32'h3ae620c6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b589256),
	.w1(32'hbbfa7be0),
	.w2(32'hbb574a22),
	.w3(32'hbc33a5b8),
	.w4(32'hbbe0e0e3),
	.w5(32'hbc2acdc2),
	.w6(32'hbbfe7b50),
	.w7(32'hbb5be0df),
	.w8(32'hbc3312eb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc028060),
	.w1(32'hbbe53e8c),
	.w2(32'hbbca48fe),
	.w3(32'hbbe367ac),
	.w4(32'hbb8447f6),
	.w5(32'hbc017de0),
	.w6(32'hb7cade88),
	.w7(32'hbab1fde9),
	.w8(32'hbb8a590d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd47623),
	.w1(32'h3bc43fbc),
	.w2(32'h3bc9c2e3),
	.w3(32'h3adeab98),
	.w4(32'hba280e06),
	.w5(32'hbb88a523),
	.w6(32'hbb914500),
	.w7(32'h3b50a299),
	.w8(32'h3b42a702),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc67879),
	.w1(32'h3c94b5d6),
	.w2(32'h3c4b77b5),
	.w3(32'h3bfce10b),
	.w4(32'h3b74ffc4),
	.w5(32'h3c7a8af4),
	.w6(32'h3bbb81de),
	.w7(32'h3c86fecd),
	.w8(32'h3c5dd9c3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9941789),
	.w1(32'hbc33db72),
	.w2(32'hbc07eb27),
	.w3(32'hba58e611),
	.w4(32'hbbb30636),
	.w5(32'h3acba2a4),
	.w6(32'hbca7c23c),
	.w7(32'hbc293010),
	.w8(32'hba327219),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fed8f1),
	.w1(32'hba3d1ab0),
	.w2(32'h3a55021d),
	.w3(32'h3a5ceab4),
	.w4(32'h3b28c6f6),
	.w5(32'hbac94ede),
	.w6(32'h37dd6e11),
	.w7(32'h3b65544b),
	.w8(32'hbbacd0b6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab8313),
	.w1(32'hbbea989a),
	.w2(32'h3ad21954),
	.w3(32'hbbf978e3),
	.w4(32'hb963b4fc),
	.w5(32'hbb691e19),
	.w6(32'hbbe2bcb5),
	.w7(32'h3a1ab8ed),
	.w8(32'hbc0685eb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d81d0),
	.w1(32'h3abdb073),
	.w2(32'hba69c9f2),
	.w3(32'hba4d1792),
	.w4(32'h3b47de15),
	.w5(32'hbb226043),
	.w6(32'hbb35e3e8),
	.w7(32'h3b65fc34),
	.w8(32'h3b1b2afa),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac40b10),
	.w1(32'hbb5fb285),
	.w2(32'hba81be60),
	.w3(32'h39a99a8e),
	.w4(32'hbb9b5ded),
	.w5(32'hba50a6ff),
	.w6(32'h3b07d08a),
	.w7(32'hbba49d4f),
	.w8(32'h3ae36ae5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52ea70),
	.w1(32'hbba1b0cc),
	.w2(32'hbad199c5),
	.w3(32'hbb73df39),
	.w4(32'h3ac084c2),
	.w5(32'h3b34d8fc),
	.w6(32'hbb921532),
	.w7(32'h3b707014),
	.w8(32'hbb3bd799),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadf92b),
	.w1(32'h3b7e8e93),
	.w2(32'h3b6b2594),
	.w3(32'h3b0952dc),
	.w4(32'h3bbe76b3),
	.w5(32'hba83b62a),
	.w6(32'h3b4bfa19),
	.w7(32'h3a84914a),
	.w8(32'hba85d717),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4bd88),
	.w1(32'hbc0027e9),
	.w2(32'hbbeb6e5b),
	.w3(32'hbc150dc4),
	.w4(32'hbbcf5696),
	.w5(32'hb9c98a2d),
	.w6(32'hbbd5f546),
	.w7(32'hbbcf3177),
	.w8(32'hbb645517),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaaacda),
	.w1(32'h3b4db25a),
	.w2(32'hbaf06899),
	.w3(32'h3b8adfa8),
	.w4(32'hb98afdd2),
	.w5(32'h3c045a1e),
	.w6(32'hba1448ab),
	.w7(32'hbb286db6),
	.w8(32'h39d25cef),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803595),
	.w1(32'hbb3e3492),
	.w2(32'h3b0de054),
	.w3(32'h3bbbfdea),
	.w4(32'h3b5c98ca),
	.w5(32'hbae193bb),
	.w6(32'h3ad2aa6d),
	.w7(32'h3b5ec15c),
	.w8(32'hbb774001),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7064b2),
	.w1(32'hb9eedf9b),
	.w2(32'h3bae8bc7),
	.w3(32'h3b3e863f),
	.w4(32'h3c3c375a),
	.w5(32'h3ba910ec),
	.w6(32'h3a4ad523),
	.w7(32'h3c130be4),
	.w8(32'h3b5990d7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3283d9),
	.w1(32'h3a85bd8f),
	.w2(32'h395b9354),
	.w3(32'h3bb60674),
	.w4(32'h3bb64bf9),
	.w5(32'hb909374d),
	.w6(32'h3ac5a5cc),
	.w7(32'h3be310f2),
	.w8(32'h3b567989),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9287820),
	.w1(32'hbb1f9ca8),
	.w2(32'hbb15e377),
	.w3(32'h3b3a83f2),
	.w4(32'hbb1974d1),
	.w5(32'h3afc53fe),
	.w6(32'h3baa83bb),
	.w7(32'h3ba77fa0),
	.w8(32'h3b58b5bc),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381d8228),
	.w1(32'h3a323580),
	.w2(32'h3bafb08c),
	.w3(32'hb967af52),
	.w4(32'hbabb5627),
	.w5(32'hbb601aee),
	.w6(32'h3b6d30cb),
	.w7(32'h3aa27191),
	.w8(32'hbae588dd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72a390),
	.w1(32'hbb870a6e),
	.w2(32'hbb309f5e),
	.w3(32'hbaa3eb1b),
	.w4(32'hbab1d71e),
	.w5(32'hba09b6e1),
	.w6(32'h3aba55c5),
	.w7(32'hbaf23242),
	.w8(32'h3b6969a5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf9cfd),
	.w1(32'hbb1f3e54),
	.w2(32'hbb3877ce),
	.w3(32'hbb63abeb),
	.w4(32'hbbc1f44e),
	.w5(32'h3a2b19fe),
	.w6(32'hbb022c7e),
	.w7(32'hbb3eb9ae),
	.w8(32'h3b30ebbb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18db4d),
	.w1(32'h3b053843),
	.w2(32'h3ae74f50),
	.w3(32'hbaa862ff),
	.w4(32'hbb050d18),
	.w5(32'hbb6e1b2b),
	.w6(32'hba32ef05),
	.w7(32'h3af8ab22),
	.w8(32'hbb9fd032),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc2053),
	.w1(32'hbbb3a69f),
	.w2(32'hbb1bfafa),
	.w3(32'hbc20eecb),
	.w4(32'h3c233bf2),
	.w5(32'hbac0c2ba),
	.w6(32'hbc400046),
	.w7(32'h3b9ad871),
	.w8(32'hbaed262f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84f049),
	.w1(32'hbb55ed02),
	.w2(32'hbaae5e88),
	.w3(32'hb6f737de),
	.w4(32'hbb1a032e),
	.w5(32'h3a5fdda8),
	.w6(32'h3b37d151),
	.w7(32'hbb1786c4),
	.w8(32'h3ba3347f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2f9f5),
	.w1(32'h3bd87fe4),
	.w2(32'h3afefb33),
	.w3(32'h3ad0ac12),
	.w4(32'hbba81cb1),
	.w5(32'hbb5b0e57),
	.w6(32'h3b213cf1),
	.w7(32'hbb029e41),
	.w8(32'hbb828eb4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47b06e),
	.w1(32'hbbbd0655),
	.w2(32'hbb9f4e95),
	.w3(32'hbbafe96e),
	.w4(32'hb9253a6f),
	.w5(32'h3b023243),
	.w6(32'hbb3b99ae),
	.w7(32'hbc0205c6),
	.w8(32'h3b25249f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990e169),
	.w1(32'hbb3487a9),
	.w2(32'hbb896924),
	.w3(32'hbabd720c),
	.w4(32'hbb42c528),
	.w5(32'hbae2f303),
	.w6(32'hb7b961c7),
	.w7(32'h392283a7),
	.w8(32'hbb960f59),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85d2ff),
	.w1(32'hbb883579),
	.w2(32'hbbd4aa44),
	.w3(32'hbb8e494c),
	.w4(32'hbbd46e6b),
	.w5(32'h3a2d4c2c),
	.w6(32'hbbbeb21d),
	.w7(32'hbba11c13),
	.w8(32'h3aa281e6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a7284),
	.w1(32'h3896dbb2),
	.w2(32'hbb26b081),
	.w3(32'hbaa33a67),
	.w4(32'hbad47dc3),
	.w5(32'hbadbf910),
	.w6(32'hba297feb),
	.w7(32'hb9fb99f5),
	.w8(32'hbaa6173c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7df838),
	.w1(32'hbb6d2e85),
	.w2(32'h3a465cc1),
	.w3(32'hbb92761c),
	.w4(32'hb9384734),
	.w5(32'h3ac6b3f1),
	.w6(32'hbb8537ad),
	.w7(32'hbb3561a8),
	.w8(32'h38fe52a7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2da11d),
	.w1(32'hbae95436),
	.w2(32'h3aa5167b),
	.w3(32'h3c07df1b),
	.w4(32'hb914f722),
	.w5(32'hbae6b984),
	.w6(32'h3c0667fb),
	.w7(32'h394fcaa3),
	.w8(32'h3ab22bdf),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39212bab),
	.w1(32'h3bab3bab),
	.w2(32'h3bb79a15),
	.w3(32'h3b797c6c),
	.w4(32'h3ac8df94),
	.w5(32'hba76c50d),
	.w6(32'h3a637fee),
	.w7(32'h3b536a1e),
	.w8(32'h3a9b9987),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb9658),
	.w1(32'h3a325d2f),
	.w2(32'h3a84200b),
	.w3(32'hbb018236),
	.w4(32'hbb5df208),
	.w5(32'h3ab0f912),
	.w6(32'h3bb3e508),
	.w7(32'hbaf66f34),
	.w8(32'h3a977833),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29a3ef),
	.w1(32'hb9258ead),
	.w2(32'h3a8b53a2),
	.w3(32'hb8f072b8),
	.w4(32'hba35d3f5),
	.w5(32'hbb2a3c30),
	.w6(32'h3b088d62),
	.w7(32'hbb154733),
	.w8(32'hbad32f47),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacba81d),
	.w1(32'h3b04200a),
	.w2(32'h3bdb4bcb),
	.w3(32'h3b05dc15),
	.w4(32'h3bcf078f),
	.w5(32'hba0677cc),
	.w6(32'h3bd8008c),
	.w7(32'h3c3acd90),
	.w8(32'h3ac5a2bc),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a483243),
	.w1(32'hbae9d5e4),
	.w2(32'h3a80ed73),
	.w3(32'hba223a9b),
	.w4(32'h3a2da49d),
	.w5(32'hbc31bdf9),
	.w6(32'hbbd6fe08),
	.w7(32'hb9f0a5c2),
	.w8(32'hbc393d71),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34e5c0),
	.w1(32'hbc7f3c65),
	.w2(32'hbc84772d),
	.w3(32'hbc10c8a2),
	.w4(32'hbc3f9e97),
	.w5(32'hbb85ebe9),
	.w6(32'hbc6c28ac),
	.w7(32'hbc47cbf5),
	.w8(32'hbb103a94),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb546b58),
	.w1(32'hbb85e181),
	.w2(32'hbbaab1e2),
	.w3(32'hbba724b2),
	.w4(32'h3acc32f8),
	.w5(32'h3b27cd0c),
	.w6(32'hbb7c1aca),
	.w7(32'h3953035d),
	.w8(32'hbbbd0b3b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb405d56),
	.w1(32'hba1ce1cb),
	.w2(32'hbb827f55),
	.w3(32'h3b4396c9),
	.w4(32'h3a5c7fa9),
	.w5(32'h3c0ddba7),
	.w6(32'hba8461d6),
	.w7(32'hbbd86b6c),
	.w8(32'h3bdd65a6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fd111),
	.w1(32'h3c168492),
	.w2(32'h3bff55f0),
	.w3(32'h3c0d62e8),
	.w4(32'h3c108daf),
	.w5(32'h3a7daa7b),
	.w6(32'h3c04f4a0),
	.w7(32'h3bef322d),
	.w8(32'h3c24bc31),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4663c),
	.w1(32'hbad3706a),
	.w2(32'hbbffbbf2),
	.w3(32'hbb24be08),
	.w4(32'hbbe9eb6f),
	.w5(32'h3b373518),
	.w6(32'h3c3759b1),
	.w7(32'h3b9fc9a7),
	.w8(32'h3b9d9752),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb037e),
	.w1(32'h3b76d127),
	.w2(32'h3bd5f6ba),
	.w3(32'h3b7a25ad),
	.w4(32'h3b9ffd44),
	.w5(32'hbadcc88f),
	.w6(32'h3c1bc78d),
	.w7(32'h3c0b583a),
	.w8(32'h3a866f67),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81eec5),
	.w1(32'h3b333851),
	.w2(32'hbada00a4),
	.w3(32'hbb83f309),
	.w4(32'hbb3f80e8),
	.w5(32'hbb549c37),
	.w6(32'hbb48d623),
	.w7(32'hba5547a6),
	.w8(32'hba8ecbd4),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba341590),
	.w1(32'hbb647b30),
	.w2(32'hbb8c95bf),
	.w3(32'hbb4c715d),
	.w4(32'hbba347f7),
	.w5(32'h39890885),
	.w6(32'h39961ef2),
	.w7(32'hbb31d8c7),
	.w8(32'h3bbf1dd5),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99800c0),
	.w1(32'hb969e890),
	.w2(32'hbb1c9910),
	.w3(32'hbaa97e11),
	.w4(32'hbb883b10),
	.w5(32'h3b228357),
	.w6(32'h3a46bb24),
	.w7(32'hbaf63821),
	.w8(32'h3b83bdc3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51ee27),
	.w1(32'h3b54261a),
	.w2(32'h3baa1f94),
	.w3(32'h3b84a76a),
	.w4(32'h3b91b1b2),
	.w5(32'h3a9e84e0),
	.w6(32'h3bd9808d),
	.w7(32'h3bf7318b),
	.w8(32'h3a8ede27),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be58af4),
	.w1(32'h3b637870),
	.w2(32'h3bb8bb1b),
	.w3(32'h3ad33387),
	.w4(32'h3bb0091b),
	.w5(32'h3abdb42e),
	.w6(32'h3bd5bfbb),
	.w7(32'h3b9aa648),
	.w8(32'h3a78b07c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6caf86),
	.w1(32'hbace9a4c),
	.w2(32'hbafec90e),
	.w3(32'h3ad16a2a),
	.w4(32'h3b086f88),
	.w5(32'hbb7826de),
	.w6(32'hbb584169),
	.w7(32'h3b1b3ea0),
	.w8(32'hbb65f8d8),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28f2de),
	.w1(32'hbb57d2d1),
	.w2(32'hbb02a852),
	.w3(32'hba673372),
	.w4(32'hbab74e5e),
	.w5(32'hbad0d161),
	.w6(32'h3b2dc8c3),
	.w7(32'h3a86048a),
	.w8(32'hbb374a61),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb977544),
	.w1(32'hbbc510e3),
	.w2(32'hbb32a396),
	.w3(32'hba8a0710),
	.w4(32'h39062a74),
	.w5(32'h3b4ff5d6),
	.w6(32'h3b517dad),
	.w7(32'h3ad2926e),
	.w8(32'h3bf38bbb),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d19d3),
	.w1(32'h3bb91f28),
	.w2(32'h3c25dca6),
	.w3(32'h3b5b5680),
	.w4(32'h3b16dfd6),
	.w5(32'h3af99b7a),
	.w6(32'h3bcf48a2),
	.w7(32'h3bc46308),
	.w8(32'h3a8ec737),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9877c),
	.w1(32'h39ee9460),
	.w2(32'hbb3d4df9),
	.w3(32'h3b87a7e4),
	.w4(32'hbab63db9),
	.w5(32'h3a2179cd),
	.w6(32'h3b0c0445),
	.w7(32'hb9596976),
	.w8(32'h3aea54cc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc925a),
	.w1(32'h3b40fd4e),
	.w2(32'h3baefaa5),
	.w3(32'h3baff8cb),
	.w4(32'h3c400f9a),
	.w5(32'h3b642785),
	.w6(32'h3bd38836),
	.w7(32'h3c6b9959),
	.w8(32'h3ab6a0d2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b302946),
	.w1(32'h3ae30c60),
	.w2(32'h3b231328),
	.w3(32'h3ab78a4e),
	.w4(32'h3b857c3a),
	.w5(32'h3acd79ab),
	.w6(32'h3aa579a0),
	.w7(32'h3ab2fed6),
	.w8(32'hbbbc2d13),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d714e),
	.w1(32'hba92fe59),
	.w2(32'h39784d15),
	.w3(32'h39d46daa),
	.w4(32'hbbabfd4f),
	.w5(32'hbb56bcee),
	.w6(32'hbb917d64),
	.w7(32'hbc1dbb5c),
	.w8(32'hbb562b17),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00e356),
	.w1(32'hbad676ce),
	.w2(32'hbb2bce91),
	.w3(32'hbb71a77e),
	.w4(32'hbb8dfeaa),
	.w5(32'h3b2e1e27),
	.w6(32'hbaaa16cc),
	.w7(32'hbbe5e366),
	.w8(32'h3ac2aa8e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4b04a),
	.w1(32'h3b27aa21),
	.w2(32'h3a99f77d),
	.w3(32'h3b7b42c8),
	.w4(32'h3b827096),
	.w5(32'h3a3a9e9b),
	.w6(32'h3adfe7f7),
	.w7(32'h3b292e74),
	.w8(32'h3aec045b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3082e5),
	.w1(32'h3b9038dd),
	.w2(32'h3acf3728),
	.w3(32'h3af666ea),
	.w4(32'hbb19a42e),
	.w5(32'hb9925402),
	.w6(32'h3b48d448),
	.w7(32'h3b15636d),
	.w8(32'hba711ed8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bfdf3),
	.w1(32'hbb01ec9a),
	.w2(32'hbb6bdd87),
	.w3(32'hbad7a278),
	.w4(32'hbb18eed5),
	.w5(32'h3a430ec3),
	.w6(32'hbaf6b8dd),
	.w7(32'h3ae2314e),
	.w8(32'h3a28d2e3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eab69),
	.w1(32'h3b35841e),
	.w2(32'hbb71f99f),
	.w3(32'h3ad5069b),
	.w4(32'hbb781956),
	.w5(32'h3aeb51bf),
	.w6(32'h3bd36495),
	.w7(32'hbb3daa51),
	.w8(32'hb8fd0636),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb495de6),
	.w1(32'hbb24b7cf),
	.w2(32'hbb1bc31f),
	.w3(32'h3b6195d6),
	.w4(32'hbaf3d323),
	.w5(32'h3b05e4f8),
	.w6(32'h3b53e9b1),
	.w7(32'hbb849a0e),
	.w8(32'h3ad6049d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad12587),
	.w1(32'h3b9016d4),
	.w2(32'h3c0b1d97),
	.w3(32'h3ba8c331),
	.w4(32'h3bc3fc07),
	.w5(32'hba34a9e0),
	.w6(32'h3a7fe2ce),
	.w7(32'h3bdf54c8),
	.w8(32'hbaa6e4e8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92ebe8),
	.w1(32'hbb8778d2),
	.w2(32'hba369a8b),
	.w3(32'hba82926f),
	.w4(32'h395ac181),
	.w5(32'hbb4cff5d),
	.w6(32'hbb7aa1d7),
	.w7(32'h38a3200e),
	.w8(32'h3a65398e),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91c2f4),
	.w1(32'hbbde4b4f),
	.w2(32'hbc08b495),
	.w3(32'hbb57fe0d),
	.w4(32'hbc112cdc),
	.w5(32'h3b2f3a79),
	.w6(32'hbaed1da5),
	.w7(32'hbb27bbe8),
	.w8(32'hb912a39b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae787f9),
	.w1(32'hbb078ac3),
	.w2(32'h3ae34f53),
	.w3(32'hbb2054a0),
	.w4(32'hbaaa1a4e),
	.w5(32'hbb2b9d21),
	.w6(32'hb9fa855e),
	.w7(32'hbb918192),
	.w8(32'hbbb86ae5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29884e),
	.w1(32'h3ab783a2),
	.w2(32'h3bccd995),
	.w3(32'h3b8d3029),
	.w4(32'h3bdde271),
	.w5(32'hbc105d1d),
	.w6(32'hb8523002),
	.w7(32'h3b6e5e80),
	.w8(32'h3aff2b6a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb753a72),
	.w1(32'hbbcaf7b4),
	.w2(32'hbb3803d7),
	.w3(32'hbc2d6ae9),
	.w4(32'hbc2a76e9),
	.w5(32'h3b1b4e79),
	.w6(32'hb9edb1a5),
	.w7(32'hbb4e64ce),
	.w8(32'h3b363625),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34d88c),
	.w1(32'h3afcfabc),
	.w2(32'hbb176c87),
	.w3(32'h38772d15),
	.w4(32'hbb937aa8),
	.w5(32'hbbce68b3),
	.w6(32'hba0e8e35),
	.w7(32'hbab46f20),
	.w8(32'hbb425f22),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8042df),
	.w1(32'hbbbd1bd6),
	.w2(32'hb9a5c70f),
	.w3(32'hbbc59e3d),
	.w4(32'hbc02d00d),
	.w5(32'h3a6e45c3),
	.w6(32'hbc069dc7),
	.w7(32'hbbaaaac8),
	.w8(32'h39db482a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d2f3a),
	.w1(32'h3b119fa4),
	.w2(32'h3b008fcf),
	.w3(32'hba2b0900),
	.w4(32'h3b845892),
	.w5(32'h3ad30c9b),
	.w6(32'h3ada0fa5),
	.w7(32'h3b6a1c79),
	.w8(32'h3b0a63ac),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac07d76),
	.w1(32'hb9fae452),
	.w2(32'h390b0bdc),
	.w3(32'hba8a190f),
	.w4(32'h3a97eb11),
	.w5(32'h3a88edc3),
	.w6(32'hbb15fa70),
	.w7(32'hba310a7f),
	.w8(32'hb9bd4132),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03ba74),
	.w1(32'h3c26ce98),
	.w2(32'h3b489817),
	.w3(32'h3b6ab306),
	.w4(32'h3a038cc8),
	.w5(32'hba294e47),
	.w6(32'h3b7e7380),
	.w7(32'h3aa4e676),
	.w8(32'h3b3c8f54),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8fa11),
	.w1(32'hba93649a),
	.w2(32'hbad5aacb),
	.w3(32'hbb23bfb0),
	.w4(32'hbb95ddf2),
	.w5(32'h3b6957f5),
	.w6(32'hba1c591f),
	.w7(32'hbbc129ef),
	.w8(32'h3aa7d998),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb4bf8),
	.w1(32'h3b948db0),
	.w2(32'hbac8a160),
	.w3(32'h3a8a0776),
	.w4(32'hbb1646d8),
	.w5(32'hbb12b8ee),
	.w6(32'h3a9c5f60),
	.w7(32'hba9cd7fe),
	.w8(32'h3add5652),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a917071),
	.w1(32'hb955e28a),
	.w2(32'hba900aed),
	.w3(32'hbbdb9005),
	.w4(32'hbb99f4b1),
	.w5(32'h3befcb97),
	.w6(32'h3bb8ccbd),
	.w7(32'h3b54acc1),
	.w8(32'h3b10d89b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafeb06),
	.w1(32'h3b7dde47),
	.w2(32'hba997e6e),
	.w3(32'h3bd07fd9),
	.w4(32'h3bb6f3a5),
	.w5(32'hb9b55b29),
	.w6(32'h3ba7fa56),
	.w7(32'hba09714a),
	.w8(32'h39e30516),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb882364),
	.w1(32'hbb8c4ab4),
	.w2(32'hbb2714f6),
	.w3(32'hbb65f7da),
	.w4(32'hbacaa710),
	.w5(32'hbace8cdb),
	.w6(32'hbc03ceb4),
	.w7(32'hba85188f),
	.w8(32'hbb9a06bc),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34a873),
	.w1(32'h3b92149a),
	.w2(32'h3bfdd8b1),
	.w3(32'h3b8b6449),
	.w4(32'h3bf126a4),
	.w5(32'h3b9231c1),
	.w6(32'h3acfac89),
	.w7(32'h3c0af295),
	.w8(32'h3b61fda9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ced76),
	.w1(32'h3b628de7),
	.w2(32'hbafed0f2),
	.w3(32'h3b7e8260),
	.w4(32'hbabb13f4),
	.w5(32'h3bb69697),
	.w6(32'h3b41b770),
	.w7(32'hbb9f732c),
	.w8(32'h3b0e5a20),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b5dc0),
	.w1(32'h3b32a036),
	.w2(32'h3bfc73d2),
	.w3(32'h3bc2c9c9),
	.w4(32'h3c63a4a9),
	.w5(32'h3aaee32c),
	.w6(32'h372ddb6c),
	.w7(32'h3c523240),
	.w8(32'hbb9f5ef1),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9b305),
	.w1(32'h3a2df2d1),
	.w2(32'h3b7a3628),
	.w3(32'h3b31db12),
	.w4(32'h3bb1f3bf),
	.w5(32'hbbfcad4c),
	.w6(32'hbb9ade62),
	.w7(32'h3a716380),
	.w8(32'hbc39473f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc176872),
	.w1(32'hbbb82fda),
	.w2(32'hbaf4a7f1),
	.w3(32'hbb67a6a1),
	.w4(32'h3b33cc3a),
	.w5(32'hbb766ec0),
	.w6(32'hbae31bd7),
	.w7(32'h3b115a63),
	.w8(32'hbbee1646),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc181d0a),
	.w1(32'hbbf6d69d),
	.w2(32'hbbba9804),
	.w3(32'hbb807113),
	.w4(32'hba4eb520),
	.w5(32'hbae7b98e),
	.w6(32'hbb24409a),
	.w7(32'hb9a91e01),
	.w8(32'h3b984b6b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76777a),
	.w1(32'h3b8c75cf),
	.w2(32'h3adca297),
	.w3(32'h39ab0aff),
	.w4(32'hbbaf5569),
	.w5(32'hbb346474),
	.w6(32'h3bad6748),
	.w7(32'h3ab23c7c),
	.w8(32'hbac90575),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89ffac),
	.w1(32'hbac418d5),
	.w2(32'hbad9decf),
	.w3(32'hbabd19df),
	.w4(32'hbb01363b),
	.w5(32'h3b4ab8bd),
	.w6(32'h3ad028d1),
	.w7(32'hba4896ad),
	.w8(32'h3b92caeb),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97b37f),
	.w1(32'h3b8af81a),
	.w2(32'h3a4e264e),
	.w3(32'h3b33062e),
	.w4(32'hbb890235),
	.w5(32'h3c1b6882),
	.w6(32'h3b07aadf),
	.w7(32'h3a0d4b19),
	.w8(32'h3c23fd64),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c001a08),
	.w1(32'hb9e177b4),
	.w2(32'hba9875a1),
	.w3(32'hbb7526af),
	.w4(32'hb9e10c88),
	.w5(32'hbb772cf3),
	.w6(32'h3bbb9e7c),
	.w7(32'h393c1811),
	.w8(32'hbbc40dd4),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25e715),
	.w1(32'hbb78a9ee),
	.w2(32'hbbc4117c),
	.w3(32'hbb3b2843),
	.w4(32'h3bac86a2),
	.w5(32'h3b798dca),
	.w6(32'hbbcbc5dc),
	.w7(32'hbba1fefd),
	.w8(32'hbac23893),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a0aa6),
	.w1(32'hbbb0bb43),
	.w2(32'hbb94e5ad),
	.w3(32'hbb115b54),
	.w4(32'h3a0319c3),
	.w5(32'hbb168937),
	.w6(32'hba6c00cc),
	.w7(32'hbb1302eb),
	.w8(32'hbb8f86e6),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb556f42),
	.w1(32'hbad7335b),
	.w2(32'h3aa44b17),
	.w3(32'hbb1a11d6),
	.w4(32'hbb6e7e48),
	.w5(32'hbb41b860),
	.w6(32'hbb08b0a8),
	.w7(32'hba06fab0),
	.w8(32'hbba67f1b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb511bc5),
	.w1(32'h3aa9007a),
	.w2(32'hbb6037a8),
	.w3(32'hbae2d398),
	.w4(32'h3aabc93d),
	.w5(32'h3b8f4840),
	.w6(32'hbb188a14),
	.w7(32'hbb21e5ad),
	.w8(32'hb88ce6b6),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6eda73),
	.w1(32'hbb0b64ee),
	.w2(32'h3b1deca7),
	.w3(32'hb984250a),
	.w4(32'h3b8e25b8),
	.w5(32'hbab44154),
	.w6(32'hbabe687a),
	.w7(32'h3b5f3227),
	.w8(32'hbaa6c619),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb368711),
	.w1(32'hbad13960),
	.w2(32'h39aa3823),
	.w3(32'h39f64d6a),
	.w4(32'hba83e370),
	.w5(32'hbab91fb6),
	.w6(32'hb5892950),
	.w7(32'h39d887f7),
	.w8(32'hbc1a7ce5),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d6123),
	.w1(32'hbb92730e),
	.w2(32'h3ab019a1),
	.w3(32'hbbbb7e8e),
	.w4(32'h3a1242c4),
	.w5(32'h3b66b099),
	.w6(32'hbb8a2506),
	.w7(32'hba10e176),
	.w8(32'h3bc56b29),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d9c88),
	.w1(32'h3b8ead7b),
	.w2(32'h37c9e331),
	.w3(32'h39b9c80b),
	.w4(32'hbbddece4),
	.w5(32'hbb8cfa92),
	.w6(32'hb98ddf3c),
	.w7(32'hba84af0c),
	.w8(32'hbad59850),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb770001),
	.w1(32'h39e0aaba),
	.w2(32'h3a82dff4),
	.w3(32'hbaf70351),
	.w4(32'hbb99ee60),
	.w5(32'hbb1e41f9),
	.w6(32'h3bfcc918),
	.w7(32'h3b131513),
	.w8(32'hbad19535),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e8736c),
	.w1(32'h3ae53218),
	.w2(32'h3aefb9a6),
	.w3(32'hbb20047e),
	.w4(32'hbab9ad25),
	.w5(32'hbb5bdc78),
	.w6(32'h3c3f5378),
	.w7(32'h3bd9f609),
	.w8(32'hbac8f87e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12050d),
	.w1(32'h3a88cc4f),
	.w2(32'h3b8cdb25),
	.w3(32'hb750b711),
	.w4(32'h3b94964b),
	.w5(32'hbb351a0e),
	.w6(32'h3a67ba7d),
	.w7(32'h3c002fad),
	.w8(32'h3bcee34c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a334279),
	.w1(32'hbb140d05),
	.w2(32'hbb4e1ebc),
	.w3(32'hbab7e279),
	.w4(32'h39f25976),
	.w5(32'h3a089182),
	.w6(32'h3bb3b5f6),
	.w7(32'h3b8b0147),
	.w8(32'h3a30d4bc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f759e3),
	.w1(32'hb91dde9c),
	.w2(32'hba9ac520),
	.w3(32'hbb058773),
	.w4(32'hb9d47f22),
	.w5(32'h3acd4d02),
	.w6(32'hba057b05),
	.w7(32'h3af716f4),
	.w8(32'h3a6af70a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7050b),
	.w1(32'h3adacbe6),
	.w2(32'h3b16d777),
	.w3(32'hbb39fee9),
	.w4(32'h3bafd9da),
	.w5(32'hba79378a),
	.w6(32'hbb185d51),
	.w7(32'h3b807f9a),
	.w8(32'h3b5f2072),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a752fd1),
	.w1(32'hbac96c9a),
	.w2(32'hbb499a0b),
	.w3(32'hbb894da5),
	.w4(32'hbb551347),
	.w5(32'hba8871c3),
	.w6(32'h392c875c),
	.w7(32'hb88e4f72),
	.w8(32'h3a65656f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f1ef5),
	.w1(32'hbb83fef6),
	.w2(32'hbb00469c),
	.w3(32'hbbaa85c8),
	.w4(32'hbb1de9c0),
	.w5(32'h3c070d92),
	.w6(32'h3715fa6d),
	.w7(32'hbaaa08b4),
	.w8(32'h3b5872a0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc611ca),
	.w1(32'h3bbd2402),
	.w2(32'h3ca900bf),
	.w3(32'h3c3e76b9),
	.w4(32'h3c8dadef),
	.w5(32'h3b021a0b),
	.w6(32'h3c051b25),
	.w7(32'h3c9d8160),
	.w8(32'h3b8ec7b2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82571d),
	.w1(32'hbbc579dc),
	.w2(32'hba51aed1),
	.w3(32'hbb6c9638),
	.w4(32'h3b1a7c58),
	.w5(32'h3be1b37b),
	.w6(32'hbbbf208c),
	.w7(32'h3a1b1740),
	.w8(32'h3b0a17c2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8343d0),
	.w1(32'h3bb5d5b5),
	.w2(32'h3bb90782),
	.w3(32'h3ba3bc46),
	.w4(32'h3c06c0d3),
	.w5(32'hbad3f5ec),
	.w6(32'hba1e7f93),
	.w7(32'h3b3f0195),
	.w8(32'hbb505860),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a914687),
	.w1(32'h3b5af8b5),
	.w2(32'hba455dc9),
	.w3(32'h3acd10f3),
	.w4(32'hbb3fa3a3),
	.w5(32'h3b16d27f),
	.w6(32'hbb1c6530),
	.w7(32'hbbc3072c),
	.w8(32'h3a9b0fbe),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b470f54),
	.w1(32'h3acf6d19),
	.w2(32'h384175be),
	.w3(32'h3a2e796e),
	.w4(32'h3ae89b67),
	.w5(32'hb9e54e9c),
	.w6(32'h3b49f2fd),
	.w7(32'h3bee3484),
	.w8(32'hb8cfd85b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdb5f5),
	.w1(32'h3ba0a3cf),
	.w2(32'hbab37303),
	.w3(32'h3a70995f),
	.w4(32'hb9c7ab77),
	.w5(32'hbb80d3c9),
	.w6(32'hba943c61),
	.w7(32'h3b67bf1b),
	.w8(32'hbad8adf5),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37a678),
	.w1(32'hba817fe3),
	.w2(32'hb8cc54a6),
	.w3(32'hbb9a5a84),
	.w4(32'hbab54550),
	.w5(32'h3b18040f),
	.w6(32'hb912bb3b),
	.w7(32'hbb3e0d37),
	.w8(32'h3b13c382),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81b55f),
	.w1(32'hbb442e07),
	.w2(32'hbadb3de4),
	.w3(32'hbadc7222),
	.w4(32'h3a5735d1),
	.w5(32'hba2bcd34),
	.w6(32'h386414ca),
	.w7(32'hb959987e),
	.w8(32'hba7a0d73),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace487a),
	.w1(32'hb9d7cf24),
	.w2(32'hba403a67),
	.w3(32'hb795ebbb),
	.w4(32'h38a59ce4),
	.w5(32'hba11cc67),
	.w6(32'h3b9d7f2c),
	.w7(32'hb9f02647),
	.w8(32'h3b42988f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f7cca5),
	.w1(32'hbb82b751),
	.w2(32'hbab7e1a7),
	.w3(32'hbb24494d),
	.w4(32'hba6d9b54),
	.w5(32'hbab32d52),
	.w6(32'h3aa819f2),
	.w7(32'h3b31dafc),
	.w8(32'hbb52e7bd),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3274e1),
	.w1(32'hbb49a5ab),
	.w2(32'hbb09addf),
	.w3(32'hb95d49b1),
	.w4(32'h3b84d4c1),
	.w5(32'h3ba1b002),
	.w6(32'hbb387d40),
	.w7(32'h398f5614),
	.w8(32'h3ba89168),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e4417),
	.w1(32'h3a26c7ab),
	.w2(32'h3b49c569),
	.w3(32'h3b4e2737),
	.w4(32'h3b8f2547),
	.w5(32'hbada3c47),
	.w6(32'h3be84f70),
	.w7(32'h3b836879),
	.w8(32'h3ba9bb8f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab387ba),
	.w1(32'hba60a2ff),
	.w2(32'h3b8cfa55),
	.w3(32'hb978f298),
	.w4(32'h3b601cde),
	.w5(32'hbb31bc3c),
	.w6(32'h3bc69e85),
	.w7(32'h3c2483a4),
	.w8(32'h3a4e68cc),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39befe6a),
	.w1(32'h3b8d89e6),
	.w2(32'hbb09e999),
	.w3(32'hbb620186),
	.w4(32'hbbbe4701),
	.w5(32'h3b451122),
	.w6(32'hb835c1dc),
	.w7(32'hbbcb29d1),
	.w8(32'h3aaaf04d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa69c0f),
	.w1(32'h3af52c90),
	.w2(32'hb9954813),
	.w3(32'hba073e7b),
	.w4(32'hbb17e71e),
	.w5(32'hba06c37f),
	.w6(32'h3aa31a3e),
	.w7(32'hbb42ed2c),
	.w8(32'hb92caee4),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b035a2b),
	.w1(32'hbb66824f),
	.w2(32'hba9595c8),
	.w3(32'hbb3ec402),
	.w4(32'h3b016325),
	.w5(32'h3bd66227),
	.w6(32'hba8d9373),
	.w7(32'hba470d6e),
	.w8(32'h3b3c711a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb06b3b),
	.w1(32'h3c0aaa73),
	.w2(32'h3c81b9c6),
	.w3(32'h3c2a486e),
	.w4(32'h3c94c669),
	.w5(32'h3afc7ab9),
	.w6(32'h3c403b57),
	.w7(32'h3c56ab2f),
	.w8(32'h3a7918d5),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acde517),
	.w1(32'hbae3d650),
	.w2(32'hba855c07),
	.w3(32'h3886f73e),
	.w4(32'h3b01af5c),
	.w5(32'hbc0c2122),
	.w6(32'hbb99f0ad),
	.w7(32'hbb0e688a),
	.w8(32'hbb862c3d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbfa20),
	.w1(32'h39170cca),
	.w2(32'h3bf2b711),
	.w3(32'hbb303920),
	.w4(32'h3afcbbce),
	.w5(32'h3bc4ee44),
	.w6(32'h3baf46f4),
	.w7(32'h3c26cc28),
	.w8(32'hb975ab3e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba357a68),
	.w1(32'hb786aeec),
	.w2(32'hbb605e24),
	.w3(32'h3a090c5f),
	.w4(32'h398af4e8),
	.w5(32'h3ad2a1f4),
	.w6(32'h3a00c069),
	.w7(32'h3a43dda8),
	.w8(32'h3b3564f7),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba755ba8),
	.w1(32'hba98f567),
	.w2(32'hbaf691b5),
	.w3(32'h3a626ccd),
	.w4(32'h3b0c5fc1),
	.w5(32'hbaf6972b),
	.w6(32'h3af52742),
	.w7(32'hba982eeb),
	.w8(32'h3a5310f0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0efc71),
	.w1(32'h3aa687ae),
	.w2(32'h3a865386),
	.w3(32'hbb57636d),
	.w4(32'hbb45049e),
	.w5(32'h391165c0),
	.w6(32'h3abb3c1d),
	.w7(32'h3ac1d141),
	.w8(32'hb8e2e87f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c658f),
	.w1(32'h3b99c66f),
	.w2(32'h3bd3d3f8),
	.w3(32'h3c3a7f66),
	.w4(32'h3c368a0e),
	.w5(32'hb8ce5d46),
	.w6(32'h3ac62421),
	.w7(32'h3c033d16),
	.w8(32'hbb0be195),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5464cf),
	.w1(32'hbb00040d),
	.w2(32'hbb459283),
	.w3(32'hbbc149b6),
	.w4(32'hbb30248a),
	.w5(32'hbb1b83db),
	.w6(32'hbbca9709),
	.w7(32'hbbc6bb24),
	.w8(32'hbbd7c7ec),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85b52d),
	.w1(32'hbc00b085),
	.w2(32'h3bc3c603),
	.w3(32'hba89e56e),
	.w4(32'h3c52a99e),
	.w5(32'h3b267b9c),
	.w6(32'hbc43257d),
	.w7(32'h3b4d854a),
	.w8(32'h3b908389),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaac8fe),
	.w1(32'hbb0e1044),
	.w2(32'hbbac2897),
	.w3(32'h3b3c3cab),
	.w4(32'h3a867483),
	.w5(32'h3bf26edd),
	.w6(32'h3a7a46d8),
	.w7(32'h3b11c208),
	.w8(32'h3b8da357),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77966d),
	.w1(32'hbb842c01),
	.w2(32'hbbded5d5),
	.w3(32'h3aa3b709),
	.w4(32'hbabdc9fd),
	.w5(32'hb7f6bc36),
	.w6(32'hb958f94d),
	.w7(32'hbb24a0ac),
	.w8(32'h3b12bbd2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9560852),
	.w1(32'hbb3c37c8),
	.w2(32'hbb91e407),
	.w3(32'h3aa2a975),
	.w4(32'hbba9c838),
	.w5(32'h3bcdc440),
	.w6(32'hb9f5490e),
	.w7(32'hbac2fdbe),
	.w8(32'h3aad9abb),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81908f),
	.w1(32'h3b03dcd1),
	.w2(32'hbb6944fc),
	.w3(32'h3bca465e),
	.w4(32'h3b071232),
	.w5(32'h3be35213),
	.w6(32'hb84ba883),
	.w7(32'hbb214b89),
	.w8(32'h3bd2ab3c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab88fb6),
	.w1(32'h3a92b78e),
	.w2(32'h3a942640),
	.w3(32'h3b8f8d46),
	.w4(32'h3b693269),
	.w5(32'h391a11a1),
	.w6(32'h3c028081),
	.w7(32'h3afc854a),
	.w8(32'h3c09f0f2),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18a4c3),
	.w1(32'hbb880a03),
	.w2(32'h3b87ea9c),
	.w3(32'hba6282ce),
	.w4(32'hbb30bc8a),
	.w5(32'h3b923f03),
	.w6(32'hbae5c30c),
	.w7(32'hba2cd9b2),
	.w8(32'h3c087b4d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e060f),
	.w1(32'h3c17db12),
	.w2(32'h3b994aea),
	.w3(32'hba4fd18b),
	.w4(32'hbad697fb),
	.w5(32'h3c1485da),
	.w6(32'hba14c467),
	.w7(32'hb9085596),
	.w8(32'hbbbf4369),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d8e3e),
	.w1(32'hbc92d7bd),
	.w2(32'hbb4e02bd),
	.w3(32'h3cddd9c9),
	.w4(32'h3bf8d490),
	.w5(32'hbbe7b563),
	.w6(32'hbc062af2),
	.w7(32'hbb729dab),
	.w8(32'hbb207241),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b615af9),
	.w1(32'h3bb1639e),
	.w2(32'h3b63c60c),
	.w3(32'hbbfff109),
	.w4(32'hbba118e7),
	.w5(32'hbb0b6a68),
	.w6(32'h3c02ebb1),
	.w7(32'h3b4b442d),
	.w8(32'hbc0d7806),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90a078),
	.w1(32'hbba3fef3),
	.w2(32'hbbc94e62),
	.w3(32'h3ad89604),
	.w4(32'h3b8e6024),
	.w5(32'h3acb2533),
	.w6(32'hbb1e3763),
	.w7(32'hbb05d1ca),
	.w8(32'h3a866f84),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f6e5f),
	.w1(32'hbbcb6584),
	.w2(32'h3a84d230),
	.w3(32'h3bae92fa),
	.w4(32'h3b5a5bdf),
	.w5(32'hbbd2a4fa),
	.w6(32'hbbc152a1),
	.w7(32'hbb070942),
	.w8(32'h398264aa),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396265b5),
	.w1(32'h3b986311),
	.w2(32'h3bb95326),
	.w3(32'hbc1bc885),
	.w4(32'hbbd498d7),
	.w5(32'hbbc9effd),
	.w6(32'h3be90461),
	.w7(32'h3b8750bc),
	.w8(32'hba743d9c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb247b2),
	.w1(32'h3bc04aa0),
	.w2(32'h3b06dc77),
	.w3(32'hbb60291e),
	.w4(32'hbbad7d16),
	.w5(32'h3c94b559),
	.w6(32'hbb7be1e2),
	.w7(32'hba894d8a),
	.w8(32'h3a5308ee),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34ebfd),
	.w1(32'hbcb323e3),
	.w2(32'hbc87a14c),
	.w3(32'h3d0c2331),
	.w4(32'h3c756c30),
	.w5(32'h3c00b684),
	.w6(32'hbb76ea4b),
	.w7(32'hbc1ee18a),
	.w8(32'h3be86e51),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f7ea5),
	.w1(32'hbbee75f9),
	.w2(32'hbbc194ae),
	.w3(32'h3caef2d0),
	.w4(32'h3c55d1d2),
	.w5(32'hb98372bb),
	.w6(32'h3b8e419f),
	.w7(32'hba8e637a),
	.w8(32'h3b15274e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a2968),
	.w1(32'hbaafff2b),
	.w2(32'h3a16c3de),
	.w3(32'h3bec5f01),
	.w4(32'h3a7da42a),
	.w5(32'hb94fe57a),
	.w6(32'h3bdc0d56),
	.w7(32'h3b37fa24),
	.w8(32'h3bb0bf3c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1dd26),
	.w1(32'h3b86a8d1),
	.w2(32'hbb302388),
	.w3(32'hbbf933f5),
	.w4(32'hbbfc582b),
	.w5(32'hba5e4ec9),
	.w6(32'hbb9afa9e),
	.w7(32'hbbe2b07f),
	.w8(32'h3b85e564),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6eaa3),
	.w1(32'h3b2f98e1),
	.w2(32'h3b144cd8),
	.w3(32'hbb60a8db),
	.w4(32'hbad47fc0),
	.w5(32'h3b42d61f),
	.w6(32'h3afd6b1c),
	.w7(32'h3b884981),
	.w8(32'hbb4fb810),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe91abd),
	.w1(32'hbb14e0ce),
	.w2(32'hbbde9270),
	.w3(32'h3a4fff3d),
	.w4(32'h3b0c2304),
	.w5(32'h3abfd64d),
	.w6(32'hbb65f808),
	.w7(32'hbba73319),
	.w8(32'h3bb8cd1c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01d3a5),
	.w1(32'hbc389892),
	.w2(32'hbabe2d2a),
	.w3(32'h3b65ac7c),
	.w4(32'h3b410ba7),
	.w5(32'h3c19a4ca),
	.w6(32'hbb30ee04),
	.w7(32'h3abe887c),
	.w8(32'h3c1f4403),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a365739),
	.w1(32'hbb900e49),
	.w2(32'hbb6b5692),
	.w3(32'h3b879a81),
	.w4(32'h3b6f5ff6),
	.w5(32'h3a9bdd06),
	.w6(32'hbb7eda05),
	.w7(32'hba9c75e1),
	.w8(32'hbaf9c3b3),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa52a7),
	.w1(32'hbc02beaf),
	.w2(32'hbbf1cd09),
	.w3(32'h3b433afd),
	.w4(32'h3c0478e4),
	.w5(32'h3c540d60),
	.w6(32'h3b8a9b42),
	.w7(32'h3a372e68),
	.w8(32'hbaa34ff1),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b8f04),
	.w1(32'hbc0dccee),
	.w2(32'hbb78a2b7),
	.w3(32'h3b73d680),
	.w4(32'hbaefdd1e),
	.w5(32'h3bbd2e79),
	.w6(32'hba080fee),
	.w7(32'hbb8b7360),
	.w8(32'h3aa383d1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb32625),
	.w1(32'hbc107e6f),
	.w2(32'hbb80ddc0),
	.w3(32'h3bdd3120),
	.w4(32'h3be705bd),
	.w5(32'hbc22d2e9),
	.w6(32'hbac2a3ec),
	.w7(32'hb9e0a8ee),
	.w8(32'h3af38436),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b861d85),
	.w1(32'h3c226d32),
	.w2(32'h3bf706c0),
	.w3(32'hbc2a2873),
	.w4(32'hbb6c6096),
	.w5(32'hbc015919),
	.w6(32'h3bae752c),
	.w7(32'h3be1e721),
	.w8(32'hba0263f0),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98ef50),
	.w1(32'h3b1665b0),
	.w2(32'h3791cae2),
	.w3(32'h3b7e1146),
	.w4(32'hbc0539b0),
	.w5(32'hbb16e7b0),
	.w6(32'hbad38391),
	.w7(32'hbb3b41cf),
	.w8(32'h3b9d5432),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baad22b),
	.w1(32'h3b218e89),
	.w2(32'h3bdcd142),
	.w3(32'hbb15dc04),
	.w4(32'hbb736517),
	.w5(32'hbaecaa65),
	.w6(32'hba021a4d),
	.w7(32'h3b7fdc3f),
	.w8(32'h3a678f6f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea4c7e),
	.w1(32'h3bc0615f),
	.w2(32'hb9b2e1a8),
	.w3(32'hbb60d6c5),
	.w4(32'hbbd64b09),
	.w5(32'h3af24660),
	.w6(32'h3b73afe0),
	.w7(32'hbab5e6a4),
	.w8(32'h3b2198a2),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4cbe2),
	.w1(32'hbc1dcb54),
	.w2(32'hbbc9f171),
	.w3(32'hbacf5040),
	.w4(32'h3b6053c4),
	.w5(32'h3958ca83),
	.w6(32'h3bb5738a),
	.w7(32'h3b44e9d4),
	.w8(32'h3b887ee0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58ff03),
	.w1(32'hbbcb105e),
	.w2(32'hbbc56e26),
	.w3(32'h3b4de85f),
	.w4(32'hba64c18b),
	.w5(32'h3c40f8be),
	.w6(32'hbada271b),
	.w7(32'hbb7f43c5),
	.w8(32'hbbbd080a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c54a8),
	.w1(32'hbb883f44),
	.w2(32'hbb04d613),
	.w3(32'h3cbad13e),
	.w4(32'h3c7bc2db),
	.w5(32'h3be597e1),
	.w6(32'hbba0a172),
	.w7(32'hbb624bf2),
	.w8(32'h3aa53fa1),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a643af9),
	.w1(32'hbba6d5a8),
	.w2(32'hbb72b51d),
	.w3(32'h3c52cd4e),
	.w4(32'h3bc1ea31),
	.w5(32'h3c1473ee),
	.w6(32'hbb1bd217),
	.w7(32'hb9dec8ce),
	.w8(32'hbbdca71c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c0d82),
	.w1(32'hbc0c8724),
	.w2(32'hbb8aa624),
	.w3(32'h3c2f5d99),
	.w4(32'h3c282598),
	.w5(32'hba04195e),
	.w6(32'h3a113077),
	.w7(32'hbae9ced2),
	.w8(32'h3a41db08),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0441a),
	.w1(32'hbb8a72ae),
	.w2(32'hbb88d49f),
	.w3(32'hbaf0beff),
	.w4(32'h3a5be90a),
	.w5(32'hbc00b770),
	.w6(32'h3c344f57),
	.w7(32'h3b893b71),
	.w8(32'hbafd2943),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ab78b),
	.w1(32'h3bdc5873),
	.w2(32'h3b85eb8a),
	.w3(32'hbac1aa31),
	.w4(32'hba2d47e6),
	.w5(32'h3c4e0535),
	.w6(32'h3b6b05f5),
	.w7(32'h3b049203),
	.w8(32'hbb34be65),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc124bd8),
	.w1(32'hbc48cbe1),
	.w2(32'h3a6f8a56),
	.w3(32'h3b712dde),
	.w4(32'hba494686),
	.w5(32'h3b09c551),
	.w6(32'h3a8fc8af),
	.w7(32'h3b907939),
	.w8(32'hbb175e0f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule