module layer_10_featuremap_298(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e78ab),
	.w1(32'hbc1b4d9e),
	.w2(32'h3b800c11),
	.w3(32'h3aa482d1),
	.w4(32'h3bb902ab),
	.w5(32'h3a5f3ae3),
	.w6(32'hba051c95),
	.w7(32'h3b112edb),
	.w8(32'h3b473b72),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad66ba5),
	.w1(32'h3b406b43),
	.w2(32'hbc6cf119),
	.w3(32'h3bc0c767),
	.w4(32'h3b89110c),
	.w5(32'hbc3e199f),
	.w6(32'h3b2664c6),
	.w7(32'hbbab242b),
	.w8(32'hbc8e0aeb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb846b74),
	.w1(32'hbc60e69c),
	.w2(32'hbb222afc),
	.w3(32'hbc509779),
	.w4(32'h3b0e6f8b),
	.w5(32'hbbe7238e),
	.w6(32'hbc8f2ee0),
	.w7(32'hbc5e8c34),
	.w8(32'hbc0a5b57),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918d15b),
	.w1(32'h3c6214bb),
	.w2(32'h3c243978),
	.w3(32'hbb1dfbaa),
	.w4(32'h3bfac5b4),
	.w5(32'hb94271bf),
	.w6(32'h3c2e024a),
	.w7(32'h3c82f243),
	.w8(32'hbb20fc12),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97d625),
	.w1(32'h3c13742c),
	.w2(32'h3c057a46),
	.w3(32'h3b53944c),
	.w4(32'h3a37729b),
	.w5(32'hbc218d66),
	.w6(32'h3b9f1e21),
	.w7(32'h3b331ffc),
	.w8(32'hbbaee9cf),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f0f2b),
	.w1(32'h3c678512),
	.w2(32'h3c4c8c51),
	.w3(32'hbac2d51e),
	.w4(32'h3bd57738),
	.w5(32'hbc41ee71),
	.w6(32'h3b9ba334),
	.w7(32'h3c5b16ff),
	.w8(32'hbb9de9bd),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e0d98),
	.w1(32'h3c1b6af5),
	.w2(32'h3bd06215),
	.w3(32'hbafdcb2f),
	.w4(32'h3c1a06cb),
	.w5(32'hbc2f51eb),
	.w6(32'h3bed8dd0),
	.w7(32'h3c4fb348),
	.w8(32'hbc325019),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98cd45),
	.w1(32'h3c8cca98),
	.w2(32'h3ca65ac3),
	.w3(32'hbc5103f0),
	.w4(32'h3b8cd52a),
	.w5(32'h3b082a34),
	.w6(32'h3b922e4d),
	.w7(32'h3cac2cea),
	.w8(32'h3b0ca7de),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fcd62),
	.w1(32'h3c573dd8),
	.w2(32'h3c4387c0),
	.w3(32'h3afabd91),
	.w4(32'h3c029622),
	.w5(32'hbc67cbe3),
	.w6(32'h3bc604dc),
	.w7(32'h3c4950b9),
	.w8(32'hbc4c4b19),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf402c8),
	.w1(32'h3c27fc0e),
	.w2(32'h3c701e43),
	.w3(32'hbbb5090a),
	.w4(32'h3b5866b4),
	.w5(32'hbc0184db),
	.w6(32'hbaaa1608),
	.w7(32'h3c295d2c),
	.w8(32'hbbbe5d8d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affc01e),
	.w1(32'h3c2572bd),
	.w2(32'h3b74384b),
	.w3(32'hba38ecbb),
	.w4(32'h3c0f71fc),
	.w5(32'h3be0663a),
	.w6(32'h3c0c95f1),
	.w7(32'h3c22e4f6),
	.w8(32'hbb4ac933),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92f136),
	.w1(32'hbca64214),
	.w2(32'hbc3ac6c6),
	.w3(32'h3b932eec),
	.w4(32'hbb11b107),
	.w5(32'h3d07311b),
	.w6(32'hbbacf205),
	.w7(32'hbc9241eb),
	.w8(32'h3cb7597d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12e154),
	.w1(32'hbb74f910),
	.w2(32'hbcb4b5b6),
	.w3(32'h3ce083b5),
	.w4(32'hbba161b4),
	.w5(32'h3b880339),
	.w6(32'h3c61367e),
	.w7(32'hbc57e51e),
	.w8(32'h3bff7556),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395021ac),
	.w1(32'hbbd9686f),
	.w2(32'h3b408651),
	.w3(32'h3b5237e1),
	.w4(32'h39c5234d),
	.w5(32'hbb2a9318),
	.w6(32'hbc0838ab),
	.w7(32'hba3f0b15),
	.w8(32'hbbfdefe3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb704829),
	.w1(32'h3a8fcf63),
	.w2(32'hbba40039),
	.w3(32'hbb47b584),
	.w4(32'hbc05939b),
	.w5(32'h3ac4fdd0),
	.w6(32'h3a4f8069),
	.w7(32'h3a75391c),
	.w8(32'h3b15ce36),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb219f6d),
	.w1(32'h3b2f4b5a),
	.w2(32'h3beecb39),
	.w3(32'hbaa7c8d7),
	.w4(32'hbb988bb0),
	.w5(32'hbaa32248),
	.w6(32'h3b78e877),
	.w7(32'hbb278a19),
	.w8(32'h3bbce491),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1008a1),
	.w1(32'h3bde05a4),
	.w2(32'h3b8f434b),
	.w3(32'h3c09e928),
	.w4(32'h3c1c5723),
	.w5(32'h3c0bc1ba),
	.w6(32'h3c4e0d33),
	.w7(32'h3c87119a),
	.w8(32'h3c1c10db),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb7924),
	.w1(32'hbc667ecb),
	.w2(32'hbc23bec8),
	.w3(32'hbad5b6a9),
	.w4(32'hbb74ec7e),
	.w5(32'h3c57ed14),
	.w6(32'hbbfea9d7),
	.w7(32'hbc309a2d),
	.w8(32'h3bed3068),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba31e53),
	.w1(32'hb89478ee),
	.w2(32'hbaa58599),
	.w3(32'hb8dbfa97),
	.w4(32'hbbf1e0e0),
	.w5(32'h3bbd2a55),
	.w6(32'hbc0fdd9e),
	.w7(32'hbc089285),
	.w8(32'h3c0f937e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ae499),
	.w1(32'h398661a0),
	.w2(32'h3b96226c),
	.w3(32'hbbcf8441),
	.w4(32'hb9db2aa8),
	.w5(32'h3b0de7e5),
	.w6(32'h3b596a29),
	.w7(32'hbb763f5a),
	.w8(32'h3b52122c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b384bf9),
	.w1(32'hbb2d865c),
	.w2(32'h3ab34207),
	.w3(32'h3b1cfc7d),
	.w4(32'hbb95c90a),
	.w5(32'hbce0a9b1),
	.w6(32'h3bc79132),
	.w7(32'hbae6489d),
	.w8(32'hbc74a44a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fe7e1),
	.w1(32'h3c9ef4cc),
	.w2(32'h3cd6910f),
	.w3(32'hbc1343bf),
	.w4(32'h3c047beb),
	.w5(32'hbb401736),
	.w6(32'h3c13ebf7),
	.w7(32'h3cd2a451),
	.w8(32'hbb844c38),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ca65b),
	.w1(32'hbb582459),
	.w2(32'h3aebe3b1),
	.w3(32'hbb33491b),
	.w4(32'h3bad470b),
	.w5(32'h3c73018b),
	.w6(32'hbc1c6bc6),
	.w7(32'hba204071),
	.w8(32'h3c612c4e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baec478),
	.w1(32'h3b1f27ee),
	.w2(32'h3b18932b),
	.w3(32'h3b87d6ec),
	.w4(32'hb90cc018),
	.w5(32'h3b966b85),
	.w6(32'hbb3566b9),
	.w7(32'hbb982c0e),
	.w8(32'h3b143c16),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b512271),
	.w1(32'hbad17554),
	.w2(32'h39e5223f),
	.w3(32'h3b90f781),
	.w4(32'h3b2eedf7),
	.w5(32'hbc6ac2f8),
	.w6(32'hbbab7055),
	.w7(32'hbc1b5ec4),
	.w8(32'hbc995903),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8ca4e),
	.w1(32'h3b5b71dd),
	.w2(32'h388e0714),
	.w3(32'hbc07de40),
	.w4(32'hbbf530b6),
	.w5(32'hbca40f34),
	.w6(32'h3a55cbac),
	.w7(32'h3c1030a8),
	.w8(32'hbc541277),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15c092),
	.w1(32'h3c3c441e),
	.w2(32'h3b9cf0d8),
	.w3(32'hbc53f078),
	.w4(32'hbbc0e251),
	.w5(32'hbbe0ae24),
	.w6(32'h3bbbe206),
	.w7(32'h3affd248),
	.w8(32'hb910b15d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c54c7),
	.w1(32'hba9fd3d8),
	.w2(32'h3b2020eb),
	.w3(32'hbad91693),
	.w4(32'hbb544e7b),
	.w5(32'h3b2a6cdc),
	.w6(32'h3abd43f3),
	.w7(32'h3b0318b2),
	.w8(32'hbb97dd17),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8afaf1),
	.w1(32'hbb029fbb),
	.w2(32'h3a28070f),
	.w3(32'h3bdf0187),
	.w4(32'h3be21326),
	.w5(32'h3a337d18),
	.w6(32'h3a34083d),
	.w7(32'h3bae0a6e),
	.w8(32'h3c3e2c07),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4427c5),
	.w1(32'h3a5170f9),
	.w2(32'h3b8b228b),
	.w3(32'h3b3e0968),
	.w4(32'hbaf24271),
	.w5(32'h3bb8b7f0),
	.w6(32'h3b69931a),
	.w7(32'hbb21c958),
	.w8(32'hbc2566c7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc718bf8),
	.w1(32'hbc85d38b),
	.w2(32'hbc984e40),
	.w3(32'hbb4177e9),
	.w4(32'hbc6bb76f),
	.w5(32'hbbdc8f3e),
	.w6(32'hbb9426be),
	.w7(32'hbc7d69de),
	.w8(32'h3bd55065),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc314836),
	.w1(32'hbc43a3f8),
	.w2(32'hbc7a0d7e),
	.w3(32'hb9c29fa7),
	.w4(32'h3b87630e),
	.w5(32'hbbc8e35c),
	.w6(32'hbc41158d),
	.w7(32'hbcaa1d58),
	.w8(32'hbc97a89f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b0199),
	.w1(32'hbc353534),
	.w2(32'hbbaa3c29),
	.w3(32'hbc5830e5),
	.w4(32'hbc93ccb2),
	.w5(32'h3bfd8367),
	.w6(32'hbca78c35),
	.w7(32'hbc46c55e),
	.w8(32'h3bdfcae2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae0f2f),
	.w1(32'hbcb20c9f),
	.w2(32'hbcb49278),
	.w3(32'h3b99e586),
	.w4(32'hbc45d310),
	.w5(32'h3a033ceb),
	.w6(32'hbc0e90c7),
	.w7(32'hbc898508),
	.w8(32'hbbe6d8e8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace0398),
	.w1(32'h3ae750c9),
	.w2(32'h3b823ce1),
	.w3(32'hbafb55b9),
	.w4(32'h3bb2b7c3),
	.w5(32'h3b9a7383),
	.w6(32'h3b82576a),
	.w7(32'hb9dfd34d),
	.w8(32'h3b31f49b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e4642),
	.w1(32'hbc859f54),
	.w2(32'hbc74ba48),
	.w3(32'h3b6d94ad),
	.w4(32'hbc4370a6),
	.w5(32'h3c12bf7e),
	.w6(32'hbbcbabf4),
	.w7(32'hbc836f73),
	.w8(32'hbc3e9ec6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1dbe8),
	.w1(32'hbb2c0542),
	.w2(32'hbc367a8e),
	.w3(32'h3c2059d8),
	.w4(32'h3b46e87b),
	.w5(32'hbbfc3b7e),
	.w6(32'hbbf3c7be),
	.w7(32'hbc48ae02),
	.w8(32'hbacd699f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d9477),
	.w1(32'h3c601637),
	.w2(32'h3a8d27bb),
	.w3(32'h3aa406aa),
	.w4(32'hbbb28146),
	.w5(32'h3b6fdd6d),
	.w6(32'h3b937ed8),
	.w7(32'hb87f8fee),
	.w8(32'hbb029917),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb4fbd),
	.w1(32'h3ae71587),
	.w2(32'hbc5e5230),
	.w3(32'h3c4a1613),
	.w4(32'h3bacfadd),
	.w5(32'hbcd36511),
	.w6(32'h3aeebca5),
	.w7(32'hbb49298e),
	.w8(32'hbbb28c87),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a63f7),
	.w1(32'h3c729de0),
	.w2(32'h3ce793b9),
	.w3(32'hbb9ebafd),
	.w4(32'h3c77eb3c),
	.w5(32'h3c149631),
	.w6(32'h3c146a33),
	.w7(32'h3cdf862f),
	.w8(32'h3b9ec99f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b453b91),
	.w1(32'hbba01117),
	.w2(32'hbaf6e6f8),
	.w3(32'h3ba75543),
	.w4(32'h3a6551bf),
	.w5(32'hbccb2018),
	.w6(32'hbbed2119),
	.w7(32'h3aa26a08),
	.w8(32'hbc64ee6b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc395874),
	.w1(32'h3bf13cfb),
	.w2(32'h3bb8842c),
	.w3(32'hbbafbc1c),
	.w4(32'h3bc09ea5),
	.w5(32'h3cc649f4),
	.w6(32'h3c90a649),
	.w7(32'h3c86b251),
	.w8(32'h3cbf2bc0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafec2af),
	.w1(32'hbbd3cdb9),
	.w2(32'hbc4b5768),
	.w3(32'h3c4a984b),
	.w4(32'hba23bb51),
	.w5(32'h3adf1b78),
	.w6(32'hbb8f560d),
	.w7(32'hbc9e5d82),
	.w8(32'h3abcf707),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ac3e7),
	.w1(32'hbaf3c8b4),
	.w2(32'hbbd27433),
	.w3(32'h3c353088),
	.w4(32'h3be678e0),
	.w5(32'hbc084e5c),
	.w6(32'hbc14ec1e),
	.w7(32'hbbcd256c),
	.w8(32'h3b5c125d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b939bb5),
	.w1(32'h3c3c3d6d),
	.w2(32'h3c41eee3),
	.w3(32'h3b9bca3c),
	.w4(32'h3c3eadc0),
	.w5(32'hbc041ff0),
	.w6(32'h3c82f324),
	.w7(32'h3c860d7d),
	.w8(32'h3c160578),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc80437),
	.w1(32'hbc4c062b),
	.w2(32'hbc55783c),
	.w3(32'hba247d67),
	.w4(32'hbb539374),
	.w5(32'hbc23a7cf),
	.w6(32'h3c992699),
	.w7(32'h3b0e15a8),
	.w8(32'hbbbb7449),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e8a94),
	.w1(32'hb9adf345),
	.w2(32'h3b71d5a3),
	.w3(32'h3ac8511f),
	.w4(32'hbadbbf40),
	.w5(32'hbb33d6f6),
	.w6(32'h3b146bca),
	.w7(32'hba7a0b2d),
	.w8(32'hbbe1aa34),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5eb559),
	.w1(32'h3ca6497a),
	.w2(32'h3c940f33),
	.w3(32'hbb378841),
	.w4(32'h3c1fa7e1),
	.w5(32'h3cd29345),
	.w6(32'h3b07d1b8),
	.w7(32'h3c961fcd),
	.w8(32'h3ca37ce8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf66e75),
	.w1(32'hbbb73607),
	.w2(32'hbc7fb7e6),
	.w3(32'h3c971132),
	.w4(32'h3b279edc),
	.w5(32'hbcef6fd5),
	.w6(32'h3c00c40a),
	.w7(32'hbc0363e6),
	.w8(32'hbc3f3572),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b21ba),
	.w1(32'h3c9eec15),
	.w2(32'h3ccaae76),
	.w3(32'hbbe3a519),
	.w4(32'h3ba08057),
	.w5(32'hba6a0ab2),
	.w6(32'h3c784414),
	.w7(32'h3cc374e0),
	.w8(32'hbc0050a6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40f362),
	.w1(32'hbc07f1eb),
	.w2(32'hbc29d8ab),
	.w3(32'hbbf555c6),
	.w4(32'hbc523ed4),
	.w5(32'h3c3f915e),
	.w6(32'hbc8dadab),
	.w7(32'hbc9b2802),
	.w8(32'h3c23cdd1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3e451),
	.w1(32'hbaf7bc2b),
	.w2(32'hbbdbb275),
	.w3(32'h3c2822af),
	.w4(32'h3b7c58e6),
	.w5(32'hbba214ed),
	.w6(32'h3a958f60),
	.w7(32'hbc3216b9),
	.w8(32'hbba0834a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b086790),
	.w1(32'hba5eee2f),
	.w2(32'h3b17e664),
	.w3(32'hba0dbb28),
	.w4(32'hbb0fb1e9),
	.w5(32'hbbcb75b7),
	.w6(32'hbbab6841),
	.w7(32'hbb6c7d6c),
	.w8(32'h3ae35ff1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0018b5),
	.w1(32'hbc610e46),
	.w2(32'hbc400562),
	.w3(32'hb8096e95),
	.w4(32'hb92bad94),
	.w5(32'h3c40f5be),
	.w6(32'h3922317d),
	.w7(32'hbca2b77c),
	.w8(32'h3c59f9f0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b71fb),
	.w1(32'hbb5f4bda),
	.w2(32'h378e4e33),
	.w3(32'hbb13f9ab),
	.w4(32'h3b0791d5),
	.w5(32'h3b0a800a),
	.w6(32'h3a8ab6cc),
	.w7(32'hbc02df16),
	.w8(32'h3c407ec5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3376e),
	.w1(32'h3b109472),
	.w2(32'h3b9bb963),
	.w3(32'hbbd949ff),
	.w4(32'h3993a306),
	.w5(32'h3c0fae8e),
	.w6(32'h3c04da8b),
	.w7(32'h3ad2a577),
	.w8(32'h3b9186a6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ffd62),
	.w1(32'hbb981927),
	.w2(32'hbbd9074f),
	.w3(32'hba2ae9c8),
	.w4(32'hbacdd525),
	.w5(32'hbc755ec3),
	.w6(32'hbb9b3bce),
	.w7(32'hbb5aa1f1),
	.w8(32'hbc3ecbcd),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe69401),
	.w1(32'hbc84f34b),
	.w2(32'hbb694dc2),
	.w3(32'hbc06b30b),
	.w4(32'h39048785),
	.w5(32'hbcff864c),
	.w6(32'hbc60c00d),
	.w7(32'hbbbf9d03),
	.w8(32'hbc8b72c3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb155c7),
	.w1(32'h3c37e183),
	.w2(32'h3c84786f),
	.w3(32'hbc13b46d),
	.w4(32'h3b8319ed),
	.w5(32'hbc1a3995),
	.w6(32'h3c35998f),
	.w7(32'h3c9dc586),
	.w8(32'hbbd3e0fc),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b909e77),
	.w1(32'h3c9e2877),
	.w2(32'h3b26e182),
	.w3(32'h395867df),
	.w4(32'h3baab9d7),
	.w5(32'hbaa38ce5),
	.w6(32'h3c09f7de),
	.w7(32'h3c290711),
	.w8(32'hbae833c2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb581295),
	.w1(32'h3ac1820d),
	.w2(32'h39a14d5b),
	.w3(32'hbabb6bae),
	.w4(32'hbb21a56c),
	.w5(32'hbc3c853f),
	.w6(32'hbb0a7b89),
	.w7(32'hba686674),
	.w8(32'hbbb930b7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c03e9),
	.w1(32'hb87f3230),
	.w2(32'hba48ced6),
	.w3(32'hbb99f6dd),
	.w4(32'hba886757),
	.w5(32'hbab62234),
	.w6(32'h3c373645),
	.w7(32'h3c0cbcc7),
	.w8(32'h3a710b2f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb701b9c),
	.w1(32'h3a8ff003),
	.w2(32'h3aed36a5),
	.w3(32'h39a3f265),
	.w4(32'h3b84a7cc),
	.w5(32'h3bfdd9f9),
	.w6(32'hbb3df006),
	.w7(32'hbbc66aa0),
	.w8(32'h3bc3eb39),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98fe9f),
	.w1(32'hbb21a4df),
	.w2(32'h3b0294dd),
	.w3(32'h3a90d10d),
	.w4(32'h3b59e1d7),
	.w5(32'hbb7ba0de),
	.w6(32'h3a948558),
	.w7(32'h3a38eddd),
	.w8(32'hbb5688a0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba933370),
	.w1(32'hbb4d5fee),
	.w2(32'hbb4d2dbd),
	.w3(32'hbbf236d3),
	.w4(32'h3b0415a7),
	.w5(32'h3c047c7b),
	.w6(32'hbb7c40a8),
	.w7(32'hbc187081),
	.w8(32'h3c288e5f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab214a2),
	.w1(32'hbb6817fd),
	.w2(32'h3b0ddb37),
	.w3(32'h3b222a53),
	.w4(32'hbab2ee3a),
	.w5(32'hbc0f53f2),
	.w6(32'hbb8a64ff),
	.w7(32'hbc44e54c),
	.w8(32'hbb51716b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb140126),
	.w1(32'h3baf0232),
	.w2(32'h3bc1849e),
	.w3(32'hbc1b89d2),
	.w4(32'h3944a68f),
	.w5(32'h3c9a6f48),
	.w6(32'h3c50cd26),
	.w7(32'h3bcae166),
	.w8(32'h3c4f6732),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b11a2),
	.w1(32'h3bf329d7),
	.w2(32'hbc017c8c),
	.w3(32'h3bef1132),
	.w4(32'h3aaae072),
	.w5(32'h3aa027ae),
	.w6(32'hbbabc972),
	.w7(32'hbc047744),
	.w8(32'h3b1c06ad),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa74fd0),
	.w1(32'hbb230d25),
	.w2(32'h3b3a50aa),
	.w3(32'hbc17fe51),
	.w4(32'hbb20b239),
	.w5(32'hbbd48420),
	.w6(32'hbc2a379a),
	.w7(32'hbb83be87),
	.w8(32'h3b8dc64c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56b854),
	.w1(32'hbc71966e),
	.w2(32'hbc8f5284),
	.w3(32'h3b893288),
	.w4(32'hbc3fc4e5),
	.w5(32'hbc0e63de),
	.w6(32'hbb7cdff0),
	.w7(32'hbc6433b3),
	.w8(32'hbc9fdc2b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8394d),
	.w1(32'h3b25c4d3),
	.w2(32'h3b44e00e),
	.w3(32'h3a44f523),
	.w4(32'hbbca0bdc),
	.w5(32'h3c0e1a31),
	.w6(32'hbba6093f),
	.w7(32'hbb590e8d),
	.w8(32'h3be6b57a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc00800),
	.w1(32'hbbb407c5),
	.w2(32'h38a1ba20),
	.w3(32'h3c23e7d1),
	.w4(32'h3b0a48de),
	.w5(32'h3c7124d8),
	.w6(32'h3a5bb7e4),
	.w7(32'hbb721c2e),
	.w8(32'h3c466969),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e845d1),
	.w1(32'hbbc66249),
	.w2(32'hbb9df2f0),
	.w3(32'h3b6154b3),
	.w4(32'h39e58be4),
	.w5(32'h3c946c60),
	.w6(32'h3b1c6c41),
	.w7(32'hbb5633d7),
	.w8(32'h3c0c07c9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86bb90),
	.w1(32'hbc8735ce),
	.w2(32'hbce78b67),
	.w3(32'h3cb5037c),
	.w4(32'hbb3179f9),
	.w5(32'h3a7ca010),
	.w6(32'h3b333463),
	.w7(32'hbc32c2f4),
	.w8(32'h3bbf7702),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38344a9c),
	.w1(32'hba9885d8),
	.w2(32'hbba4bd8a),
	.w3(32'h3a3a2eb8),
	.w4(32'h3b240793),
	.w5(32'h3d397646),
	.w6(32'h3c2f6021),
	.w7(32'h3ba9b907),
	.w8(32'h3cf7a07e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c4e6c),
	.w1(32'hbcc47577),
	.w2(32'hbd1ebf79),
	.w3(32'h3cb5071b),
	.w4(32'hbbebd5f9),
	.w5(32'h3c20a299),
	.w6(32'hbbbaf5bd),
	.w7(32'hbcf03e6c),
	.w8(32'h3bad65bd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd85d0),
	.w1(32'hba309e9f),
	.w2(32'h3baecd5a),
	.w3(32'hbb5c87d5),
	.w4(32'hbb53dda8),
	.w5(32'h3b164a42),
	.w6(32'hbc385813),
	.w7(32'h3a3b7796),
	.w8(32'h3c0bc39f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b446067),
	.w1(32'hbc3c56ee),
	.w2(32'hbb72d483),
	.w3(32'hba392661),
	.w4(32'hbbb5cc03),
	.w5(32'h3c0cc89d),
	.w6(32'hbc0e836f),
	.w7(32'hbc0a179d),
	.w8(32'h3b621088),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83eaaa),
	.w1(32'h3b727673),
	.w2(32'h3b5a9fff),
	.w3(32'h3bfde838),
	.w4(32'h3ba360b1),
	.w5(32'h3a6133f1),
	.w6(32'h3bbdd02b),
	.w7(32'hbac5f4b7),
	.w8(32'hbb05848a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcf79f),
	.w1(32'h3b0dcb5c),
	.w2(32'h3b8a28e9),
	.w3(32'h3b92cd7e),
	.w4(32'h3bbea31d),
	.w5(32'h3c63897e),
	.w6(32'h3b34af61),
	.w7(32'h3bfe4ab0),
	.w8(32'h3bcf171a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34f641),
	.w1(32'h3a9bf056),
	.w2(32'hbc00c360),
	.w3(32'h3a5f7594),
	.w4(32'h3a110be2),
	.w5(32'h3cba860e),
	.w6(32'h3a7bce71),
	.w7(32'hbac6f23d),
	.w8(32'h3c9880d6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cd2b1),
	.w1(32'hbca93d02),
	.w2(32'hbcd1e6f7),
	.w3(32'h3c413ddc),
	.w4(32'hbc12b68e),
	.w5(32'h3bd28b61),
	.w6(32'hbb3a64fa),
	.w7(32'hbc8ff9a0),
	.w8(32'h3b317e35),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a2abd),
	.w1(32'hbb9cd0aa),
	.w2(32'h3b33b1f8),
	.w3(32'h3b15effb),
	.w4(32'hb8cbfd7c),
	.w5(32'hbc514297),
	.w6(32'hbc06b570),
	.w7(32'hbb850cca),
	.w8(32'hbc6429ba),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb942b3c),
	.w1(32'h3c1bf397),
	.w2(32'hbb96865d),
	.w3(32'hbc0f8eca),
	.w4(32'hbb444b66),
	.w5(32'hbb22d334),
	.w6(32'h3b27e67e),
	.w7(32'h3b3904ae),
	.w8(32'hbafc3dcf),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8634676),
	.w1(32'hbbd3cc5f),
	.w2(32'hb92587f3),
	.w3(32'h3b15f533),
	.w4(32'h3962160c),
	.w5(32'h3b34fa0d),
	.w6(32'hbb2cc341),
	.w7(32'hbb741edb),
	.w8(32'hbae778d9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c8e23),
	.w1(32'hbc428562),
	.w2(32'hbb1930d0),
	.w3(32'hbb8caaf1),
	.w4(32'hb91b371d),
	.w5(32'hbc71ab65),
	.w6(32'h3af827aa),
	.w7(32'h3a767d3d),
	.w8(32'hbc9182d2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e8f88),
	.w1(32'hbc8ef280),
	.w2(32'hbc6d6d7b),
	.w3(32'hbcb1e5ce),
	.w4(32'hbbdce0d8),
	.w5(32'hbb27f660),
	.w6(32'hbc1b8e6a),
	.w7(32'hbc23e444),
	.w8(32'hbbf2a766),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5ef70),
	.w1(32'h3aafede7),
	.w2(32'h3b68c63c),
	.w3(32'hbbb1ec0f),
	.w4(32'hbbc69fe3),
	.w5(32'hbc7576a5),
	.w6(32'hbb319a6a),
	.w7(32'hbbb40588),
	.w8(32'hbb8a87d7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb265a54),
	.w1(32'h3c5bb0b7),
	.w2(32'h3c2f0bf6),
	.w3(32'h3abe0f62),
	.w4(32'h3b99c2de),
	.w5(32'h3bd070e6),
	.w6(32'h3c34db64),
	.w7(32'h3c6230d8),
	.w8(32'h3b73b573),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8b940),
	.w1(32'h3b886422),
	.w2(32'h3bfcc437),
	.w3(32'hba892dd4),
	.w4(32'h3b8d8b1f),
	.w5(32'h3b7d3acb),
	.w6(32'hbc43911c),
	.w7(32'h3b09f066),
	.w8(32'h3b21d374),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad15229),
	.w1(32'hb98ed7a0),
	.w2(32'hbc46003b),
	.w3(32'hbbd3af3f),
	.w4(32'hbb1cecc5),
	.w5(32'hbbd689fa),
	.w6(32'h3b824053),
	.w7(32'hbbabf547),
	.w8(32'h3b41f4db),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bfec7),
	.w1(32'h3a32ad1d),
	.w2(32'h3c0395ea),
	.w3(32'hbc2a1e13),
	.w4(32'hbb8a8ca0),
	.w5(32'hbc96ff59),
	.w6(32'hbbb1555c),
	.w7(32'h3a0e8e04),
	.w8(32'hbbd9c352),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390aa40d),
	.w1(32'hbc101d29),
	.w2(32'hbb905921),
	.w3(32'hbb5dfaf2),
	.w4(32'hba8daef9),
	.w5(32'hbbb67491),
	.w6(32'hbb9250f9),
	.w7(32'hbb87501e),
	.w8(32'hbc555bae),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec826d),
	.w1(32'hbb878964),
	.w2(32'h3b9f1bd3),
	.w3(32'hbc25d76a),
	.w4(32'h3be8aec6),
	.w5(32'hbbe58956),
	.w6(32'hbc855cc2),
	.w7(32'hbb4c3dd2),
	.w8(32'hbba8623f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadf5a5),
	.w1(32'h38ee179e),
	.w2(32'h3b3e1cbb),
	.w3(32'hbad8d04f),
	.w4(32'hbbed7325),
	.w5(32'hbc99ba8f),
	.w6(32'hbb485c03),
	.w7(32'hbbe19d77),
	.w8(32'h3bf4b991),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8f4e5),
	.w1(32'hbc66431f),
	.w2(32'hbc1dab14),
	.w3(32'hbc40ef87),
	.w4(32'h3b8d5821),
	.w5(32'h3b1d9e77),
	.w6(32'hbb8a2451),
	.w7(32'hbca00504),
	.w8(32'hbaca4e78),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f6772),
	.w1(32'h3a9e8ddd),
	.w2(32'hbc0d07d7),
	.w3(32'h3ae29f98),
	.w4(32'h3b8940cb),
	.w5(32'hbb03c4bc),
	.w6(32'hba3e87d9),
	.w7(32'hbbd61f72),
	.w8(32'hbc80f068),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4697ee),
	.w1(32'hbb8a54af),
	.w2(32'h3becb411),
	.w3(32'hbc29180f),
	.w4(32'hbc6bcb1c),
	.w5(32'h3a5da61c),
	.w6(32'hbcc8d36a),
	.w7(32'hba24ce5a),
	.w8(32'h3903de64),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2dda3),
	.w1(32'h39a8bbcb),
	.w2(32'h375907b5),
	.w3(32'hba999dc7),
	.w4(32'hba954fa5),
	.w5(32'hbbbdaa78),
	.w6(32'hbba79b54),
	.w7(32'hbbcc5330),
	.w8(32'hbc0b4dfd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ba25a),
	.w1(32'h3b14a5e2),
	.w2(32'h3c33d061),
	.w3(32'hbbca3c48),
	.w4(32'h3b93433f),
	.w5(32'h3c4c0543),
	.w6(32'hbc23beaa),
	.w7(32'h3ac63482),
	.w8(32'h3c86b365),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0edeb),
	.w1(32'hbad1a316),
	.w2(32'hbacb1c37),
	.w3(32'h3bad07a6),
	.w4(32'h3bb7d3a0),
	.w5(32'hba43e43d),
	.w6(32'h3bd9f556),
	.w7(32'h3c034bd6),
	.w8(32'hbc48bb20),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87b9b1),
	.w1(32'hbaa38d20),
	.w2(32'h3b928509),
	.w3(32'h3abf1499),
	.w4(32'h3bc7b94f),
	.w5(32'hbb0d3927),
	.w6(32'hbba1ff9a),
	.w7(32'hbbc9566a),
	.w8(32'hbb64266d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61981e),
	.w1(32'h3b3f70b1),
	.w2(32'h3a98f8aa),
	.w3(32'hb8321ad2),
	.w4(32'h3b1e8a3d),
	.w5(32'h3c504b9f),
	.w6(32'h3b094359),
	.w7(32'h3abd3aaa),
	.w8(32'h3b27babd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c137714),
	.w1(32'h3bedd458),
	.w2(32'h3c250594),
	.w3(32'h3c190f14),
	.w4(32'h3c494e9b),
	.w5(32'h3c41fc9f),
	.w6(32'hbb849723),
	.w7(32'h3b508f3e),
	.w8(32'h38289c57),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05e598),
	.w1(32'h3ba53d00),
	.w2(32'h3a66a347),
	.w3(32'h3926f1a1),
	.w4(32'hba13fe3e),
	.w5(32'h3bae446c),
	.w6(32'hbc18d0cd),
	.w7(32'hbba1aebc),
	.w8(32'h3b7ec818),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18306a),
	.w1(32'hbbe5cab5),
	.w2(32'hbb225b5e),
	.w3(32'hbb72f932),
	.w4(32'hb990ec45),
	.w5(32'h3b867b7b),
	.w6(32'hbb67f25e),
	.w7(32'h3ae8661b),
	.w8(32'h3a1eb87e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e0250),
	.w1(32'h3af38149),
	.w2(32'hbbc61125),
	.w3(32'hba4c7499),
	.w4(32'hbaf1e8cf),
	.w5(32'h3b31cdad),
	.w6(32'hbc16d69b),
	.w7(32'hbba02699),
	.w8(32'h3ab18cbe),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1dea28),
	.w1(32'h3b758059),
	.w2(32'h3ad21b9f),
	.w3(32'h3beec93c),
	.w4(32'h3b31a221),
	.w5(32'hbb5c920f),
	.w6(32'h3bbc3333),
	.w7(32'h3b0f12c2),
	.w8(32'hbb80995b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1101c),
	.w1(32'hbb5e28e7),
	.w2(32'hbbd1b57b),
	.w3(32'h39b2be8c),
	.w4(32'hbadd76a9),
	.w5(32'hbae5135e),
	.w6(32'hbbf40b0d),
	.w7(32'hbc08c0f3),
	.w8(32'hbad28e79),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09fa48),
	.w1(32'h39b410ea),
	.w2(32'hbbef1f26),
	.w3(32'h3b536f5d),
	.w4(32'hbb4013ec),
	.w5(32'h3a8a90fc),
	.w6(32'h3baae3d4),
	.w7(32'hbb53c660),
	.w8(32'h3ae20930),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc82e1e),
	.w1(32'h3b763a25),
	.w2(32'hba8a2a2f),
	.w3(32'h3b3b7909),
	.w4(32'h3bb0abd3),
	.w5(32'h3a79ba8e),
	.w6(32'hb949f770),
	.w7(32'hbaaa7330),
	.w8(32'hbaef394f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d175d4),
	.w1(32'h3b4bb3e2),
	.w2(32'h3a86d698),
	.w3(32'hba4c31d8),
	.w4(32'hb9e02e9f),
	.w5(32'hbb68cbc3),
	.w6(32'hbb83abc8),
	.w7(32'hbb2588e1),
	.w8(32'h3ac0aa63),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea7d29),
	.w1(32'h3b404f42),
	.w2(32'hbbe97221),
	.w3(32'hba78ec0c),
	.w4(32'hbbafb0d5),
	.w5(32'hbb517c57),
	.w6(32'h3c4b9917),
	.w7(32'hbaae3117),
	.w8(32'h3a4357bb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e9bc6c),
	.w1(32'hba923ecd),
	.w2(32'h3b0fd9d2),
	.w3(32'hbbeda46d),
	.w4(32'hbaa6682e),
	.w5(32'hbc194420),
	.w6(32'hba65de03),
	.w7(32'h3a5e73cd),
	.w8(32'hbc3df32d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaef243),
	.w1(32'hbc19a7f5),
	.w2(32'h3a030cd9),
	.w3(32'hba8da8fe),
	.w4(32'h3be5c2fe),
	.w5(32'h3a381938),
	.w6(32'hbc2e79c2),
	.w7(32'hbbb25b1c),
	.w8(32'hbb6032e7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae386f4),
	.w1(32'h3a9ee582),
	.w2(32'h3aa10355),
	.w3(32'hbb398f47),
	.w4(32'h3aa29481),
	.w5(32'hbb61b204),
	.w6(32'hbb726cab),
	.w7(32'hbb02acd8),
	.w8(32'hba2b825d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb604dbc),
	.w1(32'hbb8a5b2b),
	.w2(32'hbbef4f01),
	.w3(32'hbbbfe97a),
	.w4(32'hbbc0d898),
	.w5(32'h3c1e7702),
	.w6(32'hbb65fe5a),
	.w7(32'hbb8f8b0c),
	.w8(32'hb9a9dfaa),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b972863),
	.w1(32'h3b82ef3a),
	.w2(32'h3b89680a),
	.w3(32'h3b82fdee),
	.w4(32'hb83130a4),
	.w5(32'h3bca0c2b),
	.w6(32'hbbd9c13c),
	.w7(32'hbbb58c62),
	.w8(32'h3b38a793),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5c031),
	.w1(32'h3bed6817),
	.w2(32'h3c2978ff),
	.w3(32'h3bd7f2e5),
	.w4(32'h3be40527),
	.w5(32'hbba1342b),
	.w6(32'h3b8fda58),
	.w7(32'h3bfebf3a),
	.w8(32'hbc89be55),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc213e73),
	.w1(32'hbc8a75df),
	.w2(32'hbc028629),
	.w3(32'hbc18b999),
	.w4(32'hba939e97),
	.w5(32'h3b99f8b1),
	.w6(32'hbcee3d54),
	.w7(32'hbc4f2576),
	.w8(32'h3b5e0ed0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedb6f2),
	.w1(32'h3b4406a7),
	.w2(32'h3b394d0d),
	.w3(32'h3bac120d),
	.w4(32'h3a6e594f),
	.w5(32'hbbd86eb4),
	.w6(32'h3ad0b279),
	.w7(32'h3aa98e6e),
	.w8(32'hbbd8e194),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1d90b),
	.w1(32'h3b0c0ee1),
	.w2(32'hba747b47),
	.w3(32'h3a66d67c),
	.w4(32'hbadde44d),
	.w5(32'h3b7087b2),
	.w6(32'h3b7d76da),
	.w7(32'hba87bcee),
	.w8(32'h3c3c4c70),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef6ddf),
	.w1(32'h3a2f3295),
	.w2(32'h3b9d49ce),
	.w3(32'hb907b295),
	.w4(32'hbb064291),
	.w5(32'hbaab6767),
	.w6(32'h3c2b880b),
	.w7(32'h3c081221),
	.w8(32'h3b6dbd20),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b186488),
	.w1(32'h3ba12924),
	.w2(32'hbb309a81),
	.w3(32'h3aa86382),
	.w4(32'hba8d2676),
	.w5(32'hbba87140),
	.w6(32'h3c2a3796),
	.w7(32'hbaca733b),
	.w8(32'h3ba32998),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad717b),
	.w1(32'h3bd51593),
	.w2(32'h3c086053),
	.w3(32'hbbb330a4),
	.w4(32'hbbdb4aba),
	.w5(32'h392d79c3),
	.w6(32'h3b710dae),
	.w7(32'h3b4c074d),
	.w8(32'h3a934659),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd05e74),
	.w1(32'h3b20cf3d),
	.w2(32'h3b031933),
	.w3(32'hbada1b4c),
	.w4(32'hba45df18),
	.w5(32'h3b96272f),
	.w6(32'hbafe50a7),
	.w7(32'hba0a355a),
	.w8(32'h3b7ac323),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa246a0),
	.w1(32'h3b50c64c),
	.w2(32'h3aaf2ba3),
	.w3(32'h3c057ea7),
	.w4(32'hba449c02),
	.w5(32'hbb53ffc8),
	.w6(32'h3c1b5a3a),
	.w7(32'hbaa30264),
	.w8(32'hbb959287),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999b870),
	.w1(32'hbb519b89),
	.w2(32'h39d07df5),
	.w3(32'hbb08bcbe),
	.w4(32'hba053306),
	.w5(32'hbad4d01f),
	.w6(32'hbba6a00e),
	.w7(32'h3a5ff4c3),
	.w8(32'hbb05185f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbca6cd),
	.w1(32'hbbeec0bc),
	.w2(32'hbbd00b6f),
	.w3(32'hbbe77cdd),
	.w4(32'hbbe1a7c3),
	.w5(32'h3b429593),
	.w6(32'hbb63c89c),
	.w7(32'hbb41884d),
	.w8(32'h3a87c1ab),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f445e2),
	.w1(32'h3b0441f2),
	.w2(32'hb999f35d),
	.w3(32'h3a9a1be0),
	.w4(32'hbb653cc3),
	.w5(32'h3b5b0702),
	.w6(32'h3b36b313),
	.w7(32'hbb2b9c1a),
	.w8(32'h3c3b37d8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6da004),
	.w1(32'h3ba53be1),
	.w2(32'h3b946cbc),
	.w3(32'h397d32fe),
	.w4(32'h3bb654d9),
	.w5(32'h3b04be1b),
	.w6(32'h3bdcb567),
	.w7(32'h3b9bfb4e),
	.w8(32'h3b9acc57),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf75457),
	.w1(32'h3c32d546),
	.w2(32'h3c0ad2c4),
	.w3(32'h3bf40c80),
	.w4(32'h3ba9b867),
	.w5(32'h3b56dc0f),
	.w6(32'h3c4559de),
	.w7(32'h3b9f1255),
	.w8(32'hbb1fe370),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20f9ca),
	.w1(32'h3b825f29),
	.w2(32'h3b2509af),
	.w3(32'h3c027c66),
	.w4(32'h3b4aa217),
	.w5(32'h3b807bc1),
	.w6(32'h3a0052df),
	.w7(32'hbc09117a),
	.w8(32'h3bdcf95b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba44d6),
	.w1(32'h3c1a48ae),
	.w2(32'h3bb4f9c7),
	.w3(32'h3b8db131),
	.w4(32'h3b3f6b91),
	.w5(32'h37987ad6),
	.w6(32'h3c1518bc),
	.w7(32'h3b046fee),
	.w8(32'hba990f99),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab8a61),
	.w1(32'hbb4b689b),
	.w2(32'hbb7e7955),
	.w3(32'hbbe23a81),
	.w4(32'hbbfe62bc),
	.w5(32'hbb5fe1b7),
	.w6(32'hbb209237),
	.w7(32'hbc0018f5),
	.w8(32'hbbc618cf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc092c27),
	.w1(32'hbc275b0d),
	.w2(32'hbc6f086b),
	.w3(32'hbbcc384c),
	.w4(32'hbbc4728d),
	.w5(32'hbb9c3c72),
	.w6(32'hbbd4a7b6),
	.w7(32'hbc193524),
	.w8(32'h3a0f1261),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f4078),
	.w1(32'h3ab6a987),
	.w2(32'hbbdfb3d8),
	.w3(32'hbac9db4b),
	.w4(32'hbbd0e20e),
	.w5(32'h3ba09376),
	.w6(32'h3beb3357),
	.w7(32'hbb99c775),
	.w8(32'h3bcbbb1d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2512a6),
	.w1(32'h3c13090e),
	.w2(32'h3bb6e6fc),
	.w3(32'h3bdd906d),
	.w4(32'h3b82eed5),
	.w5(32'h3b59dade),
	.w6(32'h3c327e83),
	.w7(32'h3b494063),
	.w8(32'h3c0eaf7a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba59000),
	.w1(32'h3be708d5),
	.w2(32'h3b2d5d3d),
	.w3(32'h3ac7e5b6),
	.w4(32'hb9a53b90),
	.w5(32'h3b01ac8e),
	.w6(32'h3c039004),
	.w7(32'h3a3a8e12),
	.w8(32'h3b095ea2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96c301),
	.w1(32'h3b2258d9),
	.w2(32'h3b535dee),
	.w3(32'h3b2b2725),
	.w4(32'h3b4f15b3),
	.w5(32'hb94e6774),
	.w6(32'h3993d69c),
	.w7(32'h3b027c3c),
	.w8(32'hbb63995c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3a993),
	.w1(32'hbaaf7d14),
	.w2(32'hbb9e664e),
	.w3(32'hba471e19),
	.w4(32'hbb5f1e6b),
	.w5(32'hba102159),
	.w6(32'hbb3e6951),
	.w7(32'hbbf1494b),
	.w8(32'hbac94acf),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a54a9),
	.w1(32'hbb46346a),
	.w2(32'hbbb6db8d),
	.w3(32'hbaf656eb),
	.w4(32'hbbbef4d7),
	.w5(32'hbb558dad),
	.w6(32'hbb4dad64),
	.w7(32'hbbd8fe73),
	.w8(32'hba2582e7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00eaac),
	.w1(32'h3bcf224b),
	.w2(32'h3b688493),
	.w3(32'h3a77546d),
	.w4(32'h3bbc6fbb),
	.w5(32'hb9a28039),
	.w6(32'h3b7a4629),
	.w7(32'h3b899f97),
	.w8(32'hb9a6c9f5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e72b1e),
	.w1(32'h3b55a7b3),
	.w2(32'h3a2caace),
	.w3(32'h3b8d2eac),
	.w4(32'h39e01c2e),
	.w5(32'h3b6a0c51),
	.w6(32'h3c30704e),
	.w7(32'h3bb5987d),
	.w8(32'h3be2d1b7),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c103803),
	.w1(32'h3b8aa28f),
	.w2(32'hbaeedb46),
	.w3(32'h3b3965b0),
	.w4(32'hbb1d3ed8),
	.w5(32'h3a8919ce),
	.w6(32'h3c1611b2),
	.w7(32'h389b3cd8),
	.w8(32'hbaf4c4b9),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97de74),
	.w1(32'hbb3e05c5),
	.w2(32'hba9de1c7),
	.w3(32'hbae44561),
	.w4(32'h3ad477d5),
	.w5(32'h3b1f9ea1),
	.w6(32'hbb909f57),
	.w7(32'hbb024875),
	.w8(32'hbbd57e5e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc46bd8),
	.w1(32'h3b8fc4f3),
	.w2(32'h3bfc6ef2),
	.w3(32'hbb76ef14),
	.w4(32'h3ab49c95),
	.w5(32'hba400446),
	.w6(32'hbc3d9f86),
	.w7(32'hbbc2f7fe),
	.w8(32'hbad1798b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c91a4),
	.w1(32'hbaf40ed9),
	.w2(32'h3a53dedc),
	.w3(32'hb995fe43),
	.w4(32'hbb37b93c),
	.w5(32'hbb7c1f82),
	.w6(32'h3ada6d3a),
	.w7(32'hbb032e18),
	.w8(32'hba535722),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73618a),
	.w1(32'h37c13313),
	.w2(32'h3b5afc1e),
	.w3(32'h3adfa9de),
	.w4(32'h3b2b8350),
	.w5(32'hbb8697dd),
	.w6(32'h3ba61615),
	.w7(32'h3bb8c725),
	.w8(32'hbb8f1259),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb33ccc),
	.w1(32'hbb4b2bdf),
	.w2(32'hbacff653),
	.w3(32'hbb9ce5ac),
	.w4(32'hbb221e0c),
	.w5(32'hbbcb8a75),
	.w6(32'hbbb08481),
	.w7(32'hbb6a81f1),
	.w8(32'hbb872d68),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ba6f2),
	.w1(32'hbb3e5e5d),
	.w2(32'hba80654f),
	.w3(32'hbc070ea9),
	.w4(32'hbb853c4d),
	.w5(32'hbbe9fe68),
	.w6(32'hbb605496),
	.w7(32'hbb331c90),
	.w8(32'hbb9a8d0d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb43cb),
	.w1(32'h3b6c816b),
	.w2(32'hbb25f122),
	.w3(32'h3bda25dc),
	.w4(32'h3b08eab4),
	.w5(32'hbb0fc4a5),
	.w6(32'h3c48c5bf),
	.w7(32'hb9f04c85),
	.w8(32'hbb90f7f9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f24de),
	.w1(32'hbb953564),
	.w2(32'h37bb34ec),
	.w3(32'hbbe3e3ed),
	.w4(32'hba8c3d34),
	.w5(32'h3b4c2217),
	.w6(32'hbb96d556),
	.w7(32'hbb6c8c22),
	.w8(32'h3b44d128),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3db1b),
	.w1(32'h3bad49ff),
	.w2(32'h3b0cd5fa),
	.w3(32'h3c0ce219),
	.w4(32'h3bd618e7),
	.w5(32'hbb511756),
	.w6(32'h3c080dda),
	.w7(32'h3c0050dd),
	.w8(32'hbbafe108),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa247cb),
	.w1(32'hbb8188e0),
	.w2(32'hbbaa8ec5),
	.w3(32'h3a6ccdb1),
	.w4(32'hbaf40897),
	.w5(32'hbb2671e0),
	.w6(32'hb921be7d),
	.w7(32'hbbaca0dd),
	.w8(32'hbb3f54a0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe760bb),
	.w1(32'hbbbd56e6),
	.w2(32'hbc2dcbfc),
	.w3(32'hba98d227),
	.w4(32'hbb9de749),
	.w5(32'hbb92aae2),
	.w6(32'h39c02f5f),
	.w7(32'hbba2501f),
	.w8(32'hbbafd8e0),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44c75e),
	.w1(32'hbb15725e),
	.w2(32'hbb5450d7),
	.w3(32'hb924e100),
	.w4(32'hba9cd405),
	.w5(32'hbaa11513),
	.w6(32'hbb151b68),
	.w7(32'hbaae439c),
	.w8(32'hbb26bab4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb354f4e),
	.w1(32'h3ba9f10b),
	.w2(32'hbaaf8d74),
	.w3(32'h3bddc03f),
	.w4(32'hba955a93),
	.w5(32'hbb2b204e),
	.w6(32'h3c2aca86),
	.w7(32'hb9f2d918),
	.w8(32'hbb8781d2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a847705),
	.w1(32'h3b1317e2),
	.w2(32'h3bc7de43),
	.w3(32'hbb9e3c29),
	.w4(32'h39f02eaa),
	.w5(32'hbb557b57),
	.w6(32'hbc073d87),
	.w7(32'hbab3c922),
	.w8(32'h3b148eba),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3884a4d2),
	.w1(32'hba24a1ce),
	.w2(32'h3b1d1e55),
	.w3(32'hbbe7728e),
	.w4(32'hbad1b1c3),
	.w5(32'hbb21c36a),
	.w6(32'hbb676a15),
	.w7(32'h3b8ff79e),
	.w8(32'hbc42bb9b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a10c2),
	.w1(32'h3a30c991),
	.w2(32'h3bcf2a5b),
	.w3(32'hb974efff),
	.w4(32'h3b0f7b19),
	.w5(32'h3b671b2c),
	.w6(32'hbc26f871),
	.w7(32'h3a5e8e84),
	.w8(32'h3b09c20a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a835b45),
	.w1(32'hbb15875d),
	.w2(32'h3a834922),
	.w3(32'hbaebfb12),
	.w4(32'hba23f9e0),
	.w5(32'h3a6c7f78),
	.w6(32'hbb5a9c3f),
	.w7(32'hbadfa585),
	.w8(32'hbbdf857d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab9af1),
	.w1(32'hbb1b6edb),
	.w2(32'hbba4eff6),
	.w3(32'h3b65e4f4),
	.w4(32'hba82fbc2),
	.w5(32'hbb17d24d),
	.w6(32'hbb802863),
	.w7(32'hba1a5526),
	.w8(32'h3bbac54f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75bad1),
	.w1(32'hba3a94c6),
	.w2(32'h3bf17880),
	.w3(32'hbb7e84a9),
	.w4(32'h3c0e6d27),
	.w5(32'h3b69fbe6),
	.w6(32'h3bf16fb1),
	.w7(32'h3c298afa),
	.w8(32'hbc02103c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf88943),
	.w1(32'h3bb7a6a0),
	.w2(32'h3affc503),
	.w3(32'hbb0752b7),
	.w4(32'hbb507826),
	.w5(32'h3b8463c8),
	.w6(32'hbbed5443),
	.w7(32'hbbb3403b),
	.w8(32'h3c06d36c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c0d15),
	.w1(32'h3ab0b9b5),
	.w2(32'h3b86d26a),
	.w3(32'hba27ab6f),
	.w4(32'h3a107775),
	.w5(32'h3b21ec9e),
	.w6(32'h3be3857f),
	.w7(32'h3b449a25),
	.w8(32'h3ba88804),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d598a),
	.w1(32'hbae378e8),
	.w2(32'hbb7ab178),
	.w3(32'hbb91720d),
	.w4(32'h3a3852ef),
	.w5(32'hbb1a3ce8),
	.w6(32'h3b5641b2),
	.w7(32'hba13a72d),
	.w8(32'hbc1dc8bc),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7a6e7),
	.w1(32'h3b505228),
	.w2(32'hbaf99726),
	.w3(32'h3b78f4f2),
	.w4(32'h3b7fd881),
	.w5(32'hbaca57a8),
	.w6(32'h394e6261),
	.w7(32'hb820ffcc),
	.w8(32'hbb556238),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49acd8),
	.w1(32'h3b56a8cc),
	.w2(32'h3a8a5904),
	.w3(32'hba48b2bf),
	.w4(32'hbb60daaf),
	.w5(32'h3bdb09fb),
	.w6(32'hbbb544d9),
	.w7(32'hba5bacb8),
	.w8(32'h3bd87e2b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb364f6),
	.w1(32'h3b815f59),
	.w2(32'h3b31a6ae),
	.w3(32'h3c18a85d),
	.w4(32'h3b8c9ce9),
	.w5(32'h3a6a342e),
	.w6(32'h3c5c14b8),
	.w7(32'h3bb87a75),
	.w8(32'hbb42b0b2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb817228),
	.w1(32'hbba3f9cd),
	.w2(32'h3a231c95),
	.w3(32'hba1e5506),
	.w4(32'hbb67a2a9),
	.w5(32'h3b8232e0),
	.w6(32'hbbd17c3c),
	.w7(32'hbbfff803),
	.w8(32'h3ba793e3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b48d2),
	.w1(32'h3bb153e6),
	.w2(32'h3c18afa2),
	.w3(32'hbac7e241),
	.w4(32'h3bd6952e),
	.w5(32'h3b155e51),
	.w6(32'h3ac7e5f3),
	.w7(32'h3b11866b),
	.w8(32'h384e7737),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b000958),
	.w1(32'h3adce968),
	.w2(32'h3bcee6fb),
	.w3(32'h3acfdb2c),
	.w4(32'h3b927a85),
	.w5(32'h3be267a4),
	.w6(32'hbadc81b4),
	.w7(32'h3b9d2a50),
	.w8(32'h3c2260ff),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13fe7c),
	.w1(32'h3baebaec),
	.w2(32'h3b8fad1f),
	.w3(32'h3bc2552b),
	.w4(32'h39481b32),
	.w5(32'h3bf132f4),
	.w6(32'h3bc42408),
	.w7(32'h3b7d44bd),
	.w8(32'h3b428279),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b969497),
	.w1(32'h3b243b64),
	.w2(32'h3b7fb396),
	.w3(32'h3b8a5d46),
	.w4(32'h3b12924d),
	.w5(32'h3ab2d053),
	.w6(32'hbbddce74),
	.w7(32'hbb58c657),
	.w8(32'h3b944b21),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381b3f66),
	.w1(32'h3b554580),
	.w2(32'hbb8a337d),
	.w3(32'h3a6d99c3),
	.w4(32'hbb20e53f),
	.w5(32'hbbed163b),
	.w6(32'h3c06b824),
	.w7(32'h3ab28e5a),
	.w8(32'hbb960651),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099398),
	.w1(32'hbbba3983),
	.w2(32'hbba25f4a),
	.w3(32'hbbbff817),
	.w4(32'hbbbd562d),
	.w5(32'h393f295f),
	.w6(32'hbb25da6e),
	.w7(32'hbbcddb55),
	.w8(32'h3a140729),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba588d1f),
	.w1(32'hb94da259),
	.w2(32'hbaffa3a4),
	.w3(32'hba9882ab),
	.w4(32'hb98a1a97),
	.w5(32'hbb18cd7d),
	.w6(32'h3b4bafd2),
	.w7(32'h3aa49d98),
	.w8(32'hbb388d3a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89113d),
	.w1(32'hbaf8dabc),
	.w2(32'h381befc6),
	.w3(32'hba965019),
	.w4(32'h3b2c9622),
	.w5(32'h3b5884fd),
	.w6(32'hbc1fa561),
	.w7(32'hbbc07339),
	.w8(32'hbaf54184),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19fed3),
	.w1(32'hbab1b2ed),
	.w2(32'h3b438c19),
	.w3(32'hb8247059),
	.w4(32'h3b42bb0b),
	.w5(32'h3a1ebfbb),
	.w6(32'hbba6b009),
	.w7(32'hbb3cfc2f),
	.w8(32'hba2d39b6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f853dd),
	.w1(32'h3b9d8659),
	.w2(32'h3b00038e),
	.w3(32'h3a60ccda),
	.w4(32'hbad8b9db),
	.w5(32'h3af0df1f),
	.w6(32'hbb3e2a22),
	.w7(32'h38a44efe),
	.w8(32'hbbab6712),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa15bb9),
	.w1(32'h3ac2efda),
	.w2(32'hbbbf33cf),
	.w3(32'h39aab00a),
	.w4(32'hbb428db4),
	.w5(32'hba502a11),
	.w6(32'hbad69084),
	.w7(32'hbb75b6d0),
	.w8(32'h399c5d0f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ce2c51),
	.w1(32'hbafe8588),
	.w2(32'h3afb5611),
	.w3(32'h3b17e425),
	.w4(32'hba453cd4),
	.w5(32'hbb17ab60),
	.w6(32'h3b506eae),
	.w7(32'hbafa87a0),
	.w8(32'hba97c67a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae37889),
	.w1(32'hbb0360f3),
	.w2(32'h3a7f853a),
	.w3(32'hbb2df08d),
	.w4(32'hbba5b0c9),
	.w5(32'hbb4948d7),
	.w6(32'hbaef8435),
	.w7(32'hbade28b0),
	.w8(32'hba13b614),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb298e70),
	.w1(32'h3abcd256),
	.w2(32'hbb291bab),
	.w3(32'hba222e82),
	.w4(32'hbb3e0e06),
	.w5(32'hba9fc542),
	.w6(32'hbb0366ac),
	.w7(32'hbabc4797),
	.w8(32'hbbf2f178),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9900b6),
	.w1(32'hbb1addd6),
	.w2(32'hbb7eae14),
	.w3(32'hbb000716),
	.w4(32'hbb979b10),
	.w5(32'hba625f95),
	.w6(32'hbb578dbd),
	.w7(32'hba81c5a1),
	.w8(32'h3a826499),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b0929),
	.w1(32'hbafa7cad),
	.w2(32'hbb5f5bfb),
	.w3(32'hbb2c7a06),
	.w4(32'hbaee7563),
	.w5(32'hb92f85a2),
	.w6(32'h3bb8c07e),
	.w7(32'h3ab84517),
	.w8(32'hb9de1c19),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2903f4),
	.w1(32'hbc37a5a4),
	.w2(32'hbb27512d),
	.w3(32'hbc0d4cd8),
	.w4(32'hbc0f3c3f),
	.w5(32'h3807793c),
	.w6(32'hbbdbb754),
	.w7(32'hbab0b9ae),
	.w8(32'h39a6d6bb),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf85ccf),
	.w1(32'hbb1895b8),
	.w2(32'hbbcfab2a),
	.w3(32'hba4ebc55),
	.w4(32'hba7a8a1d),
	.w5(32'h3b69b197),
	.w6(32'h3aaf5922),
	.w7(32'hbb4cbbde),
	.w8(32'h3b859fe1),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5be6a),
	.w1(32'h3b5567a3),
	.w2(32'hbae5e1a1),
	.w3(32'h3bf37ddf),
	.w4(32'h3a3f0d02),
	.w5(32'h3bc694da),
	.w6(32'h3c363bb6),
	.w7(32'h3b6126e7),
	.w8(32'hbb0087c0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79d33f),
	.w1(32'hbacd602b),
	.w2(32'h3b3238a4),
	.w3(32'h3b9b9d5d),
	.w4(32'h3b9c00f1),
	.w5(32'hbb329a35),
	.w6(32'hbb6c8742),
	.w7(32'h3a30dd81),
	.w8(32'hbb5f096e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae08def),
	.w1(32'h3a899578),
	.w2(32'hba8058f8),
	.w3(32'h3b59abdb),
	.w4(32'h3ab1474d),
	.w5(32'hbacb48ab),
	.w6(32'hbb31c1b6),
	.w7(32'h3aec9773),
	.w8(32'hbb1848ba),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e23cb),
	.w1(32'hbae393fe),
	.w2(32'hbb06ca1e),
	.w3(32'h3be9237e),
	.w4(32'hbb29024f),
	.w5(32'hba8eccf1),
	.w6(32'h3b0b1a0e),
	.w7(32'hbae32b67),
	.w8(32'hba56ced0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a928b91),
	.w1(32'h3ab99b50),
	.w2(32'h3b893253),
	.w3(32'hbb0648fe),
	.w4(32'hbac85644),
	.w5(32'hbb9b2131),
	.w6(32'h3a4e2a42),
	.w7(32'h3a6f09de),
	.w8(32'hbb94b7a6),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f8339),
	.w1(32'h3a430af6),
	.w2(32'hbaafea75),
	.w3(32'hba4ddf1a),
	.w4(32'h3abd6789),
	.w5(32'h3aae1b2a),
	.w6(32'h3afb68e4),
	.w7(32'h3a934c5e),
	.w8(32'h3ca14e5e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f1f2b),
	.w1(32'h3c6bde1a),
	.w2(32'h3b97a217),
	.w3(32'h3b6f27ab),
	.w4(32'h3a3674bf),
	.w5(32'hbbacc8d4),
	.w6(32'h3c95fe19),
	.w7(32'h3baebbe9),
	.w8(32'hbbf43ab6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7a100),
	.w1(32'hb9f493dd),
	.w2(32'hbb25fb68),
	.w3(32'h3b0985e3),
	.w4(32'h38f4cef8),
	.w5(32'h3bc5ea03),
	.w6(32'hb9e048ca),
	.w7(32'hbb1e8f23),
	.w8(32'h3c0d5a88),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c4eea),
	.w1(32'h3a86e2e2),
	.w2(32'h3b3718fe),
	.w3(32'hba9a6590),
	.w4(32'h3b86d23b),
	.w5(32'hbbb97ed4),
	.w6(32'h3b9be58d),
	.w7(32'h3b0e8b4b),
	.w8(32'hbc005957),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeef8d1),
	.w1(32'hbb381cd8),
	.w2(32'h3ac13f80),
	.w3(32'hbbc95862),
	.w4(32'hbb9b31db),
	.w5(32'h38bf3266),
	.w6(32'hbbfd61d3),
	.w7(32'hbb75afea),
	.w8(32'h3915d128),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a3c01),
	.w1(32'h3a2030f0),
	.w2(32'hb8200067),
	.w3(32'hbb586d5d),
	.w4(32'h3a5dd54a),
	.w5(32'hbb39b734),
	.w6(32'h3b0aebd3),
	.w7(32'h3b2187a5),
	.w8(32'h3b1972c0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3647b0),
	.w1(32'hbbdcfd4f),
	.w2(32'hbb8fd437),
	.w3(32'hbbc8893a),
	.w4(32'hbb07da4d),
	.w5(32'h37d04937),
	.w6(32'h3af8e28f),
	.w7(32'h3b42b657),
	.w8(32'hbaeee06b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb871869),
	.w1(32'hbb738971),
	.w2(32'hbb20eb98),
	.w3(32'hbb032e68),
	.w4(32'hbad2ba86),
	.w5(32'hbb889902),
	.w6(32'hbae1993e),
	.w7(32'hba8b10b8),
	.w8(32'h3b5d6f74),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32b9fa),
	.w1(32'h3bd67dea),
	.w2(32'h3b485875),
	.w3(32'h39a73f94),
	.w4(32'hbac68990),
	.w5(32'hba4ac537),
	.w6(32'h3c415633),
	.w7(32'h3bc5ca0e),
	.w8(32'hbb4cc6d7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b4e0e),
	.w1(32'hbb372ed4),
	.w2(32'hbafaecd4),
	.w3(32'hbb2dd338),
	.w4(32'hba98bd6f),
	.w5(32'hbbad7dfe),
	.w6(32'hbbe93d63),
	.w7(32'hbbf08caf),
	.w8(32'hbc158f97),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e056d),
	.w1(32'h3a6c4393),
	.w2(32'hba97f5a4),
	.w3(32'hbb89e403),
	.w4(32'hbbb0c756),
	.w5(32'h3a72afe2),
	.w6(32'hbb12a005),
	.w7(32'hbb837b3f),
	.w8(32'h3b06b211),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ea002),
	.w1(32'h3b9b54fd),
	.w2(32'h3b95d189),
	.w3(32'h3a14c21f),
	.w4(32'h3b485454),
	.w5(32'h3ba28907),
	.w6(32'h3a23448b),
	.w7(32'h3aa9006b),
	.w8(32'h3b529130),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b2f4a),
	.w1(32'h3b899cdc),
	.w2(32'h3b372280),
	.w3(32'h3b698809),
	.w4(32'h3b80b0a5),
	.w5(32'hb99fb291),
	.w6(32'h3b000a32),
	.w7(32'h3ae416c1),
	.w8(32'h3a93f14c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b6c5e),
	.w1(32'h3b5a6804),
	.w2(32'hbb68f579),
	.w3(32'h3b6f7ec4),
	.w4(32'hba111eb6),
	.w5(32'hbb95b1f7),
	.w6(32'h3bf67086),
	.w7(32'hbb26bf3a),
	.w8(32'hbc00153c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01544f),
	.w1(32'hbb50f184),
	.w2(32'hbb0ba6df),
	.w3(32'hbb40fcd7),
	.w4(32'hbb9f3676),
	.w5(32'hbad02e2f),
	.w6(32'hbb860a68),
	.w7(32'hbb6d84b1),
	.w8(32'hbb2d1184),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dcc88),
	.w1(32'hbaa71177),
	.w2(32'h3a202c54),
	.w3(32'hbb78dad3),
	.w4(32'hba5396e1),
	.w5(32'hbb058635),
	.w6(32'hbb784a63),
	.w7(32'hbb60085e),
	.w8(32'hbb362a4e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa02c7d),
	.w1(32'h3ab9498c),
	.w2(32'hbb125c56),
	.w3(32'hbb1a99e6),
	.w4(32'h3a26e1a1),
	.w5(32'hbbb22e89),
	.w6(32'hbb1a32bc),
	.w7(32'hbb11a657),
	.w8(32'h3c0b6245),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2713b),
	.w1(32'h3c9b397d),
	.w2(32'h3c1b5f4e),
	.w3(32'h3c240ce1),
	.w4(32'h3a2cd57b),
	.w5(32'hbb9627ec),
	.w6(32'h3cfd651b),
	.w7(32'h3c356c20),
	.w8(32'hbb8e9b8d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38c730),
	.w1(32'h39926129),
	.w2(32'h3b9cc74a),
	.w3(32'hbbda4db8),
	.w4(32'hbab3762b),
	.w5(32'hba131f22),
	.w6(32'hbb7204fe),
	.w7(32'hbb0f61cf),
	.w8(32'h3ac6ae69),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a926197),
	.w1(32'hbbaceeb7),
	.w2(32'h3b0db704),
	.w3(32'hbb1ce427),
	.w4(32'hb98ceb25),
	.w5(32'h3c06f23c),
	.w6(32'hbb291645),
	.w7(32'h39eab639),
	.w8(32'h3b9e8ce5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf29b21),
	.w1(32'h3b959d67),
	.w2(32'hbb4a7287),
	.w3(32'h3bb3ae5b),
	.w4(32'h3b5af394),
	.w5(32'h3b30e66c),
	.w6(32'h3bc87456),
	.w7(32'h3ab240c6),
	.w8(32'hbb17ae9c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ef953),
	.w1(32'hb9f369f7),
	.w2(32'h39c51c9b),
	.w3(32'h3a9ddbf3),
	.w4(32'h3b28a67f),
	.w5(32'hbb152bca),
	.w6(32'hbadd6591),
	.w7(32'hb9e43753),
	.w8(32'hbb2199e4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddd37a),
	.w1(32'hbb789753),
	.w2(32'hbc1cc338),
	.w3(32'hbb41a297),
	.w4(32'hbbe15393),
	.w5(32'h3b134ec4),
	.w6(32'hb9a9add7),
	.w7(32'hbc12241a),
	.w8(32'h3b3c0056),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58c900),
	.w1(32'h3bcaabff),
	.w2(32'hbb23b385),
	.w3(32'h3bc7dfde),
	.w4(32'hbb204210),
	.w5(32'hba10fa2d),
	.w6(32'h3bcf3357),
	.w7(32'hbafd32b1),
	.w8(32'h3aa1ad1e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b0bb2),
	.w1(32'h3c2690c0),
	.w2(32'h3c31f205),
	.w3(32'h3bf96477),
	.w4(32'h3b774904),
	.w5(32'h3be7d697),
	.w6(32'h3c6b67ed),
	.w7(32'h3ba39681),
	.w8(32'h3b8a1c34),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe86b5),
	.w1(32'h3b1c5bed),
	.w2(32'h3b8d1137),
	.w3(32'h3b71a477),
	.w4(32'h3a3b3d4c),
	.w5(32'hba9a36fd),
	.w6(32'h39a1b14d),
	.w7(32'h38e1710c),
	.w8(32'hbac430af),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaac5ab),
	.w1(32'hba9f01f7),
	.w2(32'hba84263f),
	.w3(32'h3b576df0),
	.w4(32'h3a68b936),
	.w5(32'h3b15e64a),
	.w6(32'h3abff7af),
	.w7(32'h3afdffde),
	.w8(32'hba68b4cd),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a461668),
	.w1(32'h3b71b036),
	.w2(32'h3bad6f33),
	.w3(32'h3bba41e7),
	.w4(32'h3b8d8ea1),
	.w5(32'h3b23be9f),
	.w6(32'h3b8b10a5),
	.w7(32'h3ba80834),
	.w8(32'h3b2c0914),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b138d),
	.w1(32'h3b93e8a0),
	.w2(32'h3b659507),
	.w3(32'h3badd7e1),
	.w4(32'h3b6b9643),
	.w5(32'h3b909aab),
	.w6(32'h3c2fd471),
	.w7(32'h3c20e2b2),
	.w8(32'h3b9de06e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58bc56),
	.w1(32'hbbebc255),
	.w2(32'hba1d75a1),
	.w3(32'h3af4a99f),
	.w4(32'h3bdedc1d),
	.w5(32'h3bcb6c1e),
	.w6(32'h3b0e365d),
	.w7(32'h3bde14a8),
	.w8(32'h3b9d9225),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f3dde),
	.w1(32'h3c0a6d4b),
	.w2(32'h3c0c56a2),
	.w3(32'h3bc73e84),
	.w4(32'h3bfda002),
	.w5(32'h3b1ef1fb),
	.w6(32'h3b30fee1),
	.w7(32'h3ba91c76),
	.w8(32'hbb8929f0),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac43635),
	.w1(32'h3a49343c),
	.w2(32'hb958185d),
	.w3(32'h3bc2f6a2),
	.w4(32'h3b8c5c14),
	.w5(32'h399bcbb5),
	.w6(32'hbb745953),
	.w7(32'h3adffbaf),
	.w8(32'h3af9de73),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a1fd0c),
	.w1(32'h3ba03296),
	.w2(32'h38b8abb6),
	.w3(32'h3baf8ffe),
	.w4(32'h3a804c7a),
	.w5(32'hbb762690),
	.w6(32'h3bacf41a),
	.w7(32'h3a97d8f1),
	.w8(32'h3b01a655),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80ce6c),
	.w1(32'h3b1f8496),
	.w2(32'hbb069fea),
	.w3(32'h3b558f6b),
	.w4(32'hbc136acd),
	.w5(32'hbc13bdec),
	.w6(32'h3b872120),
	.w7(32'hbaa3c242),
	.w8(32'hbbd95cce),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef0b21),
	.w1(32'hbaec953c),
	.w2(32'hbbe29fff),
	.w3(32'hbbb0f6ae),
	.w4(32'hbbab2c39),
	.w5(32'h3b04dc93),
	.w6(32'h3a9a010c),
	.w7(32'h3ad8d1ab),
	.w8(32'h3aef5b3d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c9815),
	.w1(32'hbaa48f51),
	.w2(32'hbb80863d),
	.w3(32'h36acf9fb),
	.w4(32'hbb9c8c95),
	.w5(32'h397faa61),
	.w6(32'hbabeb004),
	.w7(32'hbb7555ef),
	.w8(32'h38b2ea0d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c3bc1),
	.w1(32'hbb007578),
	.w2(32'h3ae83819),
	.w3(32'hbb2b9ccd),
	.w4(32'hbafbfc75),
	.w5(32'h39c44a66),
	.w6(32'hbb9ee481),
	.w7(32'h3b2198d9),
	.w8(32'h3bc062bb),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb07ae),
	.w1(32'hbb22173b),
	.w2(32'hbb728b2e),
	.w3(32'hbab7df76),
	.w4(32'hbba95108),
	.w5(32'h3c2aac5c),
	.w6(32'h3b995c20),
	.w7(32'hbb22aa20),
	.w8(32'hbbfa9aa9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d569c),
	.w1(32'hbbdcb67f),
	.w2(32'hba2c5c06),
	.w3(32'h3c04b211),
	.w4(32'h3c007300),
	.w5(32'hbb232dcf),
	.w6(32'hbb284676),
	.w7(32'hbbe08b63),
	.w8(32'h3a27bb5f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb83b12),
	.w1(32'hbaf94f99),
	.w2(32'h3a0554fa),
	.w3(32'h3b09fd8b),
	.w4(32'h39bf8d24),
	.w5(32'h3abe6de3),
	.w6(32'h3b352f6b),
	.w7(32'h3b589139),
	.w8(32'hbb9fff20),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e98ed),
	.w1(32'hbc0de345),
	.w2(32'hba06755d),
	.w3(32'hb853ed76),
	.w4(32'hbc006d08),
	.w5(32'hbb7f47ba),
	.w6(32'hbbd313e6),
	.w7(32'hbc2b6cb2),
	.w8(32'hbb8f85f2),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58a3f7),
	.w1(32'h3aac512b),
	.w2(32'h39a27120),
	.w3(32'hba25aeb4),
	.w4(32'h39d35dc9),
	.w5(32'h3bfb37b1),
	.w6(32'hba973344),
	.w7(32'h3abbb593),
	.w8(32'h3c10aaea),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b718151),
	.w1(32'h3c192f67),
	.w2(32'hbaf1eb7b),
	.w3(32'h3c63e957),
	.w4(32'h3b2d50e1),
	.w5(32'hbaa7aa18),
	.w6(32'h3c56fe2d),
	.w7(32'h3a888710),
	.w8(32'h3a8a4f90),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66b81e),
	.w1(32'h3c260ca2),
	.w2(32'h3c095f65),
	.w3(32'h3c173458),
	.w4(32'h3c0ddd72),
	.w5(32'h3b172ac2),
	.w6(32'h3c297655),
	.w7(32'h3c45b9ae),
	.w8(32'hba1a3e21),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baad4d2),
	.w1(32'hbb09a47b),
	.w2(32'h3ad2651c),
	.w3(32'hbb7d7572),
	.w4(32'hb9c58a28),
	.w5(32'hbaf5b949),
	.w6(32'hbb354a83),
	.w7(32'h3b0417d1),
	.w8(32'hbb7d237c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58c650),
	.w1(32'hbb7157a1),
	.w2(32'h3b10a158),
	.w3(32'hbbb4a68f),
	.w4(32'hbb64b607),
	.w5(32'h3b6ee600),
	.w6(32'hbbf82c10),
	.w7(32'hbb382f5b),
	.w8(32'h3abc29c9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b424316),
	.w1(32'h39297428),
	.w2(32'h3bd1c2ec),
	.w3(32'hbb077e0f),
	.w4(32'h3b7a592f),
	.w5(32'hb992a024),
	.w6(32'hbbb5d3d0),
	.w7(32'h3a4342c1),
	.w8(32'hb95dda5c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31eb7b),
	.w1(32'h3b0e3a83),
	.w2(32'hba5154c2),
	.w3(32'hba275740),
	.w4(32'hbb7f2f2e),
	.w5(32'hbb02bf73),
	.w6(32'h3a760966),
	.w7(32'hbab2ca05),
	.w8(32'hbb34ad6f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa74c8c),
	.w1(32'hbc1e9e92),
	.w2(32'hbbc0f82e),
	.w3(32'hbb79777d),
	.w4(32'hbb43c293),
	.w5(32'h3ab8a04c),
	.w6(32'hbbbf1e5d),
	.w7(32'hbb215c0c),
	.w8(32'h3a42fd77),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b877949),
	.w1(32'hbb73829d),
	.w2(32'hbb34db66),
	.w3(32'hbb25483a),
	.w4(32'hbb09cc25),
	.w5(32'hb98b2ace),
	.w6(32'hbb8bddde),
	.w7(32'hbb67b008),
	.w8(32'h3959eac2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d1928),
	.w1(32'h3aff468a),
	.w2(32'h3adc8a3f),
	.w3(32'hbaf52cad),
	.w4(32'hbad82d85),
	.w5(32'h3b27c7e2),
	.w6(32'hbb01d914),
	.w7(32'hba9cd681),
	.w8(32'h3b9a19df),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb552e84),
	.w1(32'hba473ff3),
	.w2(32'hbb5fcd00),
	.w3(32'hbaa68ddb),
	.w4(32'hb8fb6ba1),
	.w5(32'h3bcb4663),
	.w6(32'h3a572eb7),
	.w7(32'hbaf6dc42),
	.w8(32'h3c175ffb),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8dad10),
	.w1(32'h3cc3c9ce),
	.w2(32'hbc16132d),
	.w3(32'h3cd48390),
	.w4(32'hbb9fdd33),
	.w5(32'h3b2d0e26),
	.w6(32'h3cf92e73),
	.w7(32'h3c502945),
	.w8(32'h3b022dab),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992ea57),
	.w1(32'hba395f22),
	.w2(32'hbc72c59d),
	.w3(32'h3c0ebba3),
	.w4(32'hbb5e6796),
	.w5(32'h39c3aae8),
	.w6(32'h3bb4e152),
	.w7(32'hbc48134e),
	.w8(32'hba81d53d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5146c1),
	.w1(32'hba34d88b),
	.w2(32'hbaa677de),
	.w3(32'hbaadb224),
	.w4(32'hbb2abbbc),
	.w5(32'hb9dde0de),
	.w6(32'hbb8b781d),
	.w7(32'hbb49cd33),
	.w8(32'hbb368f6a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b91bc),
	.w1(32'hbb81bf42),
	.w2(32'h3b454c66),
	.w3(32'hbaafc65b),
	.w4(32'h3b03b5fc),
	.w5(32'h3ab84ee2),
	.w6(32'hbbbf750d),
	.w7(32'h3a8b01a0),
	.w8(32'h38a9ccb0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d351e),
	.w1(32'h3ad89577),
	.w2(32'hbb516ad9),
	.w3(32'h38f68038),
	.w4(32'hbb6fec29),
	.w5(32'hbb79cff6),
	.w6(32'hb96b4d1d),
	.w7(32'hbb596b04),
	.w8(32'hbb4ce881),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39dafc),
	.w1(32'hbbbe729d),
	.w2(32'hbb0252f4),
	.w3(32'hbbf04dec),
	.w4(32'hbb3285dd),
	.w5(32'hbb01fa68),
	.w6(32'hbbd14995),
	.w7(32'hbb48972d),
	.w8(32'h3ab571ef),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0655ad),
	.w1(32'hba7c6aa2),
	.w2(32'hbb66fb74),
	.w3(32'hbac7a46f),
	.w4(32'hbb0e3961),
	.w5(32'h3aea3eb5),
	.w6(32'hbb4c7abd),
	.w7(32'hbb31486d),
	.w8(32'hb8567717),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64cd91),
	.w1(32'h3acaa96f),
	.w2(32'h3b01b3cf),
	.w3(32'h3b183d5e),
	.w4(32'h3b3fb2fe),
	.w5(32'h3b8fe6e5),
	.w6(32'h3b569a42),
	.w7(32'h3b4100a7),
	.w8(32'h39bcba3d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9912b18),
	.w1(32'hbb73afa8),
	.w2(32'hbb3786b0),
	.w3(32'hbb6c9c28),
	.w4(32'h3b4db4ed),
	.w5(32'hbbc3292d),
	.w6(32'hbbe7f96f),
	.w7(32'hbb4d8f28),
	.w8(32'h3ac1f605),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f173f),
	.w1(32'h3b4904a8),
	.w2(32'hbbb6df32),
	.w3(32'h3b873cbb),
	.w4(32'hbbe4816c),
	.w5(32'hba868306),
	.w6(32'h3ba91760),
	.w7(32'hbb988ac7),
	.w8(32'hbb1cbe19),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule