module layer_10_featuremap_113(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bf61e1),
	.w1(32'h3b4e487c),
	.w2(32'h3bad92a2),
	.w3(32'h3905358a),
	.w4(32'hba6077cc),
	.w5(32'h3b3c495d),
	.w6(32'h3b1da2e5),
	.w7(32'h3baa3235),
	.w8(32'h3b153374),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab37ee),
	.w1(32'h3a2ca996),
	.w2(32'h39c52413),
	.w3(32'h3ad33117),
	.w4(32'h3abd2bb1),
	.w5(32'h3a74ea62),
	.w6(32'hb70e6901),
	.w7(32'h39abd79d),
	.w8(32'hba6305d4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3856f7b3),
	.w1(32'hba92b207),
	.w2(32'hbac950ae),
	.w3(32'h39b73769),
	.w4(32'hb9e0f1e7),
	.w5(32'hbac5e9b8),
	.w6(32'h3b0ab1bf),
	.w7(32'h3b230e65),
	.w8(32'h3b46c46b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4924e),
	.w1(32'hbb36b232),
	.w2(32'h3a22c8cc),
	.w3(32'hbae72215),
	.w4(32'hbaa8a1d0),
	.w5(32'h3a600742),
	.w6(32'h3b3ea32e),
	.w7(32'h3b09cedf),
	.w8(32'h3b1c5d42),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a4261),
	.w1(32'h3a614d8e),
	.w2(32'h3b1c2b65),
	.w3(32'h39264612),
	.w4(32'hba495927),
	.w5(32'h3ae2fbb5),
	.w6(32'h3a9b6bb6),
	.w7(32'h3ac7de83),
	.w8(32'h3b45e1d8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b407533),
	.w1(32'hbb310b8a),
	.w2(32'hbabea82b),
	.w3(32'h3b057441),
	.w4(32'hbad5a124),
	.w5(32'hbab61bfa),
	.w6(32'hba9e2f8c),
	.w7(32'hbae4af4e),
	.w8(32'hbad8ab42),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a153f),
	.w1(32'hb9f78ebf),
	.w2(32'hb9f6deb0),
	.w3(32'hbab5a443),
	.w4(32'hb996f69f),
	.w5(32'hba020f3e),
	.w6(32'hb8892901),
	.w7(32'hb84936e2),
	.w8(32'hba712ed1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99026af),
	.w1(32'hba95a248),
	.w2(32'hba5caa26),
	.w3(32'hb9184d99),
	.w4(32'hba579c0a),
	.w5(32'hba9cdcec),
	.w6(32'h3a26b829),
	.w7(32'h39b59e0e),
	.w8(32'h3981ea47),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba676f00),
	.w1(32'h3a41fb54),
	.w2(32'hbab69587),
	.w3(32'hba699495),
	.w4(32'hb8bf918b),
	.w5(32'hbaeaa49e),
	.w6(32'h3ae1a332),
	.w7(32'hba768e25),
	.w8(32'h38e57274),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c5958),
	.w1(32'h3aa1a444),
	.w2(32'hb9cf4118),
	.w3(32'hba38b586),
	.w4(32'h3b61c359),
	.w5(32'h3ab12ebc),
	.w6(32'h3a648600),
	.w7(32'hb981a135),
	.w8(32'hba29e670),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f34f82),
	.w1(32'hbb5007a8),
	.w2(32'hbaabe82f),
	.w3(32'h3a489106),
	.w4(32'hbb3cf683),
	.w5(32'hbb1dbd31),
	.w6(32'h3c01dac3),
	.w7(32'h3c17e623),
	.w8(32'h3c15e2f4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5024ce),
	.w1(32'h3a46d990),
	.w2(32'h39f280a4),
	.w3(32'hbb382fad),
	.w4(32'h3aa0b5ef),
	.w5(32'hb96a1097),
	.w6(32'hbb0da076),
	.w7(32'hba888a0f),
	.w8(32'hbb31edb2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f2fa),
	.w1(32'hba705e45),
	.w2(32'h3954a51d),
	.w3(32'hbb22c342),
	.w4(32'h39048f12),
	.w5(32'h3a9fc285),
	.w6(32'hba0e9f19),
	.w7(32'hba044e43),
	.w8(32'hba2bba80),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edf0cf),
	.w1(32'hb92e87a7),
	.w2(32'h39e788c0),
	.w3(32'h3aad721d),
	.w4(32'hb9e4fa27),
	.w5(32'hba2a8b5c),
	.w6(32'h3a64903b),
	.w7(32'h3b0067fc),
	.w8(32'h3a1b6d55),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c689e7),
	.w1(32'hba55f667),
	.w2(32'h39eb22c2),
	.w3(32'hba8c0775),
	.w4(32'h3ab0465d),
	.w5(32'hb93e74ca),
	.w6(32'hba9fcc94),
	.w7(32'hba1b821c),
	.w8(32'hb95d02f7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb76b9),
	.w1(32'h38c11dff),
	.w2(32'hba1c88a0),
	.w3(32'h39cc24e2),
	.w4(32'hb9c1e586),
	.w5(32'hb9fe7d24),
	.w6(32'h398f6103),
	.w7(32'hba7d75af),
	.w8(32'hbaaa2135),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fc7d4),
	.w1(32'h3bd6adc2),
	.w2(32'h3bb17373),
	.w3(32'hbaa310f9),
	.w4(32'h3a15bfff),
	.w5(32'hbbd575ca),
	.w6(32'h3bd4b09f),
	.w7(32'h3b64f84b),
	.w8(32'h3b51f383),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcd3ec),
	.w1(32'h3a99b0c6),
	.w2(32'h3a58ef70),
	.w3(32'hbb6ca088),
	.w4(32'h3ae66260),
	.w5(32'h3ab1be26),
	.w6(32'h3a11eaf7),
	.w7(32'h3a49e6ba),
	.w8(32'h3a64cdf7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c836e),
	.w1(32'hb9d89bf8),
	.w2(32'hbab6d10b),
	.w3(32'h3accfe3d),
	.w4(32'h39284b42),
	.w5(32'hba9706fa),
	.w6(32'hb971b306),
	.w7(32'hb889b483),
	.w8(32'h385bf1a3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca32d3),
	.w1(32'h3a033870),
	.w2(32'hbab9fbea),
	.w3(32'hb935de30),
	.w4(32'h3a228da4),
	.w5(32'hbaa03698),
	.w6(32'h3a289c96),
	.w7(32'hba7b8e09),
	.w8(32'hb99dfcf2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b64018),
	.w1(32'h39502d9e),
	.w2(32'h3b34c43e),
	.w3(32'hba165b5f),
	.w4(32'hba40f224),
	.w5(32'h3a0fca7d),
	.w6(32'h3b63ffe7),
	.w7(32'h3b1d34b7),
	.w8(32'h3990e69b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9c904),
	.w1(32'hbad1b6b3),
	.w2(32'hba9353c7),
	.w3(32'hb84a8f73),
	.w4(32'hba793fb8),
	.w5(32'h3a53b019),
	.w6(32'hba862343),
	.w7(32'h3b325cb0),
	.w8(32'h38c7a764),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ad63b),
	.w1(32'hba82f38a),
	.w2(32'h38149f5b),
	.w3(32'h3a60f082),
	.w4(32'hbaade432),
	.w5(32'hba9c3ba8),
	.w6(32'h3bc5f9bc),
	.w7(32'h3c0b329d),
	.w8(32'h3bbd0cdc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb516ccc),
	.w1(32'hba99efe4),
	.w2(32'hba801d1e),
	.w3(32'hbb493a9e),
	.w4(32'hbaaf9489),
	.w5(32'hbab56d97),
	.w6(32'h39b4e6f2),
	.w7(32'h39ad915c),
	.w8(32'h38257496),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba573cf2),
	.w1(32'h3abc14fa),
	.w2(32'hb7a0baaf),
	.w3(32'hbaa2e238),
	.w4(32'h3b2b82ed),
	.w5(32'h3a02c832),
	.w6(32'h3bd4d4d7),
	.w7(32'h3b8dd669),
	.w8(32'h3b151e72),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99e808),
	.w1(32'h3ac76a72),
	.w2(32'h3b3d802a),
	.w3(32'hbab57fad),
	.w4(32'h3baaa605),
	.w5(32'h3b6d11f4),
	.w6(32'h38f8f530),
	.w7(32'hbaf5cc9a),
	.w8(32'h398b0cd7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a401c4d),
	.w1(32'hb9da08ae),
	.w2(32'hb910d807),
	.w3(32'h3a9d5089),
	.w4(32'hb8946a62),
	.w5(32'h39ad7aa8),
	.w6(32'hb89c5f2c),
	.w7(32'h39390836),
	.w8(32'hba05b6ad),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba256090),
	.w1(32'h3a87ce43),
	.w2(32'hb97d5d59),
	.w3(32'hb9f66bef),
	.w4(32'h3b230e19),
	.w5(32'h3ac0dfe1),
	.w6(32'h3b8bebaf),
	.w7(32'h3b250b1e),
	.w8(32'h3affcd32),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3950fee7),
	.w1(32'h3bf3858b),
	.w2(32'h3b5a2fbf),
	.w3(32'h3abce817),
	.w4(32'h3b9ebc35),
	.w5(32'hbb7f68da),
	.w6(32'h3caa214c),
	.w7(32'h3c914eff),
	.w8(32'h3c82e988),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f3f7b),
	.w1(32'h3c4e99e9),
	.w2(32'h3c192472),
	.w3(32'hba57a2e3),
	.w4(32'h3bfa4774),
	.w5(32'h3b2699b7),
	.w6(32'h3c817d20),
	.w7(32'h3c2f6b05),
	.w8(32'h3badba0c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7a873),
	.w1(32'hba89e8e5),
	.w2(32'h3a20eb44),
	.w3(32'h37ac880d),
	.w4(32'hba80d584),
	.w5(32'hb8ea11c0),
	.w6(32'h3ad19702),
	.w7(32'h3af01114),
	.w8(32'h3a7433b3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac4025),
	.w1(32'hba921325),
	.w2(32'h39e9a677),
	.w3(32'hb97bcf79),
	.w4(32'hba122fa7),
	.w5(32'h3a8d5421),
	.w6(32'h397fbd41),
	.w7(32'hb839fb38),
	.w8(32'hb9ee10df),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba366351),
	.w1(32'hb981c0b9),
	.w2(32'hbb544885),
	.w3(32'h398e424d),
	.w4(32'hb9897ae5),
	.w5(32'hbaaaa88d),
	.w6(32'hba3127e8),
	.w7(32'hba9d260c),
	.w8(32'h3adf98aa),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3801b06c),
	.w1(32'hba2401a4),
	.w2(32'h3b161e91),
	.w3(32'hbaa821b2),
	.w4(32'hbac9d43e),
	.w5(32'h3a6e4c4e),
	.w6(32'hb8a3030f),
	.w7(32'hbb0a80b6),
	.w8(32'h39804667),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22a746),
	.w1(32'hbaaeba7d),
	.w2(32'hbb4ebce8),
	.w3(32'h3ac89111),
	.w4(32'h3ab17009),
	.w5(32'hba1c83cd),
	.w6(32'h3936620a),
	.w7(32'hba22860e),
	.w8(32'hba51abb0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafeceb8),
	.w1(32'hba847281),
	.w2(32'h3ad790e0),
	.w3(32'h395fc68b),
	.w4(32'hba0a5944),
	.w5(32'h3a248ce6),
	.w6(32'h3ac1210a),
	.w7(32'h3b114b18),
	.w8(32'h3a249ded),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2f4e1),
	.w1(32'h399c5401),
	.w2(32'h39040848),
	.w3(32'hba364ecd),
	.w4(32'h3afa1b74),
	.w5(32'h3a2fbe67),
	.w6(32'h38ecfc93),
	.w7(32'hba1b59fd),
	.w8(32'hbac6ab49),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e2234),
	.w1(32'h39515ec0),
	.w2(32'h38892263),
	.w3(32'h3915fc8d),
	.w4(32'h3a355303),
	.w5(32'h3a1a1aa9),
	.w6(32'h3a172539),
	.w7(32'h3a890cb1),
	.w8(32'h3987e512),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ee900),
	.w1(32'hba5ca8b1),
	.w2(32'hba64621d),
	.w3(32'h3a3471c4),
	.w4(32'hbaac4854),
	.w5(32'hbaa1a07d),
	.w6(32'h3a6eb68b),
	.w7(32'h39f18044),
	.w8(32'h3a1aa4c2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e5ef8),
	.w1(32'hb9e4765e),
	.w2(32'hb9dea9c4),
	.w3(32'hba03075c),
	.w4(32'h383cafd2),
	.w5(32'hb9ff12f7),
	.w6(32'h391b2c48),
	.w7(32'h39c4f3e3),
	.w8(32'hba4281a4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba333774),
	.w1(32'h3ba92ef9),
	.w2(32'h3c24b535),
	.w3(32'hb9f670c7),
	.w4(32'h3b7df569),
	.w5(32'h3bf3986b),
	.w6(32'h3c49e335),
	.w7(32'h3c538d68),
	.w8(32'h3bdcea23),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c5573),
	.w1(32'hba54af40),
	.w2(32'hba9a36ed),
	.w3(32'h3b4f72b0),
	.w4(32'h39f87294),
	.w5(32'hb86f664e),
	.w6(32'hb95c2c38),
	.w7(32'h3a3d7113),
	.w8(32'hbaa28fda),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f432b),
	.w1(32'hb8d29618),
	.w2(32'h3ab45ae9),
	.w3(32'hbab8c606),
	.w4(32'hb94d7a3b),
	.w5(32'h3adf310d),
	.w6(32'hb74f78d3),
	.w7(32'h39d58f51),
	.w8(32'hba571fc2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba517c20),
	.w1(32'h3b50e1a7),
	.w2(32'h3aecdb29),
	.w3(32'h384f986a),
	.w4(32'h3b4819ad),
	.w5(32'h3a9f643b),
	.w6(32'h3a786e91),
	.w7(32'h37d23854),
	.w8(32'hbadf64d7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa24cb9),
	.w1(32'h3a701b78),
	.w2(32'hba07d5f7),
	.w3(32'h39d5a126),
	.w4(32'h3a85f196),
	.w5(32'h3a4c9a33),
	.w6(32'hb9d44ed7),
	.w7(32'h3a461ad8),
	.w8(32'h3a80a741),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86457a),
	.w1(32'hba55af5c),
	.w2(32'hb9a0cfae),
	.w3(32'hb8e4d045),
	.w4(32'h397df60d),
	.w5(32'h3a1d638a),
	.w6(32'h3ab749c8),
	.w7(32'h3ac94f44),
	.w8(32'h38f6cbe6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7b819),
	.w1(32'hba1eb1a8),
	.w2(32'h3a74e4e8),
	.w3(32'h3a1304a2),
	.w4(32'hbafd53c9),
	.w5(32'hbad65638),
	.w6(32'h39915228),
	.w7(32'h3ab16d29),
	.w8(32'hb9c0fc81),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf04981),
	.w1(32'h3bc0a8cd),
	.w2(32'hbb0bf538),
	.w3(32'hbb031fea),
	.w4(32'h3a9b0f7a),
	.w5(32'hbc195158),
	.w6(32'h3c9b85a5),
	.w7(32'h3c1c1f76),
	.w8(32'h3c7929df),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98e591),
	.w1(32'hba861685),
	.w2(32'h3a3c276d),
	.w3(32'hbac536a9),
	.w4(32'hb9d4fc45),
	.w5(32'h3a99d2f9),
	.w6(32'hb95616ba),
	.w7(32'h3a0d98ac),
	.w8(32'hba32e47a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba635e1f),
	.w1(32'hba3d60a4),
	.w2(32'h3871400b),
	.w3(32'hb9060974),
	.w4(32'hba7f9bb5),
	.w5(32'hba27a048),
	.w6(32'h39abf531),
	.w7(32'h3a8f8fd6),
	.w8(32'h39b503a1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d0f1b2),
	.w1(32'h396b4795),
	.w2(32'h3a469e41),
	.w3(32'hba14067f),
	.w4(32'hba1e44d5),
	.w5(32'h391aadc1),
	.w6(32'hba1cfa93),
	.w7(32'hb8ba74a4),
	.w8(32'hbb0f2ee2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafded2),
	.w1(32'hbaa2865c),
	.w2(32'hb937457b),
	.w3(32'hbace1433),
	.w4(32'hb92d3da9),
	.w5(32'h3aee6705),
	.w6(32'h3a973727),
	.w7(32'h3b05adbe),
	.w8(32'h3a99b186),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50b0b4),
	.w1(32'hba10ac15),
	.w2(32'h3ac531c8),
	.w3(32'hbb2e7808),
	.w4(32'h39b65494),
	.w5(32'h3b0e5059),
	.w6(32'h397e8a3d),
	.w7(32'h3a513d11),
	.w8(32'hbac60829),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5730cc),
	.w1(32'hba6e7a69),
	.w2(32'h391ce1f1),
	.w3(32'hb9edd613),
	.w4(32'hb8153625),
	.w5(32'h3ae42586),
	.w6(32'hbaa60f0c),
	.w7(32'hba080328),
	.w8(32'h392a3868),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94297ee),
	.w1(32'h3b6f5c1b),
	.w2(32'h3b2b1caf),
	.w3(32'hb9d9a2c4),
	.w4(32'h3b74e446),
	.w5(32'h3ae8fe81),
	.w6(32'h3b04727c),
	.w7(32'h39d53f31),
	.w8(32'hba63e70d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a927ab5),
	.w1(32'hbb2aca76),
	.w2(32'h3c086b92),
	.w3(32'h38597873),
	.w4(32'h3b1a86ef),
	.w5(32'h3c1df952),
	.w6(32'h3bb2d53c),
	.w7(32'h3c7ab348),
	.w8(32'h3c1695ac),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c236931),
	.w1(32'h3aba5a98),
	.w2(32'h3b51d65e),
	.w3(32'h3c20f4a1),
	.w4(32'h3a2bd4af),
	.w5(32'h3b37bb34),
	.w6(32'h3a9bcf1f),
	.w7(32'h3b33d16f),
	.w8(32'h3a91c530),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11f548),
	.w1(32'hbb10acab),
	.w2(32'h3a810edc),
	.w3(32'h3ae36cf3),
	.w4(32'hbb0d6fff),
	.w5(32'hba0ce7db),
	.w6(32'hbb0725b9),
	.w7(32'hbaf7fe04),
	.w8(32'hb9f102d4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94eb353),
	.w1(32'h3807b445),
	.w2(32'hba2aa1ab),
	.w3(32'h3ad1f7fb),
	.w4(32'h38dbddda),
	.w5(32'hba941915),
	.w6(32'h39e50930),
	.w7(32'h3a3e5aa4),
	.w8(32'h3904c03b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b78331),
	.w1(32'hba603363),
	.w2(32'hba6f4109),
	.w3(32'hbacba242),
	.w4(32'hba866bac),
	.w5(32'hba8f1a88),
	.w6(32'h3a854181),
	.w7(32'h3a2ca0ae),
	.w8(32'h39ff58ff),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f1a73),
	.w1(32'hb9c04f3c),
	.w2(32'hba974f5f),
	.w3(32'hba3579df),
	.w4(32'h3a4208bd),
	.w5(32'hb9b7f67f),
	.w6(32'h38d5df03),
	.w7(32'h3a2a0f8e),
	.w8(32'hba289dcb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ed85e),
	.w1(32'hbaa2fb05),
	.w2(32'hba3c35bb),
	.w3(32'hb9d532dd),
	.w4(32'hba85d63c),
	.w5(32'hba9c73a3),
	.w6(32'h3a5e5d47),
	.w7(32'h3b216437),
	.w8(32'h3aa0091c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa2db9),
	.w1(32'h3aba4124),
	.w2(32'hbab6d26d),
	.w3(32'hba8ec4d1),
	.w4(32'h3aac283a),
	.w5(32'h3a24e406),
	.w6(32'hbb398c83),
	.w7(32'hbb14fb4c),
	.w8(32'h3a2501dc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b298d64),
	.w1(32'h3b0a5219),
	.w2(32'h3a6e7693),
	.w3(32'h3b6c66e3),
	.w4(32'h3b15433f),
	.w5(32'h3a57445f),
	.w6(32'h3a3ff7f0),
	.w7(32'hb98bda29),
	.w8(32'hbab0a42b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a141209),
	.w1(32'hb930dcc0),
	.w2(32'hba85487d),
	.w3(32'h3967384c),
	.w4(32'h3ad75b3a),
	.w5(32'hba424ba6),
	.w6(32'h39b83101),
	.w7(32'hb9217b5f),
	.w8(32'h397b575c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925d390),
	.w1(32'hba50643a),
	.w2(32'h3b4186a3),
	.w3(32'h39aeaf14),
	.w4(32'hb836d520),
	.w5(32'h3ac76cc9),
	.w6(32'hb8eed7d5),
	.w7(32'hbadeb48e),
	.w8(32'hba94a123),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ee75c),
	.w1(32'h3b421115),
	.w2(32'h3be26667),
	.w3(32'h3ad2d215),
	.w4(32'h3ad27a78),
	.w5(32'h3bab4bdc),
	.w6(32'hbadf5da8),
	.w7(32'h3b0f39e7),
	.w8(32'h3b1d2721),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bd504),
	.w1(32'h3aea0766),
	.w2(32'h3c0bf19a),
	.w3(32'h3c08d89c),
	.w4(32'hba057799),
	.w5(32'h3b356408),
	.w6(32'h3c4b2668),
	.w7(32'h3c5609be),
	.w8(32'h3bef7aa6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5dc2f),
	.w1(32'hba008593),
	.w2(32'h3a98022c),
	.w3(32'hbb781918),
	.w4(32'hbab3f1da),
	.w5(32'h3a203873),
	.w6(32'h394c56dc),
	.w7(32'h3a99d4d7),
	.w8(32'hba80f676),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba687abe),
	.w1(32'hb6bc7426),
	.w2(32'h3b041da9),
	.w3(32'hbab57f1a),
	.w4(32'hb888fa76),
	.w5(32'hba13c9ce),
	.w6(32'h3ac4b74a),
	.w7(32'h3ab13140),
	.w8(32'hb976fb3e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5eefb),
	.w1(32'hb8399dca),
	.w2(32'hb8bdc2ae),
	.w3(32'hba6f1367),
	.w4(32'h39e44cfc),
	.w5(32'hba220583),
	.w6(32'h396b750a),
	.w7(32'h39c264ff),
	.w8(32'h3936398d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11b75b),
	.w1(32'hbb0d40a3),
	.w2(32'hb92ac012),
	.w3(32'h3951239c),
	.w4(32'hbaf026f9),
	.w5(32'hba1fc6d6),
	.w6(32'hb9bdc896),
	.w7(32'h3a5a9eb5),
	.w8(32'h3967c22b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba275d9a),
	.w1(32'hba525f74),
	.w2(32'hba302eb7),
	.w3(32'hb8f5f8c7),
	.w4(32'hba9f675b),
	.w5(32'hba9d85e2),
	.w6(32'h3a898d32),
	.w7(32'h3a50ba1c),
	.w8(32'h3a4469ca),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9a761),
	.w1(32'hba94dad1),
	.w2(32'h3aab9af5),
	.w3(32'hba266692),
	.w4(32'hba90cfa3),
	.w5(32'h3a83d569),
	.w6(32'h3a707be9),
	.w7(32'h3acf1a74),
	.w8(32'h39a08644),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ff116),
	.w1(32'h39b8c9ca),
	.w2(32'hba43f450),
	.w3(32'hba05674e),
	.w4(32'h3a286e2e),
	.w5(32'hba20ec3f),
	.w6(32'h3ab5d896),
	.w7(32'h3a875e5a),
	.w8(32'h3a0ea3d0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02e13f),
	.w1(32'h388fe2ef),
	.w2(32'h3ba5882a),
	.w3(32'hba7e24f1),
	.w4(32'h3bb2aa0b),
	.w5(32'h3bd630b6),
	.w6(32'hbba4acbd),
	.w7(32'hbb49c08a),
	.w8(32'hbab5c8dc),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae64b8a),
	.w1(32'hba5fd45f),
	.w2(32'hb9e3a48c),
	.w3(32'h3acd089c),
	.w4(32'hba2b6875),
	.w5(32'hba9ba5d2),
	.w6(32'h3aafdb89),
	.w7(32'h3a760671),
	.w8(32'h3a9c35f9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954ac4f),
	.w1(32'hb9cee178),
	.w2(32'hbafd5dc3),
	.w3(32'hba002111),
	.w4(32'h39910a88),
	.w5(32'hba8262b1),
	.w6(32'hbabc6007),
	.w7(32'h38bbeabf),
	.w8(32'h3acf6740),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e5d50),
	.w1(32'h3ba62b4d),
	.w2(32'h3b3450ae),
	.w3(32'h3aa07496),
	.w4(32'h3ba1c24c),
	.w5(32'h39f67064),
	.w6(32'h38012cf2),
	.w7(32'hbb8b9335),
	.w8(32'hbacdd0a2),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393138c6),
	.w1(32'hba89b893),
	.w2(32'h39955516),
	.w3(32'hbb263cdd),
	.w4(32'hba9a2d54),
	.w5(32'hba66c849),
	.w6(32'h3b4fead3),
	.w7(32'h3abee6e9),
	.w8(32'h3a6b0651),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52b008),
	.w1(32'h39a464d1),
	.w2(32'h3ba5d279),
	.w3(32'hba203d3d),
	.w4(32'h3a84a5ee),
	.w5(32'h3b47487c),
	.w6(32'h3c227cfb),
	.w7(32'h3c331482),
	.w8(32'h3c3383c6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c026e60),
	.w1(32'h3a8484cd),
	.w2(32'hba069ffb),
	.w3(32'h3badb40c),
	.w4(32'h3aed7f2b),
	.w5(32'h3a16436d),
	.w6(32'hb9eca433),
	.w7(32'h39c977ac),
	.w8(32'hba95970c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39286b36),
	.w1(32'h3b304de2),
	.w2(32'h3b330180),
	.w3(32'hb9a1e562),
	.w4(32'h3b14e213),
	.w5(32'h39f4598a),
	.w6(32'h3c024412),
	.w7(32'h3be9e862),
	.w8(32'h3ba292bd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68c187),
	.w1(32'h39e64296),
	.w2(32'hb9f7a130),
	.w3(32'hbace1e74),
	.w4(32'h3a6ad734),
	.w5(32'h39be3185),
	.w6(32'h39581dee),
	.w7(32'h3964dcc2),
	.w8(32'hb8e1c518),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d33068),
	.w1(32'hbb13a7f7),
	.w2(32'hbbbf484b),
	.w3(32'hb9129d47),
	.w4(32'hbc090d6f),
	.w5(32'hbc56dec6),
	.w6(32'h3ba3d94c),
	.w7(32'hba08536d),
	.w8(32'h3bbca8c7),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26eab1),
	.w1(32'h3b2be399),
	.w2(32'h3b8a2946),
	.w3(32'hbbf24571),
	.w4(32'h3b213a35),
	.w5(32'h3b5a4b0a),
	.w6(32'h3aa52f09),
	.w7(32'h3b565ff6),
	.w8(32'h3b2a5289),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcae4b),
	.w1(32'hba02c0c9),
	.w2(32'hba165d21),
	.w3(32'h3b8b2caf),
	.w4(32'h388c985c),
	.w5(32'hba50ca7e),
	.w6(32'hba092294),
	.w7(32'hbaaeecbd),
	.w8(32'hbb12400f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00fabf),
	.w1(32'hba13bbdd),
	.w2(32'h3a2b0cce),
	.w3(32'hb9f2ce54),
	.w4(32'hba56b49f),
	.w5(32'h38940856),
	.w6(32'h3ac83f6c),
	.w7(32'h3ac780d1),
	.w8(32'h39e817bc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0823b9),
	.w1(32'h3af0cc51),
	.w2(32'h3a33ea88),
	.w3(32'hb9ec44e2),
	.w4(32'h3af6e14e),
	.w5(32'h39a276cd),
	.w6(32'h3aca7d06),
	.w7(32'h3a7b47a6),
	.w8(32'hbab2698f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396871c3),
	.w1(32'hbaaabef5),
	.w2(32'h3a93eb71),
	.w3(32'hb9eb6bf4),
	.w4(32'hbacf64dc),
	.w5(32'h39414ada),
	.w6(32'h3a6d55e1),
	.w7(32'h3a701f95),
	.w8(32'hb90fa7f4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba298a9a),
	.w1(32'hba8764e6),
	.w2(32'h37a3e6b9),
	.w3(32'hba1ffd20),
	.w4(32'hba7362f2),
	.w5(32'h38b0eba1),
	.w6(32'h3b374934),
	.w7(32'h3b3de280),
	.w8(32'h3b221a06),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f1edd),
	.w1(32'h39a325bd),
	.w2(32'h371865f6),
	.w3(32'hb9a9225d),
	.w4(32'h3ae967b2),
	.w5(32'h3ad598b0),
	.w6(32'hbb13de5f),
	.w7(32'hbb0ca63e),
	.w8(32'hbb34b976),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996fdf3),
	.w1(32'h3a54a3ae),
	.w2(32'hba7c43ee),
	.w3(32'h3a93ad0d),
	.w4(32'h3a934805),
	.w5(32'hba679880),
	.w6(32'hb864e8bf),
	.w7(32'hbab2b28e),
	.w8(32'hbad1314e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad19564),
	.w1(32'h3a950c97),
	.w2(32'h3bd9171a),
	.w3(32'hba735ba0),
	.w4(32'h3b2e10df),
	.w5(32'h3ba5f1a8),
	.w6(32'h3c403af8),
	.w7(32'h3c5b9d4f),
	.w8(32'h3c159ac0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2d061),
	.w1(32'hbb07bc44),
	.w2(32'hbb28fed9),
	.w3(32'h3b899767),
	.w4(32'h38889779),
	.w5(32'hba438b13),
	.w6(32'h3a9569e1),
	.w7(32'h3aca3b22),
	.w8(32'h3abdd5e9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03ac62),
	.w1(32'hba27314c),
	.w2(32'h39defc0c),
	.w3(32'hba2628b2),
	.w4(32'hba1d00da),
	.w5(32'hb9bd4c6d),
	.w6(32'hb99c317c),
	.w7(32'h3a2c9a87),
	.w8(32'h3a27c750),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e97e9),
	.w1(32'hb9bd7489),
	.w2(32'h3ade5359),
	.w3(32'h3907e9e2),
	.w4(32'hbab0828b),
	.w5(32'hb8249fee),
	.w6(32'h3b3e8208),
	.w7(32'h3bbb76c3),
	.w8(32'h3ba450e0),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af95dd2),
	.w1(32'h3afdeaa7),
	.w2(32'h39dfeab1),
	.w3(32'hba9282e3),
	.w4(32'h3afb92b1),
	.w5(32'hb8c87150),
	.w6(32'h3aaf51bc),
	.w7(32'hb9ae67be),
	.w8(32'h3a1a33b9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1a21b),
	.w1(32'hb8f0622d),
	.w2(32'hba39e876),
	.w3(32'hbaa85eb6),
	.w4(32'h398d39ff),
	.w5(32'hba651fca),
	.w6(32'hba8a4a9f),
	.w7(32'hb98f143d),
	.w8(32'hbaddaaa6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95e145),
	.w1(32'h3b410c53),
	.w2(32'h3aa55a09),
	.w3(32'hb9a270f4),
	.w4(32'h3b81289f),
	.w5(32'h3af4d7ac),
	.w6(32'h3b989b40),
	.w7(32'h3a9ce969),
	.w8(32'h3a15ed40),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cab3c6),
	.w1(32'hbb32bb8d),
	.w2(32'h3bc7734c),
	.w3(32'h39d76ade),
	.w4(32'hb9b84ea3),
	.w5(32'h3bac60cc),
	.w6(32'hbb376b55),
	.w7(32'h3b2832e8),
	.w8(32'hbac41350),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399394a1),
	.w1(32'hbb5115f2),
	.w2(32'h3ad4d46a),
	.w3(32'h39c1b48c),
	.w4(32'hb99cb51a),
	.w5(32'h3bb4f73f),
	.w6(32'hbb8ee903),
	.w7(32'hbb13f118),
	.w8(32'hbaaa9bb3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f0d39),
	.w1(32'hbabb85df),
	.w2(32'hba4b5d0e),
	.w3(32'h3b6615b6),
	.w4(32'hba9f9766),
	.w5(32'hbafecafb),
	.w6(32'h3afbd2fd),
	.w7(32'h3aa7c209),
	.w8(32'h3add3fc4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94bce45),
	.w1(32'hbb2b04e9),
	.w2(32'hb8f5f405),
	.w3(32'hba08bc5f),
	.w4(32'hbb0899dc),
	.w5(32'hba20f261),
	.w6(32'hba31c67d),
	.w7(32'h3a3e5b96),
	.w8(32'hb8f3d0df),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c16f1),
	.w1(32'hb9ffb5ac),
	.w2(32'hb986fdaf),
	.w3(32'hb9f6f303),
	.w4(32'hb9b4343d),
	.w5(32'hba67e1a1),
	.w6(32'h3a9f99ee),
	.w7(32'h3a3c869d),
	.w8(32'h3a791139),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eccbe9),
	.w1(32'hb73779c7),
	.w2(32'hba58b036),
	.w3(32'hb9bb228e),
	.w4(32'hb7b3dd3f),
	.w5(32'hba6fe038),
	.w6(32'h3914f551),
	.w7(32'hb9b5689c),
	.w8(32'h39410592),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b12540),
	.w1(32'hba8e654e),
	.w2(32'hbb28ae91),
	.w3(32'hb9fe6909),
	.w4(32'h3a29ca36),
	.w5(32'hba548df2),
	.w6(32'h3afeedeb),
	.w7(32'h3b0e6db2),
	.w8(32'h3b28bcde),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94f5ae),
	.w1(32'hb90fa475),
	.w2(32'h3af8090a),
	.w3(32'hb9f7439d),
	.w4(32'hba08a547),
	.w5(32'h39ef3ee4),
	.w6(32'h3b567540),
	.w7(32'h3b7cc4cb),
	.w8(32'h3b0b6ef4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f4ce4),
	.w1(32'hba65f8ec),
	.w2(32'hba01b198),
	.w3(32'hb9d41f18),
	.w4(32'hba37c17c),
	.w5(32'hba8851fa),
	.w6(32'h3a6897af),
	.w7(32'h3a36aec1),
	.w8(32'h3a4b6b24),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9890cd3),
	.w1(32'h3a629fe3),
	.w2(32'h3a12e543),
	.w3(32'hb9ea17e6),
	.w4(32'h3ac6cbf9),
	.w5(32'h3af603b8),
	.w6(32'hba963a42),
	.w7(32'h3a341ffe),
	.w8(32'h3a777e96),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae708d5),
	.w1(32'h38b24afa),
	.w2(32'hb9119ad6),
	.w3(32'h3ab6f0a8),
	.w4(32'hb9b380ef),
	.w5(32'h39b20d02),
	.w6(32'h3ab2ed23),
	.w7(32'h3a6b94c7),
	.w8(32'h39b8370e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38545260),
	.w1(32'h3ad3d7fb),
	.w2(32'h3a98a2a8),
	.w3(32'hb9d42784),
	.w4(32'h3acda726),
	.w5(32'h3b6e2451),
	.w6(32'hba9e9016),
	.w7(32'hb84f1cb9),
	.w8(32'h38c0d388),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13725a),
	.w1(32'h39465893),
	.w2(32'hb938b1c7),
	.w3(32'hbb012816),
	.w4(32'hb9e0f2b4),
	.w5(32'h38cdc514),
	.w6(32'h3b0b2e75),
	.w7(32'h3a59fcde),
	.w8(32'h38bb5c99),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba059e33),
	.w1(32'hba60557f),
	.w2(32'hbaf6ab1c),
	.w3(32'hba779e35),
	.w4(32'h3a95858b),
	.w5(32'h3910a45b),
	.w6(32'h3a6a2c82),
	.w7(32'h3aa9913a),
	.w8(32'h395551ae),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba829187),
	.w1(32'hb89482e9),
	.w2(32'h39849213),
	.w3(32'h39937457),
	.w4(32'hbaa61153),
	.w5(32'h3adaa64b),
	.w6(32'hba61c2e9),
	.w7(32'hba2f9de5),
	.w8(32'hba893a0e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d30bed),
	.w1(32'hba87dd02),
	.w2(32'hba1c4c77),
	.w3(32'h3aa98a15),
	.w4(32'hba588fce),
	.w5(32'hbab79cdd),
	.w6(32'h3abdf7fd),
	.w7(32'h3a85feeb),
	.w8(32'h3aab8c4d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9207ea3),
	.w1(32'hbaa46436),
	.w2(32'hba413297),
	.w3(32'hb9f6562d),
	.w4(32'hba82472a),
	.w5(32'hbaa8c287),
	.w6(32'h397cdc09),
	.w7(32'h39e498ad),
	.w8(32'h3a302d17),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbdd22),
	.w1(32'hba3885ba),
	.w2(32'hba5ddea6),
	.w3(32'hb9671907),
	.w4(32'hb99ce700),
	.w5(32'hba950057),
	.w6(32'h3a8d196f),
	.w7(32'h3a1cffdf),
	.w8(32'h3a996853),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91dab44),
	.w1(32'hbac4f6e9),
	.w2(32'hbb19725c),
	.w3(32'hb9075284),
	.w4(32'h38a3d5a4),
	.w5(32'h38c57162),
	.w6(32'hbaeec80a),
	.w7(32'h39894156),
	.w8(32'h3923d4aa),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4faaf0),
	.w1(32'hba19164b),
	.w2(32'h3a1e2884),
	.w3(32'hba2d414f),
	.w4(32'hb900fc7e),
	.w5(32'h3a175b1a),
	.w6(32'h3abbd96f),
	.w7(32'h3a99adfb),
	.w8(32'h3abe87e0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedacd9),
	.w1(32'hbad6d57b),
	.w2(32'hba31e6fb),
	.w3(32'h3a30b0c2),
	.w4(32'hb9b28846),
	.w5(32'h3a0ef701),
	.w6(32'h3911753d),
	.w7(32'h3a644689),
	.w8(32'h3822f0ff),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bf1cb),
	.w1(32'hb8184000),
	.w2(32'hbb32628a),
	.w3(32'h3a0a860f),
	.w4(32'hb8ca9a04),
	.w5(32'hbaac6b41),
	.w6(32'h3a51b0db),
	.w7(32'hba795de7),
	.w8(32'hb9d29d65),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4725fe),
	.w1(32'hbab463e0),
	.w2(32'hba81a016),
	.w3(32'hb91fcb96),
	.w4(32'hbaae1245),
	.w5(32'hba954025),
	.w6(32'h3a1b6735),
	.w7(32'h3a170cfe),
	.w8(32'h39a4d0f9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c211c),
	.w1(32'hbb12dcc3),
	.w2(32'hbb2aed42),
	.w3(32'hba5a6548),
	.w4(32'hba982990),
	.w5(32'h39f63183),
	.w6(32'hbb98976b),
	.w7(32'hbb0fd4ea),
	.w8(32'hbb20f35b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1da780),
	.w1(32'h3a113caf),
	.w2(32'h3ad7ee47),
	.w3(32'h38f50a1e),
	.w4(32'h3a4bd713),
	.w5(32'h3add9f11),
	.w6(32'h3b067eff),
	.w7(32'h38afdb94),
	.w8(32'hb9e88bd5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb882de9e),
	.w1(32'h3a82c178),
	.w2(32'h39a7b474),
	.w3(32'h3ab5f08d),
	.w4(32'h39ad6051),
	.w5(32'hba3a7e4c),
	.w6(32'h3bb05130),
	.w7(32'h3b07c786),
	.w8(32'h3abf30dc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09bded),
	.w1(32'hb6842ee9),
	.w2(32'hb699184e),
	.w3(32'hb99be254),
	.w4(32'h353d315f),
	.w5(32'hb69e10d6),
	.w6(32'hb68ae190),
	.w7(32'h367c4da7),
	.w8(32'hb7669b4d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85a30af),
	.w1(32'hb53e2c0f),
	.w2(32'h36f99033),
	.w3(32'hb8070401),
	.w4(32'hb86791fc),
	.w5(32'hb799139a),
	.w6(32'hb7153bde),
	.w7(32'hb7b73aa6),
	.w8(32'h3604c3ca),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8328a32),
	.w1(32'hb7bdc486),
	.w2(32'hb62173f3),
	.w3(32'hb84a95b5),
	.w4(32'hb829f060),
	.w5(32'hb7670eeb),
	.w6(32'hb83e71e3),
	.w7(32'hb71de3d8),
	.w8(32'hb69a8ed9),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37987acc),
	.w1(32'h36bd7b84),
	.w2(32'h3795d59e),
	.w3(32'h376d9aa6),
	.w4(32'h371e7b0c),
	.w5(32'h36eb124f),
	.w6(32'hb59ae9ee),
	.w7(32'hb73e2acf),
	.w8(32'hb4c36349),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3696c455),
	.w1(32'h3762caff),
	.w2(32'hb7651ad9),
	.w3(32'h36ad5617),
	.w4(32'h3777a2db),
	.w5(32'hb4d2c632),
	.w6(32'hb75350da),
	.w7(32'h36fd38de),
	.w8(32'hb5e3d5d7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74bc78a),
	.w1(32'hb780a5d5),
	.w2(32'hb6a91b5e),
	.w3(32'hb75e31ba),
	.w4(32'h362dc231),
	.w5(32'h362e930b),
	.w6(32'hb6acfd88),
	.w7(32'h3782bd42),
	.w8(32'h37884f24),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82a62cf),
	.w1(32'hb7eb23e8),
	.w2(32'hb7e551a6),
	.w3(32'hb759378d),
	.w4(32'hb5f82b9f),
	.w5(32'hb7c3d204),
	.w6(32'hb7af323f),
	.w7(32'hb2d26d1a),
	.w8(32'hb7ab13c9),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84a54ec),
	.w1(32'h379911fc),
	.w2(32'h3738e4c7),
	.w3(32'hb81fb6b3),
	.w4(32'h37ef844e),
	.w5(32'hb7038f80),
	.w6(32'h37d9174a),
	.w7(32'h386a1013),
	.w8(32'h37459dd5),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3775c626),
	.w1(32'h382b5b22),
	.w2(32'h381d7983),
	.w3(32'h37d44485),
	.w4(32'h37f3f87a),
	.w5(32'h37d5cfab),
	.w6(32'hb6dd5afa),
	.w7(32'hb71fb805),
	.w8(32'h37f1cc50),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886f00b),
	.w1(32'hb8470831),
	.w2(32'hb835c272),
	.w3(32'hb8224846),
	.w4(32'hb79474df),
	.w5(32'hb77ae5e1),
	.w6(32'hb7aaee80),
	.w7(32'h373ea616),
	.w8(32'hb757153d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c766b8),
	.w1(32'hb53c1607),
	.w2(32'h374cacb9),
	.w3(32'hb84b8189),
	.w4(32'hb7e5b5dd),
	.w5(32'hb807e3e5),
	.w6(32'hb7a1458d),
	.w7(32'hb79e50c5),
	.w8(32'hb6b6f715),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b9f56c),
	.w1(32'h380eded9),
	.w2(32'h37d51d91),
	.w3(32'h37e2c136),
	.w4(32'h37a57051),
	.w5(32'hb7cc986e),
	.w6(32'hb816b35b),
	.w7(32'hb87a9e9b),
	.w8(32'hb82611b6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c67ca2),
	.w1(32'hb7e47cb7),
	.w2(32'hb780ee8c),
	.w3(32'hb7471ac0),
	.w4(32'hb83013a6),
	.w5(32'hb7ef2d7d),
	.w6(32'hb655d1b0),
	.w7(32'hb7081668),
	.w8(32'hb78f691e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb766c706),
	.w1(32'hb7ac77b3),
	.w2(32'hb6867aa0),
	.w3(32'hb81a6189),
	.w4(32'hb6390b00),
	.w5(32'hb729dc06),
	.w6(32'hb7f1b7a0),
	.w7(32'h36d1f845),
	.w8(32'h37a1a36b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7abed82),
	.w1(32'hb6762832),
	.w2(32'hb6854442),
	.w3(32'hb755c3a0),
	.w4(32'hb62fe2b7),
	.w5(32'hb597c9b8),
	.w6(32'hb6cfc9f4),
	.w7(32'h372f28f1),
	.w8(32'h36b6b044),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9387a26),
	.w1(32'hb8dc8e3e),
	.w2(32'hb8ada993),
	.w3(32'hb8f1839b),
	.w4(32'hb877779d),
	.w5(32'hb717199a),
	.w6(32'hb7f5ebf5),
	.w7(32'h3828473b),
	.w8(32'h38601c34),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e39ceb),
	.w1(32'hb7bb8679),
	.w2(32'h372d4fa9),
	.w3(32'hb7ec39f7),
	.w4(32'h374f0df1),
	.w5(32'h37ee2e9e),
	.w6(32'hb7ba4f36),
	.w7(32'h3818fb4d),
	.w8(32'h38742817),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373e0aae),
	.w1(32'h367751b7),
	.w2(32'h370e8a74),
	.w3(32'hb68fc934),
	.w4(32'h3677bb4d),
	.w5(32'h366ab3f9),
	.w6(32'h34759e53),
	.w7(32'h369d802f),
	.w8(32'h35e727e7),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35bb97ae),
	.w1(32'h35aff0e9),
	.w2(32'hb5a36f51),
	.w3(32'h35b25f42),
	.w4(32'hb52a2eaf),
	.w5(32'hb6910be7),
	.w6(32'hb676a012),
	.w7(32'hb7039da2),
	.w8(32'h36a001ff),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fe0ab3),
	.w1(32'hb73fee87),
	.w2(32'hb72778d6),
	.w3(32'hb6e909de),
	.w4(32'hb794c8ba),
	.w5(32'hb7d2c2a4),
	.w6(32'h377dfd07),
	.w7(32'hb6d43218),
	.w8(32'hb719f66c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a44010),
	.w1(32'hb8868b82),
	.w2(32'hb6c2a909),
	.w3(32'hb86d7828),
	.w4(32'hb8428887),
	.w5(32'hb714454d),
	.w6(32'hb802be97),
	.w7(32'hb660b495),
	.w8(32'hb7bf8d7f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81b355a),
	.w1(32'hb7098272),
	.w2(32'hb60f2065),
	.w3(32'hb85531d3),
	.w4(32'hb698f409),
	.w5(32'h35246c42),
	.w6(32'hb83b2201),
	.w7(32'h36b7319f),
	.w8(32'h373c5f0e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3587bd37),
	.w1(32'hb6971fae),
	.w2(32'hb620ba54),
	.w3(32'hb5512988),
	.w4(32'hb6731109),
	.w5(32'hb6f05691),
	.w6(32'hb6f1d7c0),
	.w7(32'hb6088c9f),
	.w8(32'hb72c91d2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8809547),
	.w1(32'hb7db8524),
	.w2(32'hb5c62115),
	.w3(32'hb84d1768),
	.w4(32'hb81951b3),
	.w5(32'hb68c4d21),
	.w6(32'hb806a2f3),
	.w7(32'hb63fae42),
	.w8(32'h36d727f2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb791c41c),
	.w1(32'hb85b6b94),
	.w2(32'hb8614419),
	.w3(32'hb784dafd),
	.w4(32'hb86858c6),
	.w5(32'hb85e5fa1),
	.w6(32'h36a0539d),
	.w7(32'hb6a072e3),
	.w8(32'hb7c65560),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ecf98c),
	.w1(32'h385677e1),
	.w2(32'h3850bc98),
	.w3(32'h368c0fb9),
	.w4(32'hb8290807),
	.w5(32'hb855908a),
	.w6(32'hb789e9db),
	.w7(32'hb8104765),
	.w8(32'hb825ad99),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918aa8f),
	.w1(32'hb8704ce7),
	.w2(32'hb7d98b41),
	.w3(32'hb9143d79),
	.w4(32'hb88dc760),
	.w5(32'h3675b082),
	.w6(32'hb8b50563),
	.w7(32'h36d8b044),
	.w8(32'h385363f9),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80762a1),
	.w1(32'hb7d86945),
	.w2(32'hb80efd69),
	.w3(32'hb7d14cb8),
	.w4(32'hb7b7635b),
	.w5(32'hb834e0a9),
	.w6(32'hb8362eea),
	.w7(32'hb8294185),
	.w8(32'hb83c3c4f),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bba02e),
	.w1(32'h36548a70),
	.w2(32'hb80c35ed),
	.w3(32'h379e7d54),
	.w4(32'h3804d6f9),
	.w5(32'h371ecd1d),
	.w6(32'h37df896e),
	.w7(32'h380214e6),
	.w8(32'h375ebc39),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c2de49),
	.w1(32'hb8311477),
	.w2(32'hb79590c1),
	.w3(32'hb870cdd8),
	.w4(32'h372c6a2a),
	.w5(32'h373bfc33),
	.w6(32'hb8799396),
	.w7(32'hb7b5c25d),
	.w8(32'hb818b9ed),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885f102),
	.w1(32'hb8626232),
	.w2(32'hb7e3b6b0),
	.w3(32'hb8af8b21),
	.w4(32'hb88ab1b2),
	.w5(32'hb7b96881),
	.w6(32'hb7bee21e),
	.w7(32'hb5e18831),
	.w8(32'h36cea22b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d53b9f),
	.w1(32'h37509f62),
	.w2(32'hb550d640),
	.w3(32'h3733c785),
	.w4(32'h37e6bcd1),
	.w5(32'h3754a3ac),
	.w6(32'h3700c914),
	.w7(32'h37bff0a2),
	.w8(32'h380881fc),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b35d8e),
	.w1(32'h378a7c4e),
	.w2(32'h379b5c08),
	.w3(32'h371a717a),
	.w4(32'h3750ecd2),
	.w5(32'h37012ff2),
	.w6(32'h3733f45c),
	.w7(32'h375ae41c),
	.w8(32'h376e761a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365b2927),
	.w1(32'h359251a1),
	.w2(32'h36137b08),
	.w3(32'hb57e69dd),
	.w4(32'hb66c4b9f),
	.w5(32'hb6a68ac1),
	.w6(32'hb68b43da),
	.w7(32'hb707efd9),
	.w8(32'hb72312fa),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82a183e),
	.w1(32'h37714ed9),
	.w2(32'h373530ef),
	.w3(32'hb84460d3),
	.w4(32'hb79cac3f),
	.w5(32'hb7d48ed7),
	.w6(32'hb7dd08ef),
	.w7(32'hb82eb459),
	.w8(32'h3786aae4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb622c636),
	.w1(32'hb72a3651),
	.w2(32'hb61812db),
	.w3(32'hb7336ce3),
	.w4(32'hb6c8bada),
	.w5(32'h37bba03a),
	.w6(32'h357079dd),
	.w7(32'h35382f41),
	.w8(32'h37b7db20),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8adb219),
	.w1(32'hb81ff9dd),
	.w2(32'hb8045b95),
	.w3(32'hb838089c),
	.w4(32'hb719e7f8),
	.w5(32'h36da10e5),
	.w6(32'hb82f7c16),
	.w7(32'h36949b11),
	.w8(32'h37a9452f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3491e5a6),
	.w1(32'h366c6ad6),
	.w2(32'hb7a176de),
	.w3(32'h3458a18f),
	.w4(32'h370b10fb),
	.w5(32'hb785a9f0),
	.w6(32'hb70e3fb6),
	.w7(32'h35b6cf0f),
	.w8(32'hb7112150),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a9c789),
	.w1(32'h37b134ad),
	.w2(32'hb6e47da7),
	.w3(32'h385330b1),
	.w4(32'h387e36a3),
	.w5(32'h37875a5f),
	.w6(32'h37da2455),
	.w7(32'h37952a86),
	.w8(32'hb7555de4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6993c68),
	.w1(32'h33f7ba5d),
	.w2(32'hb60223ad),
	.w3(32'hb6ad6d50),
	.w4(32'h3607be82),
	.w5(32'hb5dc554f),
	.w6(32'hb7181d03),
	.w7(32'hb642c4ed),
	.w8(32'h34d4e8dc),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h351095a2),
	.w1(32'hb74ccff5),
	.w2(32'hb76615e3),
	.w3(32'h375d4529),
	.w4(32'hb71eb644),
	.w5(32'hb78f9404),
	.w6(32'hb7016e21),
	.w7(32'hb7793e0d),
	.w8(32'hb7e0d4a7),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d6e7bf),
	.w1(32'hb83bc266),
	.w2(32'hb8657acc),
	.w3(32'hb8de3b6f),
	.w4(32'hb7a0d379),
	.w5(32'hb7dab8a0),
	.w6(32'hb88611f8),
	.w7(32'h35a14e2f),
	.w8(32'hb7736768),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83f9cef),
	.w1(32'h370d3561),
	.w2(32'h38923e07),
	.w3(32'hb7e06911),
	.w4(32'h36ab69c5),
	.w5(32'h37fb9d16),
	.w6(32'hb600390f),
	.w7(32'h3773be7d),
	.w8(32'h3813e32f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b7f7d0),
	.w1(32'h3778a7a1),
	.w2(32'hb81c7baa),
	.w3(32'h38317128),
	.w4(32'h3810c4f7),
	.w5(32'hb7f03bbf),
	.w6(32'h382f0c00),
	.w7(32'h37dfba41),
	.w8(32'hb5ab64bb),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d18692),
	.w1(32'hb8885051),
	.w2(32'hb8985c6d),
	.w3(32'hb88b4db4),
	.w4(32'hb82d2323),
	.w5(32'hb836b5fc),
	.w6(32'hb80ff782),
	.w7(32'hb71481ca),
	.w8(32'hb80a38aa),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d1a290),
	.w1(32'hb732522d),
	.w2(32'h36223216),
	.w3(32'hb768573a),
	.w4(32'hb771b95e),
	.w5(32'hb71dfe3d),
	.w6(32'h373e516f),
	.w7(32'h37510ec1),
	.w8(32'h3735eef5),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb825b0d6),
	.w1(32'h370facaf),
	.w2(32'hb8289c78),
	.w3(32'hb8035e2d),
	.w4(32'hb7bd185d),
	.w5(32'hb77b1b13),
	.w6(32'hb819c47a),
	.w7(32'hb68ff3b7),
	.w8(32'h3640eb59),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87a90f2),
	.w1(32'hb8691344),
	.w2(32'hb8affeec),
	.w3(32'hb601a08f),
	.w4(32'hb7b90e43),
	.w5(32'hb8464bc2),
	.w6(32'hb7c5bcd8),
	.w7(32'hb6d374d9),
	.w8(32'hb812dca4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a6ac60),
	.w1(32'h378005c9),
	.w2(32'h377ba18f),
	.w3(32'hb7bb7e81),
	.w4(32'h38556b54),
	.w5(32'h380175c3),
	.w6(32'hb81e7e30),
	.w7(32'h381d0188),
	.w8(32'h382ad21e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb50624e9),
	.w1(32'h37a8d57d),
	.w2(32'h37923aa3),
	.w3(32'h3735acf1),
	.w4(32'h380a6cd6),
	.w5(32'h3806bc41),
	.w6(32'h37a15a21),
	.w7(32'h380a31c9),
	.w8(32'h37e762f6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb864933c),
	.w1(32'hb66109b1),
	.w2(32'h36d4d6d0),
	.w3(32'hb82d08c8),
	.w4(32'hb77129f5),
	.w5(32'hb7a3f076),
	.w6(32'hb84345cf),
	.w7(32'hb80ef50a),
	.w8(32'hb7ee1b13),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36659f98),
	.w1(32'h3593c4c0),
	.w2(32'h36719cae),
	.w3(32'hb672be3f),
	.w4(32'hb67e36c8),
	.w5(32'hb5f68f4f),
	.w6(32'hb59d7aa1),
	.w7(32'h361e3e82),
	.w8(32'hb4c2ce29),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61b2270),
	.w1(32'hb7282685),
	.w2(32'hb79a5c90),
	.w3(32'hb717a133),
	.w4(32'hb6948385),
	.w5(32'hb78ae9e3),
	.w6(32'hb6e9b23d),
	.w7(32'hb72248f7),
	.w8(32'hb7783fda),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78be35b),
	.w1(32'hb50e7cf0),
	.w2(32'hb7268fd4),
	.w3(32'hb6f71f4b),
	.w4(32'hb68d954b),
	.w5(32'h35bb50ca),
	.w6(32'hb7785816),
	.w7(32'h366914cb),
	.w8(32'h3715a1f3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8476857),
	.w1(32'hb7b9f3cc),
	.w2(32'hb80c225a),
	.w3(32'hb7a87a87),
	.w4(32'hb70b5d06),
	.w5(32'hb822f0c7),
	.w6(32'h358dcdce),
	.w7(32'h37158d2d),
	.w8(32'hb8249049),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3592f034),
	.w1(32'hb63fe06a),
	.w2(32'hb5ea33c0),
	.w3(32'hb5cb7ddc),
	.w4(32'h3612be09),
	.w5(32'h36c03fc5),
	.w6(32'hb68416fa),
	.w7(32'hb687ce6a),
	.w8(32'hb5a1636b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7589b59),
	.w1(32'hb6cfb890),
	.w2(32'hb708d63e),
	.w3(32'hb775472f),
	.w4(32'hb5ec541b),
	.w5(32'hb72d0c16),
	.w6(32'hb488a67d),
	.w7(32'hb690de2c),
	.w8(32'hb6906cc0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c162bb),
	.w1(32'hb777bb0f),
	.w2(32'hb79336da),
	.w3(32'hb80a6f55),
	.w4(32'hb7f2c26d),
	.w5(32'hb7da57c7),
	.w6(32'hb6cd6379),
	.w7(32'hb62b36f9),
	.w8(32'h36c6c166),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3769c9a2),
	.w1(32'h3680c1f7),
	.w2(32'hb7237874),
	.w3(32'h3611bfbd),
	.w4(32'hb88fc698),
	.w5(32'hb88d98e0),
	.w6(32'h35a60379),
	.w7(32'hb6f2e3af),
	.w8(32'hb7a71dfd),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e23c2),
	.w1(32'h375982a0),
	.w2(32'h3840df1a),
	.w3(32'h38816f65),
	.w4(32'h36bb4ab0),
	.w5(32'h377e6956),
	.w6(32'h37b93b6c),
	.w7(32'hb7a40d01),
	.w8(32'h3666b3dc),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3690329c),
	.w1(32'h37519a75),
	.w2(32'hb69071c0),
	.w3(32'h36b07be0),
	.w4(32'h375dd6c5),
	.w5(32'h37863c1c),
	.w6(32'h36dccb94),
	.w7(32'h37dbb8fc),
	.w8(32'h374c9705),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d1b64),
	.w1(32'h381eb831),
	.w2(32'h37f0c209),
	.w3(32'hb8a5d0c0),
	.w4(32'hb8ae3195),
	.w5(32'hb85cd631),
	.w6(32'hb8c9b168),
	.w7(32'hb8ce76e1),
	.w8(32'hb8688e02),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d2cd7),
	.w1(32'hb8bcdc9d),
	.w2(32'hb853c96d),
	.w3(32'hb9474c7d),
	.w4(32'hb903528b),
	.w5(32'hb8b0188a),
	.w6(32'hb8ad0eb3),
	.w7(32'h3759be0b),
	.w8(32'h37128082),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6164928),
	.w1(32'h3533aca0),
	.w2(32'h37c99dc0),
	.w3(32'hb632507b),
	.w4(32'h36082f82),
	.w5(32'h37bb2673),
	.w6(32'h37455fe8),
	.w7(32'h3772c2bc),
	.w8(32'h37fd9cb9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bdb36e),
	.w1(32'h36919453),
	.w2(32'hb6a67ea0),
	.w3(32'h362d6758),
	.w4(32'hb6d34f1c),
	.w5(32'h35256457),
	.w6(32'h379a10a2),
	.w7(32'hb668bb5d),
	.w8(32'h36fb20bb),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7071dd5),
	.w1(32'hb76491c3),
	.w2(32'hb7cefc8f),
	.w3(32'h36948cf0),
	.w4(32'hb634948f),
	.w5(32'hb792bd68),
	.w6(32'hb7436e2c),
	.w7(32'hb6726c50),
	.w8(32'hb7b1d887),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h351209f5),
	.w1(32'h35122abb),
	.w2(32'hb638fefa),
	.w3(32'h3682136d),
	.w4(32'hb647cf56),
	.w5(32'hb6894bb2),
	.w6(32'h367fb845),
	.w7(32'hb6b9da11),
	.w8(32'hb6e618b1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e8db34),
	.w1(32'hb79655c9),
	.w2(32'h374b3b08),
	.w3(32'hb6a36db6),
	.w4(32'hb80fb168),
	.w5(32'h3745bc7d),
	.w6(32'hb719f71b),
	.w7(32'hb7a07f0f),
	.w8(32'h37ab2289),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7269247),
	.w1(32'hb7b1ede5),
	.w2(32'hb7b14e1e),
	.w3(32'h35f35287),
	.w4(32'hb647a3ad),
	.w5(32'hb74bdc37),
	.w6(32'hb789b8d6),
	.w7(32'hb580519b),
	.w8(32'h35a97953),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb817a5f6),
	.w1(32'hb721b963),
	.w2(32'hb7bb8373),
	.w3(32'hb82a68ce),
	.w4(32'h35e7d0fb),
	.w5(32'hb2703a1c),
	.w6(32'hb5a1fc88),
	.w7(32'h384745d0),
	.w8(32'h3781446f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a65342),
	.w1(32'hb640e763),
	.w2(32'hb76c88b5),
	.w3(32'hb7f1a897),
	.w4(32'hb7451f66),
	.w5(32'hb76cd614),
	.w6(32'hb7771e2a),
	.w7(32'h36965394),
	.w8(32'hb6c6b114),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82a5a01),
	.w1(32'hb85404b9),
	.w2(32'hb88bc16c),
	.w3(32'hb84b67e5),
	.w4(32'hb842aeff),
	.w5(32'hb881dc35),
	.w6(32'hb825b5cf),
	.w7(32'hb836a202),
	.w8(32'hb825abbc),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37da0d3a),
	.w1(32'h37e7e8c9),
	.w2(32'h37e1f5a9),
	.w3(32'h37befbff),
	.w4(32'h36c55b68),
	.w5(32'hb62d2a22),
	.w6(32'h36fd9995),
	.w7(32'hb7153f58),
	.w8(32'hb747c471),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3647c762),
	.w1(32'h36a3b916),
	.w2(32'h37119b50),
	.w3(32'h36b63579),
	.w4(32'hb3542dba),
	.w5(32'h360cd7df),
	.w6(32'hb4868a6a),
	.w7(32'h36c76027),
	.w8(32'h35d567b8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38478ecf),
	.w1(32'h37c7b08c),
	.w2(32'h37ca7257),
	.w3(32'h381dc61b),
	.w4(32'h37b34549),
	.w5(32'hb7534842),
	.w6(32'h37588c82),
	.w7(32'h36ba117c),
	.w8(32'hb8355167),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c51c44),
	.w1(32'h365d423f),
	.w2(32'h3702818d),
	.w3(32'h336f75da),
	.w4(32'hb648f97a),
	.w5(32'h35d32de0),
	.w6(32'h35c40ae3),
	.w7(32'h360bd90c),
	.w8(32'hb510a880),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81ed82b),
	.w1(32'hb802b710),
	.w2(32'hb8013cf5),
	.w3(32'hb7f3adb1),
	.w4(32'hb79c90b9),
	.w5(32'hb7ddaf23),
	.w6(32'hb77634a7),
	.w7(32'hb763d470),
	.w8(32'h3648ef2a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8784bc3),
	.w1(32'hb7da2df6),
	.w2(32'hb89d159d),
	.w3(32'hb7dae2b8),
	.w4(32'h372a991c),
	.w5(32'hb8061d55),
	.w6(32'hb6b7faa2),
	.w7(32'h38138755),
	.w8(32'hb6ccfc9b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8949c43),
	.w1(32'hb844ebae),
	.w2(32'hb89fde35),
	.w3(32'hb86b28d2),
	.w4(32'hb7e9d465),
	.w5(32'hb8477465),
	.w6(32'hb7f88ee4),
	.w7(32'h372967f6),
	.w8(32'hb7ecdd71),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb675c8c3),
	.w1(32'hb629ba52),
	.w2(32'hb77a6ada),
	.w3(32'hb6db107e),
	.w4(32'hb6ff0a33),
	.w5(32'hb76d3ef0),
	.w6(32'hb62c08ca),
	.w7(32'hb722eacb),
	.w8(32'hb705c9ac),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c3b179),
	.w1(32'hb88871f9),
	.w2(32'hb85c2052),
	.w3(32'hb887b7dd),
	.w4(32'hb7eb1ed8),
	.w5(32'hb820bb64),
	.w6(32'hb7cdd3fa),
	.w7(32'h376708d2),
	.w8(32'hb63bf610),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8496300),
	.w1(32'hb7d6e6b1),
	.w2(32'hb6ceaeb1),
	.w3(32'hb85561bb),
	.w4(32'hb73ca79b),
	.w5(32'hb79f8c39),
	.w6(32'hb7757210),
	.w7(32'h37a7b0ec),
	.w8(32'h339633f0),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d23cc9),
	.w1(32'h380aa414),
	.w2(32'h371c8f41),
	.w3(32'hb8831ecc),
	.w4(32'h36d69c38),
	.w5(32'hb6a85589),
	.w6(32'hb829b545),
	.w7(32'h35e99c58),
	.w8(32'hb6ac3cd6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c9ffa0),
	.w1(32'hb4621fe4),
	.w2(32'hb6956360),
	.w3(32'hb70e2ab0),
	.w4(32'h36a32bd3),
	.w5(32'h35ef0b8c),
	.w6(32'h3613d22f),
	.w7(32'h35de92f6),
	.w8(32'h350c86ef),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb573f97f),
	.w1(32'h356c2c09),
	.w2(32'h36960552),
	.w3(32'h36f078dd),
	.w4(32'h368136e5),
	.w5(32'h360a0ffd),
	.w6(32'h3615adfa),
	.w7(32'h36e7389e),
	.w8(32'h36c70eb1),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89144f1),
	.w1(32'hb8b6a673),
	.w2(32'hb8b291a0),
	.w3(32'hb87385d1),
	.w4(32'hb87e8662),
	.w5(32'hb82e8373),
	.w6(32'hb8725809),
	.w7(32'hb8715867),
	.w8(32'hb7e4e6e9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898ac2c),
	.w1(32'hb732a113),
	.w2(32'h374d9fea),
	.w3(32'hb79001ef),
	.w4(32'h36d6f8af),
	.w5(32'h37d31490),
	.w6(32'h36cf8d04),
	.w7(32'h3899626e),
	.w8(32'h38697702),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886f359),
	.w1(32'hb7566f74),
	.w2(32'hb86866fc),
	.w3(32'hb8a77db6),
	.w4(32'hb7d2c125),
	.w5(32'hb812288e),
	.w6(32'hb83014c4),
	.w7(32'hb6afa191),
	.w8(32'hb7a39ac7),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb811d149),
	.w1(32'hb8380f8d),
	.w2(32'hb7aee7b2),
	.w3(32'h372d14ae),
	.w4(32'hb8881392),
	.w5(32'hb82bf9ae),
	.w6(32'hb7499380),
	.w7(32'hb78561e9),
	.w8(32'h37a3eeb3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6995ff2),
	.w1(32'h35c59350),
	.w2(32'hb58ff2ae),
	.w3(32'h37675159),
	.w4(32'h366a6c14),
	.w5(32'hb5d0785f),
	.w6(32'h362616bb),
	.w7(32'h36eddaae),
	.w8(32'hb5a2230c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74f550e),
	.w1(32'hb6db2725),
	.w2(32'h35fe6e6d),
	.w3(32'hb74e08da),
	.w4(32'hb557e514),
	.w5(32'hb5720920),
	.w6(32'hb502e00b),
	.w7(32'h356fc009),
	.w8(32'hb6383610),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c5a9cb),
	.w1(32'h37611f6d),
	.w2(32'h39099cfa),
	.w3(32'h3862a18a),
	.w4(32'h37a72c4c),
	.w5(32'h38e86a57),
	.w6(32'h386b5a71),
	.w7(32'hb764f65c),
	.w8(32'h387a573d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a8aa98),
	.w1(32'h38547809),
	.w2(32'h380dc131),
	.w3(32'hb7861619),
	.w4(32'hb81b217b),
	.w5(32'hb818e06a),
	.w6(32'hb8091d09),
	.w7(32'hb89427cf),
	.w8(32'hb8440453),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a20bfc),
	.w1(32'h373d69f1),
	.w2(32'h384ac43f),
	.w3(32'h3897fe71),
	.w4(32'h36e72e36),
	.w5(32'h35e8f9a6),
	.w6(32'h38526d50),
	.w7(32'hb88d9788),
	.w8(32'hb797bc41),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88192cd),
	.w1(32'hb858a035),
	.w2(32'hb863fbee),
	.w3(32'hb7b8792d),
	.w4(32'hb5432913),
	.w5(32'h36c7bf93),
	.w6(32'hb72ad5b0),
	.w7(32'h37a45aad),
	.w8(32'h377f91ed),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bbb9b0),
	.w1(32'hb8352770),
	.w2(32'hb7eaf072),
	.w3(32'hb895a669),
	.w4(32'hb7967d79),
	.w5(32'hb7155418),
	.w6(32'hb788fde0),
	.w7(32'h382148ba),
	.w8(32'h37d707cb),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6aad58b),
	.w1(32'hb61f5447),
	.w2(32'h35bd72f3),
	.w3(32'hb71a3781),
	.w4(32'hb56750bb),
	.w5(32'hb43c4ea0),
	.w6(32'hb5f95226),
	.w7(32'hb6798ff1),
	.w8(32'hb5ab6fb3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362968f8),
	.w1(32'hb63f59e0),
	.w2(32'hb6321c75),
	.w3(32'hb57ffef6),
	.w4(32'hb71bd98e),
	.w5(32'hb43a4332),
	.w6(32'h3627ad22),
	.w7(32'h36c7622c),
	.w8(32'h362bbdf8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7899382),
	.w1(32'hb79bc9ce),
	.w2(32'hb72e96f4),
	.w3(32'hb7421503),
	.w4(32'hb710fec5),
	.w5(32'h36c84209),
	.w6(32'hb7063afd),
	.w7(32'hb632c11a),
	.w8(32'h3777019b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36916cbb),
	.w1(32'h3711c5b2),
	.w2(32'hb596d835),
	.w3(32'h36983b63),
	.w4(32'h35bc3ed3),
	.w5(32'hb68c09ac),
	.w6(32'h36555932),
	.w7(32'hb61503be),
	.w8(32'hb646fa24),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66bb421),
	.w1(32'h34992762),
	.w2(32'h3684b975),
	.w3(32'hb67c9297),
	.w4(32'h37a4e830),
	.w5(32'h3793977f),
	.w6(32'hb6066374),
	.w7(32'hb6bc95ff),
	.w8(32'h36e81d5b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8adaf54),
	.w1(32'hb7f53c07),
	.w2(32'hb6d696a7),
	.w3(32'hb88ad896),
	.w4(32'hb84d0ab5),
	.w5(32'hb7b174a8),
	.w6(32'hb7eb48d4),
	.w7(32'hb78067ec),
	.w8(32'h36be7bb1),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8357e46),
	.w1(32'hb81596cc),
	.w2(32'hb7c7cc3b),
	.w3(32'hb81ba46b),
	.w4(32'hb71671d7),
	.w5(32'h3719b76e),
	.w6(32'hb7cc2eb9),
	.w7(32'hb76cc15c),
	.w8(32'hb72af6ad),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70e6139),
	.w1(32'hb7243457),
	.w2(32'hb6a0b995),
	.w3(32'hb680b6aa),
	.w4(32'hb78409d6),
	.w5(32'h36e478a0),
	.w6(32'hb5e30430),
	.w7(32'h36fdb8f8),
	.w8(32'h3725ae57),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39054c59),
	.w1(32'h3888a409),
	.w2(32'h388d578c),
	.w3(32'h3915cee0),
	.w4(32'h382c9760),
	.w5(32'h3835e829),
	.w6(32'h3875a1af),
	.w7(32'hb8356d99),
	.w8(32'hb74704fc),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a54a8d),
	.w1(32'h37499668),
	.w2(32'h370884c3),
	.w3(32'hb6cb6b7f),
	.w4(32'h37440863),
	.w5(32'h367ae34c),
	.w6(32'h36c385ba),
	.w7(32'h378c9012),
	.w8(32'h36d09a88),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a4ff61),
	.w1(32'h349705c4),
	.w2(32'h36192e75),
	.w3(32'h335b8af6),
	.w4(32'hb652c52f),
	.w5(32'hb5c277c8),
	.w6(32'hb633b08f),
	.w7(32'h36259e99),
	.w8(32'hb61fb7cb),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb717d40c),
	.w1(32'h36c96c18),
	.w2(32'h36c75458),
	.w3(32'hb791c856),
	.w4(32'hb61906ab),
	.w5(32'hb703a9c2),
	.w6(32'hb6f21026),
	.w7(32'hb70daa24),
	.w8(32'h37056636),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ccd5b5),
	.w1(32'h36c693e7),
	.w2(32'hb5c2283c),
	.w3(32'h3711ee17),
	.w4(32'h374961d9),
	.w5(32'h36788770),
	.w6(32'hb61ca3bd),
	.w7(32'hb6cd3a1c),
	.w8(32'hb72d5375),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f204f4),
	.w1(32'h3742d218),
	.w2(32'h37293639),
	.w3(32'h3649bb09),
	.w4(32'h3750f265),
	.w5(32'h36c53f42),
	.w6(32'hb6f3dc9c),
	.w7(32'h367bc08a),
	.w8(32'h363e71e1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61de0ba),
	.w1(32'hb5084974),
	.w2(32'h35f0e304),
	.w3(32'hb6a37e26),
	.w4(32'hb670b720),
	.w5(32'hb5d3fe11),
	.w6(32'hb663b85c),
	.w7(32'h36331925),
	.w8(32'hb5f18daf),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361f7a4a),
	.w1(32'h35d7d0c2),
	.w2(32'h3637c67d),
	.w3(32'hb5689d45),
	.w4(32'h3401414c),
	.w5(32'h35d78b17),
	.w6(32'h3726048b),
	.w7(32'h36c95a66),
	.w8(32'h36acd6ec),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84e7387),
	.w1(32'hb82e02a8),
	.w2(32'hb7c860b7),
	.w3(32'hb7e03d3b),
	.w4(32'hb7ba2a85),
	.w5(32'h3584e851),
	.w6(32'hb82204f8),
	.w7(32'hb7343b0b),
	.w8(32'h35d354eb),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb881d680),
	.w1(32'hb65a018b),
	.w2(32'h3801cdfc),
	.w3(32'hb88389ae),
	.w4(32'hb817b50c),
	.w5(32'hb777e4bd),
	.w6(32'hb7c4124d),
	.w7(32'h37bfb93b),
	.w8(32'h38028932),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb831a0d8),
	.w1(32'hb74f6200),
	.w2(32'hb5d42b35),
	.w3(32'hb85b0987),
	.w4(32'hb816d0d4),
	.w5(32'hb7ca726f),
	.w6(32'hb84ca1b6),
	.w7(32'hb80f4056),
	.w8(32'hb7c89160),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8200d00),
	.w1(32'h3746b156),
	.w2(32'h376c8a7c),
	.w3(32'hb80f74f4),
	.w4(32'h36ef142b),
	.w5(32'h36e6a036),
	.w6(32'hb80f0871),
	.w7(32'hb70b9f14),
	.w8(32'h37be539f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a9363d),
	.w1(32'h368bf8ad),
	.w2(32'h35fec34b),
	.w3(32'hb52c86a1),
	.w4(32'h36ab5361),
	.w5(32'hb4ad9dbf),
	.w6(32'hb538dd22),
	.w7(32'h364df7a5),
	.w8(32'h36080823),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6229255),
	.w1(32'hb589c6c5),
	.w2(32'h346f8304),
	.w3(32'h33ba39cf),
	.w4(32'hb684d198),
	.w5(32'hb6460a9d),
	.w6(32'hb60f0893),
	.w7(32'h369d7cc4),
	.w8(32'hb6cd4c3e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bcf95b),
	.w1(32'hb687e37c),
	.w2(32'h366add52),
	.w3(32'hb7018964),
	.w4(32'hb6c412c2),
	.w5(32'hb57ce9f0),
	.w6(32'hb6b518d7),
	.w7(32'h35a6d425),
	.w8(32'hb5fbd929),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34bdecc9),
	.w1(32'h34d173cf),
	.w2(32'h363ad466),
	.w3(32'hb687efc0),
	.w4(32'hb60665ef),
	.w5(32'hb49a6fec),
	.w6(32'hb663b9b9),
	.w7(32'h35b56ec1),
	.w8(32'hb68cb90c),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b1e339),
	.w1(32'h378c12f4),
	.w2(32'hb6dbfe15),
	.w3(32'hb74889e0),
	.w4(32'hb7336492),
	.w5(32'hb7f64a42),
	.w6(32'hb82b9c59),
	.w7(32'hb82ce1f8),
	.w8(32'hb84bfc09),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb768b72d),
	.w1(32'hb80a50f1),
	.w2(32'hb7e955d9),
	.w3(32'hb74d7879),
	.w4(32'hb7ed5f3b),
	.w5(32'hb7122c60),
	.w6(32'hb7d84414),
	.w7(32'hb7d5e5bf),
	.w8(32'hb7af6109),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b13eb1),
	.w1(32'h37da9aba),
	.w2(32'hb77244c7),
	.w3(32'h37e45ee3),
	.w4(32'h37cbd347),
	.w5(32'hb714500c),
	.w6(32'h37189785),
	.w7(32'h3716cbbf),
	.w8(32'hb7a21733),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a6c705),
	.w1(32'h37ad822a),
	.w2(32'hb70c0638),
	.w3(32'h37e044f5),
	.w4(32'h377178dd),
	.w5(32'hb76a0a38),
	.w6(32'h379a022f),
	.w7(32'h3595290a),
	.w8(32'hb7ea91b0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360c9e1c),
	.w1(32'hb5a3b480),
	.w2(32'h3608ef91),
	.w3(32'h3586fcfd),
	.w4(32'hb68d6c8f),
	.w5(32'hb5059f00),
	.w6(32'hb6849348),
	.w7(32'h3673da29),
	.w8(32'h322ec299),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366e2347),
	.w1(32'hb5a8fc2d),
	.w2(32'hb70117c1),
	.w3(32'hb7267c97),
	.w4(32'hb7834777),
	.w5(32'hb6a8d004),
	.w6(32'hb68df5ef),
	.w7(32'hb72e69f6),
	.w8(32'hb74879c9),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3692cc02),
	.w1(32'h378196f0),
	.w2(32'h3760fc7b),
	.w3(32'h37c0855b),
	.w4(32'h37b41d54),
	.w5(32'h37057018),
	.w6(32'h3728f1c5),
	.w7(32'h3793d9e0),
	.w8(32'h37014e4c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b9b80d),
	.w1(32'h377cb8ce),
	.w2(32'h36203c7a),
	.w3(32'hb7d02dff),
	.w4(32'hb837e7e5),
	.w5(32'hb8b764a0),
	.w6(32'hb7d1e7db),
	.w7(32'hb8023dc9),
	.w8(32'hb899d6ed),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4852cb4),
	.w1(32'hba16aad9),
	.w2(32'h38fad112),
	.w3(32'hb6ba5b5b),
	.w4(32'hba0bec13),
	.w5(32'hb8700780),
	.w6(32'hba07fd5e),
	.w7(32'hb9410750),
	.w8(32'hb8ed4dec),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8be10a9),
	.w1(32'hb9ee3a79),
	.w2(32'hb9a6a06a),
	.w3(32'hb91c95de),
	.w4(32'hb9f52b1a),
	.w5(32'hb9b8b4fc),
	.w6(32'hb9b12453),
	.w7(32'hb9b73b71),
	.w8(32'hb96d8fb9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule