module layer_6_featuremap_46(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabba52c),
	.w1(32'h3a60c8e4),
	.w2(32'hbba2c12c),
	.w3(32'h3a17136d),
	.w4(32'hbbe52e4e),
	.w5(32'hbbf54c76),
	.w6(32'h3bf236bc),
	.w7(32'hbb11e355),
	.w8(32'hbc0b65e8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd2b82),
	.w1(32'h3b88f197),
	.w2(32'hbb52d4f9),
	.w3(32'h3c25cb86),
	.w4(32'hbac91eab),
	.w5(32'hbbe4f139),
	.w6(32'h3c66b9d6),
	.w7(32'h3bb1f75e),
	.w8(32'h3ae6d97a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaf8f9),
	.w1(32'h3c87e4a5),
	.w2(32'h3d61e48a),
	.w3(32'hbc8f5cb8),
	.w4(32'h3c8f8786),
	.w5(32'hbc047936),
	.w6(32'h3acb36b6),
	.w7(32'h3d8e802c),
	.w8(32'h39b08fde),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b11ec),
	.w1(32'hbae3f7d6),
	.w2(32'hbb858ba6),
	.w3(32'hbaa39dc6),
	.w4(32'hbb660c4f),
	.w5(32'hb9920c3e),
	.w6(32'hbab331c1),
	.w7(32'hbaac99fe),
	.w8(32'h3b1eb8c3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb705e461),
	.w1(32'hba7819ba),
	.w2(32'hbb746875),
	.w3(32'h3aee200a),
	.w4(32'h3b2238a6),
	.w5(32'hbc83656f),
	.w6(32'h3c2daf64),
	.w7(32'hbb021d73),
	.w8(32'hbcbc51e6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30feae),
	.w1(32'h3ad29a71),
	.w2(32'hbabd6dfd),
	.w3(32'h3adafb96),
	.w4(32'hbb087bd1),
	.w5(32'h3a27c518),
	.w6(32'h3b7af65a),
	.w7(32'hbb7c4c22),
	.w8(32'hb9dbea02),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d03f9),
	.w1(32'h3c0c087c),
	.w2(32'hbb900ee1),
	.w3(32'h3c1525c0),
	.w4(32'hba68ce0d),
	.w5(32'hbbcf72b7),
	.w6(32'h3c0331e8),
	.w7(32'hb912c980),
	.w8(32'hbbbe30b8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda9078),
	.w1(32'hbb40d5dd),
	.w2(32'h3bc94fb3),
	.w3(32'h3b4db6c0),
	.w4(32'h3c8fa34f),
	.w5(32'h3bd953ab),
	.w6(32'hbc10276f),
	.w7(32'hbb109f69),
	.w8(32'h3c990f84),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a914ba5),
	.w1(32'hb9070b0c),
	.w2(32'hbcd35bf3),
	.w3(32'h3cbc79ab),
	.w4(32'hbc384cc1),
	.w5(32'hbc962ed4),
	.w6(32'h3c67f9f6),
	.w7(32'hbd466d1e),
	.w8(32'hbd143ab3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96f322),
	.w1(32'h3af93400),
	.w2(32'h3ad0e384),
	.w3(32'hbb4b44af),
	.w4(32'hbb90f802),
	.w5(32'hba5a61bf),
	.w6(32'hb89bd91a),
	.w7(32'hb8f0c44e),
	.w8(32'h3b9a7d46),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6c865),
	.w1(32'hbbb35cb4),
	.w2(32'h3cbd9ee5),
	.w3(32'h3b04fd61),
	.w4(32'hbc8ccb06),
	.w5(32'h3b0eb964),
	.w6(32'h3b9ce08b),
	.w7(32'h3c4767cc),
	.w8(32'h3be43d7d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbeaebc),
	.w1(32'h3bbd66f2),
	.w2(32'h3b154527),
	.w3(32'hbaae6c42),
	.w4(32'hbb695d13),
	.w5(32'h3a348109),
	.w6(32'h3ad52fce),
	.w7(32'hba5a9eea),
	.w8(32'hbaaae8f3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ee630),
	.w1(32'h3afa2b55),
	.w2(32'hbc0fc065),
	.w3(32'h3bc783d3),
	.w4(32'hbbc07884),
	.w5(32'h3c03480b),
	.w6(32'h3b9f1214),
	.w7(32'hbbeab5b2),
	.w8(32'h3c2221a4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedbc1d),
	.w1(32'h3ca68c58),
	.w2(32'hbcd91382),
	.w3(32'h3ca6864f),
	.w4(32'h3c36dc61),
	.w5(32'hbbc7dce1),
	.w6(32'h3cf92afc),
	.w7(32'hbc37a041),
	.w8(32'hbccb7867),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd165932),
	.w1(32'hb9042c2c),
	.w2(32'hb94b1480),
	.w3(32'h3c0c722b),
	.w4(32'hb9c4ba11),
	.w5(32'hbb5fedd1),
	.w6(32'hbba0cc20),
	.w7(32'h3b396ae9),
	.w8(32'hbbd08a78),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba16d06),
	.w1(32'h3a7dcd4a),
	.w2(32'h38a8547c),
	.w3(32'hbb81dbb4),
	.w4(32'hbb929de6),
	.w5(32'hbb697466),
	.w6(32'hbb8e2531),
	.w7(32'hbb1f793f),
	.w8(32'hbafb223b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae56962),
	.w1(32'hbca902eb),
	.w2(32'hbc1dfec6),
	.w3(32'hbbb4e566),
	.w4(32'h3b9eac07),
	.w5(32'h3c7855df),
	.w6(32'hbc7164e0),
	.w7(32'h38e3a83e),
	.w8(32'h3c1346af),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c070bdf),
	.w1(32'hbad4e487),
	.w2(32'hbad54d4c),
	.w3(32'hb93230d0),
	.w4(32'hb94c2772),
	.w5(32'hba54869f),
	.w6(32'h3ae5ee10),
	.w7(32'h3b0e3207),
	.w8(32'h3b532495),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b8f58),
	.w1(32'hbbde0805),
	.w2(32'h39802a03),
	.w3(32'hbc0ceabb),
	.w4(32'hbb3c0689),
	.w5(32'h3ace7695),
	.w6(32'hbc0b4d05),
	.w7(32'hba1b7b5d),
	.w8(32'h3b90888d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0e93b),
	.w1(32'hbc9c774d),
	.w2(32'hbbdd7ef0),
	.w3(32'hbbdad3f0),
	.w4(32'h3c1c5690),
	.w5(32'h3ce4276b),
	.w6(32'hbc4b8525),
	.w7(32'h3c10a64f),
	.w8(32'h3cd169d3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c9d5a),
	.w1(32'h398ddb42),
	.w2(32'hbb05326b),
	.w3(32'h3a1ae588),
	.w4(32'h3af0bfab),
	.w5(32'hb9932cfd),
	.w6(32'hbb0a3e1d),
	.w7(32'h39d2d031),
	.w8(32'hba0b8304),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8676a),
	.w1(32'hbc46c74a),
	.w2(32'hbb0ffa4b),
	.w3(32'hbbc11dd1),
	.w4(32'hbbc6f238),
	.w5(32'hbc01dba8),
	.w6(32'hbbe27895),
	.w7(32'h3965140c),
	.w8(32'h3a4e501c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcad71),
	.w1(32'hbc5b0587),
	.w2(32'hbc466cf5),
	.w3(32'hbb69574f),
	.w4(32'hbc1185a7),
	.w5(32'h3c27b2c7),
	.w6(32'hbb23e0bc),
	.w7(32'hbcd3e6b3),
	.w8(32'h3c864fd0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17bbbf),
	.w1(32'h3c60dc3f),
	.w2(32'hbc054ded),
	.w3(32'h3cae9f73),
	.w4(32'h3c86b72b),
	.w5(32'h3b9d9abe),
	.w6(32'h3c77e90a),
	.w7(32'hbac45cf8),
	.w8(32'hbbdd945e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a489f),
	.w1(32'h3cd8f58b),
	.w2(32'hbca828f4),
	.w3(32'h3ce397f9),
	.w4(32'hbb83b3de),
	.w5(32'hbd58fecf),
	.w6(32'h3d51c6d8),
	.w7(32'h3a8f051d),
	.w8(32'hbd809512),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5c3bc4),
	.w1(32'hbc1dc2dc),
	.w2(32'h3c53db2d),
	.w3(32'hbc633734),
	.w4(32'hba43bcc4),
	.w5(32'h3c3dea6e),
	.w6(32'hbb061136),
	.w7(32'h3c92719e),
	.w8(32'h3c90f25b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c161d85),
	.w1(32'h3c1ed45d),
	.w2(32'hbc7a1e19),
	.w3(32'h3aa35d22),
	.w4(32'hbc6be1f6),
	.w5(32'hbc66c8c6),
	.w6(32'h3c3c07e4),
	.w7(32'hbc25af67),
	.w8(32'hbc9175b5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cca02),
	.w1(32'h3b183c3d),
	.w2(32'hbb74ecff),
	.w3(32'h3b93061f),
	.w4(32'h39ad7c2e),
	.w5(32'hbb068f17),
	.w6(32'h3b0ee518),
	.w7(32'hba38763d),
	.w8(32'hbaf239c4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3f9d7),
	.w1(32'hbb5cb12a),
	.w2(32'hba83f782),
	.w3(32'hbb00ba93),
	.w4(32'hba249a13),
	.w5(32'hbab64c5a),
	.w6(32'hbb4728a1),
	.w7(32'hbaf24b99),
	.w8(32'hbb498335),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf05cfd),
	.w1(32'hbbb2d5da),
	.w2(32'hbcdac3a2),
	.w3(32'h3ce043d6),
	.w4(32'h3c736e8b),
	.w5(32'hbcb993d7),
	.w6(32'h3c6e3ff3),
	.w7(32'hbb9d8230),
	.w8(32'hbca9a22a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce70980),
	.w1(32'h3c2da3e7),
	.w2(32'h3c22c67a),
	.w3(32'hbbb7029f),
	.w4(32'hbc42d31b),
	.w5(32'hba887c56),
	.w6(32'h3bb78656),
	.w7(32'hbc7c01d8),
	.w8(32'hbcd150ae),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d047c),
	.w1(32'h3cf5182a),
	.w2(32'h3c966944),
	.w3(32'hba8423c0),
	.w4(32'h3bb9544b),
	.w5(32'hbc4a47e8),
	.w6(32'h3c92d0aa),
	.w7(32'h3c2566e6),
	.w8(32'hbc536c3d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb13795),
	.w1(32'hbca01d8b),
	.w2(32'h3c507ad5),
	.w3(32'hbcd1cab9),
	.w4(32'h3c1256c3),
	.w5(32'h3ca51e4a),
	.w6(32'hbc372f76),
	.w7(32'h3d1a4017),
	.w8(32'h3d34350d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0b549e),
	.w1(32'hbb98bf02),
	.w2(32'hbc9d384e),
	.w3(32'h3c496e6c),
	.w4(32'h3cb5d3f5),
	.w5(32'h3bea12f7),
	.w6(32'h3c22b8ea),
	.w7(32'h3c8e336a),
	.w8(32'h3c900802),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a26c3),
	.w1(32'hbbd7f00e),
	.w2(32'hbb82ee3c),
	.w3(32'hbaa4f4d8),
	.w4(32'hbb138991),
	.w5(32'hba2727be),
	.w6(32'h3a552fd4),
	.w7(32'hbb0c460a),
	.w8(32'hb99fe2da),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7493f9),
	.w1(32'hbbbf3517),
	.w2(32'h3a88a490),
	.w3(32'hbbcc742d),
	.w4(32'h3bf5fc55),
	.w5(32'h3bbad4b2),
	.w6(32'h3a30059d),
	.w7(32'h3b3916ae),
	.w8(32'h3b104ab7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59693e),
	.w1(32'h390ef7c7),
	.w2(32'h3b8f6640),
	.w3(32'hbbf3921a),
	.w4(32'hbc01ec64),
	.w5(32'hbb8dbe50),
	.w6(32'hbad72c4a),
	.w7(32'hbb617e93),
	.w8(32'h3ad93f60),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8aeafd),
	.w1(32'hba905594),
	.w2(32'h3a5764f5),
	.w3(32'hb9adbae8),
	.w4(32'h3a1d920c),
	.w5(32'hbacb37eb),
	.w6(32'hbaaff2ce),
	.w7(32'h3ae6bbd2),
	.w8(32'hbb7fe6aa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb158c9a),
	.w1(32'h3cc2564c),
	.w2(32'h3c065666),
	.w3(32'h3cd69413),
	.w4(32'hbc48ae62),
	.w5(32'hbd0244a8),
	.w6(32'h3cdd1a98),
	.w7(32'hbb90894f),
	.w8(32'hbd08c4cf),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a8c42),
	.w1(32'h3c3b9479),
	.w2(32'h3c8073dd),
	.w3(32'hb839c1b7),
	.w4(32'h3c0f5d48),
	.w5(32'hbb5ba2fc),
	.w6(32'h3c9890a4),
	.w7(32'h3cceeafa),
	.w8(32'hbbc50d45),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa3a15),
	.w1(32'hbadf7764),
	.w2(32'h3be32075),
	.w3(32'hbb1a0605),
	.w4(32'hbc606387),
	.w5(32'h396496d6),
	.w6(32'h3b1b1b6d),
	.w7(32'hbb90c52e),
	.w8(32'h3c2ee303),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c859e1c),
	.w1(32'hbaa0d092),
	.w2(32'hbb7a5c94),
	.w3(32'hba326a18),
	.w4(32'hbab2a7ee),
	.w5(32'h3a4763c0),
	.w6(32'hba83d258),
	.w7(32'hba814e37),
	.w8(32'h3b0cc44d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab57661),
	.w1(32'hba9b59ec),
	.w2(32'h3ab8f6ed),
	.w3(32'hbb2e01e0),
	.w4(32'hbb85d40b),
	.w5(32'hbbdcc77c),
	.w6(32'h3b2741f6),
	.w7(32'h3a480221),
	.w8(32'hbba31134),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81e11f),
	.w1(32'h3bb6cb16),
	.w2(32'hbbbc9cc5),
	.w3(32'h3ad70a2d),
	.w4(32'hbb903993),
	.w5(32'hbc301715),
	.w6(32'h3c0fc644),
	.w7(32'hbc6602db),
	.w8(32'hbc8a3366),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf91d96),
	.w1(32'h3aca90ee),
	.w2(32'h3b5e500c),
	.w3(32'hbaa7e571),
	.w4(32'hbbb120e6),
	.w5(32'hbb41af35),
	.w6(32'h3a5e6e1b),
	.w7(32'hbb0bd4de),
	.w8(32'hbb4ceee7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7a12f),
	.w1(32'h3d4c7306),
	.w2(32'h3d414795),
	.w3(32'hbc3ebf03),
	.w4(32'hbd367a74),
	.w5(32'hbd3e448b),
	.w6(32'h3d020606),
	.w7(32'hbc011981),
	.w8(32'hbd01896d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12adde),
	.w1(32'hbb8cb816),
	.w2(32'hbbf5836e),
	.w3(32'hbb8673bf),
	.w4(32'hbbd2122b),
	.w5(32'h3c3e78a8),
	.w6(32'h39e139ae),
	.w7(32'hb95fca85),
	.w8(32'h3c648059),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b7a66),
	.w1(32'hbc95dceb),
	.w2(32'hbc0917e5),
	.w3(32'hbc807a55),
	.w4(32'h3b6233d1),
	.w5(32'h3c9b51ca),
	.w6(32'hb98a28f6),
	.w7(32'h3c7ee9ad),
	.w8(32'h3ca036a5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66f31b),
	.w1(32'h3a829418),
	.w2(32'hbacb7f5f),
	.w3(32'h3b9ca14f),
	.w4(32'h3aea49d1),
	.w5(32'h3b5853a6),
	.w6(32'h3b97ecd2),
	.w7(32'hbadc1a71),
	.w8(32'h3b0dae04),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab98640),
	.w1(32'h3bc15920),
	.w2(32'h3cb31f00),
	.w3(32'h3c0defe2),
	.w4(32'h3c79854d),
	.w5(32'h3ba64426),
	.w6(32'h3c53fe62),
	.w7(32'h3cef3ed2),
	.w8(32'h3b2b2af9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7baf0c),
	.w1(32'hbb6e22dc),
	.w2(32'hbc5668d5),
	.w3(32'h3b042002),
	.w4(32'hbbd4fb0f),
	.w5(32'hbad848b4),
	.w6(32'h3a1d1f4d),
	.w7(32'hbc19090b),
	.w8(32'hb878240a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb840e5a),
	.w1(32'hbc24b27d),
	.w2(32'hbc22b7a6),
	.w3(32'hbbad8963),
	.w4(32'hbbb2afc8),
	.w5(32'hbbc61355),
	.w6(32'hbbd77658),
	.w7(32'hbbde51d6),
	.w8(32'hbbca872f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee3a59),
	.w1(32'hbc1db43a),
	.w2(32'hbc0be96a),
	.w3(32'hbba98bc6),
	.w4(32'hbb60505f),
	.w5(32'hbb7b8022),
	.w6(32'hbc32c4f2),
	.w7(32'hbbbf45c4),
	.w8(32'hbb9e812d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd975b2),
	.w1(32'h3b76e048),
	.w2(32'hb7e94857),
	.w3(32'h3c5a9b72),
	.w4(32'h3c164d0e),
	.w5(32'hba9801d3),
	.w6(32'h3c2825c4),
	.w7(32'h3b511a34),
	.w8(32'hbbffd724),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f8f2a),
	.w1(32'hbad0d6c5),
	.w2(32'hbbca601d),
	.w3(32'hba5df422),
	.w4(32'hbb8e1038),
	.w5(32'hbb33d5c7),
	.w6(32'h3b134ede),
	.w7(32'hbb04348e),
	.w8(32'h3b0e2e92),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e0e4c),
	.w1(32'hbc4d36df),
	.w2(32'h3c2be013),
	.w3(32'h3c4a815b),
	.w4(32'hbb00fdba),
	.w5(32'hbcc677a1),
	.w6(32'h3a2b784d),
	.w7(32'hbc783c0f),
	.w8(32'hbb5d1dba),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a479a),
	.w1(32'h3b57c353),
	.w2(32'h3b54d0a3),
	.w3(32'h3b0de05c),
	.w4(32'h3aff8ce2),
	.w5(32'h3b820259),
	.w6(32'h3aa68afc),
	.w7(32'h3a8f5ecc),
	.w8(32'h3b0ed01d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf8afd),
	.w1(32'h3be1237b),
	.w2(32'h3c4b10c3),
	.w3(32'hbb764e37),
	.w4(32'hbb43972c),
	.w5(32'hbafcd420),
	.w6(32'hbb612145),
	.w7(32'h3bd12857),
	.w8(32'hbc130b22),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e94e5),
	.w1(32'hbac72e22),
	.w2(32'hba4994f0),
	.w3(32'hbb046aea),
	.w4(32'hbb3169eb),
	.w5(32'hbb62cb79),
	.w6(32'hba9d2222),
	.w7(32'hbac84f68),
	.w8(32'hbb48d588),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ec98e),
	.w1(32'hbbe1b684),
	.w2(32'h3b083b71),
	.w3(32'h3c8d2f46),
	.w4(32'hbbfb1bef),
	.w5(32'hbc61130b),
	.w6(32'hbbbc326f),
	.w7(32'hbba24613),
	.w8(32'h3b154b86),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b409b92),
	.w1(32'h3bd210a3),
	.w2(32'h3c81efc0),
	.w3(32'h3b9ee496),
	.w4(32'h3b0fc59f),
	.w5(32'hbb1b269d),
	.w6(32'h3c001ad3),
	.w7(32'h3c2454e0),
	.w8(32'h3ba5a7fe),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e8253),
	.w1(32'hbbb0e174),
	.w2(32'hbca3b4ab),
	.w3(32'h3c13716d),
	.w4(32'h3bb511b0),
	.w5(32'hbbbf1c5a),
	.w6(32'h3cc969b1),
	.w7(32'h3c3b522a),
	.w8(32'h3916100e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99af994),
	.w1(32'hbbc91768),
	.w2(32'hbc83e009),
	.w3(32'h3b748317),
	.w4(32'h3baae66b),
	.w5(32'h3ac9437b),
	.w6(32'hbb5dc93e),
	.w7(32'h39bbd9f1),
	.w8(32'h3b71d647),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e7d93),
	.w1(32'hba6387b4),
	.w2(32'hba576655),
	.w3(32'h3b14c065),
	.w4(32'h3b8b00e2),
	.w5(32'h3b970c72),
	.w6(32'hbb20779b),
	.w7(32'h395285c1),
	.w8(32'h3b1471fa),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule