module layer_8_featuremap_75(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcaca7),
	.w1(32'hbb286070),
	.w2(32'h3bb15927),
	.w3(32'hba14f4df),
	.w4(32'h39f57863),
	.w5(32'h3bc0dc62),
	.w6(32'h3acd5d19),
	.w7(32'h3a88f985),
	.w8(32'h3a8169ee),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8099be),
	.w1(32'h3960070b),
	.w2(32'h3a249b65),
	.w3(32'h39cccd41),
	.w4(32'hb62c937c),
	.w5(32'hbb081385),
	.w6(32'hba864f90),
	.w7(32'hba6cb255),
	.w8(32'hbb2ce265),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80e0604),
	.w1(32'h3a1511ef),
	.w2(32'h3a856f27),
	.w3(32'h3ac74295),
	.w4(32'h3a8309d9),
	.w5(32'hba857729),
	.w6(32'hba9f3095),
	.w7(32'hbb1898f5),
	.w8(32'hbb68f91b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4d163),
	.w1(32'hba8df979),
	.w2(32'h39a29a3e),
	.w3(32'hbbbe8101),
	.w4(32'h3a2cc74e),
	.w5(32'h3b27e9b4),
	.w6(32'hba2f60c9),
	.w7(32'hbb831240),
	.w8(32'hbb606388),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82e49b),
	.w1(32'hbaa9631d),
	.w2(32'hba256459),
	.w3(32'hbaed937d),
	.w4(32'hba31d80e),
	.w5(32'hba63ff2c),
	.w6(32'hba235711),
	.w7(32'hba8544a8),
	.w8(32'hba77d713),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba42262),
	.w1(32'h3b8320e8),
	.w2(32'hbbc6b312),
	.w3(32'hb78e2a14),
	.w4(32'hba8f448d),
	.w5(32'hbb98d5aa),
	.w6(32'hbab2a8f7),
	.w7(32'hbbf02cbe),
	.w8(32'hbbabd181),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae9dbe),
	.w1(32'hba00ba05),
	.w2(32'hb947b8b0),
	.w3(32'hb9884354),
	.w4(32'hb9a70760),
	.w5(32'hb9091410),
	.w6(32'hb9e80326),
	.w7(32'hb924d5c5),
	.w8(32'hb9360bdf),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93d6c1),
	.w1(32'hbb39ea4f),
	.w2(32'h3b8e6104),
	.w3(32'hbb331f0f),
	.w4(32'hbb264802),
	.w5(32'hb96b4d9e),
	.w6(32'hbabb84b0),
	.w7(32'hbb5e6276),
	.w8(32'hbb4b9d5d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad30e7e),
	.w1(32'hba8326cd),
	.w2(32'h3aa1adcc),
	.w3(32'hb86fc348),
	.w4(32'hb7f75c24),
	.w5(32'hbaa2a831),
	.w6(32'hba8527c6),
	.w7(32'hbad953c0),
	.w8(32'hbb240e27),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd3ca8),
	.w1(32'hbb2a5723),
	.w2(32'h3b97bfee),
	.w3(32'h3a0ff184),
	.w4(32'h38b2c033),
	.w5(32'hb94568fc),
	.w6(32'hba159749),
	.w7(32'h3aae6575),
	.w8(32'hbab5d243),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6abf48),
	.w1(32'h3a6db2ea),
	.w2(32'h3c046087),
	.w3(32'hbb776db8),
	.w4(32'h3aea3a7a),
	.w5(32'h3c35f463),
	.w6(32'h3a3e7319),
	.w7(32'hba2dd3a7),
	.w8(32'h3b160e0d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1d4f8),
	.w1(32'hbb978e23),
	.w2(32'h3aabd1d1),
	.w3(32'hb9395ef5),
	.w4(32'hbaf8f076),
	.w5(32'hbaa502a2),
	.w6(32'h3b853ce6),
	.w7(32'h3b23fe58),
	.w8(32'hbac2169c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9811e),
	.w1(32'h391e89c4),
	.w2(32'hb99ca810),
	.w3(32'h3b111bba),
	.w4(32'h3a2400e9),
	.w5(32'hbb35c872),
	.w6(32'h391fb233),
	.w7(32'h39fd4113),
	.w8(32'hbb1597fb),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4eae6),
	.w1(32'hbaf818ea),
	.w2(32'hbaca3b60),
	.w3(32'hb941a124),
	.w4(32'hbae8e75f),
	.w5(32'hbab7b0f8),
	.w6(32'hba96f087),
	.w7(32'hba6ad0ae),
	.w8(32'hb9c011eb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba100b37),
	.w1(32'hba79a102),
	.w2(32'hba50319b),
	.w3(32'hb9fa716d),
	.w4(32'hba6b5795),
	.w5(32'hba2ccac7),
	.w6(32'hba49393a),
	.w7(32'hba35483d),
	.w8(32'hb9305a92),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a99e42),
	.w1(32'hb98a2ba8),
	.w2(32'h391dbe33),
	.w3(32'h36c14e32),
	.w4(32'hb91d2587),
	.w5(32'h38e2975e),
	.w6(32'hb9dbaa49),
	.w7(32'hb917d484),
	.w8(32'h3a07cf09),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac6faf),
	.w1(32'hba662431),
	.w2(32'h3a583978),
	.w3(32'hb8c6d0fa),
	.w4(32'hbb36dd66),
	.w5(32'h39742af3),
	.w6(32'hba14cd74),
	.w7(32'hb9fb5d34),
	.w8(32'hba2dbe9b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe18b7a),
	.w1(32'hbb531a75),
	.w2(32'h3b31cbbe),
	.w3(32'h3aa36d02),
	.w4(32'hbace1811),
	.w5(32'hbab23ae4),
	.w6(32'h3ad89ead),
	.w7(32'h3a48b5a3),
	.w8(32'hbb36ba68),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd3038c),
	.w1(32'hbc25c037),
	.w2(32'h3c89eb78),
	.w3(32'hbc4f03d0),
	.w4(32'h3b0e529d),
	.w5(32'h3cca2316),
	.w6(32'h3c23ac12),
	.w7(32'h3b44c46c),
	.w8(32'hbbd90189),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f44a81),
	.w1(32'hba9118bd),
	.w2(32'h39191326),
	.w3(32'h3b50eaef),
	.w4(32'h3a2da618),
	.w5(32'hbad32c48),
	.w6(32'h3b36c00c),
	.w7(32'h3bb7d6c7),
	.w8(32'h3b9577e7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2e94f),
	.w1(32'h3b56ffa0),
	.w2(32'h3b417d89),
	.w3(32'h3bd46cea),
	.w4(32'h3ab2ff75),
	.w5(32'h3af6f1a5),
	.w6(32'h3be99be6),
	.w7(32'h3bc429cd),
	.w8(32'h39ad2c9c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9e1c2),
	.w1(32'h3b33e80c),
	.w2(32'h3ab738ae),
	.w3(32'h3b2d4f54),
	.w4(32'h3adb85bd),
	.w5(32'hba9826e3),
	.w6(32'hb950e5c8),
	.w7(32'hbaa059b0),
	.w8(32'h39f48150),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb684498),
	.w1(32'hbb8ce374),
	.w2(32'h3c8ebd56),
	.w3(32'h3bc5ae2c),
	.w4(32'h3b9f22c6),
	.w5(32'h3cc8fca4),
	.w6(32'h3c4966b2),
	.w7(32'h3c475f90),
	.w8(32'h3c05ef50),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac4cb5),
	.w1(32'h3b5c9a73),
	.w2(32'h3a3b3ed8),
	.w3(32'h3ba830f6),
	.w4(32'h3b21041c),
	.w5(32'hba0f2506),
	.w6(32'h3b11f591),
	.w7(32'h3a3beec8),
	.w8(32'h3afe61ea),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44e4a3),
	.w1(32'h3a066f45),
	.w2(32'h3a973c6c),
	.w3(32'h3ac213ea),
	.w4(32'h3a7669cc),
	.w5(32'h3ab5a961),
	.w6(32'h3a24e6c1),
	.w7(32'h3aa9733f),
	.w8(32'h3b4346b6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b86a5),
	.w1(32'hbb74f41e),
	.w2(32'h3b019420),
	.w3(32'h3b804df9),
	.w4(32'h391b2f80),
	.w5(32'h3bd5851c),
	.w6(32'h3c16f477),
	.w7(32'h3b88ec91),
	.w8(32'h3affdaa6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee27f3),
	.w1(32'h3a54631a),
	.w2(32'h3a65d20b),
	.w3(32'h3af89a65),
	.w4(32'h3a474d3e),
	.w5(32'h3a4510d2),
	.w6(32'h3aac2ac2),
	.w7(32'h3ac26ba0),
	.w8(32'h39bd611d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd399e05),
	.w1(32'hbd90b8e3),
	.w2(32'h3b2539a2),
	.w3(32'hbd3011ff),
	.w4(32'hbd9a04b1),
	.w5(32'h3cdd62a2),
	.w6(32'h3cd57a7c),
	.w7(32'h3c6939d9),
	.w8(32'hbd51bb3b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e9aa0),
	.w1(32'hbb2bcf2a),
	.w2(32'h3b2c72d1),
	.w3(32'hba588f29),
	.w4(32'hba8acaba),
	.w5(32'h3b3ee610),
	.w6(32'h3b593d52),
	.w7(32'h3b904b6b),
	.w8(32'h3ae38d27),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b652e),
	.w1(32'hba42246e),
	.w2(32'hb9b2c914),
	.w3(32'hba2928a3),
	.w4(32'hba51b49c),
	.w5(32'hba2f07f9),
	.w6(32'hba1809f0),
	.w7(32'hba84d895),
	.w8(32'hba8ece52),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f893e9),
	.w1(32'hba24d2f2),
	.w2(32'h397694ec),
	.w3(32'hb8692b7b),
	.w4(32'hba3f4e07),
	.w5(32'h3a2321ea),
	.w6(32'h388e1535),
	.w7(32'hba669907),
	.w8(32'h39dcb2ea),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5f105),
	.w1(32'h3b402d11),
	.w2(32'h3a73fc58),
	.w3(32'h3b1ea7b8),
	.w4(32'h39058ac5),
	.w5(32'hbacce176),
	.w6(32'h3ad0c5fe),
	.w7(32'h3984df7b),
	.w8(32'hbb7ec151),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92b26d0),
	.w1(32'h39594cea),
	.w2(32'hb999e199),
	.w3(32'hb8fdfd0f),
	.w4(32'hb89c49c0),
	.w5(32'hb8c60751),
	.w6(32'hb985760c),
	.w7(32'hb9fbca86),
	.w8(32'h39a5f476),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b3623),
	.w1(32'hb9a10ffa),
	.w2(32'hb968872f),
	.w3(32'h39ba51d6),
	.w4(32'hb85944b4),
	.w5(32'hb936ae4f),
	.w6(32'h39dfdaae),
	.w7(32'hb9250b12),
	.w8(32'h3a01bc0d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a3d0e),
	.w1(32'h3adb93f6),
	.w2(32'hba928e28),
	.w3(32'h3bbd2509),
	.w4(32'h3b011ac3),
	.w5(32'hbb54183d),
	.w6(32'hbb626ddb),
	.w7(32'hba164906),
	.w8(32'hb9845cfe),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc9e1b),
	.w1(32'hbbcf053b),
	.w2(32'h3b7d9374),
	.w3(32'hbb9de2c1),
	.w4(32'hbb1a2333),
	.w5(32'h3b5fbd58),
	.w6(32'h39999c88),
	.w7(32'h3b395b8b),
	.w8(32'h3ac4c2fd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1c3ab),
	.w1(32'h3a88bbbe),
	.w2(32'h3ab25dd4),
	.w3(32'h3ae68280),
	.w4(32'h3ac81e5c),
	.w5(32'h3a97e4fa),
	.w6(32'h3aa83c3e),
	.w7(32'h3acd7567),
	.w8(32'hb9bfdb78),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39456e1b),
	.w1(32'h3ab1f7ca),
	.w2(32'h3b411e4e),
	.w3(32'h3946baf5),
	.w4(32'h3a44f511),
	.w5(32'h3abfe55f),
	.w6(32'h3a8a4586),
	.w7(32'h3a7917fc),
	.w8(32'hb767833d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88dd25),
	.w1(32'hbac757ad),
	.w2(32'hbab2cf9e),
	.w3(32'hba686ca8),
	.w4(32'hbac0f06b),
	.w5(32'hba8e150f),
	.w6(32'hbab68cde),
	.w7(32'hbaa712a8),
	.w8(32'h3a2b5355),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8b47f),
	.w1(32'hb6faed8d),
	.w2(32'h3aa7f8f1),
	.w3(32'h3aafb90e),
	.w4(32'h3a4163ec),
	.w5(32'h3b00d0ff),
	.w6(32'h394a87a9),
	.w7(32'h39b3d4da),
	.w8(32'h3aa2b824),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabe637),
	.w1(32'hba9cf33b),
	.w2(32'h3be3ff56),
	.w3(32'h3ae119e7),
	.w4(32'h3b943cbc),
	.w5(32'h3ba04814),
	.w6(32'h3c6027d5),
	.w7(32'h3c00683f),
	.w8(32'hbc5f0672),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb909fc9),
	.w1(32'hbb36edc0),
	.w2(32'h3984a469),
	.w3(32'h3b011fd9),
	.w4(32'hbb8e619b),
	.w5(32'h3b2721e6),
	.w6(32'hbb9a27df),
	.w7(32'hbbbd338f),
	.w8(32'hbc1ef70c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44ca0f),
	.w1(32'hbc9156e5),
	.w2(32'h3b6a707e),
	.w3(32'h3c3e984e),
	.w4(32'h3d20941e),
	.w5(32'hbc6a02ac),
	.w6(32'hbcc4d5be),
	.w7(32'h3c868131),
	.w8(32'h39e9132f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a20a8),
	.w1(32'hbb2862b6),
	.w2(32'h3b7c2c9a),
	.w3(32'hba9b9aa9),
	.w4(32'hbc51f71f),
	.w5(32'h3afcd087),
	.w6(32'h3c441ad7),
	.w7(32'h3b094ec4),
	.w8(32'hbb2058f0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5b92d),
	.w1(32'hbc1360cc),
	.w2(32'h3bc05dba),
	.w3(32'h3ac1001e),
	.w4(32'hbb360b11),
	.w5(32'h3c88605d),
	.w6(32'h3aa766c3),
	.w7(32'hbb61616c),
	.w8(32'hbc7543cf),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc325df9),
	.w1(32'hbc8ed438),
	.w2(32'hbbf9aad1),
	.w3(32'h3b24337f),
	.w4(32'hbbb2db8a),
	.w5(32'h3b859776),
	.w6(32'hbc8ead6f),
	.w7(32'hbc5c5ae5),
	.w8(32'hbcea560b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0252f7),
	.w1(32'h3bace355),
	.w2(32'hbd2fe43a),
	.w3(32'hbc8d55c0),
	.w4(32'hbc756adf),
	.w5(32'hbc1c8fc6),
	.w6(32'hbd0e4dd2),
	.w7(32'hbce590ad),
	.w8(32'h3a9a811e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0aae3),
	.w1(32'hbc7b626b),
	.w2(32'hbbc36bad),
	.w3(32'h3b4b83e6),
	.w4(32'hbbe1d22d),
	.w5(32'h3c028a46),
	.w6(32'h3b51615c),
	.w7(32'hbc8094d4),
	.w8(32'hbc967d6e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d2cd3),
	.w1(32'h39c8c1d0),
	.w2(32'hbac7f6a6),
	.w3(32'h3c104d3f),
	.w4(32'h3d3b08d4),
	.w5(32'h3c96e6bf),
	.w6(32'hbccdb956),
	.w7(32'hbba02e52),
	.w8(32'hbc153e19),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd99427),
	.w1(32'hbbd293c7),
	.w2(32'h3b84410e),
	.w3(32'h3b014fa8),
	.w4(32'hbb992d7f),
	.w5(32'h3c3ac72d),
	.w6(32'h3ad8bf08),
	.w7(32'hbbb50a9b),
	.w8(32'hba815a49),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c562f85),
	.w1(32'h3bb32bcf),
	.w2(32'hba23586b),
	.w3(32'h3c2ad964),
	.w4(32'hbb3cb843),
	.w5(32'hbc2581e3),
	.w6(32'h3c72693d),
	.w7(32'h3be26a4a),
	.w8(32'hbbb9f601),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c5d04),
	.w1(32'hbc1f8773),
	.w2(32'h3c36b757),
	.w3(32'hbca02342),
	.w4(32'hbc83b088),
	.w5(32'h3c8653d9),
	.w6(32'h3c79ca82),
	.w7(32'h3b105d28),
	.w8(32'h3bcb7d52),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5771f8),
	.w1(32'hbc1fac41),
	.w2(32'h3b616b7e),
	.w3(32'hbb9621b8),
	.w4(32'h3cc006bf),
	.w5(32'h3cbcdffb),
	.w6(32'hbc22fb53),
	.w7(32'hbc54bc2c),
	.w8(32'hbc811586),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16dc51),
	.w1(32'hba316ddc),
	.w2(32'h3bd19c02),
	.w3(32'h3c09c301),
	.w4(32'h3d0b2b22),
	.w5(32'h3ca8505a),
	.w6(32'hbcc668d9),
	.w7(32'hbbb9229a),
	.w8(32'hbbeea5cb),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77aa4d),
	.w1(32'hbc1eb421),
	.w2(32'hbb680332),
	.w3(32'h3c613a5d),
	.w4(32'hba1fb759),
	.w5(32'hbbabd8c0),
	.w6(32'hbc370953),
	.w7(32'h3c3883d5),
	.w8(32'h3c0e971f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52b96b),
	.w1(32'hbb9c6c11),
	.w2(32'h3c327a8c),
	.w3(32'h3c04bd44),
	.w4(32'hbc0da44a),
	.w5(32'h3c7e6f53),
	.w6(32'h3ca0325e),
	.w7(32'h3c8e79fb),
	.w8(32'hbc6e2d0b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f43fe),
	.w1(32'h3bc2a650),
	.w2(32'h3c192719),
	.w3(32'hbbfa716e),
	.w4(32'hbc4bd8d1),
	.w5(32'h3c20e80b),
	.w6(32'h3b957133),
	.w7(32'hbbbdd39d),
	.w8(32'hbbfaf272),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a2283),
	.w1(32'hba3d8524),
	.w2(32'hba4d0a33),
	.w3(32'hbc2e0a7c),
	.w4(32'h3d0945b5),
	.w5(32'hbb8558db),
	.w6(32'h3ce045c8),
	.w7(32'hbb515cef),
	.w8(32'h3c065c36),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f5308),
	.w1(32'hbc6c53e7),
	.w2(32'hbc48f54f),
	.w3(32'hbbc0cf27),
	.w4(32'hbaafca0a),
	.w5(32'h3b9bdafd),
	.w6(32'h3c9a17ac),
	.w7(32'h3bdf6e4a),
	.w8(32'hbbe66751),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb3b56),
	.w1(32'h3bcec43f),
	.w2(32'hbbf55c9e),
	.w3(32'hbaf11576),
	.w4(32'h3ca6c3bd),
	.w5(32'hb9fb782e),
	.w6(32'hbcfdbfe6),
	.w7(32'hbbb627da),
	.w8(32'h3be37b96),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8387ad),
	.w1(32'h3bd0e6dd),
	.w2(32'hbbdae93c),
	.w3(32'h3c593fc7),
	.w4(32'h3a4d8cd8),
	.w5(32'hbcabba7f),
	.w6(32'hbc9a1552),
	.w7(32'hbc53b9ce),
	.w8(32'hbc387ce2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22dbb2),
	.w1(32'hbc16a834),
	.w2(32'hba97ff0e),
	.w3(32'h3c083a16),
	.w4(32'h3b2af78f),
	.w5(32'h3c628b71),
	.w6(32'hbc83e493),
	.w7(32'hbc42a0c5),
	.w8(32'hbaa19599),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2691b4),
	.w1(32'hba03a38f),
	.w2(32'h3c1dcd47),
	.w3(32'h3a8abfb8),
	.w4(32'hbc2eb5f9),
	.w5(32'hb9194448),
	.w6(32'h3c42933e),
	.w7(32'h3c1d7f27),
	.w8(32'hbc8c97bf),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d6ff8),
	.w1(32'h3b2675d5),
	.w2(32'hba929d8b),
	.w3(32'hbb1a9dd2),
	.w4(32'h3c153bfe),
	.w5(32'h3c472d8e),
	.w6(32'h3c55ab07),
	.w7(32'h3b5007be),
	.w8(32'hbb2e7d89),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68b497),
	.w1(32'h3b4ed53f),
	.w2(32'h3bb2b510),
	.w3(32'h3b9a0665),
	.w4(32'hbb254d1d),
	.w5(32'h3b8dd123),
	.w6(32'h3b90f9cc),
	.w7(32'h3a2d19e6),
	.w8(32'h3a901df6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02d886),
	.w1(32'hbb2c7b41),
	.w2(32'h3af15742),
	.w3(32'hb99547c0),
	.w4(32'hbbd39233),
	.w5(32'h3a664984),
	.w6(32'h3bd215fd),
	.w7(32'h3a69bbb1),
	.w8(32'hbb3d1aa2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e36cf),
	.w1(32'hba76f46a),
	.w2(32'hba96d296),
	.w3(32'hb8c71f66),
	.w4(32'hbb8c49dc),
	.w5(32'hba9d161c),
	.w6(32'h3ac0fd8c),
	.w7(32'hbb2cf481),
	.w8(32'hbc8f5c4a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce8ecf6),
	.w1(32'hbc5a58be),
	.w2(32'hbc971bf4),
	.w3(32'h3b69f18b),
	.w4(32'h37b8b1e1),
	.w5(32'h3c08c336),
	.w6(32'h38d0793b),
	.w7(32'hbc9496ed),
	.w8(32'hbc28a19f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f4ecfa),
	.w1(32'hbb4d536b),
	.w2(32'h39f93a1a),
	.w3(32'h3bab52d7),
	.w4(32'hbb680fc6),
	.w5(32'h3b8fd323),
	.w6(32'hbae3626b),
	.w7(32'hbb87082f),
	.w8(32'h3d0fe290),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15b578),
	.w1(32'hbca8cc19),
	.w2(32'hbbc00cb0),
	.w3(32'hbccddf39),
	.w4(32'hbd5936b9),
	.w5(32'h3b20daf4),
	.w6(32'h3d6c82ba),
	.w7(32'h3ca77830),
	.w8(32'hba883d03),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cbfd9),
	.w1(32'hbafaa5ab),
	.w2(32'hb9d721dd),
	.w3(32'h3b87569e),
	.w4(32'hbba0964f),
	.w5(32'h3a68a3a5),
	.w6(32'hbb5a05de),
	.w7(32'hbb93a84d),
	.w8(32'hbbfa3419),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1354da),
	.w1(32'hbaa0c14d),
	.w2(32'h3ab8ff60),
	.w3(32'h3bb9e4c5),
	.w4(32'hbb884f77),
	.w5(32'h3bc6aa85),
	.w6(32'hba81f37b),
	.w7(32'hbb42c1ca),
	.w8(32'hbba46b51),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac20584),
	.w1(32'hbb15cfb1),
	.w2(32'hba21c3d9),
	.w3(32'h3b9dcd46),
	.w4(32'hbba9ea9e),
	.w5(32'h3b21f7c1),
	.w6(32'hbb9f474c),
	.w7(32'hbba46244),
	.w8(32'hbce7de77),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca063d0),
	.w1(32'hbc254628),
	.w2(32'hbb0ecc50),
	.w3(32'hbc86935b),
	.w4(32'hbcef2788),
	.w5(32'hbab00fa7),
	.w6(32'hbd02d56b),
	.w7(32'hbc540f5c),
	.w8(32'hbc6b2877),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4db89),
	.w1(32'hbb7e4daf),
	.w2(32'hbb588e23),
	.w3(32'h3bcc2f6f),
	.w4(32'h3aeedbd9),
	.w5(32'h3b6b38a2),
	.w6(32'hbc0f72ce),
	.w7(32'hbc1db318),
	.w8(32'hbaf9efc8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3bbc4),
	.w1(32'hbb108e67),
	.w2(32'h3b06ed41),
	.w3(32'hba9c9d30),
	.w4(32'hbbf6785b),
	.w5(32'h3ae8f8ff),
	.w6(32'h3b9490a6),
	.w7(32'h3af8b187),
	.w8(32'hbbf181ad),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ec5a7),
	.w1(32'hbb888dfa),
	.w2(32'hb9eb473c),
	.w3(32'h3b55bb51),
	.w4(32'hbb15cb44),
	.w5(32'h3b791928),
	.w6(32'hbbe3c72e),
	.w7(32'hbba6f820),
	.w8(32'h3d24ce75),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc295c1c),
	.w1(32'hbc6ad599),
	.w2(32'hbc52d79f),
	.w3(32'hbc9102dc),
	.w4(32'hbd480604),
	.w5(32'hbc542f39),
	.w6(32'h3d9e9231),
	.w7(32'h3cd30081),
	.w8(32'h3c8c0c46),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0c73c),
	.w1(32'hbc335e79),
	.w2(32'hbc04e355),
	.w3(32'hbc52be4f),
	.w4(32'hbd2f3cc2),
	.w5(32'hbc9fa5a4),
	.w6(32'h3d1712a9),
	.w7(32'h3bdef76f),
	.w8(32'hb99486ce),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7258a),
	.w1(32'hbb73ed7d),
	.w2(32'h3b9e5579),
	.w3(32'h3b3f3835),
	.w4(32'hba8d3810),
	.w5(32'h3badb224),
	.w6(32'h3c0815d6),
	.w7(32'h3ad9876a),
	.w8(32'hbc0105a0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7036b),
	.w1(32'h3c66a4d0),
	.w2(32'hbb4cf003),
	.w3(32'hbc7815f0),
	.w4(32'h3ba08012),
	.w5(32'hba41fc31),
	.w6(32'hbbab3d95),
	.w7(32'hba0fb0d9),
	.w8(32'hbbf445ed),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80d507),
	.w1(32'h3b30b088),
	.w2(32'h3ba09b84),
	.w3(32'h3b8a620b),
	.w4(32'h3acfbd42),
	.w5(32'h3c7b3d2e),
	.w6(32'hbc3fc297),
	.w7(32'hbc2b8c11),
	.w8(32'hbc05c88c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f2742),
	.w1(32'hbbaf2bcc),
	.w2(32'h3c1a0077),
	.w3(32'h3c0206ae),
	.w4(32'h3b6ee57a),
	.w5(32'h3cc55de6),
	.w6(32'hbb712aea),
	.w7(32'hba8c8f36),
	.w8(32'hbc10cb0f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc317b5),
	.w1(32'hbc168265),
	.w2(32'hbc32df09),
	.w3(32'hbc9f7108),
	.w4(32'h3cd84eda),
	.w5(32'hba93f5ab),
	.w6(32'hbc9a3db3),
	.w7(32'h389deeea),
	.w8(32'hbc6f0aba),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1526c7),
	.w1(32'hbb0d812e),
	.w2(32'h3c700d48),
	.w3(32'h3b7fd44c),
	.w4(32'h3cba0246),
	.w5(32'h3cbc56e4),
	.w6(32'hbbc7aa74),
	.w7(32'hb97d617f),
	.w8(32'hbb4db46b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0afb22),
	.w1(32'h3a1e6f42),
	.w2(32'h3b40ba2a),
	.w3(32'h3b17d91e),
	.w4(32'hbbc06bc2),
	.w5(32'h3c617ffd),
	.w6(32'h37c53bf6),
	.w7(32'hbbee4244),
	.w8(32'hbc67a669),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca117fe),
	.w1(32'hb97b8df1),
	.w2(32'hbb61990c),
	.w3(32'h3c353e13),
	.w4(32'h3d775627),
	.w5(32'h3cc839e1),
	.w6(32'hbd03e9bd),
	.w7(32'hbbb9c1a0),
	.w8(32'hbc0eed66),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f595c),
	.w1(32'hbb5abeeb),
	.w2(32'h3bad287f),
	.w3(32'h3a71b65c),
	.w4(32'hbba888b3),
	.w5(32'h3c790398),
	.w6(32'h3b3bbdb5),
	.w7(32'hbb9e62d8),
	.w8(32'hbb72aeac),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc152d54),
	.w1(32'h3aac3a73),
	.w2(32'hbb987e78),
	.w3(32'hbb5dc1b0),
	.w4(32'h3cf329f8),
	.w5(32'h3b91bb60),
	.w6(32'hbcb83b9f),
	.w7(32'hbc217b7d),
	.w8(32'hbca698a4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89e014),
	.w1(32'hb93060b0),
	.w2(32'hbb32be18),
	.w3(32'h3c21a1c6),
	.w4(32'h3d6520d2),
	.w5(32'h3cbbe1d9),
	.w6(32'hbcf06faa),
	.w7(32'hbba0e4a5),
	.w8(32'hbc854183),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8240a7),
	.w1(32'hbadbcfb2),
	.w2(32'hbb86e36e),
	.w3(32'h3c1a1b7b),
	.w4(32'h3d425d58),
	.w5(32'h3ca06f79),
	.w6(32'hbccb4b4f),
	.w7(32'hbba17279),
	.w8(32'hbc7e1299),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5751b6),
	.w1(32'h3adaa79f),
	.w2(32'hbb86fced),
	.w3(32'h3bca63b5),
	.w4(32'h3c9d6df2),
	.w5(32'h3aaa9cb4),
	.w6(32'hbca2ff76),
	.w7(32'hbc20081d),
	.w8(32'h3c5eeb0d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be10ce8),
	.w1(32'hbbb0ca6e),
	.w2(32'h3ccbc741),
	.w3(32'h3b4efa5c),
	.w4(32'h3b882c8b),
	.w5(32'h3d03ee8c),
	.w6(32'h3c8382d2),
	.w7(32'hbc314c4c),
	.w8(32'h3b036367),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a486d33),
	.w1(32'hb96afcd6),
	.w2(32'h3b3e4f78),
	.w3(32'hba44c9cb),
	.w4(32'hbba5ee57),
	.w5(32'h39f35f2b),
	.w6(32'h3ba8fb23),
	.w7(32'h3acc179b),
	.w8(32'hbc9282d2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bc9f5),
	.w1(32'h38af244f),
	.w2(32'hbc587c84),
	.w3(32'hbc5efd77),
	.w4(32'hb73a5573),
	.w5(32'hbb174ea9),
	.w6(32'hbc5fb9c3),
	.w7(32'hbc9d72bb),
	.w8(32'hbd0822f5),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49df09),
	.w1(32'h3c2f2135),
	.w2(32'h3cac1ed7),
	.w3(32'h3c08d024),
	.w4(32'h3d170cd5),
	.w5(32'h3c8df2cc),
	.w6(32'hbd0b5133),
	.w7(32'h391e8605),
	.w8(32'hbb52f9e0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82fff0),
	.w1(32'hba534802),
	.w2(32'hbbbfb9a6),
	.w3(32'hbc22143e),
	.w4(32'hba85b2c9),
	.w5(32'h3b771991),
	.w6(32'h3c838028),
	.w7(32'hbc63994f),
	.w8(32'h3b9a81e5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc024519),
	.w1(32'h3c51a1a7),
	.w2(32'hbb312934),
	.w3(32'hb8ed0e2e),
	.w4(32'hbbd095b3),
	.w5(32'h3c0fb79e),
	.w6(32'hbc2a34f0),
	.w7(32'h3ab1cec9),
	.w8(32'h3d107ce6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeb35c),
	.w1(32'hbc2e99ed),
	.w2(32'hbc87205c),
	.w3(32'hbc5263d9),
	.w4(32'hbd313e1f),
	.w5(32'hbc9c7fad),
	.w6(32'h3d805bce),
	.w7(32'h3c91b96f),
	.w8(32'hbbb9ba61),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb096fc1),
	.w1(32'hbb626c2b),
	.w2(32'h3b8e7fcb),
	.w3(32'h3ba2c75f),
	.w4(32'hbb96074d),
	.w5(32'h3c4e91d6),
	.w6(32'h39f54581),
	.w7(32'hbb4cea3e),
	.w8(32'hbcb66697),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a426a),
	.w1(32'h3c0a2abb),
	.w2(32'hbb921e38),
	.w3(32'h3ba21c7f),
	.w4(32'h3ce4f585),
	.w5(32'h3ab86570),
	.w6(32'hbce8311a),
	.w7(32'hbbb4d574),
	.w8(32'h39fe4842),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c023b),
	.w1(32'h3a561713),
	.w2(32'h3b63f695),
	.w3(32'h3ac16f6c),
	.w4(32'hbb96d7a0),
	.w5(32'h3a34c700),
	.w6(32'h3b218775),
	.w7(32'hb879eb43),
	.w8(32'h3ce29470),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba496496),
	.w1(32'hbc2308da),
	.w2(32'hbc87e16f),
	.w3(32'hbc8d4552),
	.w4(32'hbd9a7153),
	.w5(32'hbd1315fe),
	.w6(32'h3d96ae60),
	.w7(32'h3c812b9b),
	.w8(32'hbca029fe),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd7fe2),
	.w1(32'h3c288a39),
	.w2(32'hba80e3a7),
	.w3(32'h3bcd8274),
	.w4(32'h3cd910b1),
	.w5(32'h3be1ed91),
	.w6(32'hbcc9e38c),
	.w7(32'hbc1b6f8a),
	.w8(32'hbbb3fdc8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89baf7),
	.w1(32'h3b0d1fa1),
	.w2(32'h39bff717),
	.w3(32'h3bd89c08),
	.w4(32'h3cc6c917),
	.w5(32'h3c1bd52b),
	.w6(32'hbc6e5499),
	.w7(32'hbb681842),
	.w8(32'h3a1655df),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1be8bd),
	.w1(32'hbc14e660),
	.w2(32'h3a20eef9),
	.w3(32'hbc6d6b87),
	.w4(32'hbc01fdbf),
	.w5(32'h3b8c6589),
	.w6(32'hbb8a1106),
	.w7(32'hbb3c829c),
	.w8(32'h3b1f6c63),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22920b),
	.w1(32'hba41353c),
	.w2(32'hbb336994),
	.w3(32'hbc6d1a67),
	.w4(32'hbd26c3f2),
	.w5(32'hbb58fccb),
	.w6(32'h3bd9d1cb),
	.w7(32'hbccbc8a1),
	.w8(32'h3a2a5ac1),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba323bb),
	.w1(32'hbb3f74f4),
	.w2(32'hbc0b58de),
	.w3(32'hb805244d),
	.w4(32'h3bc2b06f),
	.w5(32'hbb18ea46),
	.w6(32'hbc5404d8),
	.w7(32'hbbb11124),
	.w8(32'hbb73542a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a869c0),
	.w1(32'hbb7a69a5),
	.w2(32'hbb3508cd),
	.w3(32'hbb7b0eb7),
	.w4(32'h3affc726),
	.w5(32'hb9e8e37d),
	.w6(32'hbc48f86e),
	.w7(32'hbbd99713),
	.w8(32'h3c049d0a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e24eb7),
	.w1(32'hbc06fdff),
	.w2(32'hbba57614),
	.w3(32'hbc07d740),
	.w4(32'hbaa16ea7),
	.w5(32'hbaacfdc6),
	.w6(32'h3bbde3b8),
	.w7(32'h3bfa7dcd),
	.w8(32'hbc940046),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ab8dc),
	.w1(32'hbcc5a1da),
	.w2(32'hbcec8a12),
	.w3(32'h3bb75f85),
	.w4(32'h3cc47f3b),
	.w5(32'hbc1c80b0),
	.w6(32'h3d0b68b0),
	.w7(32'h3c902c78),
	.w8(32'hbc3151ba),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc730491),
	.w1(32'hbc039b97),
	.w2(32'hbb4f387f),
	.w3(32'hbc36c6f5),
	.w4(32'hbc0725ea),
	.w5(32'hbc01de99),
	.w6(32'hbc617ba9),
	.w7(32'h3b356162),
	.w8(32'hb9ca8ad1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb618f0),
	.w1(32'h3bb50410),
	.w2(32'h3cc1f741),
	.w3(32'hbcafa3b8),
	.w4(32'hbcce01a8),
	.w5(32'h3b12fc28),
	.w6(32'h3d0bd72d),
	.w7(32'h3cbb5c46),
	.w8(32'hba2c30fc),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1b6eb),
	.w1(32'hbc0ec8f8),
	.w2(32'hbbd5c4f2),
	.w3(32'hbb79b27a),
	.w4(32'h3b2358d9),
	.w5(32'hbad16228),
	.w6(32'hbc154c9c),
	.w7(32'hbb65b07c),
	.w8(32'h3aae403a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d1a5b),
	.w1(32'hbb337980),
	.w2(32'hbb3095fe),
	.w3(32'h3a85b358),
	.w4(32'h3b497818),
	.w5(32'h3974a2d1),
	.w6(32'hbbf33f8f),
	.w7(32'hbb03ea6e),
	.w8(32'h3b351304),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be992db),
	.w1(32'hbbe49755),
	.w2(32'hbc1a40bb),
	.w3(32'h3b440714),
	.w4(32'h3bcb3c0e),
	.w5(32'hba2595a5),
	.w6(32'hbc9352d6),
	.w7(32'hbbab2784),
	.w8(32'hbc773f65),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70d43a),
	.w1(32'hbb974a6c),
	.w2(32'h3be94c7f),
	.w3(32'h3c4206b7),
	.w4(32'hbc35ae8c),
	.w5(32'hbc21cf4d),
	.w6(32'hbca86259),
	.w7(32'h3c9dfbbb),
	.w8(32'h3be496b1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5b3fe),
	.w1(32'hbbeb48d4),
	.w2(32'h3c29937d),
	.w3(32'hbcf025d1),
	.w4(32'hbcd7da46),
	.w5(32'hbc148681),
	.w6(32'h3ccf7f08),
	.w7(32'h3c806947),
	.w8(32'hbb90f001),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c7723),
	.w1(32'hbbacea35),
	.w2(32'hbc0c1319),
	.w3(32'hbca6b11b),
	.w4(32'hbc0f4799),
	.w5(32'h3c033cfa),
	.w6(32'hbb8acd05),
	.w7(32'hbbf0960e),
	.w8(32'h3b96d9a5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48128d),
	.w1(32'h3b70d7c9),
	.w2(32'hbb87fd82),
	.w3(32'hb95bfd31),
	.w4(32'h3bd80923),
	.w5(32'h3c3f81ec),
	.w6(32'h3b8babc8),
	.w7(32'h3c46bfdf),
	.w8(32'hbb91ec59),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a031d),
	.w1(32'hbb3a0570),
	.w2(32'h3c1f2744),
	.w3(32'h3c052643),
	.w4(32'hbb682522),
	.w5(32'hbc8362ab),
	.w6(32'hbc11d49f),
	.w7(32'h3b559219),
	.w8(32'hbbcc9561),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd43380b),
	.w1(32'hbc81b361),
	.w2(32'hbd256129),
	.w3(32'hbd052b43),
	.w4(32'hbd3e4b24),
	.w5(32'hbbc5047a),
	.w6(32'hbd052e07),
	.w7(32'hbcb84bfd),
	.w8(32'hbb34307e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39273101),
	.w1(32'hba8d0748),
	.w2(32'hbc183dad),
	.w3(32'h3c8336e5),
	.w4(32'h3c8e0de2),
	.w5(32'h3c0690ad),
	.w6(32'hbba3e44b),
	.w7(32'hbbfede61),
	.w8(32'hba3dc806),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc88b1f),
	.w1(32'hb915fe79),
	.w2(32'h3bbd34a5),
	.w3(32'hbc1e923b),
	.w4(32'hbc595319),
	.w5(32'hbac2d938),
	.w6(32'h3c8602f4),
	.w7(32'hbbae7596),
	.w8(32'hbc2be270),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a5df2),
	.w1(32'h3b258724),
	.w2(32'hbb85f456),
	.w3(32'hbc5561ad),
	.w4(32'h3c780a06),
	.w5(32'h3c277aa2),
	.w6(32'h3c30a23e),
	.w7(32'h3bedd183),
	.w8(32'h3c08c8a6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbffd8f),
	.w1(32'hbc84c052),
	.w2(32'hbc9dea9a),
	.w3(32'hbc60c6dd),
	.w4(32'hbbfe547b),
	.w5(32'hbbec6fb7),
	.w6(32'hbafe77d7),
	.w7(32'h3a4540b9),
	.w8(32'hbac911bb),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3405b),
	.w1(32'hbb0afc5a),
	.w2(32'hbc4fa171),
	.w3(32'h3bd96ace),
	.w4(32'h3c19310e),
	.w5(32'hbba825d8),
	.w6(32'hbc286b31),
	.w7(32'hbc77dc42),
	.w8(32'hbc85902d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd326e32),
	.w1(32'hbbbe2975),
	.w2(32'hbc949436),
	.w3(32'hbcc120a5),
	.w4(32'hbd2eaa04),
	.w5(32'hbae47cec),
	.w6(32'hbcdd12c8),
	.w7(32'hbd530945),
	.w8(32'hbb8a74b9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule