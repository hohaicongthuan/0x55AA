module layer_10_featuremap_48(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2aa495),
	.w1(32'hbb4568bc),
	.w2(32'hbc02be43),
	.w3(32'hbc4f3ea2),
	.w4(32'hbbfa7415),
	.w5(32'hbc37b7ae),
	.w6(32'hbc4393dc),
	.w7(32'hbc218c5b),
	.w8(32'hbc371a2b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45deab),
	.w1(32'hbbc8d42d),
	.w2(32'hbb6e65aa),
	.w3(32'hbc60f06b),
	.w4(32'hbc0d426d),
	.w5(32'h3b1faae5),
	.w6(32'hbc165e70),
	.w7(32'h3b40d38f),
	.w8(32'h3b2abc48),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09e8d5),
	.w1(32'h3b79b565),
	.w2(32'h3b5c6a7e),
	.w3(32'h3af45422),
	.w4(32'h3c3456fb),
	.w5(32'h3bb0a130),
	.w6(32'h3aed642a),
	.w7(32'h3b5b7df9),
	.w8(32'h3bc48a02),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba024f76),
	.w1(32'h3c1ad025),
	.w2(32'hbbbb781d),
	.w3(32'h3b1134f5),
	.w4(32'h3a08a62c),
	.w5(32'hbb3c7ed4),
	.w6(32'hbb2a74d7),
	.w7(32'h3b8076a0),
	.w8(32'hbbe80720),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5de789),
	.w1(32'hbbc2880b),
	.w2(32'h3a0d4923),
	.w3(32'hbb7e6d79),
	.w4(32'h3aeaa3c2),
	.w5(32'hbb8cff32),
	.w6(32'hbc0dcffa),
	.w7(32'h3b996b82),
	.w8(32'hbc15516a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5915c1),
	.w1(32'hba928a09),
	.w2(32'h3bc0e083),
	.w3(32'hbbee8b54),
	.w4(32'h3a48ddef),
	.w5(32'h3b38a6e2),
	.w6(32'hbae14c8a),
	.w7(32'h3b97897a),
	.w8(32'h3b74af88),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c040387),
	.w1(32'hbbeefedc),
	.w2(32'hbcb33c6e),
	.w3(32'h3b12a5d1),
	.w4(32'hbc1ddd75),
	.w5(32'hbc8cadd0),
	.w6(32'h3c2cec8b),
	.w7(32'h3a1d421f),
	.w8(32'hbc986d7d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05e004),
	.w1(32'h3bae5ea6),
	.w2(32'hbc4e1cce),
	.w3(32'h3c23b226),
	.w4(32'hbb0acacf),
	.w5(32'hbabba58f),
	.w6(32'hbbc5481e),
	.w7(32'hbcba0c73),
	.w8(32'hbc48ebb3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f62228),
	.w1(32'hba962dfe),
	.w2(32'h3bf4e71a),
	.w3(32'hb9042bf7),
	.w4(32'hbb0fb327),
	.w5(32'hba2b3d1b),
	.w6(32'h398e4c86),
	.w7(32'hba1238db),
	.w8(32'h3793d647),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f7bbb),
	.w1(32'hbc2aa3d4),
	.w2(32'hbc6e850f),
	.w3(32'hbc8c9a30),
	.w4(32'hbc49f4f2),
	.w5(32'hbc4df79c),
	.w6(32'hbbccf03a),
	.w7(32'hbbec0aa6),
	.w8(32'hbc314390),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37b03e),
	.w1(32'h39c1df7b),
	.w2(32'h38f5c9a5),
	.w3(32'h39f76288),
	.w4(32'hbb386025),
	.w5(32'h3bb6aa2b),
	.w6(32'hbad569c4),
	.w7(32'hbb2c84d2),
	.w8(32'h3a94fc37),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4912aa),
	.w1(32'h3c18cd90),
	.w2(32'hbccaddbf),
	.w3(32'h3c5208ca),
	.w4(32'h3c08e008),
	.w5(32'hbcc8ed92),
	.w6(32'h3c1408e0),
	.w7(32'h3b80a706),
	.w8(32'hbcbc1201),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d990e),
	.w1(32'hbc6659f4),
	.w2(32'hbcec7f2e),
	.w3(32'hbc3cda18),
	.w4(32'hbc8c9965),
	.w5(32'hbca9186c),
	.w6(32'hbc19197e),
	.w7(32'hbc9e3d2a),
	.w8(32'hbcac8253),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa20b7e),
	.w1(32'h3ad0d14c),
	.w2(32'hbc301233),
	.w3(32'hb8845f7c),
	.w4(32'h3aa15310),
	.w5(32'hbc0d666e),
	.w6(32'h3b80b3e9),
	.w7(32'hb8521526),
	.w8(32'hbc08fc2a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e0f96),
	.w1(32'hba6d1db3),
	.w2(32'h3c4f1478),
	.w3(32'hbc200219),
	.w4(32'h3b8de35f),
	.w5(32'h3c50a244),
	.w6(32'hbba6277a),
	.w7(32'h3b076029),
	.w8(32'h3b706274),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba87a95),
	.w1(32'hb709f206),
	.w2(32'hbcdbac2b),
	.w3(32'hbad20fc4),
	.w4(32'h3b126837),
	.w5(32'hbc82cbfb),
	.w6(32'hbc376b87),
	.w7(32'hbc3358ce),
	.w8(32'hbc902475),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b439682),
	.w1(32'hba4b20b1),
	.w2(32'h39df4b72),
	.w3(32'h3acc3c82),
	.w4(32'hbac02e59),
	.w5(32'h3be8a8fb),
	.w6(32'h390e6e95),
	.w7(32'hbad76834),
	.w8(32'h3b8d7725),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a5a5a),
	.w1(32'hbc8ea28f),
	.w2(32'hbd00a338),
	.w3(32'h3c989322),
	.w4(32'hbbf1f525),
	.w5(32'hbd2346fc),
	.w6(32'h3c0acbb7),
	.w7(32'hbb5471fa),
	.w8(32'hbce864b5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb141fbe),
	.w1(32'hbbfb124a),
	.w2(32'hbc85dd10),
	.w3(32'hbac67232),
	.w4(32'hbbafbde1),
	.w5(32'hbbd0d309),
	.w6(32'h3b63b336),
	.w7(32'hbb8d6ad9),
	.w8(32'hbc040ecf),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdefc1f),
	.w1(32'h3ba347b4),
	.w2(32'h3b818d06),
	.w3(32'h3bd9ecbc),
	.w4(32'h3c0610ec),
	.w5(32'h3be279ab),
	.w6(32'h3c290c89),
	.w7(32'h3b4d1ac6),
	.w8(32'h3b801058),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dd015),
	.w1(32'h3ad7f9ff),
	.w2(32'h3be7cf40),
	.w3(32'h3c042791),
	.w4(32'h3bf49fbc),
	.w5(32'h3c3a5b45),
	.w6(32'h3ad2332b),
	.w7(32'h3b101767),
	.w8(32'h3bf4252a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd63add),
	.w1(32'h3c526542),
	.w2(32'h3b8cfde8),
	.w3(32'h3bac265a),
	.w4(32'h3baafe33),
	.w5(32'h3bfedd1a),
	.w6(32'h3c3f05cd),
	.w7(32'h3c1b23d7),
	.w8(32'h3b8c8731),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e661b),
	.w1(32'hbc1fe7b9),
	.w2(32'hbd32a485),
	.w3(32'hbbf08549),
	.w4(32'h3b8eea50),
	.w5(32'hbceadac3),
	.w6(32'hb940c537),
	.w7(32'hbbf9e9e3),
	.w8(32'hbcdc0cfe),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04976a),
	.w1(32'hbbc75d7c),
	.w2(32'hbba38d1a),
	.w3(32'hbc7c203f),
	.w4(32'hbc287acf),
	.w5(32'hbbb1c37e),
	.w6(32'hbc45e55a),
	.w7(32'hbbca25f3),
	.w8(32'h3a47ef35),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc193134),
	.w1(32'h3c457367),
	.w2(32'h3cf175a0),
	.w3(32'hbcbe8eb9),
	.w4(32'h3c501987),
	.w5(32'h3ce6ffb7),
	.w6(32'hbc56dd8f),
	.w7(32'h3c46b744),
	.w8(32'h3cd90b6c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9da3be),
	.w1(32'h3b387c19),
	.w2(32'h3af90863),
	.w3(32'h3aabf83c),
	.w4(32'hba9f2340),
	.w5(32'hbb84292b),
	.w6(32'h3bab60b4),
	.w7(32'hba1282ea),
	.w8(32'hbbf1417f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e1344),
	.w1(32'hbbaf53a4),
	.w2(32'h3ae8a50e),
	.w3(32'hbb27968b),
	.w4(32'hbb90b9e4),
	.w5(32'h3bcf5846),
	.w6(32'hbbc60fec),
	.w7(32'h3bd04ab8),
	.w8(32'h3ae3f21b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bbe58),
	.w1(32'h3c3060e9),
	.w2(32'h3bb0bd98),
	.w3(32'hbbd228d6),
	.w4(32'h3c53ee5d),
	.w5(32'h3ca29aea),
	.w6(32'hbbc06ecf),
	.w7(32'h3cc3fddf),
	.w8(32'h3c6f5ee6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ac40c),
	.w1(32'hbc71f345),
	.w2(32'hbbb46217),
	.w3(32'h3b8ac2e7),
	.w4(32'hbb62586d),
	.w5(32'hbc540ec5),
	.w6(32'hbb6763e2),
	.w7(32'hbc28edf4),
	.w8(32'hbb4ef1cb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe14c1),
	.w1(32'h3c024e39),
	.w2(32'h3cc72c80),
	.w3(32'hbcf4841a),
	.w4(32'hbc81bc4a),
	.w5(32'h3cc74b11),
	.w6(32'hbc4d89d4),
	.w7(32'hbbbac18f),
	.w8(32'h3cadf2ad),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c8012),
	.w1(32'hbb222e8f),
	.w2(32'hbc840772),
	.w3(32'h3b4e020a),
	.w4(32'h3b921da1),
	.w5(32'hbcaa09af),
	.w6(32'hbb645e77),
	.w7(32'hbb4cf38c),
	.w8(32'h3a9ac8e8),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd017bee),
	.w1(32'hbc414ea3),
	.w2(32'hbc7b3109),
	.w3(32'hbd3c9970),
	.w4(32'hbcd09080),
	.w5(32'hbd33f417),
	.w6(32'hbc767dfc),
	.w7(32'hbade4edb),
	.w8(32'hbcc8ec7b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc148651),
	.w1(32'hbb93f72c),
	.w2(32'hbc67c85f),
	.w3(32'hbd563a53),
	.w4(32'hbcb7e6ae),
	.w5(32'hbb2288ff),
	.w6(32'hbcff24fd),
	.w7(32'hbc2b836d),
	.w8(32'h39605f8b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d2d1b),
	.w1(32'hbbce7ba7),
	.w2(32'hbbac49d9),
	.w3(32'hbbaecfc0),
	.w4(32'hba0c1c70),
	.w5(32'hbb201164),
	.w6(32'hbb27e884),
	.w7(32'h3a2542c7),
	.w8(32'hbb6a3e5a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12f270),
	.w1(32'h3bb25954),
	.w2(32'h38c92224),
	.w3(32'hba42b504),
	.w4(32'hbabf36d1),
	.w5(32'hbacdae7d),
	.w6(32'hbc1fbf47),
	.w7(32'hbb70a2a6),
	.w8(32'h3a8a303a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb68a4),
	.w1(32'h3b8b732f),
	.w2(32'hbd1705b7),
	.w3(32'h3b8a4ae3),
	.w4(32'h3a2a9de8),
	.w5(32'hbcfe319b),
	.w6(32'h3b498265),
	.w7(32'h3b7efff1),
	.w8(32'hbcb45823),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4161a8),
	.w1(32'h3c6d3821),
	.w2(32'hbd2a561b),
	.w3(32'hbd6562c3),
	.w4(32'h3cc9b0f0),
	.w5(32'hbd1728c1),
	.w6(32'hbd3f91fb),
	.w7(32'h3bb3917c),
	.w8(32'hbd213d0b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a56a6),
	.w1(32'h3cf25718),
	.w2(32'h3d291951),
	.w3(32'hbc0eb8df),
	.w4(32'h3d055512),
	.w5(32'h3d5b0641),
	.w6(32'hbb64734f),
	.w7(32'h3cfa75a6),
	.w8(32'h3d91ef39),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd31c749),
	.w1(32'hbc38d8e2),
	.w2(32'h3cfbb3be),
	.w3(32'hbcafefa1),
	.w4(32'hbb0ef1e4),
	.w5(32'h3cef76bf),
	.w6(32'h3cec15e1),
	.w7(32'h3d03bdab),
	.w8(32'h3d326956),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2535c),
	.w1(32'h3c75346e),
	.w2(32'h3c03c59a),
	.w3(32'hbba8fc94),
	.w4(32'h3c81bc38),
	.w5(32'h3c13b676),
	.w6(32'hbba93227),
	.w7(32'hba713394),
	.w8(32'h3c2a5651),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacee1f4),
	.w1(32'h38f187c3),
	.w2(32'hbbfd67bb),
	.w3(32'hbaf4d3c9),
	.w4(32'hb9a7ecc3),
	.w5(32'hbbffbc72),
	.w6(32'h3ab4a518),
	.w7(32'hb9926f48),
	.w8(32'hbbddfff2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42b7ca),
	.w1(32'hbb54e32b),
	.w2(32'hbc1fb5ec),
	.w3(32'hbc3de3fa),
	.w4(32'h3ae92c14),
	.w5(32'hbc133173),
	.w6(32'h3b000986),
	.w7(32'h3b306891),
	.w8(32'h3bd6fbb2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb4a027),
	.w1(32'h3b30e6e4),
	.w2(32'hbb62828d),
	.w3(32'hbcca5268),
	.w4(32'h39f087a5),
	.w5(32'h3ae80349),
	.w6(32'h3c67c1a9),
	.w7(32'h3c41bf4c),
	.w8(32'h3adb5fa0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc167682),
	.w1(32'hbc92bb3d),
	.w2(32'hbcf474ee),
	.w3(32'h3b851dd8),
	.w4(32'hbba6696e),
	.w5(32'hbbe5d219),
	.w6(32'hbaae6966),
	.w7(32'hba042fed),
	.w8(32'hbcab6627),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41d69f),
	.w1(32'h3c3e2f70),
	.w2(32'h3c9085dc),
	.w3(32'hbc7e1189),
	.w4(32'hbc96ce48),
	.w5(32'h3b3ccf27),
	.w6(32'hbc9ddc06),
	.w7(32'hbc40e017),
	.w8(32'hbbf42345),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf438fc),
	.w1(32'h3b81f958),
	.w2(32'h3b1cb5d7),
	.w3(32'hbced5612),
	.w4(32'hbbf3bb9a),
	.w5(32'h3ba55429),
	.w6(32'hbcb01719),
	.w7(32'hbbe364ca),
	.w8(32'hbaeaaa52),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e012b),
	.w1(32'hba89f021),
	.w2(32'h3b336bd2),
	.w3(32'hbac677eb),
	.w4(32'h3c78c008),
	.w5(32'h3c8c1f7f),
	.w6(32'h3c3e9e82),
	.w7(32'h3c92a47a),
	.w8(32'h3c68e136),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc0dce),
	.w1(32'hbc8b549b),
	.w2(32'hbd28ad7f),
	.w3(32'h3c5c2587),
	.w4(32'hbc28cd42),
	.w5(32'hbd1f3af2),
	.w6(32'h3cd2e139),
	.w7(32'h3b5e8066),
	.w8(32'hbcfbbef4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1a78e),
	.w1(32'h3b3dd004),
	.w2(32'hbcb31056),
	.w3(32'h3b31e0e3),
	.w4(32'h3b501310),
	.w5(32'hbc48b8f1),
	.w6(32'h3bc0876c),
	.w7(32'h3bb84560),
	.w8(32'hbac1d939),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7186c),
	.w1(32'hbb0205b1),
	.w2(32'hbb475b1e),
	.w3(32'hbcb4d447),
	.w4(32'hbbf8ca60),
	.w5(32'h3c5705e8),
	.w6(32'h3b8f1449),
	.w7(32'h3c09ff7d),
	.w8(32'hbb9083fa),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c940d1f),
	.w1(32'h3c740287),
	.w2(32'hbc5c3918),
	.w3(32'h3c8af09b),
	.w4(32'h3c6c992c),
	.w5(32'h3b1d002e),
	.w6(32'hbc112eac),
	.w7(32'h3a90b741),
	.w8(32'hbb2ace38),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9213f0),
	.w1(32'hbb23c10d),
	.w2(32'h3a8a7e1b),
	.w3(32'hbc15987a),
	.w4(32'h3bd9b34c),
	.w5(32'h3c7a501f),
	.w6(32'hba8a3b7e),
	.w7(32'h3bcfdcaa),
	.w8(32'hbc13f9cc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8333bc),
	.w1(32'h3cb4a545),
	.w2(32'hbc4fa3b2),
	.w3(32'h3c521f8d),
	.w4(32'h3c6c8d5e),
	.w5(32'hbc07951f),
	.w6(32'hbbac450f),
	.w7(32'hbb1bcfff),
	.w8(32'hbb485417),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc306d53),
	.w1(32'hbc7fbdf2),
	.w2(32'hbd75e6de),
	.w3(32'hbb8447b8),
	.w4(32'hbafa5eab),
	.w5(32'hbd34af0b),
	.w6(32'h3bf81faf),
	.w7(32'hbb850a72),
	.w8(32'hbbac286c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f86a8),
	.w1(32'hbb244d48),
	.w2(32'hbc8c9677),
	.w3(32'h3a6b8d14),
	.w4(32'h3b855674),
	.w5(32'hbcbe161b),
	.w6(32'h3ca97d29),
	.w7(32'h3c42b8f5),
	.w8(32'hbc919843),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83739a),
	.w1(32'hbb86ed03),
	.w2(32'hbb808391),
	.w3(32'hbd45acf3),
	.w4(32'hbd32ae0e),
	.w5(32'hbbfb2a1e),
	.w6(32'hbceebd8b),
	.w7(32'hbc8bc3d8),
	.w8(32'h3c082151),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fa912),
	.w1(32'h3c1a0f9c),
	.w2(32'hbb67a7a8),
	.w3(32'hba8720c8),
	.w4(32'h3c74fbaf),
	.w5(32'h3c0758a0),
	.w6(32'h3c0f288e),
	.w7(32'h3ba9a964),
	.w8(32'h3b7485f0),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ebffa),
	.w1(32'h388937fe),
	.w2(32'h3b3cc6f4),
	.w3(32'h3b418d7b),
	.w4(32'h3b3ffae5),
	.w5(32'h3bf368b4),
	.w6(32'hbaa74bae),
	.w7(32'h3b74dff8),
	.w8(32'h3bbadab7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a213b27),
	.w1(32'h39f34a88),
	.w2(32'hbb1536ca),
	.w3(32'h3bcdaa68),
	.w4(32'h3b864726),
	.w5(32'h3a9bbc9c),
	.w6(32'h3c0232bb),
	.w7(32'h3bb026a1),
	.w8(32'h3c19e5ee),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bfcd5),
	.w1(32'hba1c2183),
	.w2(32'hbc287de4),
	.w3(32'hbbcf5833),
	.w4(32'h392e5489),
	.w5(32'h3bbd70a9),
	.w6(32'h3b884e35),
	.w7(32'h3bbadeea),
	.w8(32'h3c2b2460),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bb689),
	.w1(32'hbc88775d),
	.w2(32'hbc964260),
	.w3(32'h3bb09a9c),
	.w4(32'h3b829343),
	.w5(32'hbc84fba3),
	.w6(32'h3c0ab233),
	.w7(32'h3afdecb5),
	.w8(32'hbc1c5c1b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53e820),
	.w1(32'h3aa613cc),
	.w2(32'hbc4511c2),
	.w3(32'hbb87ef96),
	.w4(32'h3c9d184c),
	.w5(32'hbc0602e5),
	.w6(32'h3a656997),
	.w7(32'h3b2246b7),
	.w8(32'hbbc7ce24),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b18ab),
	.w1(32'hbaa6b7e6),
	.w2(32'hbc01088a),
	.w3(32'hbb820e22),
	.w4(32'hbb46b70f),
	.w5(32'h3bff6492),
	.w6(32'h3b57da50),
	.w7(32'hb9aa8bcc),
	.w8(32'hbabb3dd6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8dc6d),
	.w1(32'hbc20dec9),
	.w2(32'h3b9ae3cb),
	.w3(32'h3b905573),
	.w4(32'h3a22573c),
	.w5(32'h3a0fb39e),
	.w6(32'hbbce9b2d),
	.w7(32'hbc2bf969),
	.w8(32'h3b9fa51c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e2d93),
	.w1(32'hbc8ef02d),
	.w2(32'h3b2fb4f6),
	.w3(32'hbc4bed1b),
	.w4(32'hbc747c19),
	.w5(32'hba13e024),
	.w6(32'hbb9270d0),
	.w7(32'h3b59b132),
	.w8(32'hba1a2e43),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda149f),
	.w1(32'h3b66b3d4),
	.w2(32'hbb12ed76),
	.w3(32'h3b20a5be),
	.w4(32'h38219712),
	.w5(32'h3bb25349),
	.w6(32'hbb975ca2),
	.w7(32'hbbbf3bf4),
	.w8(32'h3abf9cd3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca34b31),
	.w1(32'hbc2030ff),
	.w2(32'hbd5ffabf),
	.w3(32'h3c027038),
	.w4(32'h3b9c7e5b),
	.w5(32'hbd27f906),
	.w6(32'h3c39864b),
	.w7(32'hbb450ed1),
	.w8(32'hbcfce2f1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d3e7f),
	.w1(32'h3bb82b4e),
	.w2(32'hbc4ec53a),
	.w3(32'h3b48300f),
	.w4(32'h3902990b),
	.w5(32'hbb0393d0),
	.w6(32'hbd105918),
	.w7(32'hbcbd100c),
	.w8(32'hbcc488e4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47d3d9),
	.w1(32'hbaf1ac6d),
	.w2(32'hbc4c0ddc),
	.w3(32'h3cafab37),
	.w4(32'h3c002338),
	.w5(32'hbc5a0019),
	.w6(32'hbb30b218),
	.w7(32'hbca8a48a),
	.w8(32'hbcb37acd),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fcc01),
	.w1(32'h3c9ab985),
	.w2(32'h3cfd0f6c),
	.w3(32'hbcd47dac),
	.w4(32'h3c43a77d),
	.w5(32'h3d368315),
	.w6(32'hbcb91a61),
	.w7(32'h3baf2c8f),
	.w8(32'h3d126199),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78233c),
	.w1(32'hbbeeeac2),
	.w2(32'hbb4ec0aa),
	.w3(32'h3baa1893),
	.w4(32'h395fc21d),
	.w5(32'hbbb88676),
	.w6(32'h3c0410a1),
	.w7(32'hbba13c47),
	.w8(32'h39632d7d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90706d),
	.w1(32'h3afaf438),
	.w2(32'h3a64f5d5),
	.w3(32'hba3bdaa7),
	.w4(32'h3c03a639),
	.w5(32'hbb12a1d0),
	.w6(32'h3a937e38),
	.w7(32'hbaa38f72),
	.w8(32'h3b6b836e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9a982),
	.w1(32'hbb36483a),
	.w2(32'hbbfc89e7),
	.w3(32'h3c24c1aa),
	.w4(32'h3bef0315),
	.w5(32'h3c40e8f7),
	.w6(32'h3c8bb74f),
	.w7(32'h3c346adb),
	.w8(32'h3cc22085),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e95d7),
	.w1(32'h3a332c49),
	.w2(32'hbb490dd8),
	.w3(32'h3b311617),
	.w4(32'h3c10275f),
	.w5(32'hbb10ab63),
	.w6(32'h3cc2865b),
	.w7(32'h3c59eb1d),
	.w8(32'hbbf26730),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c294cba),
	.w1(32'h3c03b61e),
	.w2(32'hbc337bb1),
	.w3(32'h3c09f954),
	.w4(32'h3bcf8ac9),
	.w5(32'h3b806946),
	.w6(32'h3b9d3fbf),
	.w7(32'h3b0c6d55),
	.w8(32'h3c61a512),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc168484),
	.w1(32'hbc859d47),
	.w2(32'hbb82f342),
	.w3(32'hbb7f85b9),
	.w4(32'hbbba4b96),
	.w5(32'h3bc0fdb0),
	.w6(32'h3ca13826),
	.w7(32'h3c13ba64),
	.w8(32'h3b067792),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b35c3),
	.w1(32'h3c80fd5f),
	.w2(32'hbc98df97),
	.w3(32'h3d05abb6),
	.w4(32'h3d19e60c),
	.w5(32'hbc3504d0),
	.w6(32'h3ce71b94),
	.w7(32'h3c52ac6c),
	.w8(32'hbc06461a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19ee06),
	.w1(32'h3ace850f),
	.w2(32'h3c3dc304),
	.w3(32'hbb9c246c),
	.w4(32'h3ca0806a),
	.w5(32'h3c3c0dbd),
	.w6(32'h3c009396),
	.w7(32'h3c5f87aa),
	.w8(32'h3952588b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ad587),
	.w1(32'hbbddf497),
	.w2(32'hbc1f4440),
	.w3(32'h3c3a1602),
	.w4(32'hba395570),
	.w5(32'hbc288f3b),
	.w6(32'h3c939942),
	.w7(32'h3c374986),
	.w8(32'hbc1961af),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c490d01),
	.w1(32'h3c1997f1),
	.w2(32'hbc36f373),
	.w3(32'hbb8e1a4a),
	.w4(32'h3bf6e57f),
	.w5(32'hbbed1166),
	.w6(32'h3bf19ba9),
	.w7(32'h3c245bdd),
	.w8(32'hbc075911),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9bbac),
	.w1(32'h392473d7),
	.w2(32'hbb4a17b4),
	.w3(32'hbb56dee5),
	.w4(32'hba0e16e5),
	.w5(32'h3c292c2d),
	.w6(32'hbb0840e9),
	.w7(32'h3b1e0fda),
	.w8(32'hba34edbd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef6f9f),
	.w1(32'hbb06ecf0),
	.w2(32'hbd0d717f),
	.w3(32'h3c4afc4e),
	.w4(32'h3c16ed73),
	.w5(32'hbd19d12e),
	.w6(32'h3a1c1996),
	.w7(32'hbb3eb35b),
	.w8(32'hbc99cccd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60c804),
	.w1(32'h3b8b50e8),
	.w2(32'hbb984fc3),
	.w3(32'hbc6cb60a),
	.w4(32'h3b524510),
	.w5(32'hba615f66),
	.w6(32'hbc540e8f),
	.w7(32'hbc978565),
	.w8(32'hbbb7ca51),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4075dc),
	.w1(32'h3bdd7957),
	.w2(32'hb9546163),
	.w3(32'h3c23c368),
	.w4(32'h3c66a2be),
	.w5(32'h3bc3c8dd),
	.w6(32'h3c6efbf8),
	.w7(32'h3c43f834),
	.w8(32'h3ab38cd9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c698a),
	.w1(32'h3bc6759e),
	.w2(32'h3b608ae3),
	.w3(32'h3c2df956),
	.w4(32'h3c64aa45),
	.w5(32'h3bfedf6b),
	.w6(32'h3ba465da),
	.w7(32'h3c816da2),
	.w8(32'h3bff0d4e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a8ae4),
	.w1(32'h3b13e38e),
	.w2(32'h3b24139b),
	.w3(32'h3ba0a0a1),
	.w4(32'h3b066878),
	.w5(32'h3af6c110),
	.w6(32'hbc168641),
	.w7(32'hbc1fa646),
	.w8(32'h3bfc6281),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacb4f3),
	.w1(32'h3c21cf36),
	.w2(32'h3b3211b7),
	.w3(32'hbb8d07c5),
	.w4(32'h3c3f7174),
	.w5(32'h3c1e7016),
	.w6(32'hba0825e3),
	.w7(32'h3b661452),
	.w8(32'h3c057f7b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afebc08),
	.w1(32'hbb3a6191),
	.w2(32'h3bc47ef8),
	.w3(32'hbb2affdc),
	.w4(32'h39ca44bc),
	.w5(32'h3c0bf3b6),
	.w6(32'hbb11e832),
	.w7(32'hbaf6e24c),
	.w8(32'hba7fc36c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08058c),
	.w1(32'h3ca9eaaa),
	.w2(32'hbb1a1326),
	.w3(32'h3c049125),
	.w4(32'h3cc80c16),
	.w5(32'hba08e26a),
	.w6(32'hbcd3d76f),
	.w7(32'hbb735dcc),
	.w8(32'hbc10b674),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a2aa8),
	.w1(32'h3b0724a3),
	.w2(32'hbcd1522b),
	.w3(32'hbbc60a56),
	.w4(32'hbb9db0d8),
	.w5(32'hbc7b1115),
	.w6(32'hbb6df0fe),
	.w7(32'hbaa891cc),
	.w8(32'hbc84df1f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5d5d7),
	.w1(32'h3ae23c77),
	.w2(32'h3c8f6cf8),
	.w3(32'hbbeb7134),
	.w4(32'h3ba599a9),
	.w5(32'h3d0419a6),
	.w6(32'hbb315c2f),
	.w7(32'h3c5b6d1d),
	.w8(32'h3d00a2b7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf8a33),
	.w1(32'h3b56c3d6),
	.w2(32'hbd40c292),
	.w3(32'h3bf7c126),
	.w4(32'h3c8ca0fd),
	.w5(32'hbd14547f),
	.w6(32'h3c43f07b),
	.w7(32'h3c47419b),
	.w8(32'hbcb3814c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8531d1),
	.w1(32'h3c18cf80),
	.w2(32'h3c8ee318),
	.w3(32'hbbd48929),
	.w4(32'h3c0d7bd8),
	.w5(32'h3cb292b8),
	.w6(32'h3b6d2217),
	.w7(32'h3c6c9a08),
	.w8(32'h3cb39e36),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23abf9),
	.w1(32'hbac92aa8),
	.w2(32'hbc861565),
	.w3(32'h3ba47fe7),
	.w4(32'h3b7a868e),
	.w5(32'hbaf0347f),
	.w6(32'hbbcfc211),
	.w7(32'hbbc27b9a),
	.w8(32'hbcd1ba43),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c380837),
	.w1(32'h3c2e2310),
	.w2(32'hbac9bbc3),
	.w3(32'h3cc159c6),
	.w4(32'h3c83df0e),
	.w5(32'hbc458059),
	.w6(32'hbb446c4b),
	.w7(32'h3b273d38),
	.w8(32'hbb976e78),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe2643),
	.w1(32'hbb861040),
	.w2(32'h3c7614d2),
	.w3(32'hbd02feac),
	.w4(32'hbbbbb140),
	.w5(32'h3c99c9e9),
	.w6(32'h3aef70b3),
	.w7(32'h3c71cad6),
	.w8(32'h3cfeea9d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ee9dc),
	.w1(32'hbb9820b9),
	.w2(32'h3c2aabcc),
	.w3(32'hbc0ea281),
	.w4(32'h3b43a279),
	.w5(32'h3ab501e8),
	.w6(32'h3b14875e),
	.w7(32'h3b615364),
	.w8(32'h3b2c2040),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e64e5),
	.w1(32'hbb95ed1b),
	.w2(32'hbcbee0a7),
	.w3(32'hbc51704f),
	.w4(32'h3bae7a62),
	.w5(32'hbc749f9e),
	.w6(32'hbac3f90e),
	.w7(32'h3b526c5f),
	.w8(32'hbb734922),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70b81f),
	.w1(32'hbadd7aee),
	.w2(32'hbcec680c),
	.w3(32'hbc1df252),
	.w4(32'hba51f35a),
	.w5(32'hbc00baa2),
	.w6(32'h3cc684ff),
	.w7(32'h3c99500b),
	.w8(32'hbc6c33c2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2bff1),
	.w1(32'h3c634c20),
	.w2(32'hbd04c3b7),
	.w3(32'hbc882cba),
	.w4(32'h3d4eb4d6),
	.w5(32'hbcc39dbb),
	.w6(32'hbd301e6c),
	.w7(32'h3c019f88),
	.w8(32'hbc96b237),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd180871),
	.w1(32'hbb8a3190),
	.w2(32'h3cd0007a),
	.w3(32'hbd3da87d),
	.w4(32'h3c65899e),
	.w5(32'h3ccdce7f),
	.w6(32'h3c268adf),
	.w7(32'h3d456d50),
	.w8(32'h3d38e975),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd24854f),
	.w1(32'hbc80cb36),
	.w2(32'h3bdb203c),
	.w3(32'hbd791158),
	.w4(32'hbc5e4aac),
	.w5(32'h3c103672),
	.w6(32'hbc93c781),
	.w7(32'h3c291984),
	.w8(32'hbb13dac5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc588c89),
	.w1(32'h397a559f),
	.w2(32'hbcf04ed5),
	.w3(32'hbc2cbdf9),
	.w4(32'h3c5403fd),
	.w5(32'hbcd052a1),
	.w6(32'h3bb27f8a),
	.w7(32'h3c65510d),
	.w8(32'hbcd1f71c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b9c965),
	.w1(32'h3bd62cc7),
	.w2(32'h3b2864f1),
	.w3(32'hbb5cf576),
	.w4(32'h3bd606e9),
	.w5(32'h39e43f53),
	.w6(32'hbbcf4215),
	.w7(32'hba51514b),
	.w8(32'hbabf55e2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f186f),
	.w1(32'h3ca31c72),
	.w2(32'hbce20298),
	.w3(32'hbcd09b44),
	.w4(32'h3cdd36b1),
	.w5(32'hbc737d55),
	.w6(32'hbcff4888),
	.w7(32'hbb644092),
	.w8(32'hbcabba6a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53bd9b),
	.w1(32'h3b12f0c1),
	.w2(32'hbcbf5abf),
	.w3(32'h3c3c24d9),
	.w4(32'h3c02b301),
	.w5(32'hbc6a3d9d),
	.w6(32'h3ca81879),
	.w7(32'h3b8a01ec),
	.w8(32'hbb5cde5b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074cc1),
	.w1(32'h3b6b3b31),
	.w2(32'hbb3be1c1),
	.w3(32'hbb71bbe8),
	.w4(32'h3aed3ce1),
	.w5(32'hbb59c461),
	.w6(32'hbb30f280),
	.w7(32'hbb8721c0),
	.w8(32'h3bb67d42),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe8714),
	.w1(32'h3ab112bb),
	.w2(32'hbc234c26),
	.w3(32'hbbfa0500),
	.w4(32'h3bb2ece6),
	.w5(32'h3bb6a760),
	.w6(32'h3b8f1083),
	.w7(32'h3b1eb3c8),
	.w8(32'hbc27d894),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa301e1),
	.w1(32'h3bd7e3ab),
	.w2(32'hbd109c00),
	.w3(32'h3b9d98b2),
	.w4(32'h3bb8b00b),
	.w5(32'hbcb75797),
	.w6(32'h3c66834f),
	.w7(32'h3b98288b),
	.w8(32'hbca1ee87),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd27dbf6),
	.w1(32'hbc20e241),
	.w2(32'h3c4ac42f),
	.w3(32'hbd236219),
	.w4(32'hb9b67c70),
	.w5(32'h3c9f6eda),
	.w6(32'hbc039388),
	.w7(32'h3c4afdd6),
	.w8(32'h3c321b40),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66f11f),
	.w1(32'h3934810d),
	.w2(32'h3c962460),
	.w3(32'hbc498c56),
	.w4(32'hbbf61bb9),
	.w5(32'h3ccd2378),
	.w6(32'h3c429d6e),
	.w7(32'h3c7ddced),
	.w8(32'h3d11f73f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb221500),
	.w1(32'h3c2ef46d),
	.w2(32'hbb767515),
	.w3(32'hbb0456d9),
	.w4(32'h3bfc6f5d),
	.w5(32'hbb7dcaf7),
	.w6(32'h3bd57b34),
	.w7(32'h3b60a703),
	.w8(32'hbc1ff230),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c77bb),
	.w1(32'h3cc88925),
	.w2(32'hbc4af11d),
	.w3(32'h3b5ff256),
	.w4(32'h3cbb313d),
	.w5(32'hbc802046),
	.w6(32'hbcadeda1),
	.w7(32'hbc21604e),
	.w8(32'hb693fdf6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d26c4),
	.w1(32'hbba57fbc),
	.w2(32'hbd07a063),
	.w3(32'hbd0983e9),
	.w4(32'hbc0dcc2f),
	.w5(32'hbcdc2935),
	.w6(32'h3c02bb37),
	.w7(32'h3c08a946),
	.w8(32'hbc9ee423),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78735d),
	.w1(32'hbbc017df),
	.w2(32'h3c0cf8c6),
	.w3(32'hbd09df2f),
	.w4(32'hbc8fb4eb),
	.w5(32'h3c2bcaa4),
	.w6(32'hbc8d5675),
	.w7(32'hbc315a78),
	.w8(32'hbb3a2c27),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c049442),
	.w1(32'h3c112b49),
	.w2(32'hb9b73639),
	.w3(32'h3c447dda),
	.w4(32'h3c2a5ed7),
	.w5(32'hba8a86d6),
	.w6(32'hbb732b12),
	.w7(32'hbbcac7fb),
	.w8(32'hbb8bebec),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d84f4),
	.w1(32'hbb12fdce),
	.w2(32'hbb57a31a),
	.w3(32'h3bb14a54),
	.w4(32'h3ba4f108),
	.w5(32'hbb14cf70),
	.w6(32'hbb12f9a0),
	.w7(32'hbbf59db5),
	.w8(32'hbbb823ed),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb268d34),
	.w1(32'hbb236d7c),
	.w2(32'hbc7af00f),
	.w3(32'h3ad0c736),
	.w4(32'h39a9bb3a),
	.w5(32'hbb8ec3bc),
	.w6(32'hbb16c28b),
	.w7(32'hbb9a0e5a),
	.w8(32'h3c4ae630),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf98ed2),
	.w1(32'hbc807172),
	.w2(32'hbc80b02c),
	.w3(32'hbcb31bf2),
	.w4(32'hbc7b0852),
	.w5(32'hbcaf18e3),
	.w6(32'h3b00fb2a),
	.w7(32'h3b6e2d78),
	.w8(32'hbc0b17e5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd053564),
	.w1(32'hbce6cc92),
	.w2(32'h3bccdaa9),
	.w3(32'hbd335564),
	.w4(32'hbce04485),
	.w5(32'h3c0203e1),
	.w6(32'hbc39b80c),
	.w7(32'hbae59dbe),
	.w8(32'h39d8b8e9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01ddd6),
	.w1(32'hbbd125d8),
	.w2(32'hba46a150),
	.w3(32'hb8b5c7ac),
	.w4(32'h3b63103b),
	.w5(32'hba966a7c),
	.w6(32'h3b0d5267),
	.w7(32'hbad4792b),
	.w8(32'hbb49b62e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b018dc),
	.w1(32'h3b1aeb0c),
	.w2(32'hbc27eeb1),
	.w3(32'h3a6bbfe7),
	.w4(32'h3809635a),
	.w5(32'hbbb9f110),
	.w6(32'hbacf37d8),
	.w7(32'hbac5496b),
	.w8(32'hbc029671),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf87b1a),
	.w1(32'h3c023846),
	.w2(32'h3c8f591c),
	.w3(32'hbbbab3f5),
	.w4(32'h3b15f788),
	.w5(32'h3d08a84a),
	.w6(32'hbadc4280),
	.w7(32'h3a053075),
	.w8(32'h3cbc7491),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadb6bb),
	.w1(32'h3ba5680f),
	.w2(32'h3b664023),
	.w3(32'h3b4dac46),
	.w4(32'hbb75d2fb),
	.w5(32'h3b2a6de3),
	.w6(32'h3c039b20),
	.w7(32'hbbbe49e1),
	.w8(32'h3b8cc6e4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc461b),
	.w1(32'hbb37d286),
	.w2(32'hbaf6194b),
	.w3(32'h3b45cb39),
	.w4(32'hbb2eea6a),
	.w5(32'hb925414d),
	.w6(32'h3b23f31f),
	.w7(32'hbb319e03),
	.w8(32'hbb9fb078),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc11e7),
	.w1(32'h3bcfaae0),
	.w2(32'hbc472e28),
	.w3(32'h3c06c7b6),
	.w4(32'h3ba3d8af),
	.w5(32'hbc28e494),
	.w6(32'h3b13d65d),
	.w7(32'h3ac04a14),
	.w8(32'hbc3c93d2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea2981),
	.w1(32'h3bd71f38),
	.w2(32'hbbc0e4e6),
	.w3(32'h3a832619),
	.w4(32'h3a0740b9),
	.w5(32'hb9cb5a9d),
	.w6(32'hbbb93c06),
	.w7(32'hbc70991c),
	.w8(32'hbc67db9a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c276ade),
	.w1(32'h3c9542e9),
	.w2(32'hbca42070),
	.w3(32'h3c69b8df),
	.w4(32'h3c9cd792),
	.w5(32'hbd09ebb0),
	.w6(32'hbc2254fd),
	.w7(32'hbc4b5e6c),
	.w8(32'hbccc0844),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9cd3f),
	.w1(32'h3b0f02b2),
	.w2(32'hbd057fd5),
	.w3(32'hbb1965b2),
	.w4(32'h3c67d2fa),
	.w5(32'hbd126351),
	.w6(32'h3bc82d63),
	.w7(32'h3b1b9c7f),
	.w8(32'hbcbee43d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eef1a),
	.w1(32'hbb2a31d7),
	.w2(32'hbbcab451),
	.w3(32'hbca40959),
	.w4(32'h3bdbcc77),
	.w5(32'hbb744172),
	.w6(32'h3ac56928),
	.w7(32'h3beb17ea),
	.w8(32'h3c4cbba4),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8defc9),
	.w1(32'h3b0d6ef0),
	.w2(32'hbbd3c377),
	.w3(32'h3b1d37cd),
	.w4(32'h3bda882a),
	.w5(32'hbb0f6696),
	.w6(32'h3b6be1b4),
	.w7(32'h3b77dc3a),
	.w8(32'hbab25780),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3088c7),
	.w1(32'h3b6939e4),
	.w2(32'hbc406c0a),
	.w3(32'hbb10d81a),
	.w4(32'hbb70172d),
	.w5(32'h3a605d67),
	.w6(32'h3baf9511),
	.w7(32'h3b69f004),
	.w8(32'h3c400f84),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc613d92),
	.w1(32'h3bd81972),
	.w2(32'hbaea92ea),
	.w3(32'hbc1873b4),
	.w4(32'hbb80a8cb),
	.w5(32'h380ac5f2),
	.w6(32'h387cf815),
	.w7(32'h3a1d8432),
	.w8(32'hbc88e162),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7c84a),
	.w1(32'hbb4e1e8b),
	.w2(32'hbb77a947),
	.w3(32'hbc87d447),
	.w4(32'hbc0abaad),
	.w5(32'hbb4cce26),
	.w6(32'hbc2af484),
	.w7(32'h39ff9948),
	.w8(32'hbbeeae7d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d450a),
	.w1(32'hbbbebd90),
	.w2(32'hbcf8de4b),
	.w3(32'h3ba78b78),
	.w4(32'h3a0c517b),
	.w5(32'hbce2b477),
	.w6(32'hbb3c60e5),
	.w7(32'hbb713240),
	.w8(32'hbc8a4607),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb847d2a7),
	.w1(32'h3c48f735),
	.w2(32'h3c388996),
	.w3(32'h390eecdd),
	.w4(32'h3c0a89c4),
	.w5(32'h3b15ce2d),
	.w6(32'h3bb2775f),
	.w7(32'h3c3ff51e),
	.w8(32'h3c1cf083),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371c343b),
	.w1(32'hbaf7448f),
	.w2(32'hbc60858d),
	.w3(32'hbc0b546c),
	.w4(32'h3c360af6),
	.w5(32'h3b347b15),
	.w6(32'h3c156952),
	.w7(32'h3bb04ecd),
	.w8(32'hba0d436b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b508a4f),
	.w1(32'hbb7a4d04),
	.w2(32'hbcabf589),
	.w3(32'h3b9d7145),
	.w4(32'hb9f31880),
	.w5(32'hbc711721),
	.w6(32'h3be4b956),
	.w7(32'h3b43ea4d),
	.w8(32'hbc71e613),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b046b10),
	.w1(32'h3c23e39a),
	.w2(32'hbb20044a),
	.w3(32'h3bacb555),
	.w4(32'h3c9f854d),
	.w5(32'h3c52f874),
	.w6(32'hbb9a9bc6),
	.w7(32'h3bea071b),
	.w8(32'h3bdcb12e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad112da),
	.w1(32'h3bc24f44),
	.w2(32'hbc83f2d1),
	.w3(32'hbc92e0d6),
	.w4(32'hbbd24343),
	.w5(32'hbc688494),
	.w6(32'h3bdb59f9),
	.w7(32'hbb5be7ab),
	.w8(32'hbc3a17d6),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c0f0a),
	.w1(32'h3a2c3859),
	.w2(32'hbc309222),
	.w3(32'h3aabaa18),
	.w4(32'h3881a644),
	.w5(32'hbc551b0a),
	.w6(32'h3b8d3817),
	.w7(32'h3b17169b),
	.w8(32'hbbee90f2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaced4c),
	.w1(32'h3d1227f3),
	.w2(32'h3c2ae3ef),
	.w3(32'hbc192f58),
	.w4(32'h3c86d991),
	.w5(32'h3cee6dfc),
	.w6(32'hbc252ecc),
	.w7(32'h3c43b08f),
	.w8(32'h3d6cea45),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1c3901),
	.w1(32'hbc8b70d7),
	.w2(32'hbb56af70),
	.w3(32'hbc29ff27),
	.w4(32'hbc0b4f97),
	.w5(32'hb97f9800),
	.w6(32'h3c825e7c),
	.w7(32'h3cbcb720),
	.w8(32'h3b98307b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24c20c),
	.w1(32'hba881fa8),
	.w2(32'h3b29d3c2),
	.w3(32'hbbc2a200),
	.w4(32'hbb86d8ee),
	.w5(32'h3bb6dec6),
	.w6(32'hbadabd47),
	.w7(32'hba54572d),
	.w8(32'h3a91d66e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ff7c4),
	.w1(32'h3b90c50b),
	.w2(32'h3a947473),
	.w3(32'h3be0a2fe),
	.w4(32'h3bfcb3b0),
	.w5(32'h3b9e71f8),
	.w6(32'h3abb8992),
	.w7(32'h3b0eb809),
	.w8(32'h3c061adc),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb806046),
	.w1(32'hba0ff20e),
	.w2(32'hbb4f6278),
	.w3(32'h3b56beb0),
	.w4(32'h3a667229),
	.w5(32'hbb9379e0),
	.w6(32'h3b86c788),
	.w7(32'h3a7c3f10),
	.w8(32'hba05b43e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf49ce),
	.w1(32'h3c0f5d1e),
	.w2(32'hbbbe2a70),
	.w3(32'hbbc1cde1),
	.w4(32'h3c3eae50),
	.w5(32'h3b546c69),
	.w6(32'hbbf54d79),
	.w7(32'h3c2a3e64),
	.w8(32'h3c55afe1),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd00a6b1),
	.w1(32'hbc98b113),
	.w2(32'hbc0d15ba),
	.w3(32'hbcac7fb3),
	.w4(32'hbc369d47),
	.w5(32'hbaa29237),
	.w6(32'h3bfc58d9),
	.w7(32'h3b959935),
	.w8(32'hbc049a6e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73d55e0),
	.w1(32'h3b8b67c7),
	.w2(32'h3bacd444),
	.w3(32'hbb3fa82e),
	.w4(32'hbbb22e61),
	.w5(32'h3ac8930d),
	.w6(32'hbbc552f9),
	.w7(32'hbafdb269),
	.w8(32'h3a982f2e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8d3f0),
	.w1(32'h3c1984b3),
	.w2(32'hbc726435),
	.w3(32'hbbf22f2f),
	.w4(32'h3c089e8b),
	.w5(32'hbc3da6d7),
	.w6(32'h3b0fee92),
	.w7(32'h3be70888),
	.w8(32'hbc2a26f3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f2831),
	.w1(32'hbb283a1a),
	.w2(32'hba5bb663),
	.w3(32'hbc027d04),
	.w4(32'hba4cd0cf),
	.w5(32'h3b9d9c30),
	.w6(32'h3bda03a8),
	.w7(32'hbb3effc0),
	.w8(32'h3b42522e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e4e31),
	.w1(32'h3b2b39ad),
	.w2(32'hbce3d769),
	.w3(32'hbb0b6a2e),
	.w4(32'h3b758142),
	.w5(32'hbcc3212f),
	.w6(32'h3bedc990),
	.w7(32'h3badff68),
	.w8(32'hbc9bf9c7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0da030),
	.w1(32'h3c417630),
	.w2(32'hbaad934e),
	.w3(32'hbc18eec5),
	.w4(32'h3bee7617),
	.w5(32'h3c2056f6),
	.w6(32'hbc30f593),
	.w7(32'h3c57a5ba),
	.w8(32'h3cf63dce),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd305c24),
	.w1(32'hbc94ac9c),
	.w2(32'h3b910c0a),
	.w3(32'hbc784a3b),
	.w4(32'hbc86ec1d),
	.w5(32'h3c97932b),
	.w6(32'h3c7aafaf),
	.w7(32'h3c5370e0),
	.w8(32'h3c3d8d47),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c824eea),
	.w1(32'h3c62e135),
	.w2(32'h3aafd544),
	.w3(32'h3ccc6ec4),
	.w4(32'h3cbf8199),
	.w5(32'h3b0f8aec),
	.w6(32'h3c8a12b8),
	.w7(32'h3c871d5a),
	.w8(32'h3ae565ed),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbcf63),
	.w1(32'h3bb8908b),
	.w2(32'h3c519b7f),
	.w3(32'hbc4b5328),
	.w4(32'h3b797a27),
	.w5(32'h3b560ed2),
	.w6(32'hbc37807e),
	.w7(32'h3b8e28e5),
	.w8(32'h3b149c3a),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d5bb9),
	.w1(32'hbbd065c1),
	.w2(32'h3c715979),
	.w3(32'h3b9377c1),
	.w4(32'h3c456251),
	.w5(32'h3c32a321),
	.w6(32'hbb814a56),
	.w7(32'h3c8c5fe5),
	.w8(32'h3c476ac3),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce2153),
	.w1(32'h3c383d30),
	.w2(32'h3bf84c31),
	.w3(32'h3b410236),
	.w4(32'h3997f075),
	.w5(32'h3bf63580),
	.w6(32'h3c9e4986),
	.w7(32'h3c29358b),
	.w8(32'h3c371e37),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6092db),
	.w1(32'hbae51725),
	.w2(32'hbbd66c9c),
	.w3(32'hbc0119a5),
	.w4(32'hbb8b7f5f),
	.w5(32'hbc67b572),
	.w6(32'hbb1b1a76),
	.w7(32'hbbbbc73e),
	.w8(32'h39151992),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ece616),
	.w1(32'hbc140cb6),
	.w2(32'hbcae83af),
	.w3(32'hbc3e2f1a),
	.w4(32'hbc1114da),
	.w5(32'hbbf49739),
	.w6(32'hbc5aefe8),
	.w7(32'hbc892249),
	.w8(32'hbb560bf7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83881c),
	.w1(32'h3bfae990),
	.w2(32'hbc74e70c),
	.w3(32'hbbed6db9),
	.w4(32'hbab852a6),
	.w5(32'hbbd18a0b),
	.w6(32'hbbcbac0e),
	.w7(32'hbc866fba),
	.w8(32'hbb8fc4eb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4ee1c),
	.w1(32'h3a0c6cf5),
	.w2(32'hbb8ee839),
	.w3(32'h3ad269b1),
	.w4(32'hbadd4f44),
	.w5(32'hbac85a8c),
	.w6(32'h3bb4f427),
	.w7(32'h3bc85e36),
	.w8(32'h3c1f98ef),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3754d2),
	.w1(32'h3b181914),
	.w2(32'h3c50b6f4),
	.w3(32'hbcc6b220),
	.w4(32'hbc45e2fc),
	.w5(32'h3c71fbbf),
	.w6(32'hbc923027),
	.w7(32'hbb8c8efe),
	.w8(32'h3bb06dfe),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2e261),
	.w1(32'h3b7b313a),
	.w2(32'h3c0717e5),
	.w3(32'h3bb78a98),
	.w4(32'h3b10055a),
	.w5(32'h3ab18ba4),
	.w6(32'h3b86986e),
	.w7(32'h3bd8f72e),
	.w8(32'hbb52f551),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec688a),
	.w1(32'hbb8dfb95),
	.w2(32'hbbe539d5),
	.w3(32'h3c91c53c),
	.w4(32'hbbf0c70b),
	.w5(32'hbbd837b8),
	.w6(32'h38eebe38),
	.w7(32'hbc768956),
	.w8(32'hbc2dad78),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee6ea1),
	.w1(32'hbc0aa78c),
	.w2(32'h3c1dba2b),
	.w3(32'hbbaff197),
	.w4(32'hbc5b0c8f),
	.w5(32'h3cdede8b),
	.w6(32'hbbd22c45),
	.w7(32'hbb1360fb),
	.w8(32'hbc3a914a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c8cf1),
	.w1(32'hbb1f364b),
	.w2(32'hbc2874b9),
	.w3(32'h3d090688),
	.w4(32'hbbc9aff0),
	.w5(32'hbc5170e2),
	.w6(32'h3cc7c3b1),
	.w7(32'h3c1ef9eb),
	.w8(32'h3c9e4b8a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c591750),
	.w1(32'h3cd5366c),
	.w2(32'h3bf63f86),
	.w3(32'hbc973e0f),
	.w4(32'h3cbba62d),
	.w5(32'h3c3268ad),
	.w6(32'hbccff5d0),
	.w7(32'hb9d91d2a),
	.w8(32'h3c5ab335),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26a7bb),
	.w1(32'h3c65787e),
	.w2(32'hbc0ea854),
	.w3(32'hbb0e588f),
	.w4(32'h3c918a41),
	.w5(32'h3b70fef7),
	.w6(32'hba27f3ca),
	.w7(32'h3b3eaa7f),
	.w8(32'hbb26dd49),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc532f2b),
	.w1(32'h3c279177),
	.w2(32'h3b0d333a),
	.w3(32'hbbbb8e77),
	.w4(32'hbc2feb28),
	.w5(32'h3c59e105),
	.w6(32'h3c03a389),
	.w7(32'hbc60f52d),
	.w8(32'h3c032a81),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fc28e),
	.w1(32'h3bb247f1),
	.w2(32'h3b328d80),
	.w3(32'hbb3fccaf),
	.w4(32'hbbac6d4f),
	.w5(32'h3b80fa83),
	.w6(32'h3caf76c4),
	.w7(32'h3c016fca),
	.w8(32'hb905357f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc335cc),
	.w1(32'hbbae8106),
	.w2(32'hbb9169cb),
	.w3(32'h38f0f4b1),
	.w4(32'hbb868d85),
	.w5(32'hbbd5cf80),
	.w6(32'hb94570dd),
	.w7(32'h3b6713d6),
	.w8(32'h3bfdba91),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9466fb),
	.w1(32'hbbcde624),
	.w2(32'hbcc160be),
	.w3(32'hbc84dd99),
	.w4(32'h3b9711b6),
	.w5(32'hbcb72550),
	.w6(32'h3c0a843d),
	.w7(32'h3b292e91),
	.w8(32'hbc93a003),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8af8fe),
	.w1(32'hbc58d391),
	.w2(32'hbc433ef7),
	.w3(32'h3ac181fb),
	.w4(32'hbb00cf02),
	.w5(32'h3b9bf882),
	.w6(32'hbb0ee7df),
	.w7(32'h3b98e941),
	.w8(32'hbbfc801a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69e42a),
	.w1(32'hbc5ff6b5),
	.w2(32'hbc8b436d),
	.w3(32'h3c3e11f7),
	.w4(32'hbbf8cff2),
	.w5(32'hbb2ffe07),
	.w6(32'h3c70bcd0),
	.w7(32'h3ba630d3),
	.w8(32'hbbfe79a1),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f9743),
	.w1(32'h3c1d8c25),
	.w2(32'h3b763caa),
	.w3(32'h3c029e29),
	.w4(32'h3bc783ff),
	.w5(32'h3b1c4e5b),
	.w6(32'h3d052f4b),
	.w7(32'h3b7791ee),
	.w8(32'hba87adb4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3011b1),
	.w1(32'hba4f5cbd),
	.w2(32'hbc28676f),
	.w3(32'hbaef980c),
	.w4(32'h3a8766b0),
	.w5(32'hbc5a5d4d),
	.w6(32'hbb8ad655),
	.w7(32'hba5cdc67),
	.w8(32'hbca48801),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ecf09),
	.w1(32'hbbb1ffbe),
	.w2(32'h3c0a87d2),
	.w3(32'hbbdbe4b3),
	.w4(32'hbb880d8b),
	.w5(32'hba159831),
	.w6(32'hbb0412ed),
	.w7(32'h3a66e296),
	.w8(32'h3bca5f70),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5484b5),
	.w1(32'hbb2e4b40),
	.w2(32'h3c8dfd88),
	.w3(32'h3b09b49d),
	.w4(32'h3ad8911d),
	.w5(32'h3bb20c34),
	.w6(32'h3bfee79a),
	.w7(32'h3ba407ec),
	.w8(32'h3aa94a06),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43de26),
	.w1(32'hba540f3b),
	.w2(32'h3b8458b2),
	.w3(32'h3ba75d03),
	.w4(32'hbb9cb128),
	.w5(32'h3b9f644d),
	.w6(32'h3be826ce),
	.w7(32'h3b85d038),
	.w8(32'h3bb8c720),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62752e),
	.w1(32'hbb89be52),
	.w2(32'hbc9f97ce),
	.w3(32'hbc28b840),
	.w4(32'hbc5f1e29),
	.w5(32'hbcaa3920),
	.w6(32'h3ab415f8),
	.w7(32'hbb912ce8),
	.w8(32'hbb09e11a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd338a),
	.w1(32'h3bf790bf),
	.w2(32'hbb0ebf05),
	.w3(32'h3930858e),
	.w4(32'h3c41fa3f),
	.w5(32'h3a0cbf2a),
	.w6(32'hbb22ee71),
	.w7(32'h3c152993),
	.w8(32'h3b7c7a11),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c085729),
	.w1(32'h3bc73859),
	.w2(32'hbb44ee44),
	.w3(32'hbc39373e),
	.w4(32'h3b8f77dd),
	.w5(32'hbc1053de),
	.w6(32'hbc7111b5),
	.w7(32'h3a876582),
	.w8(32'h3ad6860d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5bf7e),
	.w1(32'h3c75c2c9),
	.w2(32'hbb4616d0),
	.w3(32'hbcb537d3),
	.w4(32'h3b561ea3),
	.w5(32'h3c48fee5),
	.w6(32'hbc9a31f6),
	.w7(32'hbc0a6bfd),
	.w8(32'h3c6ba263),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf8a79c),
	.w1(32'hbc6c2958),
	.w2(32'hbc53fd24),
	.w3(32'hbc054299),
	.w4(32'hbcd81989),
	.w5(32'hbc67ea33),
	.w6(32'h3cbd2fac),
	.w7(32'h3a62da54),
	.w8(32'hbbe882f4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09fd87),
	.w1(32'h3ab5a4e6),
	.w2(32'hbc4a9f45),
	.w3(32'hbc801bd1),
	.w4(32'h3c12c119),
	.w5(32'hbbc8d231),
	.w6(32'hbc0cc7c1),
	.w7(32'h3b3c6e64),
	.w8(32'h3abae163),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5c04b),
	.w1(32'h3ba69b06),
	.w2(32'h3a9a5391),
	.w3(32'h3b87be7b),
	.w4(32'h3bac926a),
	.w5(32'h3bb622a4),
	.w6(32'h3ab2a7a1),
	.w7(32'h3c2170c5),
	.w8(32'hbb188596),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba72ee6),
	.w1(32'hbaf2f4e1),
	.w2(32'hbd513262),
	.w3(32'h3c0772f9),
	.w4(32'hbbfc98fc),
	.w5(32'hbd28ecf9),
	.w6(32'h3bac912a),
	.w7(32'hbca0c3bf),
	.w8(32'hbd04a49a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b013b),
	.w1(32'h3cf7af5e),
	.w2(32'h3c1c0b1d),
	.w3(32'hbcf86b60),
	.w4(32'h3c9a9255),
	.w5(32'h3d066070),
	.w6(32'hbcb6b8f7),
	.w7(32'h3aa41ed6),
	.w8(32'h3cad33a8),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd9a923),
	.w1(32'hbba9e7f8),
	.w2(32'hbc4affaa),
	.w3(32'h3cf65c16),
	.w4(32'h3cb1e046),
	.w5(32'hbbb7a0f8),
	.w6(32'h3d06f711),
	.w7(32'h3d0a46b6),
	.w8(32'hbc35a0c8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc53e67),
	.w1(32'h3b5ec1e7),
	.w2(32'hbbf2a0ea),
	.w3(32'hbbf2ae4d),
	.w4(32'hbbac97bb),
	.w5(32'hbb625f8b),
	.w6(32'hbad0aff9),
	.w7(32'hbb86dcc6),
	.w8(32'hbbc65944),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f4435),
	.w1(32'hbbc5a03f),
	.w2(32'h3c595a1d),
	.w3(32'hbbb86d67),
	.w4(32'hbbe6917e),
	.w5(32'h3c7d6255),
	.w6(32'hbc250f87),
	.w7(32'hbc193a16),
	.w8(32'h3bc51b67),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35a3aa),
	.w1(32'h3c4b83a5),
	.w2(32'h3b160380),
	.w3(32'h3c972df7),
	.w4(32'h3c37834a),
	.w5(32'hbae30b31),
	.w6(32'h3c60d797),
	.w7(32'h3bf105c5),
	.w8(32'hbac41de6),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967a23),
	.w1(32'hba9edfed),
	.w2(32'hbc598542),
	.w3(32'h3ba041e9),
	.w4(32'h3b80e417),
	.w5(32'hbc1d29dd),
	.w6(32'h3b28be4b),
	.w7(32'h3bf057af),
	.w8(32'hbc05e7f4),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a6d9c),
	.w1(32'hbbb3f921),
	.w2(32'h3c11ab13),
	.w3(32'h3c57fd76),
	.w4(32'h3b88fea8),
	.w5(32'h3c6f35bf),
	.w6(32'h3bee2cc4),
	.w7(32'h3c2f9679),
	.w8(32'h3c1e793f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad05e63),
	.w1(32'h3c7ec767),
	.w2(32'h3bd96d72),
	.w3(32'hbb3e0ae8),
	.w4(32'h3c5cdd3b),
	.w5(32'h3c0eb4b3),
	.w6(32'hba1597ee),
	.w7(32'h3c03ca58),
	.w8(32'h3bb8bb66),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41e4a6),
	.w1(32'h3bcaffe6),
	.w2(32'hba855dc5),
	.w3(32'h3c171019),
	.w4(32'h3bac1c07),
	.w5(32'hba30d967),
	.w6(32'h3b0d797a),
	.w7(32'h3be8f600),
	.w8(32'h3b073860),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ac8b0),
	.w1(32'hbc0d305c),
	.w2(32'hbcc2b4a7),
	.w3(32'hbbc9545e),
	.w4(32'hbbcbbeda),
	.w5(32'hbc8f8758),
	.w6(32'hbb3218f0),
	.w7(32'hbbdf975f),
	.w8(32'hbcccc60e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28af86),
	.w1(32'h3bcdf5d8),
	.w2(32'hbbfc6442),
	.w3(32'hbc59ee3c),
	.w4(32'hbc16a45d),
	.w5(32'hbc65e367),
	.w6(32'hbb9ed938),
	.w7(32'hbca10bb5),
	.w8(32'hbbba95e2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c215e80),
	.w1(32'hbbde8562),
	.w2(32'h3b2b4ff2),
	.w3(32'h3b46342e),
	.w4(32'h3c09e14c),
	.w5(32'h3ae0bdab),
	.w6(32'hbc4a666a),
	.w7(32'h3ab95a4e),
	.w8(32'hbac88338),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc67a4),
	.w1(32'hba2ec65f),
	.w2(32'hbc9ed790),
	.w3(32'hba90f654),
	.w4(32'h3ae54ae5),
	.w5(32'hbc9c07c7),
	.w6(32'hbb512afc),
	.w7(32'hbc417aff),
	.w8(32'hbc772eca),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4cac5),
	.w1(32'hbc30ae9d),
	.w2(32'h389399d5),
	.w3(32'hbc554835),
	.w4(32'hbc8cf1dc),
	.w5(32'h3968ae03),
	.w6(32'hbbdf36aa),
	.w7(32'hbc340b9d),
	.w8(32'hba424d40),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2347e4),
	.w1(32'hbc2f6257),
	.w2(32'hbbd38bcf),
	.w3(32'hbc141a5a),
	.w4(32'hbc307c1c),
	.w5(32'hbb5148d6),
	.w6(32'hbc2eac73),
	.w7(32'hbc0f6385),
	.w8(32'hbbaf2c8f),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28e976),
	.w1(32'h3bfc3f03),
	.w2(32'h3c60dc9e),
	.w3(32'hbc027ff3),
	.w4(32'h3ba6daab),
	.w5(32'h3c0e9d60),
	.w6(32'hbbc268d2),
	.w7(32'h3b0a9dc7),
	.w8(32'h3c205a29),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb958b2f7),
	.w1(32'h3b8aec20),
	.w2(32'h3c50c56c),
	.w3(32'hbba76c43),
	.w4(32'hbb358c6d),
	.w5(32'h3ab5de5c),
	.w6(32'hbb89204e),
	.w7(32'h38c2c535),
	.w8(32'hba6cd614),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d52358),
	.w1(32'hbb6cf623),
	.w2(32'hbbb21077),
	.w3(32'hbb4244eb),
	.w4(32'h3b72ffc2),
	.w5(32'h3c1b6ff0),
	.w6(32'h3bf05aa4),
	.w7(32'h3b537bbd),
	.w8(32'h3c71ba18),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96583c),
	.w1(32'h3c821f02),
	.w2(32'h3c23bd67),
	.w3(32'hbc8ad01f),
	.w4(32'h3aed36bc),
	.w5(32'h3c1d4b1b),
	.w6(32'hbbc71c01),
	.w7(32'hbbe1acf8),
	.w8(32'h3c3df5fb),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf38c6),
	.w1(32'h3b820cb2),
	.w2(32'hbc4129c9),
	.w3(32'hbba23e0b),
	.w4(32'h3b3a5df7),
	.w5(32'hbc030721),
	.w6(32'h3b270b19),
	.w7(32'h3b74c51a),
	.w8(32'hbbfdb529),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3176f6),
	.w1(32'hbb5a3dbc),
	.w2(32'hbc189a7c),
	.w3(32'hbc0c8e74),
	.w4(32'hbc7ba1f5),
	.w5(32'hbbc81a5c),
	.w6(32'h3b408c53),
	.w7(32'hbbffca63),
	.w8(32'hbb246eed),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f7a3a),
	.w1(32'hbaacc5b4),
	.w2(32'h3b8579ef),
	.w3(32'hba20bfbb),
	.w4(32'hbac3cf79),
	.w5(32'h3a898ac5),
	.w6(32'h39fa1e1b),
	.w7(32'h3aae8c83),
	.w8(32'h3a641938),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35fe94),
	.w1(32'hbb2f5987),
	.w2(32'h3c97bfd1),
	.w3(32'hbb6524c5),
	.w4(32'hbbcc780b),
	.w5(32'h3b016af3),
	.w6(32'hbbebd1a4),
	.w7(32'hbbe45aa1),
	.w8(32'hbcc421e3),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc59f32),
	.w1(32'hbb1121ca),
	.w2(32'hbc6efea9),
	.w3(32'h3d42a1de),
	.w4(32'h3d40de64),
	.w5(32'hbb2d9177),
	.w6(32'h3aa5394e),
	.w7(32'h3d0ad9bf),
	.w8(32'hbca05011),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d38e3),
	.w1(32'hbb7a3d10),
	.w2(32'hbc9651ca),
	.w3(32'h3c1aa592),
	.w4(32'h3be5581f),
	.w5(32'hbca24dff),
	.w6(32'h3b3d7ed0),
	.w7(32'h3af9c5e0),
	.w8(32'hbc3be56f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc697433),
	.w1(32'h3bdad5df),
	.w2(32'hba193686),
	.w3(32'hbcae58c7),
	.w4(32'h3c30a582),
	.w5(32'hbafa4161),
	.w6(32'hbcb63604),
	.w7(32'h3b4bca36),
	.w8(32'h3a73ceba),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0014f7),
	.w1(32'hbb05a07f),
	.w2(32'hbd246ed4),
	.w3(32'hbc3e04ce),
	.w4(32'h3c0e325b),
	.w5(32'hbce7b365),
	.w6(32'hbbae9c3a),
	.w7(32'h3ba398f2),
	.w8(32'hbc916604),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9da199),
	.w1(32'h3a7a56e7),
	.w2(32'h3bf41416),
	.w3(32'h3935da4c),
	.w4(32'hba2f62d6),
	.w5(32'h3bbb98d9),
	.w6(32'hba4c3621),
	.w7(32'hba166640),
	.w8(32'h39934d43),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c883a3b),
	.w1(32'hbb8a4cdb),
	.w2(32'hba7c6460),
	.w3(32'h3be2ae18),
	.w4(32'h3b0a7e15),
	.w5(32'hbc240bac),
	.w6(32'h3aac69b8),
	.w7(32'hba0bfa0a),
	.w8(32'hbc19745b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d16da),
	.w1(32'h3ceb188d),
	.w2(32'hbcd3dcbf),
	.w3(32'h3c0d67eb),
	.w4(32'h3d6a7d47),
	.w5(32'hbcaad1ca),
	.w6(32'hbcae32e9),
	.w7(32'h3cafe8a0),
	.w8(32'hbbf27234),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f417a),
	.w1(32'hbc2395e8),
	.w2(32'hbd0336a9),
	.w3(32'h3c66585e),
	.w4(32'h3b5bbd7e),
	.w5(32'hbcb289cd),
	.w6(32'hbc4496e9),
	.w7(32'hbbc1bb3d),
	.w8(32'hbcb8fc6f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d1ad4),
	.w1(32'hbad29a51),
	.w2(32'hbca95a27),
	.w3(32'h3bade7b8),
	.w4(32'h3c8aa688),
	.w5(32'hbc8ddf2e),
	.w6(32'h3bc3715b),
	.w7(32'h3c4c66b5),
	.w8(32'hbc394eed),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25b309),
	.w1(32'h3c3a95fc),
	.w2(32'h3c9c9af6),
	.w3(32'hbc23ed49),
	.w4(32'h3b830693),
	.w5(32'h3ca661ce),
	.w6(32'h3a511d2d),
	.w7(32'h3c21abc7),
	.w8(32'h3ce03312),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce934f),
	.w1(32'h3c407427),
	.w2(32'h3c881e84),
	.w3(32'hbc8ed490),
	.w4(32'h3b99fd65),
	.w5(32'h3c9c2037),
	.w6(32'hbb816e18),
	.w7(32'h3af56c9a),
	.w8(32'h3c13d938),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0904bd),
	.w1(32'hba8db2b9),
	.w2(32'h3989553b),
	.w3(32'h3c344513),
	.w4(32'h3b9b460b),
	.w5(32'hbaa4d105),
	.w6(32'h3ba04639),
	.w7(32'h3a23d91e),
	.w8(32'h3b739d44),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bf478),
	.w1(32'h3bd65dec),
	.w2(32'h3b8f339c),
	.w3(32'hbc0c0187),
	.w4(32'hbb184ce4),
	.w5(32'h3b3f7386),
	.w6(32'hbb491d33),
	.w7(32'h3b4202af),
	.w8(32'h399535d5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcc54d),
	.w1(32'h3b0f4bdb),
	.w2(32'hba0a3662),
	.w3(32'hbb8c11d8),
	.w4(32'hbb28d915),
	.w5(32'h3c1f3a2e),
	.w6(32'hbc0977df),
	.w7(32'hbbb16a4c),
	.w8(32'hbbe3c9eb),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bd9a8),
	.w1(32'hbb88e741),
	.w2(32'h3c32bb96),
	.w3(32'h3c4c8c3f),
	.w4(32'h3c013ee5),
	.w5(32'h399bb717),
	.w6(32'h3ca8106e),
	.w7(32'h3bfdaf19),
	.w8(32'h3b772917),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3da4b),
	.w1(32'hba3ee10b),
	.w2(32'hbbdf1a9f),
	.w3(32'hbb1133e5),
	.w4(32'hbc3684a9),
	.w5(32'h3aa46097),
	.w6(32'hba9899c0),
	.w7(32'h3b13e611),
	.w8(32'hbc2a4c41),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc165b81),
	.w1(32'h3b0fa06f),
	.w2(32'hbc377552),
	.w3(32'h3b273eec),
	.w4(32'hbbdbb603),
	.w5(32'hbc1c5e9e),
	.w6(32'hbb0cdf0a),
	.w7(32'hbc55c806),
	.w8(32'hbc25359c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b103b05),
	.w1(32'h3bdd23dc),
	.w2(32'h3c1460db),
	.w3(32'hbc088eb7),
	.w4(32'h3ac1b919),
	.w5(32'h3bf28b79),
	.w6(32'h3b449f31),
	.w7(32'hbb8233b7),
	.w8(32'h3ba79fd1),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c217123),
	.w1(32'h3c224671),
	.w2(32'h3bb80a88),
	.w3(32'h3b033a63),
	.w4(32'hbb190495),
	.w5(32'h3bc2a101),
	.w6(32'h3adc81ef),
	.w7(32'hbad131ad),
	.w8(32'h3b9c0768),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82c318),
	.w1(32'h3bd7ce7a),
	.w2(32'hbd2ef070),
	.w3(32'hbb8737f5),
	.w4(32'h3bc8a2c3),
	.w5(32'hbd027b3c),
	.w6(32'hbc152b41),
	.w7(32'h3bf0712f),
	.w8(32'hbc88683e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb271159),
	.w1(32'h3c38ed65),
	.w2(32'hbc4f4ff2),
	.w3(32'hba57152f),
	.w4(32'h3c1bc1d5),
	.w5(32'hbbfcb11a),
	.w6(32'h3af57df0),
	.w7(32'hbba65f4f),
	.w8(32'hbc43c8c7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2dced),
	.w1(32'h3b980832),
	.w2(32'h3b40fa76),
	.w3(32'hbb7522a3),
	.w4(32'h3b39b5ca),
	.w5(32'hbafde942),
	.w6(32'h3aae1d5c),
	.w7(32'hbb8ba64f),
	.w8(32'h3bb6cb7c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61428b),
	.w1(32'h3b8c2b07),
	.w2(32'hbc826376),
	.w3(32'h3c0a5664),
	.w4(32'h3c2ced68),
	.w5(32'hbc8bbfd0),
	.w6(32'hbabadd36),
	.w7(32'h399ec7c5),
	.w8(32'hbc48b68f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed2106),
	.w1(32'h3aa0d92f),
	.w2(32'hbaebc3ae),
	.w3(32'hb9806576),
	.w4(32'h3bd797a3),
	.w5(32'h3c0f38ee),
	.w6(32'hbc396fd2),
	.w7(32'h3b00ae99),
	.w8(32'hbb47f1ae),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82ba91),
	.w1(32'hbc2a8270),
	.w2(32'hbbed963d),
	.w3(32'h3b2bfa78),
	.w4(32'hbc4eacd5),
	.w5(32'h3c18b6c5),
	.w6(32'h3bf918c3),
	.w7(32'hbab95929),
	.w8(32'h3bf372c6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee8b93),
	.w1(32'h3c849fd1),
	.w2(32'hbc4ddcd7),
	.w3(32'h3c025c5a),
	.w4(32'h3bb74c01),
	.w5(32'hbc4f3804),
	.w6(32'h3bd4432a),
	.w7(32'h3bae7327),
	.w8(32'hbc373249),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf8f59),
	.w1(32'hbb9a1539),
	.w2(32'hba4c8ebd),
	.w3(32'hbbd8a42b),
	.w4(32'h3b605701),
	.w5(32'h3b4da96b),
	.w6(32'hbc29994a),
	.w7(32'hbbea94a5),
	.w8(32'h3ae6e0e2),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25daf0),
	.w1(32'h3b06ce81),
	.w2(32'h39808ec5),
	.w3(32'h3c427098),
	.w4(32'h3b242587),
	.w5(32'h3bbff9df),
	.w6(32'h3c2b727e),
	.w7(32'h3c30984a),
	.w8(32'h3c7127b3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc829884),
	.w1(32'hbc975e8f),
	.w2(32'hbce83e35),
	.w3(32'hbcb52079),
	.w4(32'hbc93225c),
	.w5(32'hbca373f6),
	.w6(32'h3ba45cf1),
	.w7(32'hbc450bec),
	.w8(32'hbca84636),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d18cc),
	.w1(32'h3bc0e813),
	.w2(32'hbc71e4af),
	.w3(32'h3b6f9488),
	.w4(32'h3abd43a7),
	.w5(32'hbc205e75),
	.w6(32'hbb5c5685),
	.w7(32'hbb5a7328),
	.w8(32'hb8042e15),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c2fca),
	.w1(32'h3b81420a),
	.w2(32'hbb967537),
	.w3(32'h3cecb82b),
	.w4(32'h3c512094),
	.w5(32'hbc06ae34),
	.w6(32'h3cb53972),
	.w7(32'h3ca8e31a),
	.w8(32'hbc840de4),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9060316),
	.w1(32'hbc359991),
	.w2(32'hbaf4dee4),
	.w3(32'h3c07e7bc),
	.w4(32'hbb85daef),
	.w5(32'h3b89596e),
	.w6(32'h3c645e11),
	.w7(32'h3b1ebf82),
	.w8(32'hbbd54cfb),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4cd50d),
	.w1(32'hbbad4bc2),
	.w2(32'hbb6b4583),
	.w3(32'h37886e66),
	.w4(32'hbbecccc7),
	.w5(32'hbb9b84ec),
	.w6(32'hb9060922),
	.w7(32'hbba97a89),
	.w8(32'h3c514d56),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21f527),
	.w1(32'hbc9263ad),
	.w2(32'hb965dac2),
	.w3(32'hbaf84d10),
	.w4(32'h3b954b40),
	.w5(32'h3b4be92b),
	.w6(32'hbb096ea4),
	.w7(32'h3b848fc2),
	.w8(32'h3baaaea8),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97aee3),
	.w1(32'h3bc18ddf),
	.w2(32'hbc170774),
	.w3(32'h3b351c6e),
	.w4(32'h3a54c85a),
	.w5(32'h3bb48d3c),
	.w6(32'h3bdd5118),
	.w7(32'h3aac73b0),
	.w8(32'h3b14d1a0),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb463e),
	.w1(32'h3bec973f),
	.w2(32'hbc5bde2c),
	.w3(32'hbc83de0c),
	.w4(32'hbc477fcc),
	.w5(32'hbc12c602),
	.w6(32'hbc25d48c),
	.w7(32'hbc5b5b78),
	.w8(32'hbc1b6e80),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fb510),
	.w1(32'h3bf87282),
	.w2(32'hbc249879),
	.w3(32'hbbaa8851),
	.w4(32'hb9d5144f),
	.w5(32'hbc3db34a),
	.w6(32'h3bdf6f4a),
	.w7(32'hbba9b614),
	.w8(32'hbb3beae2),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90284ab),
	.w1(32'hbae4a2f7),
	.w2(32'hba0472cc),
	.w3(32'hbbe700ed),
	.w4(32'hbb5c1d6e),
	.w5(32'hb957b2c2),
	.w6(32'hbba97f36),
	.w7(32'hbc14f57f),
	.w8(32'hba9f38ff),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ae4de),
	.w1(32'hbb5f9580),
	.w2(32'hbbbc26a2),
	.w3(32'hbb2cbe5b),
	.w4(32'hbbc9eb20),
	.w5(32'hbb71cabf),
	.w6(32'hbac82eaa),
	.w7(32'hbb855119),
	.w8(32'hb8bb3383),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00faa7),
	.w1(32'hba099f7b),
	.w2(32'h3a0261ea),
	.w3(32'hbbe2cc24),
	.w4(32'hbb8835ff),
	.w5(32'hbc94e7cc),
	.w6(32'hba5d346c),
	.w7(32'hbbb5a216),
	.w8(32'hbc18e2ca),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c9d01),
	.w1(32'hba3ebf2a),
	.w2(32'hbb53b28e),
	.w3(32'hb9b1c7e4),
	.w4(32'h3c7dda94),
	.w5(32'hbbbc14ef),
	.w6(32'hbce86fd1),
	.w7(32'hbbfdcadc),
	.w8(32'hbb600269),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dfe20),
	.w1(32'h3b93848d),
	.w2(32'h3bf3ff08),
	.w3(32'h398a8d56),
	.w4(32'h3bbf7caf),
	.w5(32'hb9d8a7dd),
	.w6(32'hbb146017),
	.w7(32'h3afd8dea),
	.w8(32'h3badfa32),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84f41f),
	.w1(32'h3c138cb2),
	.w2(32'hbd270a8f),
	.w3(32'h3b2f7390),
	.w4(32'h3c8bec2f),
	.w5(32'hbc92d912),
	.w6(32'h3ba2fc29),
	.w7(32'h3bf03a01),
	.w8(32'hbc5fff2d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b387ac5),
	.w1(32'h3a1bdf1f),
	.w2(32'h3b4c9848),
	.w3(32'h3be70f0a),
	.w4(32'hb905389d),
	.w5(32'h3b89db1f),
	.w6(32'h3a6a47f7),
	.w7(32'h3878b42b),
	.w8(32'h3c0e6959),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0d504),
	.w1(32'h3c3d517b),
	.w2(32'h3bd36b87),
	.w3(32'hbca8a6c4),
	.w4(32'hbb7e8bdd),
	.w5(32'h3c06e063),
	.w6(32'hbc437625),
	.w7(32'hbc29317c),
	.w8(32'h3b693930),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule