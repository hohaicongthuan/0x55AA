module layer_10_featuremap_296(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada5cee),
	.w1(32'h3b1f7d51),
	.w2(32'h3aeef7c9),
	.w3(32'h3ae4d686),
	.w4(32'h3a4cea8d),
	.w5(32'h3a7c08b4),
	.w6(32'h3b197173),
	.w7(32'h3aa0885b),
	.w8(32'h3a3975fb),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb565df5),
	.w1(32'hbacc0c3f),
	.w2(32'hba89121e),
	.w3(32'hbb0cc84a),
	.w4(32'h3a78141f),
	.w5(32'h3920ed27),
	.w6(32'hbb62a2a1),
	.w7(32'hbaad7365),
	.w8(32'hbafaf658),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb804a997),
	.w1(32'h38bc6d89),
	.w2(32'hb9a41f1c),
	.w3(32'hb7cb1708),
	.w4(32'hb9d2e46e),
	.w5(32'hb9ef7fb7),
	.w6(32'hb98e12a9),
	.w7(32'hba087053),
	.w8(32'hba183fcc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f0569),
	.w1(32'h3a088808),
	.w2(32'h3a277faa),
	.w3(32'hba50cc47),
	.w4(32'h382e35b2),
	.w5(32'hbac27dd8),
	.w6(32'hbaa57ae2),
	.w7(32'hb8885b70),
	.w8(32'hbade164f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d77d9),
	.w1(32'hb99e805f),
	.w2(32'h3a4e6360),
	.w3(32'hbb3222ca),
	.w4(32'hba773f0d),
	.w5(32'hba1555df),
	.w6(32'hbb3f744d),
	.w7(32'hba9c36fd),
	.w8(32'hb9fa0b68),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb945b936),
	.w1(32'h380a9581),
	.w2(32'h39bec4cf),
	.w3(32'hba01e0ad),
	.w4(32'hb94b6958),
	.w5(32'h3a9de353),
	.w6(32'hba6a7b2f),
	.w7(32'hb95958e1),
	.w8(32'h3aa12353),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b287614),
	.w1(32'hbb23198d),
	.w2(32'hbb750e1e),
	.w3(32'h3ac54a00),
	.w4(32'hbb5a75e5),
	.w5(32'hbbd02f62),
	.w6(32'h3af04017),
	.w7(32'hb88ed481),
	.w8(32'hbb8d5fc3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc652068),
	.w1(32'hbc130b50),
	.w2(32'hbbd87aa2),
	.w3(32'hbc08356b),
	.w4(32'hbbdda76c),
	.w5(32'hbb2ad1dd),
	.w6(32'hbbff7905),
	.w7(32'hba7e4218),
	.w8(32'h3a2b0c63),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cc15d),
	.w1(32'hbab2f6bd),
	.w2(32'hb9eec958),
	.w3(32'hbb66e258),
	.w4(32'hbb06f3b3),
	.w5(32'hbb79a72a),
	.w6(32'hbb3f6b54),
	.w7(32'hba371a46),
	.w8(32'hbb4c2bad),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6b9f2),
	.w1(32'hbb70a7cd),
	.w2(32'hbbf3eca1),
	.w3(32'hbbe39374),
	.w4(32'hbb9a6f8c),
	.w5(32'hbba35a50),
	.w6(32'hbc3de1bb),
	.w7(32'hbc088bee),
	.w8(32'hbbf5951b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9372a86),
	.w1(32'h3897c7c5),
	.w2(32'h3a9514c0),
	.w3(32'hb907ec67),
	.w4(32'h3a7c8f65),
	.w5(32'h3a550e72),
	.w6(32'hbab6e081),
	.w7(32'h3609957e),
	.w8(32'h389f3a64),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba394a5),
	.w1(32'h3a55569a),
	.w2(32'hba9e6900),
	.w3(32'h3b683d6a),
	.w4(32'h3a2dba4a),
	.w5(32'hba5659bf),
	.w6(32'h3b1471d7),
	.w7(32'h3a809956),
	.w8(32'h3ab80cbf),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ee30d),
	.w1(32'hb9b4b4a1),
	.w2(32'hbb1ef73a),
	.w3(32'h3a9a11f3),
	.w4(32'h3a8d1d4f),
	.w5(32'hbb36eecb),
	.w6(32'hbb197fe2),
	.w7(32'hba270b86),
	.w8(32'hbb8a2272),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c6c18),
	.w1(32'hbba05dee),
	.w2(32'hbbacc8cd),
	.w3(32'hbb28fb60),
	.w4(32'hbb4da046),
	.w5(32'hbb20b553),
	.w6(32'hbb142a54),
	.w7(32'hbb0f1350),
	.w8(32'hbb1c59ba),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4db8d),
	.w1(32'hba7fad2e),
	.w2(32'hba2340ae),
	.w3(32'hbb5895b9),
	.w4(32'hb8f3dd28),
	.w5(32'h3a7179c7),
	.w6(32'hbb9eeb7d),
	.w7(32'hbb0aebeb),
	.w8(32'hbaaa1e94),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc005c07),
	.w1(32'hbbb29840),
	.w2(32'hbc0a5aac),
	.w3(32'hbc166f5d),
	.w4(32'hbb4d77f8),
	.w5(32'hbb6c9f28),
	.w6(32'hbc0c61d8),
	.w7(32'hbb5cb48f),
	.w8(32'hbba9a181),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e4a34),
	.w1(32'h3aa5c6ee),
	.w2(32'h3aa89b4b),
	.w3(32'hba49cfd5),
	.w4(32'h3a922186),
	.w5(32'h3b1a69e7),
	.w6(32'hba4372db),
	.w7(32'h3a7aef27),
	.w8(32'h3af3df18),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb67349),
	.w1(32'hbb36c256),
	.w2(32'hbb97b134),
	.w3(32'hbb69ef49),
	.w4(32'hbaed5379),
	.w5(32'hbbe1ddcd),
	.w6(32'hbbb8c15d),
	.w7(32'hba54c163),
	.w8(32'hbbf8c919),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec273b),
	.w1(32'hbacbff98),
	.w2(32'hbb6d0765),
	.w3(32'hbacac3c9),
	.w4(32'hb9dfee89),
	.w5(32'hbb7d208c),
	.w6(32'hbb2e7446),
	.w7(32'hbaf450fb),
	.w8(32'hbb987271),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d39540),
	.w1(32'hb98a4165),
	.w2(32'hb98c6e62),
	.w3(32'h38a0cb3d),
	.w4(32'h399845ea),
	.w5(32'h3a4c1a82),
	.w6(32'hb7f47f2e),
	.w7(32'h38690acf),
	.w8(32'h396ce72f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39303e01),
	.w1(32'h3a01bf53),
	.w2(32'h384ade5d),
	.w3(32'h3ab9f82e),
	.w4(32'h3ab48ddd),
	.w5(32'hb9da6183),
	.w6(32'h3a3d96ac),
	.w7(32'h38282881),
	.w8(32'hb98c06b0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3685a),
	.w1(32'h3a8abfab),
	.w2(32'h3a977190),
	.w3(32'hb939b85e),
	.w4(32'h3abcbb1a),
	.w5(32'h39389b65),
	.w6(32'hb7192b3c),
	.w7(32'h3a999108),
	.w8(32'hb90ead14),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9f195),
	.w1(32'hbbbe0466),
	.w2(32'hbbe47486),
	.w3(32'hbc17fe4d),
	.w4(32'hbb3ff2dc),
	.w5(32'hbc1758e6),
	.w6(32'hbc0f7cb2),
	.w7(32'hbb9f8fdc),
	.w8(32'hbc5fabfd),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947649),
	.w1(32'hba9e872e),
	.w2(32'hbb130a7e),
	.w3(32'hbb7b0629),
	.w4(32'h3a03f81b),
	.w5(32'hbb3e739a),
	.w6(32'hbbfd3597),
	.w7(32'hbaf9dbe9),
	.w8(32'hbbacd8f0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2392b8),
	.w1(32'h3b3294a0),
	.w2(32'h3a125032),
	.w3(32'hbb9d91bf),
	.w4(32'h3b231d60),
	.w5(32'hba8ec076),
	.w6(32'hbc0c5a4d),
	.w7(32'hbb50e6bb),
	.w8(32'hbb8e9ab3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba530072),
	.w1(32'hba5f7fa4),
	.w2(32'hba8b28d5),
	.w3(32'hbad4d0c1),
	.w4(32'hbac89b28),
	.w5(32'h383b0eae),
	.w6(32'hbab14fbe),
	.w7(32'hba9dd5db),
	.w8(32'h3a8d77a6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b797f),
	.w1(32'h3a1bd737),
	.w2(32'hb9fa76eb),
	.w3(32'h39f3683d),
	.w4(32'hb9cf1c08),
	.w5(32'h3aafbbb1),
	.w6(32'h3a67a377),
	.w7(32'hba1343d7),
	.w8(32'h3ad00636),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16385a),
	.w1(32'h3b54750a),
	.w2(32'h3afa524f),
	.w3(32'h39c1846c),
	.w4(32'h3b49cce5),
	.w5(32'hbb00f3b7),
	.w6(32'h3ac808de),
	.w7(32'h3b58eaeb),
	.w8(32'hba35699b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b284a),
	.w1(32'h3b6cbe93),
	.w2(32'h3b330071),
	.w3(32'h3bc054ef),
	.w4(32'h3bd0a7c3),
	.w5(32'h3ba6a663),
	.w6(32'h3bee5c23),
	.w7(32'h3bf93b9c),
	.w8(32'h3bdfc8dc),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8f3f3),
	.w1(32'h3a34d438),
	.w2(32'hb8d2152a),
	.w3(32'hbbfb14c4),
	.w4(32'hbb826dce),
	.w5(32'hbbab7515),
	.w6(32'hbc24a1d1),
	.w7(32'hbbcf7499),
	.w8(32'hbbd70ce5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f10d6d),
	.w1(32'h3ab7f788),
	.w2(32'h3a601f35),
	.w3(32'hba6c2dae),
	.w4(32'h39282253),
	.w5(32'h3a8cb688),
	.w6(32'h39c40dbf),
	.w7(32'h3a8b20d0),
	.w8(32'h3b02fdd6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1f712),
	.w1(32'h3ae9de7c),
	.w2(32'h3b01433f),
	.w3(32'h3ab38e62),
	.w4(32'h3b20032e),
	.w5(32'hba6530dd),
	.w6(32'h3b3544cf),
	.w7(32'h3b082eb2),
	.w8(32'hba4de208),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9edd36),
	.w1(32'hbaaca013),
	.w2(32'hbad52e03),
	.w3(32'hbb6b5d11),
	.w4(32'hba8bef72),
	.w5(32'h3aa4f480),
	.w6(32'hbb82a1e1),
	.w7(32'hba8acb81),
	.w8(32'h3a98d7b2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b91d9),
	.w1(32'hbb3845a5),
	.w2(32'hbb1c7e56),
	.w3(32'hbb46e9be),
	.w4(32'hbb455845),
	.w5(32'hbb19f4a8),
	.w6(32'hbb760ea3),
	.w7(32'hbb42b7ab),
	.w8(32'hbb79ed47),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab94b61),
	.w1(32'hbac5ba44),
	.w2(32'hba9d0c1b),
	.w3(32'h39912d4d),
	.w4(32'hb8f78505),
	.w5(32'h3a1da66b),
	.w6(32'hba4b20e8),
	.w7(32'hba2de3dc),
	.w8(32'h39f66932),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe35b5),
	.w1(32'hb9c96d53),
	.w2(32'hb990b230),
	.w3(32'h3a6a42ae),
	.w4(32'h39050551),
	.w5(32'hbaa2f52a),
	.w6(32'hba375491),
	.w7(32'hb8a81af4),
	.w8(32'hba261d2d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a6d42),
	.w1(32'hbbe5b4fd),
	.w2(32'hbb329c33),
	.w3(32'hbbdd7f0a),
	.w4(32'hbb49789e),
	.w5(32'h3b71d640),
	.w6(32'hbc31a1b5),
	.w7(32'hbb27bb41),
	.w8(32'h3bf1364c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b537f05),
	.w1(32'h3be39de3),
	.w2(32'h3bca1e21),
	.w3(32'h3aa3f998),
	.w4(32'h3bffb700),
	.w5(32'h3c2fbaab),
	.w6(32'hbbfa263d),
	.w7(32'hba6a4971),
	.w8(32'h3bca3415),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41d6e6),
	.w1(32'h3c2bb867),
	.w2(32'h3be4aca1),
	.w3(32'h3bd98008),
	.w4(32'h3bbdb6e1),
	.w5(32'hbb244dd7),
	.w6(32'h3b8171e1),
	.w7(32'h3b2f3662),
	.w8(32'hbb95423d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12ff96),
	.w1(32'hbabfd89b),
	.w2(32'hba425be8),
	.w3(32'hbadea58e),
	.w4(32'h3a7c831b),
	.w5(32'h3a4ee46f),
	.w6(32'hbb6b9a3b),
	.w7(32'hba4025dc),
	.w8(32'h393882bd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2aae16),
	.w1(32'hbb0f997a),
	.w2(32'hbaea0434),
	.w3(32'hbb1d8ad4),
	.w4(32'hbaf5eb52),
	.w5(32'hbb1fe034),
	.w6(32'hbaddc5ec),
	.w7(32'hba851e47),
	.w8(32'hbad8884f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b933f),
	.w1(32'hb6ed096e),
	.w2(32'hba231a23),
	.w3(32'hba0ae217),
	.w4(32'hba25c2b5),
	.w5(32'h398e17ca),
	.w6(32'hba03b79f),
	.w7(32'hba44514b),
	.w8(32'h36addb19),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39686688),
	.w1(32'h39727074),
	.w2(32'h3a4b692e),
	.w3(32'hb9819aa0),
	.w4(32'h3a9cc36a),
	.w5(32'h3abdb99f),
	.w6(32'hba8b65d0),
	.w7(32'h39c52faf),
	.w8(32'h3a2fc051),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cf423),
	.w1(32'h39257f33),
	.w2(32'hbc39c896),
	.w3(32'hbc1e14f9),
	.w4(32'hb9c7c521),
	.w5(32'hbc5e7985),
	.w6(32'hbc08695e),
	.w7(32'h3af9a176),
	.w8(32'hbc2691b4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc14c9),
	.w1(32'hbaff203e),
	.w2(32'hbb5b1271),
	.w3(32'hbbeab5e4),
	.w4(32'hbb037167),
	.w5(32'hbaeb5217),
	.w6(32'hbc18d98e),
	.w7(32'hbb97514e),
	.w8(32'hbb8b48b3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55d3d2),
	.w1(32'hba543f87),
	.w2(32'hbb85ab34),
	.w3(32'hbb81d9db),
	.w4(32'hbb0cedd6),
	.w5(32'hbba2230e),
	.w6(32'hbc27cadb),
	.w7(32'hbbb55373),
	.w8(32'hbbdc0b68),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc802ed8),
	.w1(32'hbc16ef20),
	.w2(32'hbc38318a),
	.w3(32'hbc8111f7),
	.w4(32'hbc2bd19d),
	.w5(32'hbbf39384),
	.w6(32'hbc75d121),
	.w7(32'hbc229020),
	.w8(32'hbbccf96f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60f2c9),
	.w1(32'hba3323d4),
	.w2(32'hbbcf66b6),
	.w3(32'hbaba55cf),
	.w4(32'hba6cce94),
	.w5(32'hbc161743),
	.w6(32'hbad089cb),
	.w7(32'h3848e7c3),
	.w8(32'hbc187f18),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15dffe),
	.w1(32'h3ab3447a),
	.w2(32'hbaaca7aa),
	.w3(32'h3a807507),
	.w4(32'h3ab78307),
	.w5(32'hbb5955cd),
	.w6(32'h3a288f9b),
	.w7(32'h3af50724),
	.w8(32'hba7b8a11),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2774aa),
	.w1(32'hba49908e),
	.w2(32'hbb1c13b8),
	.w3(32'hba81bcee),
	.w4(32'hbb0e4a3f),
	.w5(32'hbbc11d81),
	.w6(32'hbab58d5b),
	.w7(32'hba69e3e5),
	.w8(32'hbbb985c3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19c505),
	.w1(32'h3ac673b6),
	.w2(32'hbace95ab),
	.w3(32'h3a807b66),
	.w4(32'h3a6eadb5),
	.w5(32'hbae14f50),
	.w6(32'h3a36c47b),
	.w7(32'h3ac700f8),
	.w8(32'hba986752),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8503aa),
	.w1(32'hbad01fbd),
	.w2(32'hbb097479),
	.w3(32'hbb7bb0d7),
	.w4(32'hba8f8c47),
	.w5(32'hbb0e03ab),
	.w6(32'hbb913e98),
	.w7(32'hbb3ca8a0),
	.w8(32'hbb6158d1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc2016),
	.w1(32'hba156628),
	.w2(32'h3817c168),
	.w3(32'hbabc2206),
	.w4(32'hba8ed5e8),
	.w5(32'hbaf99092),
	.w6(32'hbabbf0e6),
	.w7(32'hb819da57),
	.w8(32'hba833fa7),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20fb44),
	.w1(32'hb9ebbd9a),
	.w2(32'hbc017209),
	.w3(32'hba45d925),
	.w4(32'hba8cf57c),
	.w5(32'hbbf37b69),
	.w6(32'hba732781),
	.w7(32'hbac93bd5),
	.w8(32'hbbd08b03),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf4e39),
	.w1(32'hba783854),
	.w2(32'hbb193543),
	.w3(32'h39922647),
	.w4(32'h39fcb521),
	.w5(32'hbb3804c1),
	.w6(32'h395986df),
	.w7(32'h380f1526),
	.w8(32'hbb352556),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacf43b),
	.w1(32'hba5363f5),
	.w2(32'hb885f80b),
	.w3(32'hb8b8ff8b),
	.w4(32'h3a1a459e),
	.w5(32'hb9b6f59a),
	.w6(32'hba74ef25),
	.w7(32'hb9c0d494),
	.w8(32'hb9e69b92),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b37ee),
	.w1(32'hb9c00482),
	.w2(32'hb9bf62fc),
	.w3(32'hb91c94e4),
	.w4(32'hb9e4a3c2),
	.w5(32'hb88b969f),
	.w6(32'hb8526c99),
	.w7(32'hba076a2b),
	.w8(32'h3a014e6f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9ca8a),
	.w1(32'h3abc2038),
	.w2(32'hb89edd0e),
	.w3(32'h3a5e58da),
	.w4(32'hb8886db9),
	.w5(32'hb9df1ab7),
	.w6(32'h3a6446aa),
	.w7(32'hb9fed3bc),
	.w8(32'hb96f1f76),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39822435),
	.w1(32'h3af0a726),
	.w2(32'h3aec7251),
	.w3(32'h38b9683e),
	.w4(32'h3a79f872),
	.w5(32'h39416033),
	.w6(32'h398ecef3),
	.w7(32'h398cdb1b),
	.w8(32'hb8c4d700),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf0c90),
	.w1(32'h3a312d5d),
	.w2(32'h3a8351d1),
	.w3(32'hba83204a),
	.w4(32'h39f7054a),
	.w5(32'h3a2c329a),
	.w6(32'hb9753189),
	.w7(32'h3a8e79e5),
	.w8(32'h3a567316),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc464f),
	.w1(32'h39a494e0),
	.w2(32'hba9ac171),
	.w3(32'hbaf2418a),
	.w4(32'hb809d6a4),
	.w5(32'hbb56d251),
	.w6(32'hba83a563),
	.w7(32'h39f27f44),
	.w8(32'hbb876fa9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb76162),
	.w1(32'h3ad8c5c9),
	.w2(32'hbac8bb63),
	.w3(32'hbb3cbe11),
	.w4(32'h3b0e0690),
	.w5(32'hbb70731e),
	.w6(32'h39dfc802),
	.w7(32'h3b289113),
	.w8(32'hbb8cac92),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e1b82),
	.w1(32'hb9c9bf06),
	.w2(32'h3a088823),
	.w3(32'hba6e0782),
	.w4(32'hb9c90955),
	.w5(32'h38835903),
	.w6(32'hbac19a57),
	.w7(32'hb9b11763),
	.w8(32'hb8a47d7f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cce9a5),
	.w1(32'hb97c5c8b),
	.w2(32'hb9adfd97),
	.w3(32'h39ce59a2),
	.w4(32'hb93b618a),
	.w5(32'hb8e13b72),
	.w6(32'h388cce59),
	.w7(32'hb9ac2a7a),
	.w8(32'hb8cf788f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a4ef9),
	.w1(32'h393d103e),
	.w2(32'hb9843b62),
	.w3(32'h3a02c751),
	.w4(32'hb8e56319),
	.w5(32'hb9cc408b),
	.w6(32'hb5db997d),
	.w7(32'hb9fc09ad),
	.w8(32'hba10dc4d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60faa8),
	.w1(32'hba6ab8d2),
	.w2(32'hba3d7817),
	.w3(32'hb9c77835),
	.w4(32'hb861fe55),
	.w5(32'h3ab0ff36),
	.w6(32'hba192699),
	.w7(32'h3926ec7e),
	.w8(32'h3ab9935e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b07e1),
	.w1(32'hbb3a3a14),
	.w2(32'hbbe27771),
	.w3(32'hbb2abde2),
	.w4(32'hb9ac09c1),
	.w5(32'hbb9350e9),
	.w6(32'hbb0a1486),
	.w7(32'h38a8ab90),
	.w8(32'hbb20c8c2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e5159),
	.w1(32'hbb87fa37),
	.w2(32'hbbc78ecf),
	.w3(32'hba39d322),
	.w4(32'h38c3bf92),
	.w5(32'hbb9a4880),
	.w6(32'hbc36a516),
	.w7(32'hbbe4bdac),
	.w8(32'hbc02b6eb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99f2a7),
	.w1(32'hbaa551ce),
	.w2(32'hbbbb5d80),
	.w3(32'hbb883153),
	.w4(32'h38f04440),
	.w5(32'hbbca6094),
	.w6(32'hbb476860),
	.w7(32'hbaaebb4d),
	.w8(32'hbbe784ec),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e5a7f),
	.w1(32'h39fdec95),
	.w2(32'hbb385b3a),
	.w3(32'hbc0784bf),
	.w4(32'hbabcd88d),
	.w5(32'hba62c219),
	.w6(32'hbc827d33),
	.w7(32'hbc14b745),
	.w8(32'hbbd93c00),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5823a),
	.w1(32'hb9ed6c67),
	.w2(32'hba876a3f),
	.w3(32'hba06ed68),
	.w4(32'hba24924f),
	.w5(32'h391551d8),
	.w6(32'hb9799c8b),
	.w7(32'hb9215b39),
	.w8(32'hb9aea2df),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39419fff),
	.w1(32'hb8d15162),
	.w2(32'hb9282690),
	.w3(32'h39903063),
	.w4(32'h3a0ee7b7),
	.w5(32'h3a80a5e9),
	.w6(32'h39a0407f),
	.w7(32'h39b711cc),
	.w8(32'h3ad0134a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2a205),
	.w1(32'h3a992f6a),
	.w2(32'h3abadcab),
	.w3(32'h3a542241),
	.w4(32'h3a57925b),
	.w5(32'h3acd0935),
	.w6(32'h3a71f6b0),
	.w7(32'h3a58eb8f),
	.w8(32'h3a4ed9a3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05a4a0),
	.w1(32'hb8947c0f),
	.w2(32'hb99fad6c),
	.w3(32'h3a43c82a),
	.w4(32'h3a9fde23),
	.w5(32'h3a034d4e),
	.w6(32'hba22592e),
	.w7(32'hb8b8e3d0),
	.w8(32'hba0603e4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0d0b6),
	.w1(32'h3a815ee2),
	.w2(32'h3a1b71c9),
	.w3(32'h3ab9ec1c),
	.w4(32'h39d5b314),
	.w5(32'h3ada6856),
	.w6(32'h3a4512cc),
	.w7(32'hb805c1a9),
	.w8(32'h3a06dc8b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c25fb7),
	.w1(32'hba2f0a56),
	.w2(32'h399569bb),
	.w3(32'h37f834ea),
	.w4(32'h396d1ccf),
	.w5(32'hbb37e7c2),
	.w6(32'hbb0ca963),
	.w7(32'hb9188284),
	.w8(32'hbb131690),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfa00b),
	.w1(32'hbb68688e),
	.w2(32'hbba4bc85),
	.w3(32'hbb8c11bd),
	.w4(32'hbb29db7d),
	.w5(32'hbb41e069),
	.w6(32'hbbd3cddd),
	.w7(32'hbb0bffce),
	.w8(32'hbb46e55a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac89fb7),
	.w1(32'h39967de2),
	.w2(32'hbae270b5),
	.w3(32'hbb03c78f),
	.w4(32'h39a5cf63),
	.w5(32'h3a86d0b9),
	.w6(32'hbb87af7b),
	.w7(32'hbb44240b),
	.w8(32'hbb24b3f2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2da66d),
	.w1(32'hb9664d11),
	.w2(32'hbb08dcbc),
	.w3(32'hba3aef72),
	.w4(32'h399de80f),
	.w5(32'hba9f20cb),
	.w6(32'hbb087b9c),
	.w7(32'hb9a6871d),
	.w8(32'hbb140949),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb58de),
	.w1(32'hba101622),
	.w2(32'hb9c09963),
	.w3(32'h3a816416),
	.w4(32'hb98342a7),
	.w5(32'hbb2a4588),
	.w6(32'h3897f575),
	.w7(32'h3a937378),
	.w8(32'hba1a4ad8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1ceb6),
	.w1(32'hbb5599d6),
	.w2(32'hbb289930),
	.w3(32'hbb9ea71d),
	.w4(32'hbaa8a710),
	.w5(32'hb96144fd),
	.w6(32'hbbbd20a8),
	.w7(32'hbb368fd8),
	.w8(32'hbb11b5ba),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f7933),
	.w1(32'h399b0437),
	.w2(32'h3a1baaaa),
	.w3(32'hba176471),
	.w4(32'h3911ec2c),
	.w5(32'hba90d9e3),
	.w6(32'hbaa17d1e),
	.w7(32'hb9ff7e39),
	.w8(32'hbaf6d848),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90c92d),
	.w1(32'h3a819f65),
	.w2(32'h39ccfa70),
	.w3(32'h3a2633b9),
	.w4(32'h3a12bbb3),
	.w5(32'h3a2f74ef),
	.w6(32'h39d39afa),
	.w7(32'h39d8e73c),
	.w8(32'hb99f2b1c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fea23),
	.w1(32'hbabfa80f),
	.w2(32'hba9518be),
	.w3(32'hb9810211),
	.w4(32'h393e2d0a),
	.w5(32'h39c2f650),
	.w6(32'hbb1327f6),
	.w7(32'hba87aa86),
	.w8(32'hb99c4049),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a104f07),
	.w1(32'h39c4567e),
	.w2(32'h399ef3b5),
	.w3(32'h383b8ec9),
	.w4(32'h38db9ac2),
	.w5(32'h3a6c88aa),
	.w6(32'hb9c9676d),
	.w7(32'hb84f3c87),
	.w8(32'h3a2177fc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc39ed),
	.w1(32'h3aeed51a),
	.w2(32'h3ae98f77),
	.w3(32'h3a4e88d1),
	.w4(32'h3a15eb67),
	.w5(32'hba4074e8),
	.w6(32'h3a39d992),
	.w7(32'h3a89927d),
	.w8(32'h3992c1d6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e68d5),
	.w1(32'h3a07f8f4),
	.w2(32'hbb36508e),
	.w3(32'hbb4a2de5),
	.w4(32'h3a138542),
	.w5(32'h3a30ffc5),
	.w6(32'hbb9928e3),
	.w7(32'hbb4e24bf),
	.w8(32'hbab4f221),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1e99c),
	.w1(32'h3a22bf8c),
	.w2(32'h3a05d5a2),
	.w3(32'hba0c4dae),
	.w4(32'h398d5c5a),
	.w5(32'h3afd163a),
	.w6(32'hb9e3c921),
	.w7(32'h39760d4a),
	.w8(32'h3ad17214),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ada40),
	.w1(32'h3adfc150),
	.w2(32'h3b242c91),
	.w3(32'h3a1ee780),
	.w4(32'h3b0f04a8),
	.w5(32'h3aae1677),
	.w6(32'hbb1a433c),
	.w7(32'h3a13a81d),
	.w8(32'hb9f1e4ba),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba935e1a),
	.w1(32'h3a15c5e9),
	.w2(32'hbb762c93),
	.w3(32'hba28f53e),
	.w4(32'hb93afc06),
	.w5(32'hbb612d72),
	.w6(32'hbb812e65),
	.w7(32'hba9c3aa7),
	.w8(32'hbb9989a0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4916b7),
	.w1(32'h3b65b40f),
	.w2(32'h3b290510),
	.w3(32'h3ad8ed3d),
	.w4(32'h3b06f6fc),
	.w5(32'h390d4d5e),
	.w6(32'hb99fd83d),
	.w7(32'h3a3e7759),
	.w8(32'hb94d05e4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1a136),
	.w1(32'hbbda9965),
	.w2(32'hbb74ff6b),
	.w3(32'hbbdcbcbf),
	.w4(32'hbbbdbbba),
	.w5(32'hbb25a724),
	.w6(32'hbbb677b5),
	.w7(32'hbbad049b),
	.w8(32'hbb51f61b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7eaaf6),
	.w1(32'h3bd25b78),
	.w2(32'h3bd8561b),
	.w3(32'h3b574da3),
	.w4(32'h3b84846b),
	.w5(32'h3b331588),
	.w6(32'h3a14ddd6),
	.w7(32'h3adc19f0),
	.w8(32'h3a028005),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02a84f),
	.w1(32'hbbbcffd4),
	.w2(32'hbc2054f6),
	.w3(32'hbbac5bdc),
	.w4(32'hbb8bc4c7),
	.w5(32'hbbd7d020),
	.w6(32'hbbe6adce),
	.w7(32'hbbb24e9a),
	.w8(32'hbc00180e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb003eaa),
	.w1(32'hbb282cd6),
	.w2(32'hbb810231),
	.w3(32'hbb52d53a),
	.w4(32'hbaff4844),
	.w5(32'hbb7f7f97),
	.w6(32'hbb325d37),
	.w7(32'hbb11d655),
	.w8(32'hbb4a1936),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cb625),
	.w1(32'hb915c0f1),
	.w2(32'h3910979e),
	.w3(32'hbb96841a),
	.w4(32'hba323b24),
	.w5(32'hb9b1d78c),
	.w6(32'hbbb54b33),
	.w7(32'hbb18216e),
	.w8(32'hb97ca0e1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2f141),
	.w1(32'h3aa7ffe7),
	.w2(32'h39b5a12f),
	.w3(32'h3a8d22de),
	.w4(32'h3ac60b29),
	.w5(32'hba80c627),
	.w6(32'h36c5ae05),
	.w7(32'h3bb82b50),
	.w8(32'h3af1bde5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa83214),
	.w1(32'h3b126820),
	.w2(32'hbbc41a88),
	.w3(32'hba08034c),
	.w4(32'hbad439e3),
	.w5(32'hbc01124d),
	.w6(32'hbb29a4ef),
	.w7(32'h3ad31d9a),
	.w8(32'hbbf676d6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65259e),
	.w1(32'h3b527c8f),
	.w2(32'hba095c6f),
	.w3(32'h3adffb23),
	.w4(32'hbb6bc8b6),
	.w5(32'hbc125cf6),
	.w6(32'hba45dd3a),
	.w7(32'hbb1f6db5),
	.w8(32'hbc04446f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc8b8b),
	.w1(32'hbb985f03),
	.w2(32'hbb243fd8),
	.w3(32'hbbf72880),
	.w4(32'h39886a27),
	.w5(32'h3bc9ffea),
	.w6(32'hbc0a21c5),
	.w7(32'hba84c7c0),
	.w8(32'h3ba9a234),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4ad2f),
	.w1(32'h3ba3f888),
	.w2(32'h3bef76d1),
	.w3(32'hbc5aabeb),
	.w4(32'hbb9fa71d),
	.w5(32'h3be0929b),
	.w6(32'hbc47cfbf),
	.w7(32'hba0249c6),
	.w8(32'h3c8c6251),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a4a94),
	.w1(32'h39636b02),
	.w2(32'hbba596ec),
	.w3(32'h3af12122),
	.w4(32'hbb05c4a8),
	.w5(32'hbbb7e1a2),
	.w6(32'h39b72353),
	.w7(32'h3c07afe4),
	.w8(32'hbc143816),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd80057),
	.w1(32'hbb76636d),
	.w2(32'hbb8b11db),
	.w3(32'hbc3ea115),
	.w4(32'hbaa66d95),
	.w5(32'hbb2c1e11),
	.w6(32'hbbe7832a),
	.w7(32'h3a74332d),
	.w8(32'hbaa79f5f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ec80f),
	.w1(32'h399e7058),
	.w2(32'hbbfbc703),
	.w3(32'hbbb1dc8e),
	.w4(32'hbb62820b),
	.w5(32'hbbb8e743),
	.w6(32'hb99d66ff),
	.w7(32'h3b942865),
	.w8(32'h3b08802a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b9692),
	.w1(32'hbbf1f46a),
	.w2(32'hbb982cbb),
	.w3(32'hbbf26a0b),
	.w4(32'hbabdbd56),
	.w5(32'hbb2df28b),
	.w6(32'hbbbee061),
	.w7(32'h3afe990f),
	.w8(32'h386d9cb2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d8d44),
	.w1(32'h395ad693),
	.w2(32'hbbb0eaf7),
	.w3(32'hbb19b1e5),
	.w4(32'hbb33e08c),
	.w5(32'hbbf55a15),
	.w6(32'hbabc86fe),
	.w7(32'hbb72fbc6),
	.w8(32'hbbc46adb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2e6c9),
	.w1(32'hb8878af0),
	.w2(32'hbb0a3a20),
	.w3(32'h39dc515d),
	.w4(32'hb8f768c9),
	.w5(32'hba9dc456),
	.w6(32'h39f5d4cf),
	.w7(32'h39ab8e5e),
	.w8(32'hba2499ca),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfc1c8),
	.w1(32'h39bd8dbd),
	.w2(32'h38ff58d7),
	.w3(32'hbb7d854b),
	.w4(32'h3a94e7c5),
	.w5(32'hbac21060),
	.w6(32'hbb3ad017),
	.w7(32'hb970ad90),
	.w8(32'hbb2414f0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae941b7),
	.w1(32'h3bd9a257),
	.w2(32'hbb6b8488),
	.w3(32'h3b2dac6d),
	.w4(32'h3a44bb13),
	.w5(32'hbb7276dd),
	.w6(32'h3a86dc54),
	.w7(32'h3b0eb292),
	.w8(32'hbb62e484),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a9dd3),
	.w1(32'h3b46bb2d),
	.w2(32'hbb05bf4b),
	.w3(32'hb9a0b45a),
	.w4(32'h3b20cfee),
	.w5(32'hbb85b10b),
	.w6(32'hba105f2c),
	.w7(32'h3b4db29a),
	.w8(32'hba24e2d3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9dbd8d),
	.w1(32'h3b87e86c),
	.w2(32'h3aa89379),
	.w3(32'hbb2815f3),
	.w4(32'hb8898b19),
	.w5(32'hbacec60a),
	.w6(32'hb97b3db7),
	.w7(32'h3aa8edd7),
	.w8(32'hbb0144ca),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7df04),
	.w1(32'h3b96b341),
	.w2(32'hb9f50d0a),
	.w3(32'h3b331bed),
	.w4(32'h3b2e64c0),
	.w5(32'hba220b51),
	.w6(32'h3b4a3b6f),
	.w7(32'h3a0c3cf9),
	.w8(32'hbb3f4cc8),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9949ffa),
	.w1(32'h3a918658),
	.w2(32'h3b2d2ae9),
	.w3(32'h39bf245b),
	.w4(32'h3b2ec468),
	.w5(32'h3b0655a8),
	.w6(32'hbb7f5966),
	.w7(32'h3a5a8135),
	.w8(32'hbacad685),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18d8ce),
	.w1(32'hbc0a1770),
	.w2(32'hbbe5e559),
	.w3(32'hbc22d742),
	.w4(32'hbbb60888),
	.w5(32'hbbbf9565),
	.w6(32'hbbbcd44f),
	.w7(32'hbbd83076),
	.w8(32'hbc01a84b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69e0b9),
	.w1(32'hba4062ea),
	.w2(32'hbb458105),
	.w3(32'hbb6a78c4),
	.w4(32'hbb56873e),
	.w5(32'hbb26511e),
	.w6(32'hbb9b3bab),
	.w7(32'hbb6dfad4),
	.w8(32'h398bea82),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac42ea4),
	.w1(32'h3b8920e1),
	.w2(32'hbb0515d3),
	.w3(32'h3b8854e3),
	.w4(32'h3acb504c),
	.w5(32'hba790263),
	.w6(32'h3bfa060e),
	.w7(32'h3c1906a5),
	.w8(32'hb9ed0e4d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45139a),
	.w1(32'hbaaf01e1),
	.w2(32'hba4d84b1),
	.w3(32'hbb35f730),
	.w4(32'hbacefbc6),
	.w5(32'hba19ef89),
	.w6(32'hba457172),
	.w7(32'hb9c905f6),
	.w8(32'h3a9faeee),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba914213),
	.w1(32'hba9fcdbf),
	.w2(32'h39e5034f),
	.w3(32'hbab2b40b),
	.w4(32'hba8ec8af),
	.w5(32'h3ac72f18),
	.w6(32'hb9964d9e),
	.w7(32'h3adfdb0a),
	.w8(32'h3b75b6d7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cb350),
	.w1(32'hbaab20c5),
	.w2(32'h3a935acf),
	.w3(32'hba183e5a),
	.w4(32'h3af39daa),
	.w5(32'hba218278),
	.w6(32'h3b8bd0cb),
	.w7(32'h3bce1749),
	.w8(32'h37928cae),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb245438),
	.w1(32'hba772d8a),
	.w2(32'hb9264c4a),
	.w3(32'hbab34532),
	.w4(32'hbab3b043),
	.w5(32'h3ad5f31a),
	.w6(32'hbb6a4695),
	.w7(32'hba35ec81),
	.w8(32'hbb9917fe),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fa53b),
	.w1(32'hb9ebe591),
	.w2(32'h3a0b7745),
	.w3(32'hbab93517),
	.w4(32'hbabd71fa),
	.w5(32'hbb122404),
	.w6(32'hbb611103),
	.w7(32'hb975379d),
	.w8(32'hbb102610),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87bf90),
	.w1(32'h38891dfd),
	.w2(32'hbb12d1c3),
	.w3(32'hbb128be3),
	.w4(32'hbb1ba738),
	.w5(32'hba02ea12),
	.w6(32'hbb1b1611),
	.w7(32'hba3952d7),
	.w8(32'hbb9372a7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc31678),
	.w1(32'hbb20417f),
	.w2(32'hbb524352),
	.w3(32'hbb9fad79),
	.w4(32'hba8df915),
	.w5(32'hbab9128e),
	.w6(32'hbc22cb4e),
	.w7(32'hbba2a5cf),
	.w8(32'hbbb53298),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41eaee),
	.w1(32'h3adb47ca),
	.w2(32'hb8231f01),
	.w3(32'h3ac2d854),
	.w4(32'h3a880694),
	.w5(32'hbae344f4),
	.w6(32'hbb048fd3),
	.w7(32'hbb190778),
	.w8(32'h39f96935),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d1692),
	.w1(32'hbad69f25),
	.w2(32'hba78b3a0),
	.w3(32'hbb9a58ba),
	.w4(32'hbb1d1d7f),
	.w5(32'hbab1a82f),
	.w6(32'hba82244a),
	.w7(32'h391ef52e),
	.w8(32'hba8dedd4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71ddc9),
	.w1(32'hbadf0e32),
	.w2(32'hb9a66d85),
	.w3(32'hbb093c7d),
	.w4(32'hbb8e3400),
	.w5(32'h39499ee5),
	.w6(32'hb9a7a59e),
	.w7(32'hbaaa9b1a),
	.w8(32'h3a8a8f86),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bebd51),
	.w1(32'hba2f5f56),
	.w2(32'hba727372),
	.w3(32'h399cdc8e),
	.w4(32'h3a4d61e6),
	.w5(32'h39790fc7),
	.w6(32'h3ae4e353),
	.w7(32'h3b0d592b),
	.w8(32'hbb127399),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb371643),
	.w1(32'hbbd35102),
	.w2(32'hbba72f8f),
	.w3(32'h37bff3e0),
	.w4(32'hbb9865b1),
	.w5(32'hbb821f1e),
	.w6(32'hbb876fe1),
	.w7(32'hbb974184),
	.w8(32'hbb9a2f36),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4de8f),
	.w1(32'hbb3c671e),
	.w2(32'hbb08e372),
	.w3(32'hba21d1c3),
	.w4(32'h3ae756bf),
	.w5(32'hbb56a1c8),
	.w6(32'hbb48112e),
	.w7(32'hba240278),
	.w8(32'hbb3ac62f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba643b92),
	.w1(32'hb928b9d7),
	.w2(32'hb9a98bfa),
	.w3(32'h3a049c07),
	.w4(32'h38ae2923),
	.w5(32'hbb90b1e5),
	.w6(32'hb7ece8d0),
	.w7(32'h38a688ef),
	.w8(32'h3bc4d7c6),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa30145),
	.w1(32'h3c1a1a66),
	.w2(32'h3b7b1055),
	.w3(32'hb80b86d8),
	.w4(32'hbaa2244d),
	.w5(32'hba81fc31),
	.w6(32'h3bb9a90a),
	.w7(32'h3c5a37e0),
	.w8(32'h3924e0dc),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06723e),
	.w1(32'h3ae54a4d),
	.w2(32'h36b6881f),
	.w3(32'h39e2e1a4),
	.w4(32'h3ab2850e),
	.w5(32'h3b5b4767),
	.w6(32'h39efd2d9),
	.w7(32'h3a24a67c),
	.w8(32'h3bb15a01),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c1163),
	.w1(32'h3a3c5062),
	.w2(32'hbb068520),
	.w3(32'h3af3d7e5),
	.w4(32'hba1788c5),
	.w5(32'hbaa8e6c8),
	.w6(32'h3b9ee4e9),
	.w7(32'h3ba28fba),
	.w8(32'hbb211c03),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb42f92),
	.w1(32'hbb52223a),
	.w2(32'hbb8cc88b),
	.w3(32'hbb7a159e),
	.w4(32'hb995cffe),
	.w5(32'hbb81a67a),
	.w6(32'hbb071adf),
	.w7(32'hb9e63b74),
	.w8(32'hbb5e632b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccbe9b),
	.w1(32'hba9476a5),
	.w2(32'hbb8e6250),
	.w3(32'hbb80dd49),
	.w4(32'hbb2bf85e),
	.w5(32'hbb936b3a),
	.w6(32'hbb0b0b2b),
	.w7(32'hb9d46354),
	.w8(32'hbb63db75),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdabcb),
	.w1(32'hbabf39ff),
	.w2(32'hb921dedc),
	.w3(32'hbb484bb1),
	.w4(32'hba381414),
	.w5(32'h39f15b29),
	.w6(32'hbba0d1bc),
	.w7(32'hba7f275a),
	.w8(32'hb8b45e00),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a81189),
	.w1(32'hb907fea1),
	.w2(32'hba98af31),
	.w3(32'hbae13bc6),
	.w4(32'h38b142a3),
	.w5(32'h39af0bce),
	.w6(32'hba86b2fd),
	.w7(32'h3aecaa60),
	.w8(32'hbb3a2d85),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3cf97),
	.w1(32'hba60b2e0),
	.w2(32'hba914148),
	.w3(32'hba38f0a2),
	.w4(32'h3a50abfe),
	.w5(32'hbb3b13ee),
	.w6(32'hbacc530b),
	.w7(32'h3a719b56),
	.w8(32'hbb6dd273),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb080298),
	.w1(32'h3ae61f8e),
	.w2(32'h3ac89905),
	.w3(32'hbacc459e),
	.w4(32'h3b1e1e8e),
	.w5(32'h3a6e3aea),
	.w6(32'hbb8d5809),
	.w7(32'h39ef8922),
	.w8(32'hba4b0700),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6c973),
	.w1(32'hbb5460b7),
	.w2(32'hbb7fc4d3),
	.w3(32'hbb2aaea7),
	.w4(32'hba433efd),
	.w5(32'hbb21c778),
	.w6(32'hbb7bf917),
	.w7(32'hbb493252),
	.w8(32'hbbb239e7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3a9d7),
	.w1(32'h3acd8808),
	.w2(32'hb9e7616d),
	.w3(32'h3a215cfb),
	.w4(32'hb88512dc),
	.w5(32'hbbc082d2),
	.w6(32'hbb68acd3),
	.w7(32'hbb074874),
	.w8(32'hbbb12e3c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb182e10),
	.w1(32'hb9950ace),
	.w2(32'h3b172ac2),
	.w3(32'hbbe824e5),
	.w4(32'hbb0b7d78),
	.w5(32'hbb5b0fa0),
	.w6(32'hbbfcf6a9),
	.w7(32'hbbee96ba),
	.w8(32'hbb88ea5e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d849a4),
	.w1(32'h3af2a774),
	.w2(32'h3a4ac960),
	.w3(32'hba7f232e),
	.w4(32'h3a27e543),
	.w5(32'h3a576b68),
	.w6(32'h3aa00ee1),
	.w7(32'h3b0bf9db),
	.w8(32'hba78bd7d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbc1fd),
	.w1(32'hbb152d3c),
	.w2(32'hb9a3958f),
	.w3(32'hba2fa942),
	.w4(32'hbadd3663),
	.w5(32'hba0061de),
	.w6(32'hbb205fbc),
	.w7(32'hbb18e34e),
	.w8(32'h3ac7fff7),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcef47),
	.w1(32'h3b1d35c5),
	.w2(32'h3ac7655c),
	.w3(32'hb9372788),
	.w4(32'hba40559d),
	.w5(32'hbb0218a9),
	.w6(32'h3b0a9340),
	.w7(32'h3ac29931),
	.w8(32'h3a3906ec),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38051cd6),
	.w1(32'h3a10655d),
	.w2(32'h399139f3),
	.w3(32'hba8ae45a),
	.w4(32'hba341e80),
	.w5(32'hba6f4884),
	.w6(32'h39a8e940),
	.w7(32'h3aa28aa1),
	.w8(32'h3b55f842),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f1b62),
	.w1(32'hb768b240),
	.w2(32'hba91588f),
	.w3(32'hbb2ab583),
	.w4(32'hbaa45080),
	.w5(32'hbaf493f2),
	.w6(32'hba812ba8),
	.w7(32'hb9b0a899),
	.w8(32'hbb691531),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7c00d),
	.w1(32'hba9430fe),
	.w2(32'hbb802658),
	.w3(32'hbac04596),
	.w4(32'hbab39efa),
	.w5(32'hbb2555ac),
	.w6(32'hbb724cc6),
	.w7(32'hbbd5741b),
	.w8(32'hbb8f9ed3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3948f6cc),
	.w1(32'h398e27b4),
	.w2(32'h3a7e496e),
	.w3(32'hbb1d2fe2),
	.w4(32'hbb007d06),
	.w5(32'h3979d889),
	.w6(32'hbaab5d16),
	.w7(32'hb92eb3a1),
	.w8(32'h3a5d44a6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac153de),
	.w1(32'hb906d5c1),
	.w2(32'hbb1b9a08),
	.w3(32'hbba0704d),
	.w4(32'hbad5451a),
	.w5(32'hbb9cfeee),
	.w6(32'hbb69cc29),
	.w7(32'hbaac53de),
	.w8(32'hbc02683a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82e7cc),
	.w1(32'hbbc4dd99),
	.w2(32'hbbbe6842),
	.w3(32'hbb078c88),
	.w4(32'h39f5efaf),
	.w5(32'hbb4c2df1),
	.w6(32'hbb390349),
	.w7(32'hbb2d5063),
	.w8(32'hbb498312),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5c9fc),
	.w1(32'hbbb3aafe),
	.w2(32'hba98d647),
	.w3(32'hbc0dba2a),
	.w4(32'hbbb132cf),
	.w5(32'hbc1682b1),
	.w6(32'hbc096dac),
	.w7(32'hbb61c2c7),
	.w8(32'h3bef57d2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f30da),
	.w1(32'h3a3a8acf),
	.w2(32'hba9ca27b),
	.w3(32'hbbe96d5c),
	.w4(32'hbba9b54a),
	.w5(32'hba8afa92),
	.w6(32'h3aa19855),
	.w7(32'h3c4ab7c4),
	.w8(32'hbb4d6380),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1625f1),
	.w1(32'h3b0bf2b5),
	.w2(32'hbad71861),
	.w3(32'h3b0ab175),
	.w4(32'h3a8aee47),
	.w5(32'hbb1a3e50),
	.w6(32'h3b4f675a),
	.w7(32'h3af7688a),
	.w8(32'h3b1d7419),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c161116),
	.w1(32'h3be77662),
	.w2(32'h3b603446),
	.w3(32'h3be7c579),
	.w4(32'h3b25f811),
	.w5(32'h3a7a60e0),
	.w6(32'h3bfd08d3),
	.w7(32'h3bfb5505),
	.w8(32'h3b8c1316),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38b359),
	.w1(32'hbbc0531e),
	.w2(32'hbb77a920),
	.w3(32'hbc2687ee),
	.w4(32'hbb6434a4),
	.w5(32'hbb753bfa),
	.w6(32'hbc0c7bb4),
	.w7(32'hbba158e8),
	.w8(32'hba975ccc),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb938f80a),
	.w1(32'h3b03fe0d),
	.w2(32'h3b2bd9c1),
	.w3(32'h3ab9bc56),
	.w4(32'h3af64604),
	.w5(32'h3aa2e9a1),
	.w6(32'h3aff9b98),
	.w7(32'h3b60c436),
	.w8(32'hbaa293fa),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d1cbd),
	.w1(32'h3bb014f0),
	.w2(32'h3a77484a),
	.w3(32'h3b055d1f),
	.w4(32'h3add4da4),
	.w5(32'h3b2a54f4),
	.w6(32'hba93ec42),
	.w7(32'h39abd67e),
	.w8(32'h38597b11),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71f27c),
	.w1(32'hb88bbb8f),
	.w2(32'h3a965b8a),
	.w3(32'hba37b81e),
	.w4(32'hbb055102),
	.w5(32'hbb83d60a),
	.w6(32'hbab284cc),
	.w7(32'hbb8027f6),
	.w8(32'hba9d3d6d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1622c),
	.w1(32'hbb3839d5),
	.w2(32'hbb1e4512),
	.w3(32'hbbcffddc),
	.w4(32'hbb115e79),
	.w5(32'hb9b2ea0f),
	.w6(32'hbb443f66),
	.w7(32'h3ad42c6a),
	.w8(32'h39873478),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90be46),
	.w1(32'hbba3cb07),
	.w2(32'hbb8219f3),
	.w3(32'h3aaca09b),
	.w4(32'hbb79e3fc),
	.w5(32'hbb298336),
	.w6(32'hbb76eaec),
	.w7(32'hbb8c7070),
	.w8(32'hbab63b66),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3d60c),
	.w1(32'hbacdb85f),
	.w2(32'hbab90846),
	.w3(32'hb9d1df01),
	.w4(32'hb986bed7),
	.w5(32'hba28fded),
	.w6(32'h39ab1fa7),
	.w7(32'h3a2d582b),
	.w8(32'h3b9a1a61),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb889601),
	.w1(32'h3993c4c0),
	.w2(32'hbb3b4f8e),
	.w3(32'hbb92c193),
	.w4(32'hbb607f7b),
	.w5(32'hbb4702b5),
	.w6(32'hba8a1586),
	.w7(32'h3a45279f),
	.w8(32'hba48df85),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a685d),
	.w1(32'h3b343177),
	.w2(32'h3ac5fd05),
	.w3(32'hb91ce44c),
	.w4(32'h3a96381a),
	.w5(32'h38a32bee),
	.w6(32'h3b5996df),
	.w7(32'h3a84cb8f),
	.w8(32'h3a9bb939),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39363f71),
	.w1(32'hbaf39b8d),
	.w2(32'hbafeb7a3),
	.w3(32'h3aa5404a),
	.w4(32'hbaee04f2),
	.w5(32'hbac4b8b3),
	.w6(32'hbb15f655),
	.w7(32'hbb1a4b27),
	.w8(32'hba8d1c36),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67951b),
	.w1(32'h3a4260d8),
	.w2(32'h3b7564dd),
	.w3(32'hba932ffd),
	.w4(32'hb9002700),
	.w5(32'h3a14a7c4),
	.w6(32'h391acb1b),
	.w7(32'h3b1d2cc6),
	.w8(32'hbabce776),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae164d8),
	.w1(32'h3ae52696),
	.w2(32'h3ae3cb00),
	.w3(32'h3b35bcea),
	.w4(32'h3b2248f9),
	.w5(32'h3abfaa1e),
	.w6(32'h3a358e6c),
	.w7(32'hbb19f07a),
	.w8(32'h3a2abf8d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c9bb3),
	.w1(32'h39d7492f),
	.w2(32'h391b8782),
	.w3(32'hbb3af9f2),
	.w4(32'h3a3335c6),
	.w5(32'hb9f80dea),
	.w6(32'hbb3b07ac),
	.w7(32'h39864801),
	.w8(32'h3aab6836),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9b16e),
	.w1(32'hbab39cb6),
	.w2(32'hbb9dcfab),
	.w3(32'hbc0cf659),
	.w4(32'hba86186f),
	.w5(32'hbb753cea),
	.w6(32'hbc2d8959),
	.w7(32'hbba2ec52),
	.w8(32'hbb5edc6a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49045d),
	.w1(32'h3b6bd882),
	.w2(32'h3afe7926),
	.w3(32'h3b854950),
	.w4(32'h3baf36dd),
	.w5(32'hbac13544),
	.w6(32'h3bdcf838),
	.w7(32'h3bcd7596),
	.w8(32'h3b1b3b84),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c56b2),
	.w1(32'h3ae74150),
	.w2(32'h399f2c0f),
	.w3(32'hbb8c4a35),
	.w4(32'hba0850e4),
	.w5(32'h3980ddd6),
	.w6(32'hbb7925cb),
	.w7(32'hbb2e21ea),
	.w8(32'h3b1e8be5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2e95f),
	.w1(32'h3ab9e674),
	.w2(32'hb88faf1b),
	.w3(32'hba4e65cf),
	.w4(32'hbabd77d9),
	.w5(32'hbac8f04b),
	.w6(32'h3b970eaa),
	.w7(32'h3af22658),
	.w8(32'h3a7afaf9),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6cfd4),
	.w1(32'hba89e420),
	.w2(32'hbc042ceb),
	.w3(32'hbb86a06e),
	.w4(32'h39f80384),
	.w5(32'hbb86e9c5),
	.w6(32'hbb03bcb2),
	.w7(32'hb8b22542),
	.w8(32'hbbe565a9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9960ccb),
	.w1(32'hbafe406a),
	.w2(32'hbb839499),
	.w3(32'hbb78d6d7),
	.w4(32'hbac8c081),
	.w5(32'hbb0c6a2d),
	.w6(32'hbb876163),
	.w7(32'hbae647ca),
	.w8(32'hbae82acf),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb726eb4),
	.w1(32'h39ab9818),
	.w2(32'hbbb14a66),
	.w3(32'hbb8e69c3),
	.w4(32'hbb6c6ff4),
	.w5(32'hbbf0edc4),
	.w6(32'hbbe253b3),
	.w7(32'hbb2ea955),
	.w8(32'hbbd00ec4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4044a4),
	.w1(32'h3b60de8e),
	.w2(32'h3b43375e),
	.w3(32'h39ad1526),
	.w4(32'h3b2d6538),
	.w5(32'h3b29c7b3),
	.w6(32'h3b35aae3),
	.w7(32'h3b9f56e7),
	.w8(32'h3b97ba62),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd4459),
	.w1(32'hbb28dbfb),
	.w2(32'hbb2eb949),
	.w3(32'hbb7fbf19),
	.w4(32'hba77a9ce),
	.w5(32'hbb1f9d33),
	.w6(32'hbb4cd057),
	.w7(32'hb99b96a2),
	.w8(32'hbab531e5),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb854441d),
	.w1(32'hb9129d3d),
	.w2(32'h39ff66a9),
	.w3(32'hbb0beb60),
	.w4(32'hbb1ea517),
	.w5(32'h3a4c3461),
	.w6(32'hba2888e6),
	.w7(32'h398287e8),
	.w8(32'h3ac1cf9c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39971235),
	.w1(32'h3b04f506),
	.w2(32'h398f069e),
	.w3(32'hba9db5e7),
	.w4(32'hb8864893),
	.w5(32'hbb17d00e),
	.w6(32'h3b41b297),
	.w7(32'h3b5f3b43),
	.w8(32'hb9971f14),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa03d50),
	.w1(32'hb9ac1dc0),
	.w2(32'h3a502e07),
	.w3(32'hbb1fa31d),
	.w4(32'hbafc3ede),
	.w5(32'h3b326c73),
	.w6(32'h39c93383),
	.w7(32'hbab172ab),
	.w8(32'hbb2886f6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc35ba5),
	.w1(32'hbbf3010c),
	.w2(32'hbbc803e9),
	.w3(32'hbbc9792f),
	.w4(32'hbadc6508),
	.w5(32'hbbcb421e),
	.w6(32'hbbf6daef),
	.w7(32'hbb87e951),
	.w8(32'hbb92c387),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2a89b),
	.w1(32'hbac7f4f1),
	.w2(32'hbb0a1c39),
	.w3(32'hbaf9b4a9),
	.w4(32'h3835df80),
	.w5(32'hbb245e66),
	.w6(32'hb92e48cc),
	.w7(32'hb9264b81),
	.w8(32'hbbb186b5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc5097),
	.w1(32'hbb5fbff0),
	.w2(32'hbb520d48),
	.w3(32'hba936814),
	.w4(32'hba3018a0),
	.w5(32'h3ab68bac),
	.w6(32'hbb4bb8ee),
	.w7(32'hbba05199),
	.w8(32'h3c42b1ab),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eb3ca),
	.w1(32'h3be55c81),
	.w2(32'h3b7f21bd),
	.w3(32'hb9dcfe85),
	.w4(32'hba5547f6),
	.w5(32'h3af86665),
	.w6(32'h3be81d1e),
	.w7(32'h3bc9afd6),
	.w8(32'h3b745c09),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b005fdb),
	.w1(32'hb89078cb),
	.w2(32'hbb3fb26a),
	.w3(32'hbb17c6d9),
	.w4(32'hba0eb92d),
	.w5(32'hbba0b9ee),
	.w6(32'h3a5f0b87),
	.w7(32'hbad0c115),
	.w8(32'hbb99992d),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd44497),
	.w1(32'h3a8e44d7),
	.w2(32'h3a324e25),
	.w3(32'hbb399121),
	.w4(32'h3abd1ac4),
	.w5(32'hba44099c),
	.w6(32'h3aa59d92),
	.w7(32'h3b7593d3),
	.w8(32'h3b070be7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b82e3),
	.w1(32'hb93b335f),
	.w2(32'h3a030a9e),
	.w3(32'hbb3f6a5c),
	.w4(32'hbb12bc9c),
	.w5(32'h3af64848),
	.w6(32'hb9e25362),
	.w7(32'hb975df5c),
	.w8(32'h3bd5dc7a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fb8a9),
	.w1(32'hbab8331b),
	.w2(32'hbba19045),
	.w3(32'hbb3e44a7),
	.w4(32'hbb70c4b6),
	.w5(32'hbc2ef392),
	.w6(32'h38a4ed97),
	.w7(32'h3b935071),
	.w8(32'hbc6215e6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0016ea),
	.w1(32'h392de77a),
	.w2(32'hbbd7a389),
	.w3(32'hbbcc472f),
	.w4(32'h3b4bf25a),
	.w5(32'hbb440984),
	.w6(32'hbbd2e730),
	.w7(32'hba412b9b),
	.w8(32'hbbf551b1),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39265ff7),
	.w1(32'hbaa396db),
	.w2(32'hbb365e3a),
	.w3(32'h39ba3127),
	.w4(32'hba49629d),
	.w5(32'hbb9c6fd0),
	.w6(32'hba023c62),
	.w7(32'hba37890a),
	.w8(32'h3bb186d8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5cd24),
	.w1(32'h3a22aee2),
	.w2(32'hbb0fb68d),
	.w3(32'hbb1fbdf5),
	.w4(32'hbad59f73),
	.w5(32'h3a8b660d),
	.w6(32'h3b94d9a1),
	.w7(32'h3b5e09b0),
	.w8(32'h3ab1eca0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff855b),
	.w1(32'hb9d6cf94),
	.w2(32'hbb4c7822),
	.w3(32'hb9ff1782),
	.w4(32'h397dd864),
	.w5(32'hbb09ccab),
	.w6(32'h39d8ab10),
	.w7(32'hbb1191c1),
	.w8(32'hbac99d38),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bb1e0),
	.w1(32'h38f65c90),
	.w2(32'hbb512e00),
	.w3(32'hb9e20c94),
	.w4(32'h3a64ca0c),
	.w5(32'h3a8e52ab),
	.w6(32'hba53b8bc),
	.w7(32'hba95b50a),
	.w8(32'hbc3e97f9),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb909e292),
	.w1(32'hbbfb73fe),
	.w2(32'hbbe1e665),
	.w3(32'h3aff8283),
	.w4(32'hba38d0fd),
	.w5(32'hbb4bc6af),
	.w6(32'hbbf37415),
	.w7(32'hbc33ef14),
	.w8(32'hbb1fcb2b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd1fc7),
	.w1(32'h39dd2f03),
	.w2(32'hbaaeb6bc),
	.w3(32'h3ac42844),
	.w4(32'h3adb401c),
	.w5(32'h3b122085),
	.w6(32'h38a3e915),
	.w7(32'h3b51a328),
	.w8(32'hb99791e2),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6016b2),
	.w1(32'hbae3badc),
	.w2(32'hbb35b766),
	.w3(32'hba772ea8),
	.w4(32'h3a8c11f9),
	.w5(32'hbadf78fa),
	.w6(32'hbb3b6292),
	.w7(32'hbad4d8ec),
	.w8(32'hbb9ba530),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38647f),
	.w1(32'h38d31129),
	.w2(32'hba5dfd48),
	.w3(32'h3b95ebc4),
	.w4(32'h397c6001),
	.w5(32'h3b003aa5),
	.w6(32'h3a7e19d6),
	.w7(32'hbaa1da71),
	.w8(32'h3b0b635e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38451e19),
	.w1(32'h39f7db6d),
	.w2(32'hbbbbb1ce),
	.w3(32'h3a75e07b),
	.w4(32'h384b2d91),
	.w5(32'hbba8237b),
	.w6(32'hb80ccbeb),
	.w7(32'hbad63a4a),
	.w8(32'hbb70e2d0),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba348ed4),
	.w1(32'hba44c2ba),
	.w2(32'hba9c8956),
	.w3(32'hbad1a9bd),
	.w4(32'hbb0a82f1),
	.w5(32'hba488c6f),
	.w6(32'hb9503409),
	.w7(32'hba971f51),
	.w8(32'hba7201ac),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89dfc7),
	.w1(32'h3a304c28),
	.w2(32'h3acc0129),
	.w3(32'hbaa4574a),
	.w4(32'hbae2c3b8),
	.w5(32'h3ae05dea),
	.w6(32'hba5e53b1),
	.w7(32'hba7da3da),
	.w8(32'hba9be2cf),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93ce8c),
	.w1(32'hbb9f00a5),
	.w2(32'hbb65f79f),
	.w3(32'h39b34e0a),
	.w4(32'hbae797a7),
	.w5(32'hbb50eeb4),
	.w6(32'hbb64d24e),
	.w7(32'hbb34f396),
	.w8(32'hbb04df72),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbe591),
	.w1(32'hba3c8126),
	.w2(32'hbafe44a8),
	.w3(32'hbb22125e),
	.w4(32'hbabd0a4e),
	.w5(32'hbab084b8),
	.w6(32'hbaa463e5),
	.w7(32'hbb094e34),
	.w8(32'hbb1cb085),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb250036),
	.w1(32'hba3e0c45),
	.w2(32'hbac936da),
	.w3(32'hba9fa8de),
	.w4(32'h3914fd70),
	.w5(32'hbb337f4f),
	.w6(32'hbb7fe005),
	.w7(32'hba4d9798),
	.w8(32'hbb342517),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1c2b9),
	.w1(32'h3b04ab4b),
	.w2(32'hb92b974a),
	.w3(32'hbb764c41),
	.w4(32'hb99e7915),
	.w5(32'h3941b188),
	.w6(32'hbb8970e0),
	.w7(32'hbacb5a83),
	.w8(32'hbc2016dd),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a184cbb),
	.w1(32'hba9644c8),
	.w2(32'hbacc7b3a),
	.w3(32'hbb91cafa),
	.w4(32'h39478bb1),
	.w5(32'hbab31252),
	.w6(32'hbc04867e),
	.w7(32'hbbc6103f),
	.w8(32'hbba0fda0),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68da14),
	.w1(32'hbac823a6),
	.w2(32'hba56f0c7),
	.w3(32'hba04bf30),
	.w4(32'hba1a670d),
	.w5(32'hb8815aa9),
	.w6(32'h3a09f407),
	.w7(32'hbafe9289),
	.w8(32'hbb1a639c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a5803),
	.w1(32'h3a1905d3),
	.w2(32'hbb8e050c),
	.w3(32'hbbac6ff3),
	.w4(32'hba790c7c),
	.w5(32'hb97b3db6),
	.w6(32'hbbdd572a),
	.w7(32'hbb731bb6),
	.w8(32'hbb322984),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99e5f3),
	.w1(32'hbb16a496),
	.w2(32'hbb986da8),
	.w3(32'hbb214a36),
	.w4(32'hba397e4d),
	.w5(32'hbbd29c63),
	.w6(32'hbaaad8c1),
	.w7(32'h3852d867),
	.w8(32'hbb0bd8fb),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bba67),
	.w1(32'hbb201a4d),
	.w2(32'hbb7ee759),
	.w3(32'hbc0734ea),
	.w4(32'hbb8b69a5),
	.w5(32'hbac8a3f4),
	.w6(32'hbc09bb9a),
	.w7(32'hbbdf5282),
	.w8(32'hbb9cbe0f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a827c),
	.w1(32'hbaa24d00),
	.w2(32'hbb210834),
	.w3(32'hba072de2),
	.w4(32'hba24b570),
	.w5(32'hbae3ab1d),
	.w6(32'h3a032aeb),
	.w7(32'hba3a7836),
	.w8(32'hbab91c91),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cd387),
	.w1(32'h3b0c817c),
	.w2(32'h3a90b17f),
	.w3(32'h3ac27963),
	.w4(32'h395a0735),
	.w5(32'h382e0ac2),
	.w6(32'h3abdac6b),
	.w7(32'hbaae5200),
	.w8(32'hbb33e671),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee267b),
	.w1(32'h3b593069),
	.w2(32'h3b1bbf77),
	.w3(32'h3a8e3f00),
	.w4(32'h3ae1d0a7),
	.w5(32'hbb4611d6),
	.w6(32'hbbead165),
	.w7(32'hbaab9850),
	.w8(32'hbbbad1e8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea3085),
	.w1(32'hbb2c31c4),
	.w2(32'hbb7781d5),
	.w3(32'hbbceaa86),
	.w4(32'hbaf9188a),
	.w5(32'hbb359f37),
	.w6(32'hbc0deab6),
	.w7(32'hbb8b2f70),
	.w8(32'hbb919cd6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a4a5a),
	.w1(32'hbb6988ea),
	.w2(32'hbb6694f6),
	.w3(32'hbb8aa74d),
	.w4(32'hbab99e43),
	.w5(32'hbc032f5f),
	.w6(32'hbc07d66b),
	.w7(32'hbb84084b),
	.w8(32'hbbc98547),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91bc01),
	.w1(32'h3aecd93c),
	.w2(32'hbadfbf0b),
	.w3(32'hbada0fdf),
	.w4(32'hbb81ff8d),
	.w5(32'hbbbe2228),
	.w6(32'h3b67f0d5),
	.w7(32'h3b000098),
	.w8(32'hbbd5d854),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cf806),
	.w1(32'hbb5a4840),
	.w2(32'hbaa4ac33),
	.w3(32'hbb3ffd5a),
	.w4(32'hbb14556e),
	.w5(32'hbad0ec37),
	.w6(32'hbb4ced9c),
	.w7(32'hbbe07a65),
	.w8(32'h3a93e934),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c54d7),
	.w1(32'hbaed7bd6),
	.w2(32'hbacca4ba),
	.w3(32'hbb0e490c),
	.w4(32'hbb002c2d),
	.w5(32'hba8c82e9),
	.w6(32'h3a778a62),
	.w7(32'h3a1b51a4),
	.w8(32'hbb206eab),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44291b),
	.w1(32'h3b1be71c),
	.w2(32'hbb80da83),
	.w3(32'hbb2035d4),
	.w4(32'hb8cd0352),
	.w5(32'hba988418),
	.w6(32'hbba457ee),
	.w7(32'hbb109ae5),
	.w8(32'hba8548ea),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb885380),
	.w1(32'hba69dda0),
	.w2(32'hbb1ce8df),
	.w3(32'hbb18d006),
	.w4(32'h3962b67d),
	.w5(32'hbb409416),
	.w6(32'hbbb41f44),
	.w7(32'hbb0d0e26),
	.w8(32'hbbedd3c1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3678d1),
	.w1(32'h3a5407d2),
	.w2(32'hbaf00bc8),
	.w3(32'h3aaef0b9),
	.w4(32'h38e955da),
	.w5(32'hbac85021),
	.w6(32'hbaa317da),
	.w7(32'h39e7b5a8),
	.w8(32'h3ba0d403),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3da9c5),
	.w1(32'h3b9a95e6),
	.w2(32'h3a1a313b),
	.w3(32'hbb878f22),
	.w4(32'hbab74af5),
	.w5(32'hbaa460f5),
	.w6(32'hbb4a24d3),
	.w7(32'h3a146913),
	.w8(32'h3c1651e7),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c7d14),
	.w1(32'h3a9e955e),
	.w2(32'h3ad788ac),
	.w3(32'hbb8266b7),
	.w4(32'h3a47bf72),
	.w5(32'hbabc7d80),
	.w6(32'h3c03d39f),
	.w7(32'h3c5f905e),
	.w8(32'hbbb5b52c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1ddd6),
	.w1(32'hbb413eee),
	.w2(32'hba43fddf),
	.w3(32'hb97aa248),
	.w4(32'hb9a0fe82),
	.w5(32'hbb520e95),
	.w6(32'hbb048b62),
	.w7(32'hba97312c),
	.w8(32'h3a9466f5),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f61c74),
	.w1(32'hbace8c5a),
	.w2(32'hb9105b1f),
	.w3(32'hbb4bf91c),
	.w4(32'hbb60b00a),
	.w5(32'hba69c50b),
	.w6(32'hba8c674a),
	.w7(32'hbabc49fa),
	.w8(32'hbae1d535),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0e859),
	.w1(32'hb9b698a5),
	.w2(32'hbabe3114),
	.w3(32'hba80671d),
	.w4(32'hbb01ec63),
	.w5(32'hbb243ffe),
	.w6(32'hb8d485b4),
	.w7(32'hbaa8a119),
	.w8(32'hbb1041d9),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae093f),
	.w1(32'h3b31ce96),
	.w2(32'h3b5ea73d),
	.w3(32'hbbdeb968),
	.w4(32'hba1f5aac),
	.w5(32'h3a2f1ffa),
	.w6(32'hb9eeb58a),
	.w7(32'h3b0a7fb3),
	.w8(32'h3aadf1e2),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9d570),
	.w1(32'hba03c106),
	.w2(32'hbb221bac),
	.w3(32'h3ac82a53),
	.w4(32'hbab139eb),
	.w5(32'hbb3d26df),
	.w6(32'h3aa5ec66),
	.w7(32'hb97adbd3),
	.w8(32'hbaf306c2),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b7269),
	.w1(32'hbbb6ed3b),
	.w2(32'hbb8868e3),
	.w3(32'hbb9cbf19),
	.w4(32'hbb811a9e),
	.w5(32'hbb27a996),
	.w6(32'hbbfca9d8),
	.w7(32'hbbeb6193),
	.w8(32'hbb974413),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99a565),
	.w1(32'h3b2e8da7),
	.w2(32'h3ac37867),
	.w3(32'hbaabb7b1),
	.w4(32'h3a3ec26a),
	.w5(32'hbb1c6855),
	.w6(32'hbb18e1ba),
	.w7(32'hb9b1e5ce),
	.w8(32'hbb13b8d2),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0495b8),
	.w1(32'hb88097e3),
	.w2(32'hba550fcf),
	.w3(32'hb9f085b4),
	.w4(32'h3a19a823),
	.w5(32'hbaba7e1d),
	.w6(32'h3aa77b12),
	.w7(32'h3a153870),
	.w8(32'hbab94ed5),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefb788),
	.w1(32'hbbc401d5),
	.w2(32'hbbce4fb4),
	.w3(32'hbbd7d0c2),
	.w4(32'hbb84475e),
	.w5(32'hbb47e28a),
	.w6(32'hbbff04bf),
	.w7(32'hbb029ffc),
	.w8(32'hbb02ab3d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97bbd9d),
	.w1(32'h383c9926),
	.w2(32'h390f0cf9),
	.w3(32'hbab8e4d7),
	.w4(32'hba091c81),
	.w5(32'hb9f1d2d4),
	.w6(32'hba26c8ac),
	.w7(32'h38a7ad25),
	.w8(32'hbb0ba423),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986e0b6),
	.w1(32'hb9bef2ac),
	.w2(32'hb9670b30),
	.w3(32'hb9f62e62),
	.w4(32'h3a11b302),
	.w5(32'hb9aebee0),
	.w6(32'hb9b80773),
	.w7(32'h3974683e),
	.w8(32'hba478f68),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0afe28),
	.w1(32'hba838be0),
	.w2(32'hba8b8e2e),
	.w3(32'hba6c97ea),
	.w4(32'h3925be56),
	.w5(32'hbaa01647),
	.w6(32'hba988e7c),
	.w7(32'h3a32d4de),
	.w8(32'hba8c1b15),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f731b),
	.w1(32'hba1559c7),
	.w2(32'h39244ec0),
	.w3(32'h3a11d444),
	.w4(32'h396d8a42),
	.w5(32'hb981b8ca),
	.w6(32'h3a22c2c9),
	.w7(32'hb607352b),
	.w8(32'hb9248e0f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80a815),
	.w1(32'hb8a39aea),
	.w2(32'hba398e28),
	.w3(32'hba8acbe0),
	.w4(32'hba20f4b6),
	.w5(32'h3a4f2f1e),
	.w6(32'hba4afff2),
	.w7(32'hb9823236),
	.w8(32'h3b03b84d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24e4d9),
	.w1(32'h3b1d892d),
	.w2(32'h3b1f50c5),
	.w3(32'h3b07dc12),
	.w4(32'h3ae4ae94),
	.w5(32'h372052fd),
	.w6(32'h3b2b9077),
	.w7(32'h3b19eb71),
	.w8(32'h39ec696c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb737d0be),
	.w1(32'h3a1873ac),
	.w2(32'hb95b865e),
	.w3(32'h3a42db85),
	.w4(32'hb9900e19),
	.w5(32'hb83dd590),
	.w6(32'h3a43b5e7),
	.w7(32'h38c77fe7),
	.w8(32'h3977a7d1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa78a1a),
	.w1(32'h3ab8f176),
	.w2(32'h39bcba98),
	.w3(32'hba4e0fab),
	.w4(32'h3a8bf360),
	.w5(32'hba3da17c),
	.w6(32'hbaecf964),
	.w7(32'hba415da4),
	.w8(32'hba57ed28),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ac7dc),
	.w1(32'hbb758fb3),
	.w2(32'hbc025bfc),
	.w3(32'hbbdc2d01),
	.w4(32'hbba5ab01),
	.w5(32'hbbe96865),
	.w6(32'hbbb05f6f),
	.w7(32'hbb938ef1),
	.w8(32'hbbd0c6b1),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cb4e1),
	.w1(32'hbae4f466),
	.w2(32'hbb5614a9),
	.w3(32'hbb1e450e),
	.w4(32'hba69df12),
	.w5(32'hbb118b54),
	.w6(32'hbb0a9d24),
	.w7(32'hba1469e3),
	.w8(32'hbb13777c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba861e1),
	.w1(32'hbb6f83df),
	.w2(32'hbb84e689),
	.w3(32'hbb84cb42),
	.w4(32'hbb05d63e),
	.w5(32'hbb253c29),
	.w6(32'hbb77b91a),
	.w7(32'hbada278c),
	.w8(32'hbb638d4f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c34df0),
	.w1(32'h387e7dc2),
	.w2(32'h3ac513a5),
	.w3(32'h3ad044b1),
	.w4(32'h3b0888ff),
	.w5(32'hba428eec),
	.w6(32'h3af359ce),
	.w7(32'h3ada3aff),
	.w8(32'h39fabeb3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ce038),
	.w1(32'hbab96209),
	.w2(32'hbb17a2c4),
	.w3(32'hb99314bb),
	.w4(32'hb9d83bb1),
	.w5(32'h3a04d2b0),
	.w6(32'h3a3b1680),
	.w7(32'hba435164),
	.w8(32'h39fb850a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a601253),
	.w1(32'h3a849542),
	.w2(32'h3a873063),
	.w3(32'h3a0b1276),
	.w4(32'h398becff),
	.w5(32'h3ab8d63b),
	.w6(32'h39ddbbd3),
	.w7(32'h3a0c2e49),
	.w8(32'h3a9d3ee6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b334d),
	.w1(32'h3a47bcb4),
	.w2(32'h3adf83db),
	.w3(32'h3a819d22),
	.w4(32'h3a4a7a96),
	.w5(32'h3abc874b),
	.w6(32'h38bbce94),
	.w7(32'h3a7443da),
	.w8(32'h3aeeac2d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb390b60),
	.w1(32'hbab391a5),
	.w2(32'hbba46cd3),
	.w3(32'hb9dd4a47),
	.w4(32'hb90bbde7),
	.w5(32'hbb0ffe39),
	.w6(32'hba48a829),
	.w7(32'hb9a59154),
	.w8(32'hbb320c88),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a027b2),
	.w1(32'h3a7de743),
	.w2(32'h37f253d6),
	.w3(32'h3a02932b),
	.w4(32'hb9a9cead),
	.w5(32'hbb6a216a),
	.w6(32'h3af37025),
	.w7(32'h3a33d3d7),
	.w8(32'hbb8296ab),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97d7e26),
	.w1(32'hb9ce69e4),
	.w2(32'hbabd792a),
	.w3(32'h3a441eff),
	.w4(32'hb876239d),
	.w5(32'h39e97c9d),
	.w6(32'h3a8c1e03),
	.w7(32'hb7b4ee13),
	.w8(32'h3961a09f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfc582),
	.w1(32'hbace27c9),
	.w2(32'hbaff5ec8),
	.w3(32'hbb2bd9df),
	.w4(32'hbaddde25),
	.w5(32'hbb0173c4),
	.w6(32'hbab827fe),
	.w7(32'hb9c9a5ba),
	.w8(32'hbadaca33),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba335f9c),
	.w1(32'hbac91d9d),
	.w2(32'hba9b3352),
	.w3(32'hba94ed8d),
	.w4(32'hb9b1f539),
	.w5(32'hbac3f7a6),
	.w6(32'hb9cf65d8),
	.w7(32'hba3d541f),
	.w8(32'hbaab54b5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c06226),
	.w1(32'hb9e4eb8f),
	.w2(32'hbb0714c3),
	.w3(32'hba84a650),
	.w4(32'h396ada1d),
	.w5(32'hbadf00b7),
	.w6(32'hbae18365),
	.w7(32'hba8cc16a),
	.w8(32'hbb29d80e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae052d),
	.w1(32'hba695fdf),
	.w2(32'hba6bc488),
	.w3(32'hbabd222a),
	.w4(32'hba12b67a),
	.w5(32'hb9558bc2),
	.w6(32'hba7fdbdb),
	.w7(32'hba55820a),
	.w8(32'hba26cdbc),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09fb4c),
	.w1(32'hbb96f2cd),
	.w2(32'hbbf109dc),
	.w3(32'hbbf19c4c),
	.w4(32'hba62cda3),
	.w5(32'hbb850f35),
	.w6(32'hbb041a64),
	.w7(32'h3b1177ab),
	.w8(32'hbb416954),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396124e9),
	.w1(32'h39a14dd3),
	.w2(32'h399a783d),
	.w3(32'h3a84d68e),
	.w4(32'h39c33f20),
	.w5(32'hb9c24ee9),
	.w6(32'h3aab5baa),
	.w7(32'h3a3277ab),
	.w8(32'hba6f3e01),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fe957),
	.w1(32'h3a2b4b55),
	.w2(32'hba42d189),
	.w3(32'hbb110237),
	.w4(32'hb848d39d),
	.w5(32'h3a6cfef2),
	.w6(32'hbb535829),
	.w7(32'hbaba19c0),
	.w8(32'h3aa83d48),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule