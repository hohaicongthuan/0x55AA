module layer_10_featuremap_486(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07e39d),
	.w1(32'h39af4324),
	.w2(32'h3a727047),
	.w3(32'hbc02ac59),
	.w4(32'h38c429e0),
	.w5(32'h3a9791a7),
	.w6(32'hbbcfcabe),
	.w7(32'hbb05e21f),
	.w8(32'hbb555dcb),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc180f60),
	.w1(32'hbc0025c1),
	.w2(32'hbc3f96e3),
	.w3(32'hbb12f37c),
	.w4(32'h3bf22a8c),
	.w5(32'hb837081d),
	.w6(32'hbbf432bb),
	.w7(32'hbb80b6ba),
	.w8(32'hbbbaccd9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb827350),
	.w1(32'h3bcbf156),
	.w2(32'h3b6f01fc),
	.w3(32'h3a19e234),
	.w4(32'hbb3c6b08),
	.w5(32'hbbf95f61),
	.w6(32'h3b54ad2c),
	.w7(32'h3b2af634),
	.w8(32'h3c2054c5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08dcca),
	.w1(32'hbbc9c935),
	.w2(32'hba6dfa5a),
	.w3(32'hbb74162b),
	.w4(32'hbbb11054),
	.w5(32'hbbbd9852),
	.w6(32'h3beb2bcd),
	.w7(32'hbba77961),
	.w8(32'hbb8261d9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30f849),
	.w1(32'h3a857804),
	.w2(32'hba805bb9),
	.w3(32'hbb9b9840),
	.w4(32'h3b49238f),
	.w5(32'h3b3673ff),
	.w6(32'h3bb0ab4a),
	.w7(32'h3ae192b6),
	.w8(32'h3b97d2af),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94c713),
	.w1(32'hbb45e84d),
	.w2(32'h3a32da2c),
	.w3(32'h3a211093),
	.w4(32'h3b665720),
	.w5(32'hbafb0fcb),
	.w6(32'hba3172ee),
	.w7(32'hbb96c8e1),
	.w8(32'hbc010580),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada1e40),
	.w1(32'hbc2550f6),
	.w2(32'hbc46f087),
	.w3(32'h3ae3caa0),
	.w4(32'hbbb779a9),
	.w5(32'h3b3e4942),
	.w6(32'h3a53be97),
	.w7(32'hbbc3c61e),
	.w8(32'hbc63b6bc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc893dfc),
	.w1(32'hbc261c4b),
	.w2(32'hbc4b09c7),
	.w3(32'hbc686da4),
	.w4(32'h3a9a5bec),
	.w5(32'h3c17aae9),
	.w6(32'hbc51c897),
	.w7(32'h3973d9f0),
	.w8(32'hbc18f998),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda52c7),
	.w1(32'hba0c552d),
	.w2(32'hbb355e58),
	.w3(32'h3c3fe1ea),
	.w4(32'hb856336e),
	.w5(32'hbaacbc6d),
	.w6(32'h3b66b519),
	.w7(32'hbaaa21f1),
	.w8(32'h3acd05e4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97c763),
	.w1(32'hb95c9d1d),
	.w2(32'hbb90ca70),
	.w3(32'hbc240321),
	.w4(32'hbc07b32d),
	.w5(32'hbc8e1497),
	.w6(32'hbbcb852d),
	.w7(32'hbbedbc61),
	.w8(32'hbc6845a3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46ee73),
	.w1(32'hbb36d712),
	.w2(32'h3a5aa390),
	.w3(32'hbbed8509),
	.w4(32'hbbc841ec),
	.w5(32'hbaa3ca80),
	.w6(32'hbbfde4da),
	.w7(32'hb90ed819),
	.w8(32'h3b8d597c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77bc25),
	.w1(32'h3afa4b81),
	.w2(32'hba1c8a5d),
	.w3(32'hbc052ce4),
	.w4(32'h3b23f33a),
	.w5(32'hb8c136f5),
	.w6(32'hbacaa92d),
	.w7(32'h3b41a8f3),
	.w8(32'hbb00b197),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62a1dc),
	.w1(32'hbbd74b5d),
	.w2(32'hbc9681d6),
	.w3(32'hbbc4de16),
	.w4(32'h3a252565),
	.w5(32'hbc8da42c),
	.w6(32'hbb7e9310),
	.w7(32'hbb83163b),
	.w8(32'hbc1923c7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4a39),
	.w1(32'hba32088c),
	.w2(32'hbb089d85),
	.w3(32'hbc083dbb),
	.w4(32'hbb6d137d),
	.w5(32'hbbed1d4e),
	.w6(32'h3bdc2fa6),
	.w7(32'hba843d4c),
	.w8(32'h3b93391e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4323e2),
	.w1(32'h38d2a46a),
	.w2(32'hba603f65),
	.w3(32'hbb2f0cbd),
	.w4(32'hbbd62a03),
	.w5(32'hbc1b47ec),
	.w6(32'hba809c3e),
	.w7(32'h3b135ff9),
	.w8(32'h3a052b0e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10148f),
	.w1(32'hbc2dbddb),
	.w2(32'hbc5b47e1),
	.w3(32'hbb8718a4),
	.w4(32'hbb9e0b94),
	.w5(32'hbc3335a9),
	.w6(32'hbc0dfa1a),
	.w7(32'hbba92f44),
	.w8(32'hbbe70c7a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6e8c8),
	.w1(32'h3b87bdeb),
	.w2(32'h3b71e32c),
	.w3(32'hbb3ff113),
	.w4(32'hbab9c95f),
	.w5(32'hbb0eea25),
	.w6(32'hbb3ee714),
	.w7(32'hbb911623),
	.w8(32'hba84da8f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dca54),
	.w1(32'h3ad37582),
	.w2(32'hbacf6486),
	.w3(32'hbba5dc33),
	.w4(32'hbb0d85c9),
	.w5(32'hbc20e454),
	.w6(32'hbbb040d3),
	.w7(32'hbbd5efd2),
	.w8(32'hbc4d0a10),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad23ebd),
	.w1(32'hbaf6a794),
	.w2(32'hbbfa9203),
	.w3(32'hbb41ebcf),
	.w4(32'hbbc77dd8),
	.w5(32'hbc6bc03e),
	.w6(32'hb9ecaf98),
	.w7(32'h398f8109),
	.w8(32'hbbddfc23),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb566fdb),
	.w1(32'h3b89e059),
	.w2(32'h3b87518e),
	.w3(32'hbb757e0c),
	.w4(32'hbbbb685b),
	.w5(32'hbb3dab4a),
	.w6(32'hbbcfd8d0),
	.w7(32'hb968d231),
	.w8(32'hbba1fea3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d4aef),
	.w1(32'h3a71fb2c),
	.w2(32'h3b4356f9),
	.w3(32'hbc30fb33),
	.w4(32'h3b132dce),
	.w5(32'h3a1d10c4),
	.w6(32'hba6cdd93),
	.w7(32'h3b04f1e5),
	.w8(32'hba08a60e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12e2a4),
	.w1(32'h3bd817f6),
	.w2(32'h3b872d41),
	.w3(32'hb974d34f),
	.w4(32'h3bfc8b05),
	.w5(32'h3a6739a2),
	.w6(32'hb987deae),
	.w7(32'h3c3d7d0a),
	.w8(32'h3ae7a81d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f5136),
	.w1(32'hbab432f2),
	.w2(32'hb9ec0c91),
	.w3(32'hbc0bc7ee),
	.w4(32'h3b187b3b),
	.w5(32'hbb9d318e),
	.w6(32'hb9a02b8e),
	.w7(32'hbb2452a9),
	.w8(32'hbc7a167f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a9122),
	.w1(32'hbb9a33e0),
	.w2(32'hbc4bdd16),
	.w3(32'hbb19065b),
	.w4(32'hbb16f338),
	.w5(32'hbc20d6b6),
	.w6(32'hbbb40f4d),
	.w7(32'hba7a991d),
	.w8(32'hbbe29617),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6dbbe7),
	.w1(32'hbba92de7),
	.w2(32'hbbbbec1d),
	.w3(32'hbc4aa681),
	.w4(32'hbb5830a3),
	.w5(32'hbc1fefad),
	.w6(32'hbc67ec1d),
	.w7(32'h3bd0b1a0),
	.w8(32'hb9ca1713),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb834433),
	.w1(32'h3b4f7a96),
	.w2(32'h3b2311c8),
	.w3(32'hbb03a100),
	.w4(32'h3b05daa2),
	.w5(32'h39ade511),
	.w6(32'h3a8dbea3),
	.w7(32'h3b77169d),
	.w8(32'h3ad03eab),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b809ef9),
	.w1(32'h3a71ef66),
	.w2(32'h3aaefd10),
	.w3(32'hb82fbb12),
	.w4(32'hbb4d193e),
	.w5(32'hba31b152),
	.w6(32'h3aff3433),
	.w7(32'hba5bdfaf),
	.w8(32'hbbcb6629),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c44e0),
	.w1(32'hb955bfe6),
	.w2(32'hbabf8244),
	.w3(32'h3af5b143),
	.w4(32'hbabd0e80),
	.w5(32'h39f1b714),
	.w6(32'hbbe67b45),
	.w7(32'hbb421458),
	.w8(32'h3ac7541d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19de1b),
	.w1(32'h3bae43be),
	.w2(32'hba87aab2),
	.w3(32'hbbd632d7),
	.w4(32'hba818720),
	.w5(32'hba9ad871),
	.w6(32'hbc2ae954),
	.w7(32'hbba47bfd),
	.w8(32'hbba53bea),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f875d2),
	.w1(32'h3bfa518f),
	.w2(32'hb9c96b0b),
	.w3(32'hba9587b1),
	.w4(32'h3b588aa5),
	.w5(32'h3b0efb16),
	.w6(32'hbc116f04),
	.w7(32'h3a9140ee),
	.w8(32'hbba51799),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ec8b1),
	.w1(32'h3af9757d),
	.w2(32'h3945bf73),
	.w3(32'h3b71d182),
	.w4(32'hbb5e7dd7),
	.w5(32'hbb3c64fe),
	.w6(32'h3ac9b772),
	.w7(32'hbb87de9b),
	.w8(32'hbb6fb051),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c1fc3),
	.w1(32'hbc1e0915),
	.w2(32'hbc0ec7b3),
	.w3(32'h3ae25843),
	.w4(32'hba6fb733),
	.w5(32'hba3f8f39),
	.w6(32'hbb89603e),
	.w7(32'hbb4bacc6),
	.w8(32'h3a54fc9e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9264f),
	.w1(32'hbc0f0ba7),
	.w2(32'hbc403233),
	.w3(32'hbb027571),
	.w4(32'hba29ccad),
	.w5(32'hbc0d0e5e),
	.w6(32'h3b31024a),
	.w7(32'h3a84dc1a),
	.w8(32'h3c37e7b2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15b339),
	.w1(32'hbb3e65a0),
	.w2(32'hbb426398),
	.w3(32'hbc68574d),
	.w4(32'hba2b4f79),
	.w5(32'hbab9a7a3),
	.w6(32'h3be4b26a),
	.w7(32'h3bbd1919),
	.w8(32'h3c15767b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae3e7a),
	.w1(32'h3b4fc5fa),
	.w2(32'h3b313450),
	.w3(32'hbb608793),
	.w4(32'hbabfe472),
	.w5(32'hbb71c227),
	.w6(32'h3bd24913),
	.w7(32'hb8bc72ee),
	.w8(32'h3a0764c9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbf3ff),
	.w1(32'hbb3a7940),
	.w2(32'hbb72bf5b),
	.w3(32'h3aef477f),
	.w4(32'hbb4990e4),
	.w5(32'hbc297920),
	.w6(32'hba50ee22),
	.w7(32'hbb077393),
	.w8(32'hbbc994c9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e04ef),
	.w1(32'h3bd393b3),
	.w2(32'hbbd88416),
	.w3(32'hbb80bb4c),
	.w4(32'h3b9e22a5),
	.w5(32'hbbec9fd7),
	.w6(32'h3b94bb4e),
	.w7(32'h3c39132b),
	.w8(32'hbab579cb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba65d9),
	.w1(32'hbb1518c2),
	.w2(32'hbc040ec6),
	.w3(32'hbc94a423),
	.w4(32'h3ca88772),
	.w5(32'h3c5f1bcb),
	.w6(32'hbcb6cd18),
	.w7(32'hba86816f),
	.w8(32'hba5e1600),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bef30),
	.w1(32'h3c95fbe4),
	.w2(32'h3c91aef5),
	.w3(32'hbc8a4baf),
	.w4(32'h3bbd038b),
	.w5(32'h3b9c7505),
	.w6(32'hbc81c901),
	.w7(32'h3b86136e),
	.w8(32'h3bcb405c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac0220),
	.w1(32'hbbc133a6),
	.w2(32'hbb3d9c5f),
	.w3(32'hbae24cfc),
	.w4(32'h3b16f002),
	.w5(32'h3c26421a),
	.w6(32'hbbac2d07),
	.w7(32'hbbc0dca2),
	.w8(32'hbb9d3035),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f8e09),
	.w1(32'hbbaf6941),
	.w2(32'hbbd50d7e),
	.w3(32'h3bcdc18e),
	.w4(32'hb99edbb9),
	.w5(32'hbbbf3886),
	.w6(32'h38bb3826),
	.w7(32'hbac16041),
	.w8(32'hba5c817b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde4681),
	.w1(32'hbb827372),
	.w2(32'hbbc87f8d),
	.w3(32'h3ae1c54f),
	.w4(32'hbbd21a2d),
	.w5(32'hbc192b80),
	.w6(32'h3b39ab89),
	.w7(32'h3b71d1ad),
	.w8(32'h3b82076e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d627d),
	.w1(32'hbb9da8bf),
	.w2(32'hbb63e8ad),
	.w3(32'hbb6bf46f),
	.w4(32'h3bf661e8),
	.w5(32'hba1521ee),
	.w6(32'hbc07977e),
	.w7(32'hb9ead575),
	.w8(32'hbb102f2e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc442b77),
	.w1(32'hb9a6d417),
	.w2(32'hbbcc7bbb),
	.w3(32'hbc1d9567),
	.w4(32'hbb04d373),
	.w5(32'hbbe8c1fb),
	.w6(32'hbb82c378),
	.w7(32'hbc101304),
	.w8(32'hbc5718cc),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14d16a),
	.w1(32'hba4dd22a),
	.w2(32'hbc5c503c),
	.w3(32'hbbb1dfaa),
	.w4(32'h3bd1e585),
	.w5(32'hbb432d9a),
	.w6(32'hbb47acd9),
	.w7(32'h3c2e3b61),
	.w8(32'h3a4c0682),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95c654),
	.w1(32'hbb03f3f2),
	.w2(32'hbc2b5f05),
	.w3(32'hba80b72c),
	.w4(32'h3b44c848),
	.w5(32'hbbd6ee3c),
	.w6(32'hbc27e354),
	.w7(32'h3ab4e1a8),
	.w8(32'hbc0c2cbd),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a63fc),
	.w1(32'h3c0c4853),
	.w2(32'h3bc003a4),
	.w3(32'hbc007726),
	.w4(32'hbc24b6e3),
	.w5(32'hbc495ec2),
	.w6(32'hbbdbc0eb),
	.w7(32'hbb8ec34c),
	.w8(32'hbc52e0b2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbadeb6),
	.w1(32'h3b40b9ee),
	.w2(32'hbbb8af9f),
	.w3(32'hbc349b20),
	.w4(32'hbb218378),
	.w5(32'hbc243c28),
	.w6(32'hbc309854),
	.w7(32'h397970e9),
	.w8(32'hbbd5a048),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e51e6),
	.w1(32'h3b4b20a3),
	.w2(32'h34fc7280),
	.w3(32'h3afa8474),
	.w4(32'hba1b7802),
	.w5(32'hbb0854e9),
	.w6(32'h3a28579e),
	.w7(32'hbbf3642b),
	.w8(32'hbc3f6e30),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb406f4b),
	.w1(32'h3b2200ac),
	.w2(32'h3aa3d1c3),
	.w3(32'hba27d886),
	.w4(32'h3af1f20a),
	.w5(32'hba35ef85),
	.w6(32'hbc31bd71),
	.w7(32'h39d1d9b8),
	.w8(32'hbbada04c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba161b1),
	.w1(32'hbb049c1c),
	.w2(32'hbc04852e),
	.w3(32'h3be97bb8),
	.w4(32'hbb55fc7b),
	.w5(32'hbbe243f1),
	.w6(32'hbba35d81),
	.w7(32'h3accc034),
	.w8(32'h3ae2cf6f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6411d),
	.w1(32'hbba244cf),
	.w2(32'hbc0ee4dc),
	.w3(32'hbb47da99),
	.w4(32'h39837730),
	.w5(32'hbba20b76),
	.w6(32'hbb9a1c58),
	.w7(32'hbbc06a38),
	.w8(32'hbbabf098),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb004881),
	.w1(32'hbb2f43e8),
	.w2(32'hbbf09232),
	.w3(32'hbacc9328),
	.w4(32'h3bc4b904),
	.w5(32'h3c1585be),
	.w6(32'h3a12d4f3),
	.w7(32'h3b6c4b66),
	.w8(32'h3ae97790),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e7bc2),
	.w1(32'hbc6e5d05),
	.w2(32'hbcab80d2),
	.w3(32'h3ad89712),
	.w4(32'h3c10c6c7),
	.w5(32'h3c3f4493),
	.w6(32'hbb04e64e),
	.w7(32'hbb6c6cf0),
	.w8(32'hbc038cea),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27da44),
	.w1(32'h3abc1d01),
	.w2(32'hba602928),
	.w3(32'h3baaf12a),
	.w4(32'h3bf34353),
	.w5(32'h3c067adc),
	.w6(32'h3bb9f849),
	.w7(32'hbb869e83),
	.w8(32'hbab4440d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf57b8),
	.w1(32'hbc3b6a4b),
	.w2(32'hbbf4a34b),
	.w3(32'hbae0ad58),
	.w4(32'h3c8a9a5c),
	.w5(32'h3c3cf70b),
	.w6(32'hb9826853),
	.w7(32'hbc2ea72e),
	.w8(32'hbba8cd2f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba23c83),
	.w1(32'hbb88f5f3),
	.w2(32'hbbbe64ca),
	.w3(32'hbaf3d578),
	.w4(32'hbba2baab),
	.w5(32'hbbba3a9f),
	.w6(32'h3bdf6239),
	.w7(32'hbb0a8f36),
	.w8(32'hbba498ea),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb540a44),
	.w1(32'hbb5021c1),
	.w2(32'hbb296cb3),
	.w3(32'hbb5fc652),
	.w4(32'hbb964e8e),
	.w5(32'hbb52e9b4),
	.w6(32'hbbc1e46e),
	.w7(32'hb7988ba8),
	.w8(32'h3b31024e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1011e1),
	.w1(32'h3a9e8482),
	.w2(32'hbb735177),
	.w3(32'hbb9aea66),
	.w4(32'h3bb4b6f1),
	.w5(32'hbb37602f),
	.w6(32'h3a9de7a2),
	.w7(32'hbab33610),
	.w8(32'hbac7c21c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b007cb2),
	.w1(32'h3b243262),
	.w2(32'h3b3cd5db),
	.w3(32'h3ad1e34b),
	.w4(32'h3b16b4e7),
	.w5(32'h3ae05112),
	.w6(32'hbafa7493),
	.w7(32'hb9a633e3),
	.w8(32'hbc278d31),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad2020),
	.w1(32'h3a9dfca5),
	.w2(32'h3b556877),
	.w3(32'hbb294ff6),
	.w4(32'hbb59a13a),
	.w5(32'h3b79641b),
	.w6(32'hbbd9c8f4),
	.w7(32'hb9877fec),
	.w8(32'h3aba82f4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f50a1),
	.w1(32'h3a044177),
	.w2(32'hbb643e72),
	.w3(32'h3b1d30a4),
	.w4(32'hbb61dce1),
	.w5(32'hbc1accbd),
	.w6(32'h3acdad05),
	.w7(32'hba022575),
	.w8(32'hbb98d725),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66b3f9),
	.w1(32'hbc082fb8),
	.w2(32'hbb44d3ed),
	.w3(32'hbab44805),
	.w4(32'hbb7324ee),
	.w5(32'hbbf74622),
	.w6(32'hbbb3a5e9),
	.w7(32'hbbb76acb),
	.w8(32'hbbbdcfbf),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38daa3d0),
	.w1(32'hbad2a25e),
	.w2(32'hbb03f8da),
	.w3(32'hbb9a92f4),
	.w4(32'h3aa97cab),
	.w5(32'h3a56a60a),
	.w6(32'hbb7b3f65),
	.w7(32'hbb0c45b9),
	.w8(32'hbaa7d393),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52447d),
	.w1(32'h3b78ec74),
	.w2(32'h3aa33fef),
	.w3(32'hbab4ad80),
	.w4(32'h3bce8c2f),
	.w5(32'h3b8183db),
	.w6(32'hbb58eb46),
	.w7(32'h3b180477),
	.w8(32'hbb1117bd),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00c8ff),
	.w1(32'hba90a9fa),
	.w2(32'hba595bd5),
	.w3(32'h3b19f1ef),
	.w4(32'h3a9d2ebd),
	.w5(32'hbb861430),
	.w6(32'h3b320ff6),
	.w7(32'h3b854665),
	.w8(32'h3b0fbfb0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc643674),
	.w1(32'hbbbe4f66),
	.w2(32'hbc2ccd68),
	.w3(32'hbc060419),
	.w4(32'hbbea9b24),
	.w5(32'hbbd72cf8),
	.w6(32'hbc0b3daa),
	.w7(32'hbc0ecdda),
	.w8(32'hbc43ccd4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79da2b),
	.w1(32'h3b43bbac),
	.w2(32'hbc0759d0),
	.w3(32'hbc3d114d),
	.w4(32'hb9a8dbc8),
	.w5(32'hbc4fceaa),
	.w6(32'hbc1b7601),
	.w7(32'hbb0f318b),
	.w8(32'hbc7895e8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fe624),
	.w1(32'h3bb7e098),
	.w2(32'hbb9b4bc2),
	.w3(32'hbc3daeb2),
	.w4(32'h3c0dadfb),
	.w5(32'hbb638fca),
	.w6(32'hbcac16d9),
	.w7(32'h3b09a15f),
	.w8(32'h3b82fa8e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84a7a6),
	.w1(32'h3ba691dd),
	.w2(32'hbc2a001b),
	.w3(32'hbc71b788),
	.w4(32'h3c26b575),
	.w5(32'hbaa81e39),
	.w6(32'hbc9d76a1),
	.w7(32'h3c492ed8),
	.w8(32'hbae05a55),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39856f94),
	.w1(32'h3794e5b6),
	.w2(32'h381daf4e),
	.w3(32'h3975eddb),
	.w4(32'hb7e85094),
	.w5(32'hb702f2ae),
	.w6(32'h39911f19),
	.w7(32'h37d7dcfd),
	.w8(32'h387fb213),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da8ee3),
	.w1(32'h388bb55b),
	.w2(32'h3919c747),
	.w3(32'h39be3b62),
	.w4(32'h35bf7338),
	.w5(32'h38c32a78),
	.w6(32'h39eacb8d),
	.w7(32'h38f8b079),
	.w8(32'h396fe48a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad2820),
	.w1(32'hb827df3a),
	.w2(32'h3805ef86),
	.w3(32'h39acaf81),
	.w4(32'hb91106a1),
	.w5(32'hb7e48476),
	.w6(32'h39d8c360),
	.w7(32'hb8217327),
	.w8(32'h38a2e336),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae94939),
	.w1(32'h3a5f6a25),
	.w2(32'hb834f14e),
	.w3(32'hbad18cd8),
	.w4(32'hb9053247),
	.w5(32'hba1fd85c),
	.w6(32'hbb09a150),
	.w7(32'hba12c045),
	.w8(32'hba3cddcc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a64d18),
	.w1(32'h38a353a3),
	.w2(32'h38e5ae22),
	.w3(32'h398f0ed3),
	.w4(32'h379052a8),
	.w5(32'h388f9356),
	.w6(32'h39bb3260),
	.w7(32'h38b4e16e),
	.w8(32'h39069474),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7e575),
	.w1(32'hba99f8f4),
	.w2(32'hbaf94307),
	.w3(32'hbab0db1c),
	.w4(32'hbb09187b),
	.w5(32'hbb0f384b),
	.w6(32'h39e02c25),
	.w7(32'hb982912c),
	.w8(32'hbaad029d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a2738),
	.w1(32'hbb5ddd66),
	.w2(32'hbbeb40f9),
	.w3(32'hbbd0467b),
	.w4(32'hbb55a147),
	.w5(32'hbb8e66f5),
	.w6(32'hbbc93900),
	.w7(32'hbb0f06b4),
	.w8(32'hbbeb87be),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a6373),
	.w1(32'hbb87289c),
	.w2(32'hbc102cdb),
	.w3(32'hbbe20b62),
	.w4(32'hbaa270c1),
	.w5(32'hbbccea99),
	.w6(32'hbb8e19a1),
	.w7(32'h3ad6fa77),
	.w8(32'hbb51c1c2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dbfc6),
	.w1(32'h38ca1b18),
	.w2(32'hbb86b545),
	.w3(32'hbb72519a),
	.w4(32'h3a353eb1),
	.w5(32'hbb22dc1a),
	.w6(32'hbb849fd6),
	.w7(32'h3a231ba7),
	.w8(32'hbb1c5429),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b56dc),
	.w1(32'h3a1bb70e),
	.w2(32'hbb8894d3),
	.w3(32'hba605815),
	.w4(32'hbb0001f2),
	.w5(32'hbb781c22),
	.w6(32'h3a07535e),
	.w7(32'h39aa3e0e),
	.w8(32'hbb87824a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a527a),
	.w1(32'hb98bcd78),
	.w2(32'hbb661a02),
	.w3(32'hbb3d4533),
	.w4(32'h3a13a56b),
	.w5(32'hbb002432),
	.w6(32'hbb3b0df9),
	.w7(32'h3a19b425),
	.w8(32'hbac96d5d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba848496),
	.w1(32'hb903420d),
	.w2(32'hbb7afa11),
	.w3(32'hba0fd91c),
	.w4(32'hba854b24),
	.w5(32'hbb9b9750),
	.w6(32'h39de5a0f),
	.w7(32'h397f3ff0),
	.w8(32'hbb866328),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3842b41c),
	.w1(32'h36fca2d8),
	.w2(32'h37b4a201),
	.w3(32'h383d9fa0),
	.w4(32'h35272a54),
	.w5(32'h37a38260),
	.w6(32'h3856bef9),
	.w7(32'hb722db7c),
	.w8(32'h37bf0972),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381daff6),
	.w1(32'h3803c256),
	.w2(32'h38089b88),
	.w3(32'h380ccb38),
	.w4(32'h38099dcc),
	.w5(32'h36bcb2f0),
	.w6(32'h388ddee8),
	.w7(32'h37f6b94e),
	.w8(32'h36053109),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38797430),
	.w1(32'h3809accf),
	.w2(32'h38b0ba63),
	.w3(32'hb8689e45),
	.w4(32'hb8055eb4),
	.w5(32'h3814f25d),
	.w6(32'h37fc8d69),
	.w7(32'h37d69ac4),
	.w8(32'h380737c6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396dbc80),
	.w1(32'h3a28e891),
	.w2(32'h39f28896),
	.w3(32'h3921c26f),
	.w4(32'h3a017eb6),
	.w5(32'h3987410f),
	.w6(32'hb8a325c3),
	.w7(32'h39d5e162),
	.w8(32'h392cb359),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1be7bf),
	.w1(32'h39d27c34),
	.w2(32'hba23aa68),
	.w3(32'hbc06c2aa),
	.w4(32'h3b171811),
	.w5(32'h3b36c879),
	.w6(32'hbc0ea3f6),
	.w7(32'h3b6a1186),
	.w8(32'h3a84f2eb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8d35b),
	.w1(32'h39b5e54f),
	.w2(32'h3a15a495),
	.w3(32'h3a8cc8a9),
	.w4(32'h3aa41eaf),
	.w5(32'h3a8f50c5),
	.w6(32'hba42c577),
	.w7(32'h38320fe7),
	.w8(32'h39b28bec),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7682b),
	.w1(32'hba7415c3),
	.w2(32'hbbcd02a2),
	.w3(32'hbb18da6b),
	.w4(32'h39400753),
	.w5(32'hbba77fb7),
	.w6(32'hbb416ec8),
	.w7(32'h3ac6ae85),
	.w8(32'hbb9a7581),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17aeef),
	.w1(32'hbb242b0e),
	.w2(32'hbb99ec88),
	.w3(32'hbc2c60e2),
	.w4(32'hbab912c1),
	.w5(32'hbb499fe4),
	.w6(32'hbc2e3b64),
	.w7(32'hbbb14e5b),
	.w8(32'hbbb1e9a9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66134b),
	.w1(32'h3b632655),
	.w2(32'h3ad81c01),
	.w3(32'hbba520bc),
	.w4(32'h3b4568d3),
	.w5(32'h3b332ee3),
	.w6(32'hbbd8b326),
	.w7(32'h3ad2e19f),
	.w8(32'h3a00a9fd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb394ead),
	.w1(32'hba1a938f),
	.w2(32'hbb62a9a5),
	.w3(32'hbba7f5aa),
	.w4(32'hb9d8793e),
	.w5(32'h3af6935e),
	.w6(32'hbaea6647),
	.w7(32'hbab06f50),
	.w8(32'hbbd0d7e7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ab97c),
	.w1(32'h3bc01fde),
	.w2(32'h3a9df592),
	.w3(32'hb96d9648),
	.w4(32'h3b993ac6),
	.w5(32'h3a2fb449),
	.w6(32'h39f36efe),
	.w7(32'h3ba3001d),
	.w8(32'h3b1521c0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc326173),
	.w1(32'hbb641e9a),
	.w2(32'hbc0ec310),
	.w3(32'hbc1452cd),
	.w4(32'hba3e930e),
	.w5(32'hbb3b5b26),
	.w6(32'hbc2aa463),
	.w7(32'hba9ad3b6),
	.w8(32'hbbc35f8f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3679b),
	.w1(32'h393a4d6f),
	.w2(32'hbb039656),
	.w3(32'hbb819810),
	.w4(32'h3b3a96b9),
	.w5(32'h3ab7b926),
	.w6(32'hbb8b8198),
	.w7(32'h3b0dbaf3),
	.w8(32'hb91bba32),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8a6d9),
	.w1(32'h3b2452e7),
	.w2(32'hbb43c733),
	.w3(32'hbbc2b6fd),
	.w4(32'h3b4a630b),
	.w5(32'hbb1f26df),
	.w6(32'hbbf2421b),
	.w7(32'h3b80aa00),
	.w8(32'hbad3a1f0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11b3de),
	.w1(32'h3a02718d),
	.w2(32'hb7c3e299),
	.w3(32'h3a586956),
	.w4(32'h3a3885af),
	.w5(32'h38be02b5),
	.w6(32'h3a719a48),
	.w7(32'h3a1bc6f3),
	.w8(32'h3a19f871),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1a2df),
	.w1(32'hba5b33b1),
	.w2(32'hbc07aaf6),
	.w3(32'hbb857548),
	.w4(32'h3b1d30f3),
	.w5(32'hbbabf456),
	.w6(32'hbb781eb0),
	.w7(32'h3a4119a8),
	.w8(32'hbbd68c11),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54d845),
	.w1(32'h3adbf7bb),
	.w2(32'hbb4c250c),
	.w3(32'hbb4f3e07),
	.w4(32'h3b6dec6c),
	.w5(32'h3ad605db),
	.w6(32'hbac94cd2),
	.w7(32'h3b1bfc15),
	.w8(32'hbb0b9867),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee94a4),
	.w1(32'h39e20a93),
	.w2(32'hbc026826),
	.w3(32'hbad90963),
	.w4(32'h3b65e3ec),
	.w5(32'hbba3f73b),
	.w6(32'h3a859018),
	.w7(32'h3bd1be8d),
	.w8(32'hbbe17efa),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc938ce5),
	.w1(32'h3c42b5de),
	.w2(32'h3c4fd564),
	.w3(32'hbc69494c),
	.w4(32'h3c9e36cd),
	.w5(32'h3c9e9872),
	.w6(32'hbc8823b3),
	.w7(32'h3c46662b),
	.w8(32'h3bc8fcee),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8ec0f),
	.w1(32'h393267b1),
	.w2(32'hbc2f1850),
	.w3(32'hbb58a167),
	.w4(32'h3b145dbb),
	.w5(32'hbc114448),
	.w6(32'hbb3c779f),
	.w7(32'h3b7d62c0),
	.w8(32'hbbc79328),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9335c6),
	.w1(32'hb6fae761),
	.w2(32'hbba7c3cc),
	.w3(32'hb95b7b49),
	.w4(32'h39ae6b68),
	.w5(32'hbb23d0df),
	.w6(32'h3bb28465),
	.w7(32'h3bab308f),
	.w8(32'hbb98a29e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d5924),
	.w1(32'h39a7c286),
	.w2(32'h391edd78),
	.w3(32'h391d515e),
	.w4(32'h39cf6435),
	.w5(32'h39954c76),
	.w6(32'h3a04801d),
	.w7(32'h38cec5a2),
	.w8(32'h39a8168d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84a3c7),
	.w1(32'hbc2d243a),
	.w2(32'hbc61943d),
	.w3(32'hbc0d59b0),
	.w4(32'hbb6e7693),
	.w5(32'hbc328c91),
	.w6(32'hba92c33e),
	.w7(32'h3b6853fb),
	.w8(32'hbb8d341a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c06ff),
	.w1(32'h392fc70d),
	.w2(32'hbb63e4a4),
	.w3(32'hbb55bc4f),
	.w4(32'hba7bccf1),
	.w5(32'hbba96eb3),
	.w6(32'hb98185fc),
	.w7(32'h3af57057),
	.w8(32'hbb8993da),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939f22b),
	.w1(32'h398e0f14),
	.w2(32'hb806a06f),
	.w3(32'h38c39201),
	.w4(32'h39fba61c),
	.w5(32'h39a16950),
	.w6(32'hb97968b3),
	.w7(32'h395b9a8c),
	.w8(32'hb79410da),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bcf68),
	.w1(32'hbaa7210c),
	.w2(32'hbb1efb53),
	.w3(32'hba97b487),
	.w4(32'hb9f3de30),
	.w5(32'hba471d45),
	.w6(32'hbb0362af),
	.w7(32'hba67e631),
	.w8(32'hba4308a7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96a074),
	.w1(32'hbb3bc305),
	.w2(32'hbbef6673),
	.w3(32'hbb34ccb9),
	.w4(32'hbb0da69e),
	.w5(32'hbbe6ff6a),
	.w6(32'hbb036437),
	.w7(32'hbb667868),
	.w8(32'hbc0ec97b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6af900),
	.w1(32'h3ad8341f),
	.w2(32'hbbada5fb),
	.w3(32'hbaf2a9c9),
	.w4(32'h3b1cff67),
	.w5(32'hbb987167),
	.w6(32'hbad503c1),
	.w7(32'h3b3a58b3),
	.w8(32'hbb18991a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb767b3),
	.w1(32'hba4b166c),
	.w2(32'hbafee082),
	.w3(32'hbbac95c0),
	.w4(32'h3a49f133),
	.w5(32'hba4082fc),
	.w6(32'hbbb5147b),
	.w7(32'hba9a173b),
	.w8(32'hbb3d2cb2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba70300),
	.w1(32'h3a91d967),
	.w2(32'hbb744114),
	.w3(32'hbb7bbc2f),
	.w4(32'h3b129778),
	.w5(32'hbaf286b7),
	.w6(32'hbb2b5b2b),
	.w7(32'h3b2ba613),
	.w8(32'hbadaa8c2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb395272),
	.w1(32'h3b49e926),
	.w2(32'h3a8fd689),
	.w3(32'hbb12e227),
	.w4(32'h3b120986),
	.w5(32'h3986fe57),
	.w6(32'hbbc07c78),
	.w7(32'h3a844d42),
	.w8(32'hbb1d6f4a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ec8a5),
	.w1(32'hbaf24873),
	.w2(32'hbbe0d24e),
	.w3(32'hbb7b88eb),
	.w4(32'hb98bd95e),
	.w5(32'hbb31b210),
	.w6(32'hbb705382),
	.w7(32'hb9fe160a),
	.w8(32'hbb86141f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e041d),
	.w1(32'h3a5903df),
	.w2(32'hbb35d6d4),
	.w3(32'hbb1b01c9),
	.w4(32'h3abb3ac5),
	.w5(32'hbb116305),
	.w6(32'hbb153718),
	.w7(32'h3ad92351),
	.w8(32'hbb0212a4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80fa322),
	.w1(32'hb8005d10),
	.w2(32'hb85a6f45),
	.w3(32'hb790e612),
	.w4(32'hb7aa558e),
	.w5(32'h387d6c8d),
	.w6(32'hb6db209a),
	.w7(32'hb841a210),
	.w8(32'h3696ddaf),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00027e),
	.w1(32'hb98bcbb5),
	.w2(32'hb9711c5e),
	.w3(32'hb97a62d3),
	.w4(32'hb901b975),
	.w5(32'hb7a88434),
	.w6(32'hb9f92907),
	.w7(32'hb9060c81),
	.w8(32'hb92156f2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3832d0f9),
	.w1(32'h39a5815a),
	.w2(32'h394ad148),
	.w3(32'hb8f1deaa),
	.w4(32'h397f496b),
	.w5(32'h3927b667),
	.w6(32'hb8cac907),
	.w7(32'h39406c5a),
	.w8(32'h38eb6d27),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9163e38),
	.w1(32'h39f94676),
	.w2(32'h3a73b468),
	.w3(32'h39436c0d),
	.w4(32'h39ced3ec),
	.w5(32'h3a0fc090),
	.w6(32'h38393948),
	.w7(32'h39bd037d),
	.w8(32'h39400a81),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc65d92),
	.w1(32'h3a28efad),
	.w2(32'hbb768bf2),
	.w3(32'hbb5e3d1a),
	.w4(32'h3ad65575),
	.w5(32'hbb502644),
	.w6(32'hbb6c24f1),
	.w7(32'h3b24b23a),
	.w8(32'hbb2fc5c6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b99bb),
	.w1(32'hb8673d2e),
	.w2(32'h391022c7),
	.w3(32'hba38a62d),
	.w4(32'hb88928ce),
	.w5(32'h390cd39b),
	.w6(32'hba32ff08),
	.w7(32'h38bdbac1),
	.w8(32'hb7f07f33),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaed131),
	.w1(32'hba453e2a),
	.w2(32'hbb76d390),
	.w3(32'hba3efa26),
	.w4(32'hba2a42c4),
	.w5(32'hbb3de1ea),
	.w6(32'h3b0f1e81),
	.w7(32'h39d2c368),
	.w8(32'hbb13fe0b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d78f6),
	.w1(32'h39d96d62),
	.w2(32'hbb16ebee),
	.w3(32'hbc0fa6c9),
	.w4(32'h3a9e54da),
	.w5(32'hb90b2bcc),
	.w6(32'hbc1893ca),
	.w7(32'h3a8ac320),
	.w8(32'hbb068985),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ae238),
	.w1(32'h3756f8b6),
	.w2(32'hb8df0127),
	.w3(32'h398429a4),
	.w4(32'h39066f79),
	.w5(32'h39152feb),
	.w6(32'h39b3a4b7),
	.w7(32'h39a5bc07),
	.w8(32'h394ff3cb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917b731),
	.w1(32'h39a55977),
	.w2(32'hb90a487b),
	.w3(32'h39b37d22),
	.w4(32'h3a1e4f81),
	.w5(32'h3a068f21),
	.w6(32'h38155a50),
	.w7(32'h39acbcbc),
	.w8(32'h377226c6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c367fd),
	.w1(32'h3860fea5),
	.w2(32'h3895a346),
	.w3(32'h38a2f96e),
	.w4(32'h379d4c3a),
	.w5(32'h38722d7e),
	.w6(32'h388fdcef),
	.w7(32'h37b36be8),
	.w8(32'h38762fe5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa09eb6),
	.w1(32'hba5d978c),
	.w2(32'hba633644),
	.w3(32'hba9034fa),
	.w4(32'h37dbcaa0),
	.w5(32'hb9692305),
	.w6(32'hba9b4bb9),
	.w7(32'hba3e2855),
	.w8(32'hbaa178c6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44afcd),
	.w1(32'hbb51feff),
	.w2(32'hbb6d7317),
	.w3(32'h3ae0cc4d),
	.w4(32'hbb7c3546),
	.w5(32'hbbeb9d68),
	.w6(32'hb9b8545b),
	.w7(32'hbb65deed),
	.w8(32'hbbbd9c77),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99435b),
	.w1(32'hbb188bdf),
	.w2(32'hbc22f138),
	.w3(32'hbb6047d8),
	.w4(32'hbac58017),
	.w5(32'hbbe72f74),
	.w6(32'hbb5a2bf6),
	.w7(32'hbaf9711b),
	.w8(32'hbbf87742),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e96cb8),
	.w1(32'hba163294),
	.w2(32'hba3b541e),
	.w3(32'hb99ed930),
	.w4(32'hb97f5a9b),
	.w5(32'h38b683fd),
	.w6(32'h39c06aa9),
	.w7(32'h394269ca),
	.w8(32'hb9dac04b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02bf5e),
	.w1(32'hb9af149a),
	.w2(32'hbaa46ed8),
	.w3(32'hbb3e5369),
	.w4(32'hba45afa1),
	.w5(32'hba62bce8),
	.w6(32'hbb8075b7),
	.w7(32'hba80aef6),
	.w8(32'hba9ea8b5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf521d0),
	.w1(32'h3a87de78),
	.w2(32'hb9f28e74),
	.w3(32'hbb042fc1),
	.w4(32'h3a50bf2f),
	.w5(32'hba16c178),
	.w6(32'hbb18061c),
	.w7(32'h3aa9b0ad),
	.w8(32'hba35545a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ac744),
	.w1(32'h3984e3cf),
	.w2(32'hbb26cf31),
	.w3(32'hbadb53b0),
	.w4(32'h39f7ba24),
	.w5(32'hba8ffb9f),
	.w6(32'hbb2a2ff1),
	.w7(32'hb9a74f1a),
	.w8(32'hbad8a7a6),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94e2c1),
	.w1(32'hbaf70c07),
	.w2(32'hbbb1586a),
	.w3(32'hbb4a43ce),
	.w4(32'h3a857796),
	.w5(32'hba032da1),
	.w6(32'hbb32b092),
	.w7(32'h3a83082c),
	.w8(32'hb9f786c2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e238b),
	.w1(32'hbaabcbb2),
	.w2(32'hbbd7485a),
	.w3(32'hbb680f0b),
	.w4(32'hba91abc6),
	.w5(32'hbbd6bcf1),
	.w6(32'hbac4f079),
	.w7(32'hbadb0a28),
	.w8(32'hbc0de426),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95b95c),
	.w1(32'h3a104144),
	.w2(32'hbb68ac8e),
	.w3(32'hbb85298a),
	.w4(32'h3acc2335),
	.w5(32'hbaf40b05),
	.w6(32'hbb6c1787),
	.w7(32'h3b161179),
	.w8(32'hbb24d21e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1407a),
	.w1(32'hbaf6a28f),
	.w2(32'hbb8a5b28),
	.w3(32'hbb3c912e),
	.w4(32'h3abbbefa),
	.w5(32'hba8267f9),
	.w6(32'hba9853b6),
	.w7(32'h3aa07042),
	.w8(32'hbb1e4e13),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba58b26),
	.w1(32'hbac621b8),
	.w2(32'hbb9d14de),
	.w3(32'hbb66c770),
	.w4(32'hb90cee73),
	.w5(32'hbbacf7d5),
	.w6(32'hbb246499),
	.w7(32'hb92c0d82),
	.w8(32'hbbaa1668),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc28736),
	.w1(32'hb93caab8),
	.w2(32'hb9b79b7f),
	.w3(32'hbb777699),
	.w4(32'h3a8f7162),
	.w5(32'h3a4fc0dc),
	.w6(32'hbb7acd8d),
	.w7(32'h3ac48c27),
	.w8(32'hb9bc52d8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb664471),
	.w1(32'hbaa97ccb),
	.w2(32'hbbb1b1f9),
	.w3(32'hbb13f695),
	.w4(32'hb955702a),
	.w5(32'hbb749896),
	.w6(32'hba9b3bef),
	.w7(32'hb9eb057d),
	.w8(32'hbbb23037),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefd1c3),
	.w1(32'h389525be),
	.w2(32'hbab93d50),
	.w3(32'hba7bd1f1),
	.w4(32'h3a3c953c),
	.w5(32'hba892239),
	.w6(32'hba87a4c9),
	.w7(32'h3a3d6240),
	.w8(32'hba50efd5),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be49c),
	.w1(32'h3bdcb908),
	.w2(32'hb7d37cda),
	.w3(32'hbc0ce882),
	.w4(32'h3b86bd2a),
	.w5(32'hb8898b1d),
	.w6(32'hbbf7e93e),
	.w7(32'h3baa746e),
	.w8(32'hbb14df9a),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1c72f),
	.w1(32'h39c8c0be),
	.w2(32'h3a958693),
	.w3(32'hbb84c436),
	.w4(32'h3a285ff7),
	.w5(32'h3a5aebd4),
	.w6(32'hbb8e5109),
	.w7(32'h3a26be3d),
	.w8(32'hba8d335e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3703959c),
	.w1(32'hb7655c31),
	.w2(32'hb825428d),
	.w3(32'hb88cc494),
	.w4(32'hb8d68274),
	.w5(32'hb9127dbb),
	.w6(32'hb8317534),
	.w7(32'hb8b6ad9a),
	.w8(32'hb8a2bf50),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3851bfb7),
	.w1(32'h38234363),
	.w2(32'h3809b42f),
	.w3(32'h3731c578),
	.w4(32'hb6adecaa),
	.w5(32'h37c807a1),
	.w6(32'h377c1cfd),
	.w7(32'h376dbff5),
	.w8(32'h3892ebd8),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb277053),
	.w1(32'hba0e69c6),
	.w2(32'hbaf1a791),
	.w3(32'hbb3b182c),
	.w4(32'h3a56887f),
	.w5(32'h3a29db23),
	.w6(32'hbad18252),
	.w7(32'h3a39b66e),
	.w8(32'hb9a90499),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc072af3),
	.w1(32'hb9a8db4f),
	.w2(32'hbb269aca),
	.w3(32'hbb89f2b4),
	.w4(32'h3b1740fc),
	.w5(32'hba9b69a5),
	.w6(32'hbb805f86),
	.w7(32'h3b343687),
	.w8(32'hbb5b3f80),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc130d2f),
	.w1(32'hbb2a4f45),
	.w2(32'hbbf59b7f),
	.w3(32'hbc1e7ea8),
	.w4(32'hbb0b95c0),
	.w5(32'hbbf99f52),
	.w6(32'hbbfa2495),
	.w7(32'hbb07c900),
	.w8(32'hbba19774),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ffa655),
	.w1(32'h379777d7),
	.w2(32'hb7080d3b),
	.w3(32'h381ebc64),
	.w4(32'h37abf566),
	.w5(32'h3780d442),
	.w6(32'h3830a3d2),
	.w7(32'h37ad9902),
	.w8(32'h37cf697c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb31df0),
	.w1(32'hbaf17c0d),
	.w2(32'hbc03a919),
	.w3(32'hbb908ad4),
	.w4(32'hbab4c200),
	.w5(32'hbbec1b94),
	.w6(32'hbb6892e5),
	.w7(32'hb9874b9e),
	.w8(32'hbbc80d7c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d231c),
	.w1(32'hba763b99),
	.w2(32'hbb8e4737),
	.w3(32'hbb02138a),
	.w4(32'h3a2f54fe),
	.w5(32'hbb8496e1),
	.w6(32'hbb0b3e8c),
	.w7(32'h3a932774),
	.w8(32'hbb8af54d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25fc18),
	.w1(32'hbb52d79d),
	.w2(32'hbc15c70a),
	.w3(32'hba9f86c3),
	.w4(32'hbaf6e6a5),
	.w5(32'hbbac3326),
	.w6(32'h3b539b02),
	.w7(32'h3ab45870),
	.w8(32'hbb91536d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb003102),
	.w1(32'h3b2f60ca),
	.w2(32'hbbc43316),
	.w3(32'hbb1c3c19),
	.w4(32'h3b38c65d),
	.w5(32'hbb89ea84),
	.w6(32'hbb57981c),
	.w7(32'h3ba50aa0),
	.w8(32'hbadc91e2),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ffa30),
	.w1(32'h3a06dcfe),
	.w2(32'hb87a0be3),
	.w3(32'hbb1401cb),
	.w4(32'h3a0bbe3a),
	.w5(32'h39acb47a),
	.w6(32'hbb80ac19),
	.w7(32'hba0731cf),
	.w8(32'hbb04c40f),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1731ae),
	.w1(32'h39dd4638),
	.w2(32'h3a0c8921),
	.w3(32'h39a00ebd),
	.w4(32'h39a8de35),
	.w5(32'h3a2f29f1),
	.w6(32'h39aa0c9c),
	.w7(32'h3a0e5e87),
	.w8(32'h3a20159c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2a0c),
	.w1(32'h3b1fd090),
	.w2(32'h3a3f480d),
	.w3(32'hbb2e61e7),
	.w4(32'h3b61870d),
	.w5(32'h3ab9086c),
	.w6(32'hbb95db6f),
	.w7(32'h3b36feda),
	.w8(32'hb965e2a7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1330d3),
	.w1(32'h3b3a0150),
	.w2(32'h3a90b37f),
	.w3(32'hbbc69961),
	.w4(32'h3bba0414),
	.w5(32'h3b9fece2),
	.w6(32'hbc04e097),
	.w7(32'h3ae5bf89),
	.w8(32'hbb7db68b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5da3ae),
	.w1(32'h3b509530),
	.w2(32'h3a79ae1a),
	.w3(32'hbb43d26e),
	.w4(32'h3b8f5419),
	.w5(32'h3b15b96b),
	.w6(32'hbbb6605a),
	.w7(32'h3b53802c),
	.w8(32'h3a602845),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cada8),
	.w1(32'hba2be2f9),
	.w2(32'hba8229fa),
	.w3(32'hba8ae1c5),
	.w4(32'hbac60bdb),
	.w5(32'hbaaebdb9),
	.w6(32'hb65978f6),
	.w7(32'hba1d70e6),
	.w8(32'hbad501df),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7faf2),
	.w1(32'hb9f1d8db),
	.w2(32'hba116720),
	.w3(32'hb98a1030),
	.w4(32'hb9a97d05),
	.w5(32'hb953ec74),
	.w6(32'hba035c1f),
	.w7(32'hba1bd390),
	.w8(32'hba216c25),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccccfb),
	.w1(32'hbb64d4dc),
	.w2(32'hbbb59284),
	.w3(32'hbb64f792),
	.w4(32'hbae33e4e),
	.w5(32'hbb6e2599),
	.w6(32'hbb85377b),
	.w7(32'hbaa9b47d),
	.w8(32'hbb8b09e4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d0606),
	.w1(32'hb79fbcf9),
	.w2(32'hba39862e),
	.w3(32'h39241aa9),
	.w4(32'h377414a1),
	.w5(32'hb9a47480),
	.w6(32'h3a7735f1),
	.w7(32'h3a17c932),
	.w8(32'hb90e2a02),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb309ec4),
	.w1(32'h3b04dc86),
	.w2(32'hb9c7b336),
	.w3(32'hba94f4ae),
	.w4(32'h3acd5e0d),
	.w5(32'hba9f82d7),
	.w6(32'hbaeb4e4c),
	.w7(32'h3addbf64),
	.w8(32'hb9bbd276),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386df43d),
	.w1(32'h39d8cf86),
	.w2(32'h39ce90c5),
	.w3(32'hb8e209ad),
	.w4(32'h394e8767),
	.w5(32'h39bc4cd8),
	.w6(32'hb9f30355),
	.w7(32'hb91e839b),
	.w8(32'h391797d2),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb955578),
	.w1(32'h3a1b49f4),
	.w2(32'hba17ddf1),
	.w3(32'hbbb9421d),
	.w4(32'hbaaa699a),
	.w5(32'hbabc6475),
	.w6(32'hbbd5c23f),
	.w7(32'hba970815),
	.w8(32'hba803538),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f20c0a),
	.w1(32'hb748175e),
	.w2(32'h387c4a61),
	.w3(32'h38d10f88),
	.w4(32'h36b653d2),
	.w5(32'h37ed592e),
	.w6(32'h3934203c),
	.w7(32'h38ba2bf9),
	.w8(32'h385d9f1b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83c0cf5),
	.w1(32'h39ae466d),
	.w2(32'h39d746be),
	.w3(32'hb7cd22cc),
	.w4(32'h38f77928),
	.w5(32'h39bcfb63),
	.w6(32'hb8efc23f),
	.w7(32'h380f3e3c),
	.w8(32'hb6daf54c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83281a),
	.w1(32'hba85897e),
	.w2(32'hbb6b31d6),
	.w3(32'hbb0aa0c6),
	.w4(32'h3ad27888),
	.w5(32'hbad51a72),
	.w6(32'hbb0e8e75),
	.w7(32'h3a8f6cc3),
	.w8(32'hbb4528fe),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39a332),
	.w1(32'hb9ee0408),
	.w2(32'hbbf8fd91),
	.w3(32'hbbf9212f),
	.w4(32'hbb334bb3),
	.w5(32'hbc46ad0c),
	.w6(32'hbbadcc85),
	.w7(32'h3acd80e9),
	.w8(32'hbc35ade2),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb425468),
	.w1(32'h3b1ded35),
	.w2(32'h3ad4526b),
	.w3(32'hbb54a2a3),
	.w4(32'h3af0d5d6),
	.w5(32'h3acdd0e0),
	.w6(32'hbbb4f977),
	.w7(32'h3a66eb8a),
	.w8(32'h386f316a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb412737),
	.w1(32'h3ac75ce8),
	.w2(32'hbbc0f1a6),
	.w3(32'hbac040d9),
	.w4(32'h3b4340bb),
	.w5(32'hbb99c1d3),
	.w6(32'hba8986a9),
	.w7(32'h3b6c4c76),
	.w8(32'hbb786bc8),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76ecbdb),
	.w1(32'h3819e9ea),
	.w2(32'hbaa77c3d),
	.w3(32'hba50508d),
	.w4(32'hb6e2568b),
	.w5(32'hb92d3f20),
	.w6(32'hb9949b7e),
	.w7(32'h3909bc43),
	.w8(32'hb9e1b2bb),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc437af8),
	.w1(32'h3818f429),
	.w2(32'hbc3516a5),
	.w3(32'hbc1cf48f),
	.w4(32'h3b2145fd),
	.w5(32'hbc04c228),
	.w6(32'hbc1636e0),
	.w7(32'hba9e9bc6),
	.w8(32'hbc0dd8c3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe80ba2),
	.w1(32'hba20d9fd),
	.w2(32'hbb9ad93a),
	.w3(32'hbba9f03d),
	.w4(32'h3ae3cb0d),
	.w5(32'hba976490),
	.w6(32'hbbc30d97),
	.w7(32'h3afb2c84),
	.w8(32'hbb1937f0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f68a8),
	.w1(32'hba4d89b6),
	.w2(32'hbbf7c350),
	.w3(32'hbb29d469),
	.w4(32'h3a067a0f),
	.w5(32'hbc075fd6),
	.w6(32'hbad1eb2a),
	.w7(32'h3a50deeb),
	.w8(32'hbbd8e282),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd8a66),
	.w1(32'hb9d3e474),
	.w2(32'h384baa85),
	.w3(32'hba0819de),
	.w4(32'hb99f858b),
	.w5(32'h3784c207),
	.w6(32'hb99c2cfc),
	.w7(32'hb8b93ef4),
	.w8(32'h3949fc2f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf13c4d),
	.w1(32'hba3dc4f5),
	.w2(32'hbb96e364),
	.w3(32'hba9a6cad),
	.w4(32'hb9fafa64),
	.w5(32'hbb2ff081),
	.w6(32'h38c1480e),
	.w7(32'h3abb0368),
	.w8(32'hbb1a0432),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d0b1f),
	.w1(32'h382fdeee),
	.w2(32'h382b9b44),
	.w3(32'h391c56bb),
	.w4(32'h34ee05ba),
	.w5(32'h36f760b9),
	.w6(32'h393d51ca),
	.w7(32'h37b6bdb3),
	.w8(32'h38877273),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11a43e),
	.w1(32'hba345b7a),
	.w2(32'hbb612141),
	.w3(32'hb99774d1),
	.w4(32'hb98dc248),
	.w5(32'hbabef9ca),
	.w6(32'hb99a81f6),
	.w7(32'hb6bd77b2),
	.w8(32'hbad9125b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa83908),
	.w1(32'h3a0a841e),
	.w2(32'hba8cd8ee),
	.w3(32'hbab0569a),
	.w4(32'h39749fb7),
	.w5(32'hba03c86e),
	.w6(32'hbac876c4),
	.w7(32'h363c911b),
	.w8(32'hba68b974),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba653a8),
	.w1(32'hb92cd00d),
	.w2(32'hbba8bd32),
	.w3(32'hbb9fdc48),
	.w4(32'h3a534e52),
	.w5(32'hbadc76c7),
	.w6(32'hbba773de),
	.w7(32'hb9e07431),
	.w8(32'hbb8dfaec),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bfa267),
	.w1(32'h378fe006),
	.w2(32'h374170cb),
	.w3(32'h388fac64),
	.w4(32'hb5ef1e63),
	.w5(32'hb669612a),
	.w6(32'h38aba2f2),
	.w7(32'h37dde7b3),
	.w8(32'h38248d2c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38034df7),
	.w1(32'h38d7281d),
	.w2(32'hb7eaf0b0),
	.w3(32'hb81af0dc),
	.w4(32'h37835031),
	.w5(32'h37a80b8f),
	.w6(32'hb90a017c),
	.w7(32'h38ca26a8),
	.w8(32'h390967e8),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53df1c),
	.w1(32'h39c10f59),
	.w2(32'hb7d4c86b),
	.w3(32'hbb05d381),
	.w4(32'h3aa5d0da),
	.w5(32'h3a7434a8),
	.w6(32'hbb1b8630),
	.w7(32'h3a70c463),
	.w8(32'h39d21809),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae23c5),
	.w1(32'h3a7e629b),
	.w2(32'hbb070329),
	.w3(32'hbbacef6b),
	.w4(32'h3a74c5d6),
	.w5(32'hb8b57fec),
	.w6(32'hbb98c6ed),
	.w7(32'hb9aca07b),
	.w8(32'hbae597b5),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba986977),
	.w1(32'h3b07c3cf),
	.w2(32'hbaa56719),
	.w3(32'hbb122cf7),
	.w4(32'h39aa43c7),
	.w5(32'hbad39686),
	.w6(32'h3a81ed90),
	.w7(32'h3b73473a),
	.w8(32'hbb0ca5fd),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba609a0c),
	.w1(32'h395b21f7),
	.w2(32'hba1b2711),
	.w3(32'hba9c99cd),
	.w4(32'hb7ab48c1),
	.w5(32'hb9ee4413),
	.w6(32'hbab7b661),
	.w7(32'h38e0840c),
	.w8(32'hba964d4c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f6eee),
	.w1(32'hbc1087a2),
	.w2(32'hbcb3f140),
	.w3(32'hbc5eb684),
	.w4(32'hbc0fcb06),
	.w5(32'hbcab943f),
	.w6(32'hbb9c8665),
	.w7(32'hbb859351),
	.w8(32'hbc48c731),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83a90a),
	.w1(32'hba8cc060),
	.w2(32'hbbd3c97e),
	.w3(32'hbc506ebb),
	.w4(32'h3b36e1c5),
	.w5(32'h3b208eb6),
	.w6(32'hbc3f0de1),
	.w7(32'h3b8f2304),
	.w8(32'hba8ebfef),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e5192),
	.w1(32'hb99ff5a5),
	.w2(32'hba5bf728),
	.w3(32'h391b2d30),
	.w4(32'hbaa261a8),
	.w5(32'hbab1d457),
	.w6(32'h3a4c4f55),
	.w7(32'hba132f15),
	.w8(32'hbac1765a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384073fe),
	.w1(32'hb7c7eba8),
	.w2(32'hb80e2365),
	.w3(32'h38292622),
	.w4(32'hb858f106),
	.w5(32'hb7bc75d3),
	.w6(32'h381a6715),
	.w7(32'h37602782),
	.w8(32'hb76933bc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ff51bb),
	.w1(32'h370cabba),
	.w2(32'h38e5441e),
	.w3(32'h3933d569),
	.w4(32'h38c8ec18),
	.w5(32'h38dbfacd),
	.w6(32'h39b66e8b),
	.w7(32'h38c9123e),
	.w8(32'h38fd61dc),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914d9eb),
	.w1(32'h381c2bf1),
	.w2(32'h38496e72),
	.w3(32'h38f267a9),
	.w4(32'h371fbe31),
	.w5(32'h37ceb300),
	.w6(32'h39175112),
	.w7(32'h38138612),
	.w8(32'h387eba45),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a496d43),
	.w1(32'hba31da24),
	.w2(32'hbb335137),
	.w3(32'h3a2dae14),
	.w4(32'hbad2bad2),
	.w5(32'hbb6503bc),
	.w6(32'h3a3e6aa9),
	.w7(32'hba9ac284),
	.w8(32'hbb6cd217),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1a4b6),
	.w1(32'hb90a1849),
	.w2(32'hbaacc9dc),
	.w3(32'hbb900a42),
	.w4(32'h39a7067a),
	.w5(32'hbb41c36b),
	.w6(32'hbb9c1942),
	.w7(32'hb9f1c8fa),
	.w8(32'hbbcd62a1),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1db3da),
	.w1(32'hbb4cae00),
	.w2(32'hbc0e893c),
	.w3(32'hbbfec10c),
	.w4(32'hba01b04e),
	.w5(32'hbbbee7f2),
	.w6(32'hbbdfc414),
	.w7(32'h3ad68bd2),
	.w8(32'hbb27ef79),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc51d7),
	.w1(32'h3a6d2902),
	.w2(32'hb7a85bc4),
	.w3(32'hbad037b0),
	.w4(32'h39dc4bd5),
	.w5(32'h3a339f91),
	.w6(32'hbb19f95e),
	.w7(32'hb93a1211),
	.w8(32'hba31545c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba25091),
	.w1(32'hbb275f7c),
	.w2(32'hbbf79a63),
	.w3(32'hbb051fbb),
	.w4(32'h389d11c7),
	.w5(32'hbbf04e51),
	.w6(32'hbb2c8fbf),
	.w7(32'h39c05a0b),
	.w8(32'hbbd0de23),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33fb52),
	.w1(32'hb9a11ef9),
	.w2(32'hba837e4f),
	.w3(32'hb9a63a9c),
	.w4(32'h3a788be8),
	.w5(32'h387ea803),
	.w6(32'h3a04320a),
	.w7(32'h39fd5e9a),
	.w8(32'hba91b4fa),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73544d),
	.w1(32'hba0e453d),
	.w2(32'h39df0159),
	.w3(32'h3ab12acb),
	.w4(32'hba2056a3),
	.w5(32'h3a5c7094),
	.w6(32'h393d0419),
	.w7(32'h3a39c5fd),
	.w8(32'h39895acc),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa611c0),
	.w1(32'hbaf28844),
	.w2(32'hba8575bc),
	.w3(32'hbb1dd0df),
	.w4(32'hbac734b5),
	.w5(32'hb9a0c96d),
	.w6(32'hba0ba740),
	.w7(32'hb9802847),
	.w8(32'h390a7225),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30163c),
	.w1(32'hb8d025c7),
	.w2(32'hb996178d),
	.w3(32'h39b46e6b),
	.w4(32'hb9f5a239),
	.w5(32'h3a065090),
	.w6(32'h39d8ab74),
	.w7(32'h3981a7e4),
	.w8(32'h39d6c28e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2a8ec),
	.w1(32'h3ac0a7c0),
	.w2(32'h39f236ed),
	.w3(32'hbb8f4e7c),
	.w4(32'hb8e595df),
	.w5(32'hbb009d01),
	.w6(32'hbb6adb86),
	.w7(32'hb9efb5fc),
	.w8(32'hbae34bbe),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a3e9d),
	.w1(32'h3a68d4c8),
	.w2(32'hb963f247),
	.w3(32'hbc00f79a),
	.w4(32'h3bb44b49),
	.w5(32'h3bc775f9),
	.w6(32'hbc44d451),
	.w7(32'h3b70daf7),
	.w8(32'h3ab5bd81),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba735e9),
	.w1(32'hb86b1092),
	.w2(32'hbb83586a),
	.w3(32'hbb43339e),
	.w4(32'h3aa56530),
	.w5(32'hbaf8ca77),
	.w6(32'hbb6ccfd2),
	.w7(32'h39b50499),
	.w8(32'hbb50c8b6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e7041),
	.w1(32'h3a03f210),
	.w2(32'h3a862831),
	.w3(32'hbac676ab),
	.w4(32'hba6b2fe1),
	.w5(32'hb9d258e8),
	.w6(32'hba934439),
	.w7(32'hbb1c5bbc),
	.w8(32'hba8d0ae0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cf25c),
	.w1(32'h3aab4bba),
	.w2(32'hbba3f3cb),
	.w3(32'hbba3f310),
	.w4(32'h3b729190),
	.w5(32'hba84c72f),
	.w6(32'hbbc16cc7),
	.w7(32'h3b3121f4),
	.w8(32'hbb4d1d5d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb339dc6),
	.w1(32'hbad20c22),
	.w2(32'hbb572804),
	.w3(32'hbb0c9de8),
	.w4(32'hbab20980),
	.w5(32'hbb8c17c5),
	.w6(32'hbaf3659d),
	.w7(32'hba596900),
	.w8(32'hbb4c069c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69c4c8),
	.w1(32'h3ae19853),
	.w2(32'hbb80cd92),
	.w3(32'hbc4461b2),
	.w4(32'h3b9d182c),
	.w5(32'hbae50acc),
	.w6(32'hbc49b6c8),
	.w7(32'h3b99385f),
	.w8(32'hbb0a2e96),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7703a9),
	.w1(32'hba5a3f41),
	.w2(32'h3a190ee6),
	.w3(32'h3b74e1e5),
	.w4(32'hba8c9f10),
	.w5(32'hb8c43e42),
	.w6(32'h3baeb03d),
	.w7(32'hba9397a2),
	.w8(32'hba3c02b0),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25cc11),
	.w1(32'hb9410b99),
	.w2(32'h3a34cffe),
	.w3(32'hba578f3b),
	.w4(32'hba7b2b21),
	.w5(32'h39bc8f37),
	.w6(32'hba83a492),
	.w7(32'hb829b00f),
	.w8(32'hb9a3acb8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca81d0),
	.w1(32'h3b056936),
	.w2(32'hbade2e58),
	.w3(32'hbb7641d4),
	.w4(32'h3b53e883),
	.w5(32'hb8eeb34a),
	.w6(32'hbbb99a5b),
	.w7(32'h3b004c71),
	.w8(32'hbb0eb9db),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc188ee1),
	.w1(32'h3b2f7652),
	.w2(32'hbbb47f94),
	.w3(32'hbbb4cf99),
	.w4(32'h3aa15df1),
	.w5(32'hbc303488),
	.w6(32'hbb8bff62),
	.w7(32'h3b7dd3e1),
	.w8(32'hbb9d0e7f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1251be),
	.w1(32'h39c47cae),
	.w2(32'hbb591064),
	.w3(32'hbbb5ba3e),
	.w4(32'h3a366da5),
	.w5(32'hba1cb6b1),
	.w6(32'hbbaecaf7),
	.w7(32'h3af69540),
	.w8(32'hbb5499e9),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e59a2),
	.w1(32'hba28a9b7),
	.w2(32'hbb36f842),
	.w3(32'hbb16d6c7),
	.w4(32'hbb9fdfbd),
	.w5(32'hbb2a7a29),
	.w6(32'h3a9bf4ce),
	.w7(32'hbaf36e11),
	.w8(32'hbb44c0f9),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37bfef),
	.w1(32'hba817509),
	.w2(32'hbb127bea),
	.w3(32'hba25cef6),
	.w4(32'hba1c143a),
	.w5(32'hba107e90),
	.w6(32'h38ba6aa7),
	.w7(32'hba4f8f05),
	.w8(32'hba66cae5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb161394),
	.w1(32'hbb02b909),
	.w2(32'hb9954721),
	.w3(32'hbb18aa50),
	.w4(32'hbabca83a),
	.w5(32'h3a23bc76),
	.w6(32'hbb3357b6),
	.w7(32'hbac8634c),
	.w8(32'h3a237803),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4a89c),
	.w1(32'h3a872902),
	.w2(32'hbb906adb),
	.w3(32'h3b0ee3c7),
	.w4(32'hbbeb638b),
	.w5(32'hbc25ba50),
	.w6(32'h3b3827dd),
	.w7(32'hbb795fb3),
	.w8(32'hbc138d35),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fd554),
	.w1(32'hbbcd33b7),
	.w2(32'hbc1cd6d2),
	.w3(32'hbbe9cb13),
	.w4(32'hbbb85a55),
	.w5(32'hbc14f721),
	.w6(32'hbbf799cc),
	.w7(32'hbb8faf04),
	.w8(32'hbbe92857),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5eaa7),
	.w1(32'hbafe1947),
	.w2(32'hbbbfac15),
	.w3(32'hbaa31eed),
	.w4(32'hbb61b845),
	.w5(32'hbbcd612d),
	.w6(32'h3b493303),
	.w7(32'hba2c6f43),
	.w8(32'hbc02d6e6),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96a68c),
	.w1(32'h3bc920d4),
	.w2(32'h3b37057a),
	.w3(32'hbbabea1a),
	.w4(32'h3ba89fc9),
	.w5(32'h3b320ced),
	.w6(32'hbc09e585),
	.w7(32'h3b9c671a),
	.w8(32'h3a12a6cf),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc93e1),
	.w1(32'h3a0e1656),
	.w2(32'hbb75dca7),
	.w3(32'hbbb33934),
	.w4(32'h3b6fc459),
	.w5(32'h3a1d15ba),
	.w6(32'hbba4a6dd),
	.w7(32'h3bac949b),
	.w8(32'hb7e995be),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae148d4),
	.w1(32'hba640885),
	.w2(32'hb9a3d701),
	.w3(32'h3b078553),
	.w4(32'hbaef1925),
	.w5(32'hba4774f2),
	.w6(32'h3ad1db37),
	.w7(32'hbb00aa3f),
	.w8(32'hbb8a3978),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98a47f),
	.w1(32'h39a63ac5),
	.w2(32'hbabebd0b),
	.w3(32'hba5297cf),
	.w4(32'h37af94ea),
	.w5(32'h3a36f246),
	.w6(32'hbab54586),
	.w7(32'hb99e8cfe),
	.w8(32'h3ad45ebc),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f04ef7),
	.w1(32'hb966bc14),
	.w2(32'hb928d7f6),
	.w3(32'h37b8cfa9),
	.w4(32'hba489d30),
	.w5(32'h39e28e8c),
	.w6(32'hbaa82c77),
	.w7(32'hba9d9cb7),
	.w8(32'hba822f19),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44d4af),
	.w1(32'h3628c497),
	.w2(32'h3aa6c1c8),
	.w3(32'hba75109d),
	.w4(32'h3a6d4200),
	.w5(32'h3a39e29a),
	.w6(32'hbb0257fd),
	.w7(32'h3aa10d19),
	.w8(32'h3af090d9),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09636a),
	.w1(32'hbb2717c5),
	.w2(32'hbb72c2bd),
	.w3(32'h3ad3b95e),
	.w4(32'hbb7dd2a3),
	.w5(32'hbb912942),
	.w6(32'h39d2d119),
	.w7(32'hba880416),
	.w8(32'hbb5345c5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc215a1d),
	.w1(32'hbae3a55a),
	.w2(32'hbb906c01),
	.w3(32'hbbd4c68f),
	.w4(32'hbaf025d6),
	.w5(32'hbc081589),
	.w6(32'hbb5950b1),
	.w7(32'hba2258c4),
	.w8(32'hbbea0e53),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2e496),
	.w1(32'hbad27393),
	.w2(32'hbbb0e46f),
	.w3(32'hbba846dc),
	.w4(32'hb9233efe),
	.w5(32'hbada324f),
	.w6(32'hbbdf97a4),
	.w7(32'hba5d8ea9),
	.w8(32'hbb854e0e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cb301),
	.w1(32'hb8c6c46d),
	.w2(32'hba0a84e0),
	.w3(32'h39d22462),
	.w4(32'h388e6ba1),
	.w5(32'hba944b4f),
	.w6(32'h39900732),
	.w7(32'hba6da7e4),
	.w8(32'h39139570),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dfdb7),
	.w1(32'hb9f2953c),
	.w2(32'hbbee4b95),
	.w3(32'hba84e91d),
	.w4(32'hbb148580),
	.w5(32'hbb9d39a5),
	.w6(32'h3b01de0b),
	.w7(32'h3ad64509),
	.w8(32'hbc1e73da),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fc428),
	.w1(32'h3afaf410),
	.w2(32'hbaed24be),
	.w3(32'hbb388c6b),
	.w4(32'h3a67634b),
	.w5(32'hbb7d641d),
	.w6(32'hbb3c75db),
	.w7(32'h39d26dd9),
	.w8(32'hbb860483),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cab18f),
	.w1(32'hbabb72cf),
	.w2(32'hba334456),
	.w3(32'hb9d515b7),
	.w4(32'hba95049f),
	.w5(32'hba1a66cb),
	.w6(32'hbaa4f2ab),
	.w7(32'hba33ac98),
	.w8(32'hbb226cc5),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6da6f),
	.w1(32'hb97e1061),
	.w2(32'hbb042538),
	.w3(32'hba597308),
	.w4(32'hbae7b04c),
	.w5(32'hbb325e89),
	.w6(32'hba648b12),
	.w7(32'hbae50bf1),
	.w8(32'hbb87af61),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1fac1),
	.w1(32'h3a677e38),
	.w2(32'h3aaae894),
	.w3(32'hb9f44399),
	.w4(32'h3a21e6d7),
	.w5(32'h3a065ccc),
	.w6(32'hba67a2e9),
	.w7(32'h3a16d271),
	.w8(32'h381c744c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387e2997),
	.w1(32'hb920fdb5),
	.w2(32'hbad2ecfc),
	.w3(32'hb991c699),
	.w4(32'hb9f18cdd),
	.w5(32'hbb63d66f),
	.w6(32'h394a03f6),
	.w7(32'h3a03f247),
	.w8(32'hbb2b0629),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba595053),
	.w1(32'h3a81cc1b),
	.w2(32'h3a6d2a8b),
	.w3(32'hbb1305ae),
	.w4(32'h3af98a15),
	.w5(32'h3ad24057),
	.w6(32'hb749c59c),
	.w7(32'h3ae96fa9),
	.w8(32'h3a8696bd),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38037695),
	.w1(32'hbac0eeae),
	.w2(32'hbb1e707c),
	.w3(32'h3a30404d),
	.w4(32'hba1c5b26),
	.w5(32'hbb5b75b0),
	.w6(32'h3a9598d1),
	.w7(32'h39b9eed1),
	.w8(32'hba1e793d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb787798),
	.w1(32'h3b47a854),
	.w2(32'h3aaa315e),
	.w3(32'hbb8183c0),
	.w4(32'h3ad2dd00),
	.w5(32'h3af6dc1c),
	.w6(32'hbbbd2931),
	.w7(32'h3a5e9319),
	.w8(32'hb7f96008),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb997aeb),
	.w1(32'hba398b30),
	.w2(32'hbc31cc34),
	.w3(32'hbb815091),
	.w4(32'hbb52a19e),
	.w5(32'hbbe1cc72),
	.w6(32'hbb53a2cc),
	.w7(32'hbb542d0b),
	.w8(32'hbc1306fe),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ec527),
	.w1(32'hba7605e8),
	.w2(32'hbba17ced),
	.w3(32'hbb192cf3),
	.w4(32'h39b990f1),
	.w5(32'hbb1705be),
	.w6(32'hbb3faf6c),
	.w7(32'h3a870ef7),
	.w8(32'hbb452063),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d96f9),
	.w1(32'hbb891298),
	.w2(32'hbc2b29ab),
	.w3(32'hbb9885c3),
	.w4(32'hbb5a8841),
	.w5(32'hbc054d3c),
	.w6(32'hbb6b3065),
	.w7(32'hbb6a06ab),
	.w8(32'hbc03eb26),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23a070),
	.w1(32'h3ab8a038),
	.w2(32'h3a80d5b3),
	.w3(32'hbac79827),
	.w4(32'h3a122dc3),
	.w5(32'hb961b7eb),
	.w6(32'h398a13bb),
	.w7(32'h395df9a5),
	.w8(32'hbace6c14),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396bd1a2),
	.w1(32'h39e3cf71),
	.w2(32'hba23850c),
	.w3(32'h38a5d9c1),
	.w4(32'h39c0a80a),
	.w5(32'hba583078),
	.w6(32'hba8997cc),
	.w7(32'h3a0938f1),
	.w8(32'hba045453),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0bee9),
	.w1(32'hbad71396),
	.w2(32'hba78b47d),
	.w3(32'hba34f3b8),
	.w4(32'hb9846da6),
	.w5(32'hbb051202),
	.w6(32'hb91e4d81),
	.w7(32'h3a877f1a),
	.w8(32'h3a916f5a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ae551),
	.w1(32'h3a828383),
	.w2(32'h3a118208),
	.w3(32'h3aa2f04a),
	.w4(32'hb9c313be),
	.w5(32'hb954a016),
	.w6(32'h3aea9fdb),
	.w7(32'hb9717a5c),
	.w8(32'hb9a5b867),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb510f8),
	.w1(32'hbb20c665),
	.w2(32'hbbd35b2d),
	.w3(32'hbb158e77),
	.w4(32'hb8c60e18),
	.w5(32'hbb18c784),
	.w6(32'hbb0ebaa2),
	.w7(32'hbb4f0acd),
	.w8(32'hbbaf3a06),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d0231),
	.w1(32'hb9890447),
	.w2(32'hba89909f),
	.w3(32'hb9dd341f),
	.w4(32'hba108bd7),
	.w5(32'hba6908d6),
	.w6(32'hb97551fe),
	.w7(32'hb9f90c9d),
	.w8(32'hba249dc0),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb525c1b),
	.w1(32'h3b78038f),
	.w2(32'h3b81bcaf),
	.w3(32'hbb27310b),
	.w4(32'h3b466df9),
	.w5(32'h3b959ec7),
	.w6(32'hbb6f8b36),
	.w7(32'h3aabccce),
	.w8(32'h3af726bc),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8704ac),
	.w1(32'h3a9e66f5),
	.w2(32'h3a96449f),
	.w3(32'hb9dbe82e),
	.w4(32'h3b284e7d),
	.w5(32'h3b1cdcf9),
	.w6(32'h39d853fc),
	.w7(32'h3b18bb9f),
	.w8(32'h3a8c6b9a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b7b1a),
	.w1(32'hb9b827e3),
	.w2(32'h39a74ac2),
	.w3(32'h3a2dcf2a),
	.w4(32'h3aa6622c),
	.w5(32'h3b2a252e),
	.w6(32'h3ad552db),
	.w7(32'h3a8b05d4),
	.w8(32'h39dfd28e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaab0c5),
	.w1(32'h39e45de0),
	.w2(32'hba0d7267),
	.w3(32'hba6e8dea),
	.w4(32'h3a0e5c41),
	.w5(32'hba176b1b),
	.w6(32'hba8fac16),
	.w7(32'hbab3ab29),
	.w8(32'hbb042cd3),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5e909),
	.w1(32'hba3dbcc8),
	.w2(32'hbab418d3),
	.w3(32'h3a1a6f59),
	.w4(32'h39807578),
	.w5(32'hba370cc1),
	.w6(32'hb9b61adc),
	.w7(32'h3abaa7eb),
	.w8(32'h3aa8c528),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad4262),
	.w1(32'hbbc058ce),
	.w2(32'hbc4e81a8),
	.w3(32'hbb5d11aa),
	.w4(32'hbb30ff84),
	.w5(32'hbad03e22),
	.w6(32'hbb812198),
	.w7(32'hbb3ce129),
	.w8(32'hbbec2fbd),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb7614),
	.w1(32'hbb4e87e9),
	.w2(32'hbb0575fb),
	.w3(32'hbb126e4c),
	.w4(32'hbb8c2524),
	.w5(32'hbb532def),
	.w6(32'hbab8c803),
	.w7(32'hbb80220e),
	.w8(32'hbb6e593f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75b58b),
	.w1(32'h3bb4fed2),
	.w2(32'h3bb5e0d9),
	.w3(32'hbb5d3224),
	.w4(32'h3b91958e),
	.w5(32'h3bc4eb2b),
	.w6(32'hbc358ad4),
	.w7(32'h3a81478c),
	.w8(32'h3ba053d0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule