module layer_8_featuremap_225(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98cee2),
	.w1(32'h3c927889),
	.w2(32'h3cbbfb47),
	.w3(32'hbb08974b),
	.w4(32'h3ca34189),
	.w5(32'h3c032f86),
	.w6(32'hbc85a38d),
	.w7(32'hbb721e0e),
	.w8(32'h3abb1ac7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6fdaa2),
	.w1(32'h3b4ded66),
	.w2(32'hb8bbb932),
	.w3(32'h3b52bd10),
	.w4(32'h39ce4e3d),
	.w5(32'hbb28aeb9),
	.w6(32'h3a89e434),
	.w7(32'hbaa498ec),
	.w8(32'hbb05470b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ff7f1),
	.w1(32'h3c074d86),
	.w2(32'h3c44a1d2),
	.w3(32'h39b38143),
	.w4(32'hbb6c5426),
	.w5(32'hbc2bc6f9),
	.w6(32'h3aad9131),
	.w7(32'h3b99b093),
	.w8(32'hba3357bc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7d120),
	.w1(32'hb8caade5),
	.w2(32'h3aa32cb2),
	.w3(32'hbc352b7e),
	.w4(32'h3be805ab),
	.w5(32'h3ac5a97f),
	.w6(32'hbc072736),
	.w7(32'hbc4692ae),
	.w8(32'hbad43c87),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9382c),
	.w1(32'h3bbf231c),
	.w2(32'hba4d93ed),
	.w3(32'hbc0f10fa),
	.w4(32'h3ad51596),
	.w5(32'hbaffea7f),
	.w6(32'h3b66784a),
	.w7(32'h3b3f7b1f),
	.w8(32'h3b8fa214),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27cd7e),
	.w1(32'hbacf18b0),
	.w2(32'hbc462f9d),
	.w3(32'hbaa09beb),
	.w4(32'hbc328024),
	.w5(32'hbc6ce8c6),
	.w6(32'h3abe73b9),
	.w7(32'h3c027637),
	.w8(32'h3b94d8ed),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc528197),
	.w1(32'hbbd0e4fd),
	.w2(32'hbba77f67),
	.w3(32'hbbd65c75),
	.w4(32'hba6f9c72),
	.w5(32'h391b8a57),
	.w6(32'hbbcd98a8),
	.w7(32'hbc01dcca),
	.w8(32'hbb7ff693),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d2266),
	.w1(32'h3ce5f0f7),
	.w2(32'h3d404a74),
	.w3(32'hbb593339),
	.w4(32'hbb84c110),
	.w5(32'hbcdd86c2),
	.w6(32'h3cf409f8),
	.w7(32'h3c5a3560),
	.w8(32'h3bbcc848),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b8469),
	.w1(32'h3b3bc639),
	.w2(32'hba66819c),
	.w3(32'hbca8caca),
	.w4(32'h3bce9448),
	.w5(32'h3afa813e),
	.w6(32'h3a896e2b),
	.w7(32'hba1f82d4),
	.w8(32'h39cb543c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f72a6),
	.w1(32'hbc36c182),
	.w2(32'hbcb05f05),
	.w3(32'h3a9aacb0),
	.w4(32'hbbf86868),
	.w5(32'hbb855b29),
	.w6(32'hbaa7baf6),
	.w7(32'h3c3e4ed4),
	.w8(32'h3c2bd38a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc280c49),
	.w1(32'h3b817b10),
	.w2(32'hbbe4c563),
	.w3(32'h3bacb146),
	.w4(32'h3c4e770b),
	.w5(32'h3c0ebb1c),
	.w6(32'hbc89be6d),
	.w7(32'hbbe812ae),
	.w8(32'hbc56b036),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8961c),
	.w1(32'hbb0deed2),
	.w2(32'hbb9d4328),
	.w3(32'hbb905633),
	.w4(32'hbb318ec3),
	.w5(32'hbb14e184),
	.w6(32'hbaa87fde),
	.w7(32'hbb330ef7),
	.w8(32'hbb63487d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadec10c),
	.w1(32'hbc9184dc),
	.w2(32'hbc581628),
	.w3(32'hbaf66818),
	.w4(32'h3a59c20d),
	.w5(32'h3abbd13e),
	.w6(32'hbc9b3e1a),
	.w7(32'hbace9078),
	.w8(32'h3b896ea8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae000f6),
	.w1(32'h3c056289),
	.w2(32'hbb885771),
	.w3(32'h3c01d929),
	.w4(32'hbb6c5fdf),
	.w5(32'hbccfd064),
	.w6(32'h3bf1bc92),
	.w7(32'hba63da22),
	.w8(32'h3af31d63),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ba747),
	.w1(32'hbb222cf5),
	.w2(32'h3b5fc7d0),
	.w3(32'hbca8a1ee),
	.w4(32'h3b5eb095),
	.w5(32'h3bc5889f),
	.w6(32'h393ee2e4),
	.w7(32'h3a658c5d),
	.w8(32'h3b78633f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0f55c),
	.w1(32'h3a6eb38d),
	.w2(32'h3b374a06),
	.w3(32'h3ba0f5b7),
	.w4(32'h3cbe47eb),
	.w5(32'h3d00f5e3),
	.w6(32'hbc495fec),
	.w7(32'hbc1bcd34),
	.w8(32'hbaad3a3e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e15f3),
	.w1(32'h3bb2bdec),
	.w2(32'h3caae476),
	.w3(32'h3c6fc957),
	.w4(32'h3caed2e3),
	.w5(32'h3cc764ed),
	.w6(32'hbba7b399),
	.w7(32'h3c4574d8),
	.w8(32'h3c615bd1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfb6d25),
	.w1(32'h3a1355ca),
	.w2(32'h3bc1aec2),
	.w3(32'h3c561d8e),
	.w4(32'h3c20443c),
	.w5(32'h3c940897),
	.w6(32'hbccfb498),
	.w7(32'hbcf61d8b),
	.w8(32'hbc00b735),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb7996),
	.w1(32'h3bc2688d),
	.w2(32'h3c6bc496),
	.w3(32'h3c395559),
	.w4(32'hbbf92c4a),
	.w5(32'hbc811828),
	.w6(32'h3ae207f7),
	.w7(32'h3a70107c),
	.w8(32'h3b88420a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca03899),
	.w1(32'hba25b64c),
	.w2(32'h3a37d76f),
	.w3(32'h3bea7037),
	.w4(32'h3bb1f1e4),
	.w5(32'h3b6f33b4),
	.w6(32'hbb83e02c),
	.w7(32'hbace3b97),
	.w8(32'hba7959f0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b991182),
	.w1(32'hbc81537b),
	.w2(32'hbcac345e),
	.w3(32'h3aa5e6a5),
	.w4(32'hbc128bf3),
	.w5(32'hbbdb550a),
	.w6(32'h3bc69aaf),
	.w7(32'h3c0577ba),
	.w8(32'hbbfa9142),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49fed9),
	.w1(32'hbc9900b3),
	.w2(32'hbcdcf183),
	.w3(32'hba2b869c),
	.w4(32'hb880c5cb),
	.w5(32'hbc272312),
	.w6(32'hbb06ab68),
	.w7(32'h3a9557a4),
	.w8(32'hbb32abcf),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b8411),
	.w1(32'hbc6ed721),
	.w2(32'hbc3f1fc7),
	.w3(32'h3bacc0f6),
	.w4(32'h3b95030b),
	.w5(32'h3b3fdfd0),
	.w6(32'hbbca6434),
	.w7(32'hbc0bbeaa),
	.w8(32'hbc1d4e7f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe793fc),
	.w1(32'hbc65118d),
	.w2(32'hbcb9294c),
	.w3(32'h3b8d2869),
	.w4(32'h3b46f0f5),
	.w5(32'h3a737ba0),
	.w6(32'hbb9f6354),
	.w7(32'h3bd2170b),
	.w8(32'h39b4a107),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65b529),
	.w1(32'hbb882d08),
	.w2(32'hb9f539e0),
	.w3(32'hbaf983cb),
	.w4(32'hba0c0865),
	.w5(32'hbb187fa0),
	.w6(32'hba93126d),
	.w7(32'h3b3cb3e9),
	.w8(32'h3b603dcf),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4757ee),
	.w1(32'h3c60f1f8),
	.w2(32'h3c45f9e5),
	.w3(32'h3a37a2e7),
	.w4(32'hbbd06be5),
	.w5(32'hbc2843d5),
	.w6(32'h3c54a449),
	.w7(32'h3c723594),
	.w8(32'h3c578cef),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d3c6d),
	.w1(32'h3c7300fb),
	.w2(32'h3cf235e3),
	.w3(32'hbc4d7cd4),
	.w4(32'h3ca7c103),
	.w5(32'h3b090591),
	.w6(32'h387f182f),
	.w7(32'hbc03618f),
	.w8(32'h3a11bbe9),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc0893d),
	.w1(32'h3aa8adda),
	.w2(32'h3b3d70f7),
	.w3(32'h3ac3c5eb),
	.w4(32'h3c042bff),
	.w5(32'h3b2ac859),
	.w6(32'hbcb10fc1),
	.w7(32'hbc2fe35e),
	.w8(32'hbadd2e58),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dea964),
	.w1(32'h3b95a31b),
	.w2(32'hbb721f46),
	.w3(32'hbaf8df31),
	.w4(32'h3a8b2eb8),
	.w5(32'h3b1be1b2),
	.w6(32'hbb8f4d17),
	.w7(32'hbba89fba),
	.w8(32'hbbcd96fb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb298f06),
	.w1(32'hba965ad5),
	.w2(32'hbb8db2a6),
	.w3(32'h3b60676b),
	.w4(32'h3bf1ea96),
	.w5(32'h3b4afbf3),
	.w6(32'h3a170005),
	.w7(32'hba335a0a),
	.w8(32'hbc473a6e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5dbc6b),
	.w1(32'h3c02e0e5),
	.w2(32'h3b01f347),
	.w3(32'hbb905a7e),
	.w4(32'h3ae2aa27),
	.w5(32'hbb1112dd),
	.w6(32'h3b046b81),
	.w7(32'h3b07e290),
	.w8(32'hbbab2b14),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa318c),
	.w1(32'hbb429224),
	.w2(32'hbc1bec09),
	.w3(32'hb9ba816c),
	.w4(32'hbbee6c0d),
	.w5(32'h3b80ce48),
	.w6(32'h3b0f1d37),
	.w7(32'hbac97f1e),
	.w8(32'hbbc0b62d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a48c1),
	.w1(32'h3bd9ff90),
	.w2(32'h3ccc88fa),
	.w3(32'h3bcdb2cb),
	.w4(32'hba28bd0b),
	.w5(32'h3b6d82ef),
	.w6(32'hbcab30c7),
	.w7(32'hbc0af0bc),
	.w8(32'h3b04139d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71d4f1),
	.w1(32'h3c176ca5),
	.w2(32'h3cd1cba3),
	.w3(32'hbaa452d0),
	.w4(32'h3bcf87cd),
	.w5(32'h3c6a4f0e),
	.w6(32'hbc35f294),
	.w7(32'hbb677749),
	.w8(32'h3aab9ff7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22689b),
	.w1(32'hbc063fbe),
	.w2(32'hbc2b970d),
	.w3(32'hbb818f1b),
	.w4(32'hbb87a8da),
	.w5(32'hba6cc856),
	.w6(32'hba7ebe5a),
	.w7(32'hbb7a1e02),
	.w8(32'hbb9e9393),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dcd51),
	.w1(32'h3c9893f2),
	.w2(32'h3c88431e),
	.w3(32'h3b2053d0),
	.w4(32'hbbbc6340),
	.w5(32'hbc8600fb),
	.w6(32'h3c2f2e2f),
	.w7(32'h3bee8821),
	.w8(32'h3c19e693),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c739aa3),
	.w1(32'hbb278d23),
	.w2(32'hbae806a9),
	.w3(32'hbbca9689),
	.w4(32'h3a41e474),
	.w5(32'hba31f082),
	.w6(32'hbab1d593),
	.w7(32'hba9b477b),
	.w8(32'h39da97d7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0dff1),
	.w1(32'hb8a5fdc5),
	.w2(32'h3bd56a8e),
	.w3(32'h3b2c8b2d),
	.w4(32'h3ac0b4f0),
	.w5(32'h3b7fe899),
	.w6(32'h3afc200d),
	.w7(32'h3bc7f8e9),
	.w8(32'h3c310eaf),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ffb1b),
	.w1(32'hbca7e230),
	.w2(32'hbd0b2673),
	.w3(32'h3c115f3d),
	.w4(32'hbab73b91),
	.w5(32'hb895a3dc),
	.w6(32'h3aca6303),
	.w7(32'hbc34d8fc),
	.w8(32'hbc269af0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc455558),
	.w1(32'hbb68c9c5),
	.w2(32'hbb7f70e3),
	.w3(32'hbac4e428),
	.w4(32'hbb31ca74),
	.w5(32'h3ba93f4a),
	.w6(32'hbb00a47c),
	.w7(32'h3bab7239),
	.w8(32'h3c384bea),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb682edd),
	.w1(32'h3aec7dc4),
	.w2(32'h3a767c18),
	.w3(32'hbb8e216b),
	.w4(32'h3a06f964),
	.w5(32'hba11815a),
	.w6(32'h3b21bda8),
	.w7(32'h3a4b341c),
	.w8(32'h39cd6680),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ae722),
	.w1(32'h39f18ac9),
	.w2(32'h3ab420fe),
	.w3(32'h3a395b5d),
	.w4(32'hbb4c9882),
	.w5(32'hbc29532a),
	.w6(32'hbb683e52),
	.w7(32'hb9925a23),
	.w8(32'hbb959fe3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9381c0),
	.w1(32'hbb5b4839),
	.w2(32'hbb0025a9),
	.w3(32'hbbf8c3c6),
	.w4(32'hbb568962),
	.w5(32'hbbe96036),
	.w6(32'hb79824ec),
	.w7(32'hbb4e9b6e),
	.w8(32'hbb31a853),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac4435),
	.w1(32'hbc405610),
	.w2(32'hbc7ba290),
	.w3(32'hbbd0192c),
	.w4(32'hbb0bfde0),
	.w5(32'h3c919921),
	.w6(32'hbceed737),
	.w7(32'hbd28d2d8),
	.w8(32'hbc987c68),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31eb1e),
	.w1(32'h3be38cfe),
	.w2(32'h39cd3237),
	.w3(32'h3c70c156),
	.w4(32'hbc54f63d),
	.w5(32'hbd1585e9),
	.w6(32'h3ca1a4f7),
	.w7(32'h3d4e830c),
	.w8(32'h3cf3b6ae),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4465fb),
	.w1(32'h3a5fbf2e),
	.w2(32'hbb35b1ae),
	.w3(32'hbccd8d61),
	.w4(32'h3be7e7c5),
	.w5(32'h3ac3fbef),
	.w6(32'hbb466e53),
	.w7(32'hbbd7400b),
	.w8(32'hbb889415),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0104d8),
	.w1(32'hbb4a0f8e),
	.w2(32'hbbe8b9a1),
	.w3(32'hbb806bd9),
	.w4(32'hbb852ef0),
	.w5(32'h3aff4aad),
	.w6(32'hbb4c8348),
	.w7(32'hbb85166c),
	.w8(32'hbb8dfdfd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2af44c),
	.w1(32'h3be22810),
	.w2(32'h3b944c0a),
	.w3(32'h3a36d7a4),
	.w4(32'hba06b140),
	.w5(32'hbbae07ad),
	.w6(32'h3c005577),
	.w7(32'h3baf8a97),
	.w8(32'h3c3905ab),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f6821),
	.w1(32'h3bc0d9f3),
	.w2(32'hbc1bc2b7),
	.w3(32'hbb5e22b3),
	.w4(32'hbc11452f),
	.w5(32'hbc5483de),
	.w6(32'h3b430700),
	.w7(32'h3bff124f),
	.w8(32'hbb23ae93),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2be8ae),
	.w1(32'h3bed04fd),
	.w2(32'h3c3fe879),
	.w3(32'hbb892b31),
	.w4(32'hbb655973),
	.w5(32'h3b76c53d),
	.w6(32'hbc31ef73),
	.w7(32'hbc2fceb5),
	.w8(32'hbc3accc6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e8b26),
	.w1(32'h3b22b5f2),
	.w2(32'h3a69ff74),
	.w3(32'hb994fd3a),
	.w4(32'hbab5c2f5),
	.w5(32'h389090e4),
	.w6(32'h3b15d2d2),
	.w7(32'h3a5adbf0),
	.w8(32'h3b3e5a2f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26e856),
	.w1(32'h3b140c5a),
	.w2(32'h3a54541e),
	.w3(32'h39f67825),
	.w4(32'hbaab3f46),
	.w5(32'hbbebca09),
	.w6(32'h3c225b55),
	.w7(32'h3c27faab),
	.w8(32'hb8938d2b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef2f56),
	.w1(32'hba1ed674),
	.w2(32'hbb9035f3),
	.w3(32'hbb940fb5),
	.w4(32'hbb7291e7),
	.w5(32'hbbbad7e5),
	.w6(32'hbb475781),
	.w7(32'hbbb507fb),
	.w8(32'hbb87b3ad),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98379d),
	.w1(32'hbba25bc6),
	.w2(32'hbc802632),
	.w3(32'hb99c3fa8),
	.w4(32'hbc9e82c1),
	.w5(32'hbcb1b56a),
	.w6(32'h3c045f9d),
	.w7(32'hbbd0ecaa),
	.w8(32'hbbf5b00b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2994dc),
	.w1(32'h3b0d73c1),
	.w2(32'h3c2ae172),
	.w3(32'hbb37d445),
	.w4(32'hbbef4c6e),
	.w5(32'hbbd2cc69),
	.w6(32'hbc236fa3),
	.w7(32'hbc29f18b),
	.w8(32'hbc5f75a4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf51c59),
	.w1(32'hbbb6c727),
	.w2(32'h3c80273b),
	.w3(32'h3b939b0f),
	.w4(32'h3c3cf396),
	.w5(32'h3cd47107),
	.w6(32'hbd11dfcc),
	.w7(32'hbd1ece69),
	.w8(32'hbc9c8a6b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db9de),
	.w1(32'hbc253c43),
	.w2(32'hba859011),
	.w3(32'h3cc46dac),
	.w4(32'hbb209bfb),
	.w5(32'hbb72ef84),
	.w6(32'hbbe97f2a),
	.w7(32'hbbc223da),
	.w8(32'hbbfa94c5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba845339),
	.w1(32'h3921452a),
	.w2(32'hbb31d91f),
	.w3(32'h3a1e12f7),
	.w4(32'h3b29b483),
	.w5(32'hbbca47ff),
	.w6(32'h3afb22b8),
	.w7(32'h3ad7d174),
	.w8(32'h3ab6f2eb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0981a6),
	.w1(32'hbb742e0a),
	.w2(32'h3ac1a122),
	.w3(32'hba34c386),
	.w4(32'hbb4a2420),
	.w5(32'h394fb6a0),
	.w6(32'hbb59a3db),
	.w7(32'hbaf62b82),
	.w8(32'h3b6c234b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab9c57),
	.w1(32'hbc3a53c1),
	.w2(32'hbce92674),
	.w3(32'h3bbbb735),
	.w4(32'h3b53aeb2),
	.w5(32'hbab6d5cb),
	.w6(32'h3ac0a7fd),
	.w7(32'h3b48c81a),
	.w8(32'hbc0a366c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91b393),
	.w1(32'hbc1a4023),
	.w2(32'hbbab1ac0),
	.w3(32'hbb9832e2),
	.w4(32'h3b473240),
	.w5(32'hba97c619),
	.w6(32'hbc868d7b),
	.w7(32'hbc60f0f9),
	.w8(32'hbab941ab),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52920b),
	.w1(32'h3b9eab6a),
	.w2(32'h3b9ec5c9),
	.w3(32'hbb294e39),
	.w4(32'h3c38c4ad),
	.w5(32'h3bd79833),
	.w6(32'hbc037ba6),
	.w7(32'hbc0e1c51),
	.w8(32'hbc221eab),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb782f4b),
	.w1(32'h395871f3),
	.w2(32'hb99e4abe),
	.w3(32'h3a7ae42b),
	.w4(32'hbb7dd963),
	.w5(32'hbb29c6e2),
	.w6(32'h3b820dcb),
	.w7(32'h3b27aa6e),
	.w8(32'hbaa743c1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc5ebd),
	.w1(32'h3a982c99),
	.w2(32'h3a977c51),
	.w3(32'hbac6eb0b),
	.w4(32'h3a05a012),
	.w5(32'h3aa7eb7b),
	.w6(32'h389985b8),
	.w7(32'hbac4f8bb),
	.w8(32'hbb0aa481),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52b7d4),
	.w1(32'hbb525b00),
	.w2(32'hbb0f7e93),
	.w3(32'hbb177188),
	.w4(32'hbb8d30c9),
	.w5(32'hbb30d49e),
	.w6(32'hbab51f02),
	.w7(32'hbb3317be),
	.w8(32'hbb8e2f55),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9768ace),
	.w1(32'hbbfb64ca),
	.w2(32'hbbd163bd),
	.w3(32'hba0fdbb0),
	.w4(32'h3aae9e52),
	.w5(32'h39d90ca2),
	.w6(32'h3ae809d5),
	.w7(32'h3bf142b1),
	.w8(32'h3aa3decf),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7627b),
	.w1(32'hbcc27d8f),
	.w2(32'hbd248e6e),
	.w3(32'h3c191bdc),
	.w4(32'h3c1f93ce),
	.w5(32'h3c3de193),
	.w6(32'h3c264e9b),
	.w7(32'h3c0dc442),
	.w8(32'h3ba5048b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf07ea),
	.w1(32'hbb14dd53),
	.w2(32'hbad634e4),
	.w3(32'h3c8f5672),
	.w4(32'h39a46f83),
	.w5(32'hbbf30334),
	.w6(32'hbc007577),
	.w7(32'hbc089f88),
	.w8(32'hbbbacec5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cf2dd),
	.w1(32'h3cd271b7),
	.w2(32'h3d3c9782),
	.w3(32'hbc08e14b),
	.w4(32'h3c809eb5),
	.w5(32'h3c576f12),
	.w6(32'hbc696ddf),
	.w7(32'hbb85509c),
	.w8(32'hb9dce9c8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3383f),
	.w1(32'hbb809752),
	.w2(32'hbc70cc46),
	.w3(32'h3c424553),
	.w4(32'hbc4ccb44),
	.w5(32'hbc7fc401),
	.w6(32'h3c795b67),
	.w7(32'h3c51d197),
	.w8(32'h3be41d40),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed7c63),
	.w1(32'h3ac749f5),
	.w2(32'h3ac58778),
	.w3(32'hbbe090a8),
	.w4(32'h3bb87c0c),
	.w5(32'hb78b079a),
	.w6(32'h3b7e3879),
	.w7(32'h3b9d5d86),
	.w8(32'hbac341ad),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d1c9f),
	.w1(32'h3b62aaa4),
	.w2(32'hbc301c05),
	.w3(32'hbc0f2299),
	.w4(32'hbbfdf120),
	.w5(32'hbcc45de7),
	.w6(32'h3c579414),
	.w7(32'h3c63411e),
	.w8(32'h3a7789d3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35bcc4),
	.w1(32'h3bfaf551),
	.w2(32'h3a8c4621),
	.w3(32'hbc82d1ff),
	.w4(32'hbbedbb51),
	.w5(32'hbc953c2d),
	.w6(32'h3c3c7203),
	.w7(32'h3c1cf0f1),
	.w8(32'h3bf1e067),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc026105),
	.w1(32'hbb62bb00),
	.w2(32'hbc105b68),
	.w3(32'hbc194bd1),
	.w4(32'h3ba9fb3d),
	.w5(32'hbafa68a7),
	.w6(32'hbbddf3b6),
	.w7(32'hbc1d9b12),
	.w8(32'hbbf02cb2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5da5c2),
	.w1(32'hbae9b4e7),
	.w2(32'hbad7cd27),
	.w3(32'hba7277bb),
	.w4(32'hb98f7901),
	.w5(32'hbb25d5be),
	.w6(32'hbba0b44d),
	.w7(32'hbaf6e585),
	.w8(32'hbbedbdb8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe031c0),
	.w1(32'hbb22d403),
	.w2(32'hbc987781),
	.w3(32'hbb2a6c11),
	.w4(32'h3bd7522a),
	.w5(32'h3b35a506),
	.w6(32'h3a8d8501),
	.w7(32'hbc86d14e),
	.w8(32'hbc286cf3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ed0c7),
	.w1(32'hba93be4e),
	.w2(32'hb988e837),
	.w3(32'hbb311e83),
	.w4(32'hbb94c8f5),
	.w5(32'hbc2850e6),
	.w6(32'h3bdd820a),
	.w7(32'h3bdcb348),
	.w8(32'hb9868de0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12d81a),
	.w1(32'h3b69a12c),
	.w2(32'h3b832284),
	.w3(32'hbbeebc50),
	.w4(32'hb99cdf85),
	.w5(32'hbad0741b),
	.w6(32'h3bc48ccc),
	.w7(32'h3b43f962),
	.w8(32'hb79bb7d2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b1dc4e),
	.w1(32'h3ae7436e),
	.w2(32'h39f8b097),
	.w3(32'h3a49b6af),
	.w4(32'h3b83e78e),
	.w5(32'hbbc77d00),
	.w6(32'hb92c1320),
	.w7(32'hba9f91e2),
	.w8(32'hbb0414f2),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ccd46),
	.w1(32'h3b549b6f),
	.w2(32'h3c45a286),
	.w3(32'hbbac6d68),
	.w4(32'h3ca12cb4),
	.w5(32'h3cb6a669),
	.w6(32'hbd0da3cd),
	.w7(32'hbcf0c553),
	.w8(32'hbc3383a9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ca5d7),
	.w1(32'h3c2a3ded),
	.w2(32'h3c4f2a27),
	.w3(32'h3a2d02cb),
	.w4(32'hbb8fb2ca),
	.w5(32'hbc0549dd),
	.w6(32'h3b68faf1),
	.w7(32'h38e439a0),
	.w8(32'h39e45b4e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7bc21),
	.w1(32'h3cd6fc1c),
	.w2(32'h3cf8cdfe),
	.w3(32'hbc23c815),
	.w4(32'h3c463786),
	.w5(32'h39460346),
	.w6(32'h3af216e5),
	.w7(32'h3c5523a0),
	.w8(32'h3bd93221),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c255717),
	.w1(32'hb97edb23),
	.w2(32'hbb7eb8cf),
	.w3(32'hbc1c02c4),
	.w4(32'h3b1b1894),
	.w5(32'hbba130b8),
	.w6(32'h3bb8e280),
	.w7(32'hbaff6e4f),
	.w8(32'hba0c4fc0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08cf0a),
	.w1(32'h3a0282e3),
	.w2(32'hbc34b900),
	.w3(32'hbbbcc131),
	.w4(32'hbc0d8ab4),
	.w5(32'hbc4380fa),
	.w6(32'h3aead5bc),
	.w7(32'hba8a586a),
	.w8(32'h3c18ff6b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fb509),
	.w1(32'h3c39ecef),
	.w2(32'h3c6bebcd),
	.w3(32'hbc680980),
	.w4(32'h3c138099),
	.w5(32'hbad71fbd),
	.w6(32'hb997fd41),
	.w7(32'h3b9e5efc),
	.w8(32'hbaabb54f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f2eeb),
	.w1(32'h3b3cf92c),
	.w2(32'h3c012264),
	.w3(32'hbb92f606),
	.w4(32'h3c44430f),
	.w5(32'h3b1e28a2),
	.w6(32'hbbe30757),
	.w7(32'h3c74913a),
	.w8(32'h3be49374),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b454b),
	.w1(32'hbb7c0519),
	.w2(32'hbad0d3fc),
	.w3(32'hbb0900c5),
	.w4(32'hb9f1415e),
	.w5(32'h3b303584),
	.w6(32'hbac0eef2),
	.w7(32'h3a1533a9),
	.w8(32'h3ad4b4e4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2df81a),
	.w1(32'h3be0d3ab),
	.w2(32'h3c0be907),
	.w3(32'h3b8b0175),
	.w4(32'h3bdfddb5),
	.w5(32'h3b3884c6),
	.w6(32'h3b002d49),
	.w7(32'hbae3d9e9),
	.w8(32'hbae36343),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6d616),
	.w1(32'hbb9e1316),
	.w2(32'hbba0519b),
	.w3(32'h3ac7abfc),
	.w4(32'h3ba919bb),
	.w5(32'h3b128827),
	.w6(32'hbb990c8f),
	.w7(32'hbb9b6422),
	.w8(32'hbbb0d9e6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb242a4c),
	.w1(32'h3b91d201),
	.w2(32'hbb29f15a),
	.w3(32'h3bb5f82b),
	.w4(32'hbc13dcf0),
	.w5(32'hbcb436a0),
	.w6(32'h3b375053),
	.w7(32'h3bcf0c1b),
	.w8(32'h3b867291),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61d789),
	.w1(32'h3b9fd3b7),
	.w2(32'h3bd74dae),
	.w3(32'hbc033b55),
	.w4(32'hba82f704),
	.w5(32'hbc9ee8b4),
	.w6(32'h3c3a1333),
	.w7(32'h3c3a863e),
	.w8(32'h3a2a0523),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdeaf44),
	.w1(32'h3b58a322),
	.w2(32'h3c4ca074),
	.w3(32'hbc865a24),
	.w4(32'h3bcfd2ff),
	.w5(32'hbb324957),
	.w6(32'hbc2f25ec),
	.w7(32'hbb9f15fd),
	.w8(32'hbafb228a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e7e95),
	.w1(32'hbb037244),
	.w2(32'hbb7681e6),
	.w3(32'hbb87a048),
	.w4(32'hbb0e254b),
	.w5(32'hbb6484d5),
	.w6(32'hbb37c888),
	.w7(32'hba4f3315),
	.w8(32'hb9f1403f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3d757),
	.w1(32'h3aa1c3ac),
	.w2(32'hb99aa082),
	.w3(32'hb945ade0),
	.w4(32'hbb1950c6),
	.w5(32'h3a1fa119),
	.w6(32'hbb07d41e),
	.w7(32'hbb603494),
	.w8(32'hbb8c03b1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8be9f3),
	.w1(32'h3b081147),
	.w2(32'hbbb6eb62),
	.w3(32'h3ac1b3e5),
	.w4(32'hbc649fd2),
	.w5(32'hbbc42f2a),
	.w6(32'h3c01b779),
	.w7(32'hbb20aba5),
	.w8(32'hbc405356),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c269ea2),
	.w1(32'h3b2e4a8c),
	.w2(32'h3b9362d3),
	.w3(32'h3bea0817),
	.w4(32'hba188331),
	.w5(32'hbbda0540),
	.w6(32'hba39aa20),
	.w7(32'hb9d63db6),
	.w8(32'h371c0265),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c99e6),
	.w1(32'hbbfc02d7),
	.w2(32'hbcc8b1af),
	.w3(32'hbb82a327),
	.w4(32'h371d34e9),
	.w5(32'hbbb86173),
	.w6(32'h3b8cfa92),
	.w7(32'h3b8587b6),
	.w8(32'hbb5117a1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc807e64),
	.w1(32'hbc60d0aa),
	.w2(32'hbcf30582),
	.w3(32'hbba57503),
	.w4(32'h3bbc0e50),
	.w5(32'h3b76163c),
	.w6(32'hbb282bea),
	.w7(32'hbc8f7678),
	.w8(32'hbc134261),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1d5eb),
	.w1(32'hbc964ab0),
	.w2(32'hbcf18084),
	.w3(32'h3bfa4cff),
	.w4(32'hbb6aad4c),
	.w5(32'h3be48c84),
	.w6(32'hbc42cdfd),
	.w7(32'hbcbaff37),
	.w8(32'hbc59ed6b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d1191),
	.w1(32'h3bd008a4),
	.w2(32'h3c0fbe5b),
	.w3(32'h3c3d1b01),
	.w4(32'hb9db0c19),
	.w5(32'h3b28204c),
	.w6(32'hbc2011b7),
	.w7(32'hbc35cf36),
	.w8(32'h399e0eec),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c074528),
	.w1(32'h3c08b0e9),
	.w2(32'h3c6d7046),
	.w3(32'h3bd0c6dc),
	.w4(32'hbc9d3da9),
	.w5(32'hbc404a6d),
	.w6(32'h3c85daea),
	.w7(32'h3c8889ee),
	.w8(32'h3c9a6a08),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb780e6),
	.w1(32'hbb9e9c40),
	.w2(32'hbaf9a85a),
	.w3(32'h3bbc9c75),
	.w4(32'hbc6ce549),
	.w5(32'hbcacec23),
	.w6(32'h3ab6ec12),
	.w7(32'h3b99d321),
	.w8(32'h3b4473d4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c1a66),
	.w1(32'h3c4fdd81),
	.w2(32'h3c9923f7),
	.w3(32'hbc6ea31d),
	.w4(32'h3b18b9b2),
	.w5(32'hbc52905c),
	.w6(32'h3c4a3cad),
	.w7(32'h3c9bef2e),
	.w8(32'h3b618729),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a932e13),
	.w1(32'hbccb8679),
	.w2(32'hbc8d211d),
	.w3(32'hbc95df50),
	.w4(32'h3bede85b),
	.w5(32'h3bdfa5a8),
	.w6(32'hbc107861),
	.w7(32'hb9aeece8),
	.w8(32'hb9a59a41),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb083e82),
	.w1(32'hbc9fdf78),
	.w2(32'hbc8da3d7),
	.w3(32'h3c85d866),
	.w4(32'h3ca92906),
	.w5(32'h3b92123a),
	.w6(32'hbc28ac5d),
	.w7(32'hbca1463a),
	.w8(32'hbc2e6d43),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb02de8),
	.w1(32'hbb79fc6d),
	.w2(32'hbb115c05),
	.w3(32'hbb844213),
	.w4(32'h3b1e0c94),
	.w5(32'h3ac9a404),
	.w6(32'hbba9ad8d),
	.w7(32'hbb819b51),
	.w8(32'hbb615ea9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b411881),
	.w1(32'hbba919e9),
	.w2(32'hbc3e17c8),
	.w3(32'hba8f5f15),
	.w4(32'h3bd58ecb),
	.w5(32'h3bb1b246),
	.w6(32'h3b2652c4),
	.w7(32'h3b1dfd7e),
	.w8(32'hbb1b2d4e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc176603),
	.w1(32'h3bff6ced),
	.w2(32'h3baedf39),
	.w3(32'h3bc1366a),
	.w4(32'h3c1566c9),
	.w5(32'h3ae398a2),
	.w6(32'hbab2a2db),
	.w7(32'h3b07641f),
	.w8(32'h3bb55373),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b371e2a),
	.w1(32'h3bc2e35f),
	.w2(32'hbb18de4a),
	.w3(32'hbb3c80f5),
	.w4(32'hbbaeeb21),
	.w5(32'hbb7d60a5),
	.w6(32'h3b05fae1),
	.w7(32'hbb2a4557),
	.w8(32'hbb18d31e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe33320),
	.w1(32'h3b68bef1),
	.w2(32'h39b0dc27),
	.w3(32'hbba65e7e),
	.w4(32'h3b0b11dd),
	.w5(32'hb81e8bf4),
	.w6(32'h3a7d3e20),
	.w7(32'h399b009a),
	.w8(32'h37b93ba9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40c234),
	.w1(32'h3bcd6ff7),
	.w2(32'h3c423411),
	.w3(32'h3829c40a),
	.w4(32'hbb81e943),
	.w5(32'hbc3fb2c6),
	.w6(32'h3b78e067),
	.w7(32'h39e047bc),
	.w8(32'hb99cb930),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1c2e1),
	.w1(32'h3ac09197),
	.w2(32'hbac36949),
	.w3(32'hbcb426ea),
	.w4(32'hbb7daf34),
	.w5(32'hbbe8c0ce),
	.w6(32'hbabca0fc),
	.w7(32'hbb89c92c),
	.w8(32'hbb3111a2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb051d29),
	.w1(32'hbaf3fc8c),
	.w2(32'hba28103b),
	.w3(32'hbbe1b432),
	.w4(32'h3a31c439),
	.w5(32'hbba590f4),
	.w6(32'h3b2bf932),
	.w7(32'hb9e8a6dd),
	.w8(32'hbb059562),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa69a61),
	.w1(32'hbc01182f),
	.w2(32'hbcf5d345),
	.w3(32'h3b98d134),
	.w4(32'h3b54c7e6),
	.w5(32'h3be97e00),
	.w6(32'h3acf52ae),
	.w7(32'hbbaf9b18),
	.w8(32'hbb861004),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1a32a),
	.w1(32'hbbcad79b),
	.w2(32'hba0443c4),
	.w3(32'h3c76514e),
	.w4(32'h3949e536),
	.w5(32'hbb360423),
	.w6(32'hbb5ce6db),
	.w7(32'h3a266743),
	.w8(32'hba4f5827),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03214c),
	.w1(32'h38b6b7c1),
	.w2(32'hba3d70e8),
	.w3(32'hbb0ce836),
	.w4(32'hbabfae52),
	.w5(32'hbabe7ced),
	.w6(32'hba6dda3f),
	.w7(32'hbb271542),
	.w8(32'hbb72ec57),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb311610),
	.w1(32'hbbe05281),
	.w2(32'hbb3bdf35),
	.w3(32'hba01d5ce),
	.w4(32'hba3a44af),
	.w5(32'hbad37c63),
	.w6(32'hbb129ac3),
	.w7(32'h3b2053be),
	.w8(32'h3a8e5200),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba638ba0),
	.w1(32'h3b35f7ce),
	.w2(32'h3ba4b5f7),
	.w3(32'hbb1aabc7),
	.w4(32'h3bacd99a),
	.w5(32'h3aed9724),
	.w6(32'hbba7af9f),
	.w7(32'hbbe0b26d),
	.w8(32'hbb2ef552),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7a46a),
	.w1(32'h3b36baa4),
	.w2(32'h3c3b5111),
	.w3(32'h3b28af91),
	.w4(32'hbc451ac6),
	.w5(32'hbcb0b84c),
	.w6(32'hbb6d9c91),
	.w7(32'h3bbe29b8),
	.w8(32'h3c2c3117),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca88dc),
	.w1(32'hbaa7e2f1),
	.w2(32'h3ac7117b),
	.w3(32'hbc4a7747),
	.w4(32'hba2d9f4b),
	.w5(32'hba2dc421),
	.w6(32'hba63ffbb),
	.w7(32'h3ac63089),
	.w8(32'hbbecbbca),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf0266),
	.w1(32'h3c870216),
	.w2(32'h3d35e78b),
	.w3(32'h3adef6d9),
	.w4(32'h3c5e9a78),
	.w5(32'h3cb4593b),
	.w6(32'hbc8d5ee7),
	.w7(32'hbc0c9570),
	.w8(32'h3a2a3e21),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc71036),
	.w1(32'h3af17d74),
	.w2(32'h3c34f32f),
	.w3(32'h3c8805b6),
	.w4(32'h3a6935ba),
	.w5(32'hba18af66),
	.w6(32'hbba0057e),
	.w7(32'hbb21245a),
	.w8(32'hbad53365),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11441a),
	.w1(32'h3aa2b9d5),
	.w2(32'hbb3bc87c),
	.w3(32'h3adb7922),
	.w4(32'hbb0f8201),
	.w5(32'hbb8eaf6e),
	.w6(32'h39858a00),
	.w7(32'hbb59a843),
	.w8(32'hbb1d0205),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb482743),
	.w1(32'hba8eefca),
	.w2(32'hbba9fe34),
	.w3(32'hbb54afb7),
	.w4(32'h3abf39cd),
	.w5(32'hbb307426),
	.w6(32'hb71c8383),
	.w7(32'h3b8f9598),
	.w8(32'h3b41893c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b031993),
	.w1(32'hbbf06266),
	.w2(32'hbc1fd80c),
	.w3(32'h3be2d4d6),
	.w4(32'hbc85a713),
	.w5(32'hbcfd6914),
	.w6(32'h3c7a089a),
	.w7(32'h3cc78610),
	.w8(32'h3c6186d5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc805bd9),
	.w1(32'hbb39d545),
	.w2(32'hbbc718b6),
	.w3(32'hbcc5ff02),
	.w4(32'hbb6a1ff2),
	.w5(32'hbb67a5e8),
	.w6(32'hbbb5ae48),
	.w7(32'h3b8ebd77),
	.w8(32'h3bdb60d8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf69e7e),
	.w1(32'hbaa45317),
	.w2(32'hbc10f6b0),
	.w3(32'hba93bd1d),
	.w4(32'hb9a7904e),
	.w5(32'hbc12bdcc),
	.w6(32'h3a393265),
	.w7(32'hbbefd464),
	.w8(32'hb8c03227),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dc5e5),
	.w1(32'hbc25afd8),
	.w2(32'hbbadfc12),
	.w3(32'hba8f98c4),
	.w4(32'hba8bef33),
	.w5(32'h3b8a48ba),
	.w6(32'hbc249c56),
	.w7(32'hbbd38a55),
	.w8(32'h3c240a6b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule