module layer_10_featuremap_379(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf37b2f),
	.w1(32'hbb14b2db),
	.w2(32'hba84d25f),
	.w3(32'hbbe23606),
	.w4(32'hbbe0b921),
	.w5(32'hbaab99ea),
	.w6(32'hbb3fd5d5),
	.w7(32'hba588411),
	.w8(32'h3b0d3a9c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb054b3c),
	.w1(32'h3ad6795f),
	.w2(32'h3aa726c2),
	.w3(32'hbb11c240),
	.w4(32'hbb077892),
	.w5(32'hb9e034ff),
	.w6(32'h3b873364),
	.w7(32'h3a893f6e),
	.w8(32'h398bca05),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9a29d),
	.w1(32'h398d9f60),
	.w2(32'h3b7ff336),
	.w3(32'h3ab738ba),
	.w4(32'h3b6577a7),
	.w5(32'hbb09daef),
	.w6(32'hb9ad6560),
	.w7(32'hbb92bb3d),
	.w8(32'h38b20e51),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a39d9),
	.w1(32'hbb690cb1),
	.w2(32'h3b240015),
	.w3(32'h3b9bac46),
	.w4(32'hbc18c009),
	.w5(32'hbba4cf3f),
	.w6(32'hba9b50c6),
	.w7(32'h3ab7f757),
	.w8(32'h3c28d119),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82389a),
	.w1(32'hbbe33827),
	.w2(32'hba8ea3c5),
	.w3(32'hb9c3568d),
	.w4(32'hbb10bc3f),
	.w5(32'hbb60e647),
	.w6(32'h3bd0799c),
	.w7(32'hba8c91ab),
	.w8(32'h3bb1fc15),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ee97e),
	.w1(32'h3b725f24),
	.w2(32'h3ae7a12a),
	.w3(32'hbbe81f25),
	.w4(32'h3ca97ca0),
	.w5(32'h3c0eb2cc),
	.w6(32'h3b4c8ca1),
	.w7(32'hbc055cb2),
	.w8(32'hbb83ce31),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2af03e),
	.w1(32'h3aae877b),
	.w2(32'hbb92cdf2),
	.w3(32'h3bd9acee),
	.w4(32'h3bdd6abb),
	.w5(32'h3ce96d1c),
	.w6(32'h3c59b36d),
	.w7(32'hba54cd82),
	.w8(32'hbc8390f1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7af355),
	.w1(32'h3bdcc0b0),
	.w2(32'h3c027ebb),
	.w3(32'hbc2ebe03),
	.w4(32'hbc5304d2),
	.w5(32'hbbfe8a1a),
	.w6(32'hbc255976),
	.w7(32'hbb3a7edb),
	.w8(32'hbb9e1ce4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49a268),
	.w1(32'hbb6bfd9e),
	.w2(32'hbb872c1b),
	.w3(32'h3ba63f26),
	.w4(32'hbc126599),
	.w5(32'hbbcd0c72),
	.w6(32'h3b3b630f),
	.w7(32'hbbb4ea04),
	.w8(32'hbc3654ea),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a06c3),
	.w1(32'hbc93b7d9),
	.w2(32'hbcbc134d),
	.w3(32'hbc06a56a),
	.w4(32'hbb928dcc),
	.w5(32'hbbc03bda),
	.w6(32'hbba64261),
	.w7(32'hbb43fac1),
	.w8(32'hbbb878eb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6488fc),
	.w1(32'hbc09660b),
	.w2(32'hbb89202a),
	.w3(32'hbc03862f),
	.w4(32'h3baf79ea),
	.w5(32'h3c287f4c),
	.w6(32'hbb8d3297),
	.w7(32'hbbd71597),
	.w8(32'hbc44fbfa),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf89092),
	.w1(32'h3a128268),
	.w2(32'hbaa59412),
	.w3(32'h3babc35e),
	.w4(32'hbbb0b138),
	.w5(32'hbb6aaafc),
	.w6(32'hb9afa6a5),
	.w7(32'hbb4e6d6f),
	.w8(32'hbbf7abfc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc805347),
	.w1(32'hbba8295a),
	.w2(32'hbc1d6cb2),
	.w3(32'hbba3cda7),
	.w4(32'hbc5124e4),
	.w5(32'hbc707678),
	.w6(32'hbc00065b),
	.w7(32'hbb8d89a5),
	.w8(32'hba73935a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5a0ca),
	.w1(32'h3aa5d620),
	.w2(32'h3b1ef600),
	.w3(32'hbaf58724),
	.w4(32'h3bd99736),
	.w5(32'h3bac50a8),
	.w6(32'h3bdcf9f7),
	.w7(32'h3b8d66d8),
	.w8(32'hbb024aa2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10ad4c),
	.w1(32'hbb6d89ee),
	.w2(32'hbbf0c48d),
	.w3(32'h3b7ba398),
	.w4(32'h3c16e9fe),
	.w5(32'h3c91fd6d),
	.w6(32'hbbaf9975),
	.w7(32'h3bbb013e),
	.w8(32'h3b72a1ad),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc110204),
	.w1(32'hbbc0c02a),
	.w2(32'hbbea20e1),
	.w3(32'h3ae5e629),
	.w4(32'hbbc4a6b0),
	.w5(32'hbacecd4a),
	.w6(32'h3b854db5),
	.w7(32'hbb845e70),
	.w8(32'h39c00d04),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e5ae2),
	.w1(32'hbb9186c3),
	.w2(32'hbb5591d9),
	.w3(32'hbb700af3),
	.w4(32'hbb86a25c),
	.w5(32'hbbca54c4),
	.w6(32'hbaa93eb4),
	.w7(32'h3b51c76d),
	.w8(32'hbc170191),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f9e7e),
	.w1(32'hbb2b658a),
	.w2(32'hbb62016f),
	.w3(32'hbc06304a),
	.w4(32'hbbb336e1),
	.w5(32'hbb53308e),
	.w6(32'hbc46e8a4),
	.w7(32'hbb802151),
	.w8(32'hbc46aad9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a588196),
	.w1(32'hbbbef4b0),
	.w2(32'hbbed3616),
	.w3(32'h3c098a7d),
	.w4(32'hba33fe0b),
	.w5(32'hbbe19147),
	.w6(32'h3a1cae51),
	.w7(32'h3b289e15),
	.w8(32'hbb62fd4f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba089ebc),
	.w1(32'h3b8c49bf),
	.w2(32'hbc92fd33),
	.w3(32'h3b2bdf24),
	.w4(32'h3aa222f8),
	.w5(32'h3d308ae6),
	.w6(32'hba35085d),
	.w7(32'hb9ff12d3),
	.w8(32'hbcb56f44),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf17c4),
	.w1(32'hba314787),
	.w2(32'h3b5b5c13),
	.w3(32'h3bb9db17),
	.w4(32'hbb4f8c9b),
	.w5(32'hbbd94326),
	.w6(32'h3bdb05a0),
	.w7(32'hba9cdca0),
	.w8(32'h3aeae7b6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab054c3),
	.w1(32'h3b8a90e6),
	.w2(32'h3abfa9ac),
	.w3(32'hbb784e75),
	.w4(32'hbbbbdd05),
	.w5(32'hbc04bb9e),
	.w6(32'h3b3ca5ed),
	.w7(32'hbb2fbca1),
	.w8(32'h393d04e0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe33d8),
	.w1(32'hbb5153a3),
	.w2(32'hbc043bc4),
	.w3(32'hbb986d37),
	.w4(32'h3c4fe06d),
	.w5(32'h3d2ad995),
	.w6(32'hbba42905),
	.w7(32'h3c447ed8),
	.w8(32'hbc15bbee),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1289a),
	.w1(32'hbb90ba7e),
	.w2(32'hbbf69ac4),
	.w3(32'h3c84c888),
	.w4(32'hbc214d0e),
	.w5(32'hbc8a44ac),
	.w6(32'h3bb02b87),
	.w7(32'h3a2bb73c),
	.w8(32'h3aedbe84),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93d79b),
	.w1(32'hbc0094af),
	.w2(32'hbc500cd8),
	.w3(32'hbc974ef3),
	.w4(32'hbb4e9eb8),
	.w5(32'h39be09d5),
	.w6(32'hbc6cc085),
	.w7(32'h3bcb3f2a),
	.w8(32'hbbc1951b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74d24d),
	.w1(32'h3bbfe727),
	.w2(32'h3c14eb68),
	.w3(32'h3c850ccb),
	.w4(32'h38e73a70),
	.w5(32'hbc8c0787),
	.w6(32'h3b55ac4a),
	.w7(32'h3b83a347),
	.w8(32'h3bff9b39),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b5e43),
	.w1(32'hbc2bdb62),
	.w2(32'h39cbe2a5),
	.w3(32'h3ab4551c),
	.w4(32'hbb188c2c),
	.w5(32'h3ab09a45),
	.w6(32'h3b21b563),
	.w7(32'hbb605cfa),
	.w8(32'hbb8b9f69),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8f20c),
	.w1(32'h3b9ff302),
	.w2(32'hbb36b9a3),
	.w3(32'hbbbc8485),
	.w4(32'hba195ab7),
	.w5(32'hbb2dc55c),
	.w6(32'hbc020b80),
	.w7(32'hbaf6dddc),
	.w8(32'hbb54de0f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02082e),
	.w1(32'hbc5c6ce3),
	.w2(32'hbccf38bb),
	.w3(32'hbb1e43a4),
	.w4(32'h3c4817a0),
	.w5(32'h3c7d4483),
	.w6(32'hbbb1bb03),
	.w7(32'h3bafbbe0),
	.w8(32'hbc4c445a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ded09),
	.w1(32'hbb160c55),
	.w2(32'hbc1e6c2c),
	.w3(32'hbc26c5d7),
	.w4(32'h3ab2154c),
	.w5(32'hbba28ab7),
	.w6(32'hbc294c85),
	.w7(32'hbbfd8871),
	.w8(32'hbc08b324),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2522f9),
	.w1(32'h3c3fe8a6),
	.w2(32'h3bcd64ed),
	.w3(32'h3aca43f5),
	.w4(32'h3c8bf23b),
	.w5(32'h3d7d6a88),
	.w6(32'hbb4094c2),
	.w7(32'h3bdfb394),
	.w8(32'hbc330fe8),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42643f),
	.w1(32'hbb443a9e),
	.w2(32'hbb93aca2),
	.w3(32'h3c809be2),
	.w4(32'hbb3092f1),
	.w5(32'hbbb52413),
	.w6(32'h3ba3e978),
	.w7(32'hbbfc019e),
	.w8(32'hbc17ae0c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01a288),
	.w1(32'hbc023205),
	.w2(32'hbbab4e40),
	.w3(32'hb9121d72),
	.w4(32'hba30e5d4),
	.w5(32'hbbd992b6),
	.w6(32'hb9740a98),
	.w7(32'hbb8dc49e),
	.w8(32'hbbc96a20),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba914e8),
	.w1(32'hbb624adc),
	.w2(32'hbb618de2),
	.w3(32'hbc227474),
	.w4(32'hba896576),
	.w5(32'h3b93510d),
	.w6(32'hbc4ef44b),
	.w7(32'h3bd52546),
	.w8(32'hbb77353a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae71d23),
	.w1(32'h3c04c1b3),
	.w2(32'h3b9225ea),
	.w3(32'h3b0aa04d),
	.w4(32'h3c1f5581),
	.w5(32'h3bc6d419),
	.w6(32'h3b35551c),
	.w7(32'h3b56aab3),
	.w8(32'h3c071e32),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7aab65),
	.w1(32'h399c2eee),
	.w2(32'h3ae2f543),
	.w3(32'h3c085744),
	.w4(32'hba82099e),
	.w5(32'hbabb1426),
	.w6(32'hbb6881d4),
	.w7(32'h3c05539b),
	.w8(32'h3b8c4753),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1265b6),
	.w1(32'hbbb85236),
	.w2(32'hbbcf3c0f),
	.w3(32'h3a483ac8),
	.w4(32'h3b82239b),
	.w5(32'h3b2fe423),
	.w6(32'h3bcba63a),
	.w7(32'h3b82541b),
	.w8(32'hbc53a93a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0feabc),
	.w1(32'h3c2adad7),
	.w2(32'h3c0dc00d),
	.w3(32'hbc2f439e),
	.w4(32'h3ba93938),
	.w5(32'h3c8ac417),
	.w6(32'hbbf536ee),
	.w7(32'h3ba20af3),
	.w8(32'hbae8e289),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba7d7c),
	.w1(32'h3b85dfc6),
	.w2(32'h3a4dcaa3),
	.w3(32'hbc0478cf),
	.w4(32'hb8fd0083),
	.w5(32'h3aa0cd60),
	.w6(32'hbbc482c5),
	.w7(32'h3be06d1d),
	.w8(32'h3b96ca0f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39417eaa),
	.w1(32'h3b3fa59e),
	.w2(32'h3b5c79b7),
	.w3(32'h3b428402),
	.w4(32'hbb15354a),
	.w5(32'hbb278a54),
	.w6(32'h3b6b9492),
	.w7(32'h3b3c3212),
	.w8(32'h3b3d92b5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b219521),
	.w1(32'hbb201869),
	.w2(32'hba81fa60),
	.w3(32'h3bf4d65d),
	.w4(32'hbc11df78),
	.w5(32'hbbb210d3),
	.w6(32'hbb27289b),
	.w7(32'h3b21a6aa),
	.w8(32'h3c7495d9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba754d),
	.w1(32'h3b244700),
	.w2(32'h3bc3b065),
	.w3(32'hbb1ad4c4),
	.w4(32'hbb0f894d),
	.w5(32'h3ad1a953),
	.w6(32'h3c0667c2),
	.w7(32'hbc08b16e),
	.w8(32'hbbf03f36),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a557154),
	.w1(32'hbabc5cae),
	.w2(32'h3b6c70a5),
	.w3(32'hbb100547),
	.w4(32'h3ada581d),
	.w5(32'hbab8974f),
	.w6(32'hbb735fe9),
	.w7(32'h3af26ae4),
	.w8(32'h388dd6e0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28d825),
	.w1(32'hbbbc9f3c),
	.w2(32'hbc5b4961),
	.w3(32'hbbc71f80),
	.w4(32'hbc4fd6a3),
	.w5(32'hbc676568),
	.w6(32'hbc4c2475),
	.w7(32'hbc55590c),
	.w8(32'hbc395aed),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35d4e9),
	.w1(32'hbbb0b42f),
	.w2(32'hbc3f098b),
	.w3(32'hbbdab7a4),
	.w4(32'hbb621475),
	.w5(32'hbc349048),
	.w6(32'h3ac2d001),
	.w7(32'h3b17c7f1),
	.w8(32'hbb50ad7e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44dbdc),
	.w1(32'hba3b9abb),
	.w2(32'hbbfd2d3e),
	.w3(32'hbbe4d369),
	.w4(32'hbbc405b6),
	.w5(32'hbadd20a9),
	.w6(32'hba8c058a),
	.w7(32'hb8420f89),
	.w8(32'h3c5166d2),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59a839),
	.w1(32'h3afecce5),
	.w2(32'h3c2dae27),
	.w3(32'hbb4f756f),
	.w4(32'hbba17803),
	.w5(32'hba245888),
	.w6(32'h3be17f8b),
	.w7(32'hba61f422),
	.w8(32'h3b23dee7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba197b7),
	.w1(32'hbc00540e),
	.w2(32'hbc816c2b),
	.w3(32'hba27bef5),
	.w4(32'hbbff1ac4),
	.w5(32'hbbf3dc38),
	.w6(32'hbb91286d),
	.w7(32'hba776ff9),
	.w8(32'hbba57bb6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf22334),
	.w1(32'h3b0f0bc3),
	.w2(32'h3bc3f427),
	.w3(32'hbbded441),
	.w4(32'h3babcf70),
	.w5(32'hbb027699),
	.w6(32'h3a1493ef),
	.w7(32'h3b7cd2a1),
	.w8(32'h3b6eb8f9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad06a4b),
	.w1(32'h3b446393),
	.w2(32'h3bd221aa),
	.w3(32'h3a4a97cc),
	.w4(32'h3b0592e9),
	.w5(32'hbb266584),
	.w6(32'h3b4d0395),
	.w7(32'h3b0c80de),
	.w8(32'h3ab7c1a9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ee002),
	.w1(32'hbb2296a6),
	.w2(32'hbc0bc116),
	.w3(32'h3ad4c353),
	.w4(32'hbb18d871),
	.w5(32'hbc0691e8),
	.w6(32'h3b1ac170),
	.w7(32'h3c203b1f),
	.w8(32'h3a12d403),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbe98e),
	.w1(32'hbc2147e0),
	.w2(32'hbc1c7676),
	.w3(32'h3bc8f796),
	.w4(32'hbbf6ba38),
	.w5(32'hbbdad671),
	.w6(32'h39899d27),
	.w7(32'h3a777e89),
	.w8(32'h3b2ac015),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc152b40),
	.w1(32'h3ba156f4),
	.w2(32'h3b0be561),
	.w3(32'hbbd93f67),
	.w4(32'h3bde92e6),
	.w5(32'h3bbffc7e),
	.w6(32'hbc12003a),
	.w7(32'hbb7b8a33),
	.w8(32'hbb5c1195),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2465e),
	.w1(32'hbb82267b),
	.w2(32'hbc013c4c),
	.w3(32'h3a2fb6df),
	.w4(32'h3b0b8d56),
	.w5(32'hbb204b58),
	.w6(32'h3b31c43d),
	.w7(32'h3b3ddd9d),
	.w8(32'hb917fcc9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba876538),
	.w1(32'hbba1b67f),
	.w2(32'hbac75ad0),
	.w3(32'h3c28893a),
	.w4(32'hbc144d74),
	.w5(32'hbaf036db),
	.w6(32'hbb5e45a7),
	.w7(32'hbbe75673),
	.w8(32'hbbdd25f7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86ba5e),
	.w1(32'hba85e91a),
	.w2(32'hba34c9a4),
	.w3(32'h3b84877e),
	.w4(32'hbb548892),
	.w5(32'h3bf192a7),
	.w6(32'hbb6d5de0),
	.w7(32'hbbb72f28),
	.w8(32'hbb837a24),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23a0a7),
	.w1(32'hbbf62935),
	.w2(32'hbb9a9121),
	.w3(32'h39091589),
	.w4(32'h3b966199),
	.w5(32'h3c087c48),
	.w6(32'hbb81989d),
	.w7(32'h3bf96a22),
	.w8(32'h3b8a25aa),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2a26a),
	.w1(32'hba030f5c),
	.w2(32'hbb33f562),
	.w3(32'h3bb9a1ea),
	.w4(32'h3c03b8d2),
	.w5(32'hbc0d0621),
	.w6(32'h3a9c6d3d),
	.w7(32'hbc28d363),
	.w8(32'h3be24375),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb749fad),
	.w1(32'hb9011502),
	.w2(32'h3a27c6b7),
	.w3(32'hbba21365),
	.w4(32'hbc05ac4a),
	.w5(32'hbbf0eff1),
	.w6(32'h3a9f872d),
	.w7(32'hbc73a136),
	.w8(32'hbc56996e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf6d5b),
	.w1(32'hbafa49dd),
	.w2(32'h3aac546b),
	.w3(32'hbb556951),
	.w4(32'h3ab62c7c),
	.w5(32'hbc3c3811),
	.w6(32'hbc27d999),
	.w7(32'hbb04aca2),
	.w8(32'h3b8b559e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc788c),
	.w1(32'hbb9c788c),
	.w2(32'hbb806b9e),
	.w3(32'hbb9b892e),
	.w4(32'hbc906566),
	.w5(32'hbc17e61e),
	.w6(32'hbc5ad9d5),
	.w7(32'hbafae76d),
	.w8(32'h3b8d2fa2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb177a7d),
	.w1(32'hbb221d8e),
	.w2(32'hbb281545),
	.w3(32'hbc18db01),
	.w4(32'hbb92ffb6),
	.w5(32'h3acf58d6),
	.w6(32'hb892e202),
	.w7(32'hbc197ea1),
	.w8(32'hbc2cc386),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb031626),
	.w1(32'hbb8dda38),
	.w2(32'hbb8bca50),
	.w3(32'hbb120866),
	.w4(32'hbb688c51),
	.w5(32'hbb9b6c4f),
	.w6(32'hba95753a),
	.w7(32'hba0b1983),
	.w8(32'h3b3523f1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6062b),
	.w1(32'h3c1385f7),
	.w2(32'h3b015346),
	.w3(32'h3a4bb7ee),
	.w4(32'hbb296823),
	.w5(32'h3b062db1),
	.w6(32'hba2f091a),
	.w7(32'h3b0199d8),
	.w8(32'hbb0272ed),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f7da8),
	.w1(32'h3b66834c),
	.w2(32'h3b637e55),
	.w3(32'h3b447653),
	.w4(32'h3b4723d6),
	.w5(32'hba4ff35b),
	.w6(32'h39fdb6ec),
	.w7(32'h3b723665),
	.w8(32'h3b714dc1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab92ef0),
	.w1(32'h3b870304),
	.w2(32'h3b37e0df),
	.w3(32'h3b27a872),
	.w4(32'hb99b2614),
	.w5(32'h3bbbd27d),
	.w6(32'h3c07e5b2),
	.w7(32'hbb8f7002),
	.w8(32'hba8a21fe),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a10ad),
	.w1(32'h3a17bf92),
	.w2(32'hba928ac8),
	.w3(32'h3c01a1c5),
	.w4(32'hba9e3f40),
	.w5(32'hbb899c5f),
	.w6(32'h3b2a58e5),
	.w7(32'h3b9dc4bb),
	.w8(32'hba40e7b3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f1c95),
	.w1(32'h3bf6d810),
	.w2(32'hbb87f29f),
	.w3(32'h3c2a150e),
	.w4(32'hbbbbfa69),
	.w5(32'hbc9aa7e9),
	.w6(32'h3be08c9a),
	.w7(32'h3bd60ceb),
	.w8(32'h3bf4a46a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc355e4c),
	.w1(32'hbc461d38),
	.w2(32'hbc5f0772),
	.w3(32'hbbff87e5),
	.w4(32'hbc08ea4b),
	.w5(32'hbc15c1d3),
	.w6(32'hbb16f5b0),
	.w7(32'hb90d4863),
	.w8(32'hbbc2a3c2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc7b45),
	.w1(32'hbbd909ad),
	.w2(32'hbc8a8cb3),
	.w3(32'hbc0e95d5),
	.w4(32'h3b4240f0),
	.w5(32'hbbad6b6f),
	.w6(32'hbc365f66),
	.w7(32'hb99534f8),
	.w8(32'hbbc617a2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c9a88),
	.w1(32'h3772d9a3),
	.w2(32'h3b94984a),
	.w3(32'hbbb43023),
	.w4(32'h39b5f8c9),
	.w5(32'hbb2ea332),
	.w6(32'hbba7615e),
	.w7(32'hba9c41d6),
	.w8(32'h3a94c720),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a37c40),
	.w1(32'hb81a619d),
	.w2(32'hbadfcc1d),
	.w3(32'h3c1017f1),
	.w4(32'hbb3acd02),
	.w5(32'hbc2b1759),
	.w6(32'h3c60ec9a),
	.w7(32'h3a78b6e9),
	.w8(32'h3af1580e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c436979),
	.w1(32'h3a1e6c83),
	.w2(32'hbb3fb121),
	.w3(32'h3ba7d064),
	.w4(32'hbb513de7),
	.w5(32'hbb94e74b),
	.w6(32'hbc159378),
	.w7(32'hbb77dc52),
	.w8(32'hbb317d56),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3909552f),
	.w1(32'h3bbd700c),
	.w2(32'h3b1992bd),
	.w3(32'h3b7936f7),
	.w4(32'h3bcc72fb),
	.w5(32'h3b82e5d5),
	.w6(32'hbb0e2a5f),
	.w7(32'h3b7c5ae9),
	.w8(32'hba955cf2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03f5e3),
	.w1(32'hb9eca3c9),
	.w2(32'hbba68709),
	.w3(32'hbbcf2e13),
	.w4(32'h3b42b3bd),
	.w5(32'hb930f191),
	.w6(32'hbbf01366),
	.w7(32'hbb226b14),
	.w8(32'hbba84b87),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb991685),
	.w1(32'hbb2feba1),
	.w2(32'hbb66480f),
	.w3(32'hbb59119b),
	.w4(32'h39de6b07),
	.w5(32'hbbdcab74),
	.w6(32'hbb0d4874),
	.w7(32'h3b1d0230),
	.w8(32'hbb525be7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54ccca),
	.w1(32'h3abdbe5d),
	.w2(32'hbb03242a),
	.w3(32'hbbee2c07),
	.w4(32'h3a984105),
	.w5(32'h3b7a5067),
	.w6(32'hbc16c90f),
	.w7(32'h3a29fc9c),
	.w8(32'hbaefce30),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ff885),
	.w1(32'hbc94a5ed),
	.w2(32'hbc7258ad),
	.w3(32'h3a54b0bd),
	.w4(32'hbc68d2d3),
	.w5(32'hbc5209c4),
	.w6(32'h3a9a56eb),
	.w7(32'hbc2ab59a),
	.w8(32'hbc0f5a55),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c8150),
	.w1(32'hbc3141de),
	.w2(32'hbaf4ff2b),
	.w3(32'h3cf97064),
	.w4(32'hbc29d7c4),
	.w5(32'h3a8ac767),
	.w6(32'h3c3590c1),
	.w7(32'hbb49f71e),
	.w8(32'h3b1dcbee),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d7a0a),
	.w1(32'hbba756fb),
	.w2(32'hbb75c2d1),
	.w3(32'h3c84bbc0),
	.w4(32'h3a7ce702),
	.w5(32'h3b98fe9a),
	.w6(32'h3c7a08c4),
	.w7(32'hb9d76d7a),
	.w8(32'h3c193b0c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdfaf1),
	.w1(32'hbb583158),
	.w2(32'hbb52a6f8),
	.w3(32'hbb5eb0bf),
	.w4(32'hbb68c073),
	.w5(32'h3b470c5f),
	.w6(32'h3b478d17),
	.w7(32'h39f5fcea),
	.w8(32'hbb8b7f67),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaaaa24),
	.w1(32'hbbf99b6d),
	.w2(32'hbc02615b),
	.w3(32'h39ccfcae),
	.w4(32'hbc117add),
	.w5(32'hbc252c68),
	.w6(32'hbb374f8b),
	.w7(32'hbbe1d16e),
	.w8(32'hbbdf9df3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3db55f),
	.w1(32'hbc3758be),
	.w2(32'hbb537e10),
	.w3(32'h3c38397e),
	.w4(32'hbba4c2af),
	.w5(32'hba013439),
	.w6(32'h3c449f30),
	.w7(32'hbaa812fe),
	.w8(32'h3c2a07cf),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c2129),
	.w1(32'h3a8dd0d0),
	.w2(32'h3beea980),
	.w3(32'h3c1a12b6),
	.w4(32'h3ae0b853),
	.w5(32'hbbdf1f39),
	.w6(32'h3c18c652),
	.w7(32'hbb28eb15),
	.w8(32'hbc0ad410),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba78f65),
	.w1(32'h3b966de6),
	.w2(32'h3a0a37f5),
	.w3(32'h3bf81d34),
	.w4(32'h3b90f517),
	.w5(32'hbb6bf772),
	.w6(32'h3c851feb),
	.w7(32'h3b48eb9f),
	.w8(32'h3ac89881),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03bf1e),
	.w1(32'hbb529dd6),
	.w2(32'hbbf4af45),
	.w3(32'hba192184),
	.w4(32'hbb97bf88),
	.w5(32'hbc6a544c),
	.w6(32'hbb12e0bb),
	.w7(32'hbbe512b8),
	.w8(32'hbb121efa),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafeae54),
	.w1(32'h3bbc7daf),
	.w2(32'h3c2a4b91),
	.w3(32'h3b591476),
	.w4(32'h3c3b802b),
	.w5(32'h3c665a2c),
	.w6(32'hbba29a56),
	.w7(32'h3c475314),
	.w8(32'h3c23f00e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ffaf9f),
	.w1(32'hba44bedb),
	.w2(32'h3bbc0aa4),
	.w3(32'h3b396a0c),
	.w4(32'h3ac1fcb4),
	.w5(32'h3c08ef32),
	.w6(32'h3c0bbaf3),
	.w7(32'h3bd54c49),
	.w8(32'hbb9e5e8d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe1b63),
	.w1(32'hbb3cd467),
	.w2(32'hbbec6fb0),
	.w3(32'hbb1ac3d2),
	.w4(32'h3a8908dd),
	.w5(32'hbb420f6e),
	.w6(32'h3b108077),
	.w7(32'hbadf60c8),
	.w8(32'hbb140f31),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc147dd6),
	.w1(32'hbbcaac8c),
	.w2(32'hbc24ef32),
	.w3(32'hbc13ee8f),
	.w4(32'hbbb74997),
	.w5(32'hbc4b9e24),
	.w6(32'hbb0aa7a3),
	.w7(32'hbb20f0e7),
	.w8(32'hbb8e2b23),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba288dd),
	.w1(32'hbc430924),
	.w2(32'hbc1d5059),
	.w3(32'h3c81bdba),
	.w4(32'hbc0c6b8b),
	.w5(32'hbc2f8214),
	.w6(32'h3c21cc6e),
	.w7(32'hbc51304d),
	.w8(32'hbc3a97bb),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e10d7),
	.w1(32'h3bad1156),
	.w2(32'hbb6d4184),
	.w3(32'h39d9721e),
	.w4(32'h3b0884aa),
	.w5(32'hbc020d3c),
	.w6(32'hb91df5c7),
	.w7(32'h3a38ae2a),
	.w8(32'hb8d4f44e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6098a9),
	.w1(32'h39dfdc50),
	.w2(32'hb90dd862),
	.w3(32'hbb2a55ac),
	.w4(32'h3c144891),
	.w5(32'h3beaaa08),
	.w6(32'h3be7318c),
	.w7(32'h3c7f9676),
	.w8(32'h3c814bdb),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a9383),
	.w1(32'hbb102190),
	.w2(32'hbbbbbde0),
	.w3(32'h3bbe3b55),
	.w4(32'h39fc70e0),
	.w5(32'h3b04855d),
	.w6(32'h3bd810dd),
	.w7(32'hbaa30b10),
	.w8(32'hbb9e4f9c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f3eb0),
	.w1(32'h3b4d354f),
	.w2(32'hbb9d39c1),
	.w3(32'h395f0521),
	.w4(32'hb603af6e),
	.w5(32'hbc704a14),
	.w6(32'h3bd846bb),
	.w7(32'hbbfb69c4),
	.w8(32'h3bbf5a3d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61e57f),
	.w1(32'hbc562963),
	.w2(32'hbc195219),
	.w3(32'hbbc06d58),
	.w4(32'h3b6c6d36),
	.w5(32'h3c30ab72),
	.w6(32'h3a1f1a74),
	.w7(32'hbb5bd958),
	.w8(32'hba6e3e87),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8fb8f),
	.w1(32'h3aad64b5),
	.w2(32'h3af4b84f),
	.w3(32'hbbbfd8e5),
	.w4(32'h3b57c48f),
	.w5(32'hba8874c1),
	.w6(32'hbc447326),
	.w7(32'h3a74106f),
	.w8(32'hb9d8b7b7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcafdfb),
	.w1(32'hbbb0129f),
	.w2(32'hbc480310),
	.w3(32'hbb3a0c49),
	.w4(32'h3b738bce),
	.w5(32'hbc2fb07f),
	.w6(32'hbbfe5195),
	.w7(32'h3bb87a98),
	.w8(32'hba6a2524),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3838b656),
	.w1(32'h3b8cdaec),
	.w2(32'hbbbbb710),
	.w3(32'h3ba60c27),
	.w4(32'h3c0e2cdb),
	.w5(32'hb8bd88cf),
	.w6(32'h3bf1bfb0),
	.w7(32'h3c4a2a5f),
	.w8(32'h3bf6d835),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f8ab3),
	.w1(32'hb9d6647d),
	.w2(32'hbc7cfb16),
	.w3(32'h3ba598c7),
	.w4(32'hba8999c9),
	.w5(32'hbc88d4c8),
	.w6(32'hbbbeabd9),
	.w7(32'h3be0dbec),
	.w8(32'hbb76ca85),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b3da6),
	.w1(32'h3b9e7473),
	.w2(32'h3c2d42de),
	.w3(32'hbc36970e),
	.w4(32'h3c1ff06d),
	.w5(32'h3bce790e),
	.w6(32'hbb1253fa),
	.w7(32'h3c325feb),
	.w8(32'h3bac9620),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc133152),
	.w1(32'hbb302fce),
	.w2(32'hbc007221),
	.w3(32'hbbe7edeb),
	.w4(32'hba8be519),
	.w5(32'h3b17448b),
	.w6(32'hbb323283),
	.w7(32'hb97b1769),
	.w8(32'hbb19dce5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae831f2),
	.w1(32'hbb06df47),
	.w2(32'h3ab133f3),
	.w3(32'hb9e52027),
	.w4(32'h3bab56a8),
	.w5(32'h3977900b),
	.w6(32'h3b99de1a),
	.w7(32'h3bc3aff1),
	.w8(32'h396129e6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bbf5d),
	.w1(32'hbc06acc5),
	.w2(32'hbbcee829),
	.w3(32'hbaa66529),
	.w4(32'hbc3e4ae4),
	.w5(32'hbc56f544),
	.w6(32'hbba31fd6),
	.w7(32'hbc3f2985),
	.w8(32'hbbe7bf70),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11729c),
	.w1(32'hbc86965a),
	.w2(32'hbc2d49be),
	.w3(32'h3b14021a),
	.w4(32'h3b8f3eaf),
	.w5(32'hba96669b),
	.w6(32'hbc0dac08),
	.w7(32'hbb655f7a),
	.w8(32'h3c4bc039),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeac54e),
	.w1(32'hbadb7fab),
	.w2(32'hbba962eb),
	.w3(32'h3c6b3206),
	.w4(32'h3a27ba69),
	.w5(32'hbbd91d8b),
	.w6(32'h3c86b1e2),
	.w7(32'h3bae808c),
	.w8(32'h3b7ceac7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a3d9c),
	.w1(32'hbc24a211),
	.w2(32'hbb1f5498),
	.w3(32'h3b97854a),
	.w4(32'hbc261413),
	.w5(32'hbbb03763),
	.w6(32'h3be29471),
	.w7(32'hbbdd330d),
	.w8(32'hbb091d8c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6ca5f),
	.w1(32'hbb9fe689),
	.w2(32'hbc23fcb0),
	.w3(32'h3c755b20),
	.w4(32'hbbd695b5),
	.w5(32'hbc006205),
	.w6(32'h3c5dd500),
	.w7(32'hbb7d2ec5),
	.w8(32'hbb28a9ac),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd4863),
	.w1(32'hbb0a24c5),
	.w2(32'hbc1cd92b),
	.w3(32'hbbd60912),
	.w4(32'h3ba98dd6),
	.w5(32'hbbcf5ef9),
	.w6(32'hbc338962),
	.w7(32'hba77eb02),
	.w8(32'hbb06ac31),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e77a9),
	.w1(32'hbc25a3b8),
	.w2(32'hbc1368a6),
	.w3(32'hbbd91157),
	.w4(32'hb8fcd766),
	.w5(32'h3af6b7a9),
	.w6(32'hbb85ade7),
	.w7(32'hbb996b2e),
	.w8(32'h3c8905c9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca199f),
	.w1(32'hbb43470f),
	.w2(32'hbc5fdb26),
	.w3(32'hbbb5a498),
	.w4(32'hbb467e12),
	.w5(32'hbc4b1957),
	.w6(32'hbae12ed5),
	.w7(32'h3aad52c7),
	.w8(32'h3c3fea49),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe60ec),
	.w1(32'h3a93146f),
	.w2(32'hbb876419),
	.w3(32'h3b0b8972),
	.w4(32'h3b084303),
	.w5(32'hbc21106c),
	.w6(32'h3c3891e4),
	.w7(32'h3a9982cc),
	.w8(32'hba8bf6f0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959a5ad),
	.w1(32'h3bc80129),
	.w2(32'h3b873092),
	.w3(32'h3ba0292c),
	.w4(32'h3c049def),
	.w5(32'h3bcc8b5e),
	.w6(32'h3b2fe270),
	.w7(32'h3acdf5ab),
	.w8(32'hbbee1465),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc257a07),
	.w1(32'hbc3c7d91),
	.w2(32'hbbcc05d1),
	.w3(32'hbc60c229),
	.w4(32'hbc45604f),
	.w5(32'hbb990ef9),
	.w6(32'hbc9a67aa),
	.w7(32'hbc0406be),
	.w8(32'h3abc7fd4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc08564),
	.w1(32'hbb20f5eb),
	.w2(32'hbb61266e),
	.w3(32'h3ad0a343),
	.w4(32'h3a7169c3),
	.w5(32'h3b4abf44),
	.w6(32'h3bde3aaa),
	.w7(32'h3b659310),
	.w8(32'h3b350f55),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b685fa5),
	.w1(32'hbb0f0bda),
	.w2(32'h3ad1aada),
	.w3(32'hbae27e74),
	.w4(32'hbb3cf176),
	.w5(32'hbb24a592),
	.w6(32'hbb684075),
	.w7(32'hba5af2c9),
	.w8(32'h3992bda3),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b152156),
	.w1(32'hbaaa7e6f),
	.w2(32'hba51b8e9),
	.w3(32'h3b9026ff),
	.w4(32'hb9a25af7),
	.w5(32'h3af84201),
	.w6(32'h3b023088),
	.w7(32'h3b5b45b0),
	.w8(32'h3abbd774),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba220688),
	.w1(32'hbbd23bbe),
	.w2(32'hbb4d2e09),
	.w3(32'hbbfb0d6b),
	.w4(32'hbb9c5d33),
	.w5(32'h3b518e8c),
	.w6(32'hbc5b21c0),
	.w7(32'hbbc53a37),
	.w8(32'h3b2464b2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0edbf2),
	.w1(32'hb78e4b59),
	.w2(32'h3af80756),
	.w3(32'h3b93f671),
	.w4(32'h3bb4b042),
	.w5(32'h3c477397),
	.w6(32'h3bbccc46),
	.w7(32'hba5a0c8a),
	.w8(32'h3b9a298a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba068a5),
	.w1(32'hbc51980d),
	.w2(32'hbc1f7718),
	.w3(32'h3bbce740),
	.w4(32'hbbed1895),
	.w5(32'hbc3761c6),
	.w6(32'hba9d6e84),
	.w7(32'hbb414ef7),
	.w8(32'hbb251291),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64a473),
	.w1(32'hbb7baed8),
	.w2(32'hba84f7ec),
	.w3(32'h3a558953),
	.w4(32'hbba43651),
	.w5(32'h39b9d35b),
	.w6(32'hbae0841f),
	.w7(32'hbbab1e56),
	.w8(32'hbbdd0213),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8886d4),
	.w1(32'hbb7465a2),
	.w2(32'h39766347),
	.w3(32'h3a4f629f),
	.w4(32'h3a73fb52),
	.w5(32'hbad973ef),
	.w6(32'h3b5a3291),
	.w7(32'hbb16b4b6),
	.w8(32'hbc674429),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb2198),
	.w1(32'hb9cf179f),
	.w2(32'h3a93ba12),
	.w3(32'hbc5fedf8),
	.w4(32'hbb95b2c4),
	.w5(32'h3b066e45),
	.w6(32'hbc05ace2),
	.w7(32'hb9bf6e95),
	.w8(32'hba95e664),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad362cc),
	.w1(32'h3c749ace),
	.w2(32'hb98e7eec),
	.w3(32'hb9dc5d9b),
	.w4(32'h3c36055f),
	.w5(32'h3c21e7e5),
	.w6(32'h3b43e206),
	.w7(32'h3c632666),
	.w8(32'h3a9f5273),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3731d),
	.w1(32'h3c007502),
	.w2(32'h3bb03ca7),
	.w3(32'hbcd8a2bf),
	.w4(32'h3bd68ff9),
	.w5(32'h3ac21418),
	.w6(32'hbcb3e3e3),
	.w7(32'h3acafe45),
	.w8(32'h3b38b745),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bdb5d),
	.w1(32'hbc19e2f5),
	.w2(32'hbbca9e09),
	.w3(32'h3b7349e2),
	.w4(32'hbbdf3b19),
	.w5(32'hbc3acc5f),
	.w6(32'hbc13061a),
	.w7(32'hbc097408),
	.w8(32'h394980c4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0655db),
	.w1(32'hbb2a8d3c),
	.w2(32'hbb9d9837),
	.w3(32'h3c018bb3),
	.w4(32'h3b2a9bae),
	.w5(32'hbb5bcb0f),
	.w6(32'h3c066368),
	.w7(32'hba5c2a09),
	.w8(32'hba22987f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47b585),
	.w1(32'hba1a8dff),
	.w2(32'hbae4c893),
	.w3(32'hba89b2ec),
	.w4(32'h3ad83741),
	.w5(32'hbbf5e789),
	.w6(32'hbba54233),
	.w7(32'h3a8c426a),
	.w8(32'hbbbaf4bf),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc142037),
	.w1(32'h3b2f204c),
	.w2(32'hbc0750db),
	.w3(32'hbbb19926),
	.w4(32'h3c00a9dd),
	.w5(32'h3af66a5d),
	.w6(32'hb861a18e),
	.w7(32'h3b9f16a4),
	.w8(32'h3b809c1b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7f952),
	.w1(32'hbbf7fbec),
	.w2(32'hbc0769c8),
	.w3(32'hbbd3cc82),
	.w4(32'hbba95531),
	.w5(32'hbc295f29),
	.w6(32'hbb040b09),
	.w7(32'hbba951c9),
	.w8(32'hbb83efcc),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec22f9),
	.w1(32'hbbfe1d23),
	.w2(32'hbae5acaf),
	.w3(32'h3b3c59c7),
	.w4(32'hbbf5f72d),
	.w5(32'hbb51a448),
	.w6(32'h3b046b02),
	.w7(32'hbbf828bf),
	.w8(32'hbbe8d4ed),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc819958),
	.w1(32'h3bd3fac5),
	.w2(32'h3c4f0c58),
	.w3(32'hbc76ddf0),
	.w4(32'h3c1fc02c),
	.w5(32'h3c1b1283),
	.w6(32'hbc32de36),
	.w7(32'h3c0f049d),
	.w8(32'h3c630459),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3afb2d),
	.w1(32'h3b773218),
	.w2(32'hbb6c7d98),
	.w3(32'h3c8c5f2a),
	.w4(32'h3ba1172e),
	.w5(32'h3b169eb8),
	.w6(32'h3c1da054),
	.w7(32'h3b3c5d0a),
	.w8(32'h3b0c29d7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb825fdc),
	.w1(32'hbba8f2cc),
	.w2(32'hbba85f9d),
	.w3(32'hbc07ef68),
	.w4(32'hbb601ae9),
	.w5(32'h3afb322a),
	.w6(32'hbc1698d6),
	.w7(32'h3a9802ba),
	.w8(32'h3b38cef0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cc633),
	.w1(32'hbbd3f565),
	.w2(32'hbb738349),
	.w3(32'hb9576b89),
	.w4(32'h3bfa7cf2),
	.w5(32'h3beeb15e),
	.w6(32'h3b14d8c4),
	.w7(32'h3ac1bbe9),
	.w8(32'hbba76738),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd16d58),
	.w1(32'h3a4fa526),
	.w2(32'hb98cee3b),
	.w3(32'h3a837918),
	.w4(32'h3acb32f8),
	.w5(32'h3b48bd99),
	.w6(32'hbb1acc2b),
	.w7(32'hbc2526ce),
	.w8(32'hbc774227),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eb8ab),
	.w1(32'h39cff0ae),
	.w2(32'hbb8b3338),
	.w3(32'h3ae00337),
	.w4(32'h3b2715e3),
	.w5(32'hb81140ec),
	.w6(32'hbb70713d),
	.w7(32'h3b940930),
	.w8(32'h3bc4031b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0b63f),
	.w1(32'h3b630f90),
	.w2(32'hbae43658),
	.w3(32'hbb40a236),
	.w4(32'h3c41fa02),
	.w5(32'hbb0b11ae),
	.w6(32'h3b5487f6),
	.w7(32'h3b98d845),
	.w8(32'h38f73844),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baca9da),
	.w1(32'hbb97c826),
	.w2(32'hbbe8577c),
	.w3(32'h3bf4d46b),
	.w4(32'hbb4a4854),
	.w5(32'hbb2d22a1),
	.w6(32'hbbdbe053),
	.w7(32'hbc1a9ae7),
	.w8(32'hba9dfa95),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc48df7),
	.w1(32'hbbc36858),
	.w2(32'hbc168cd5),
	.w3(32'hbbea08d6),
	.w4(32'hbbdcca67),
	.w5(32'hbbb8a2b1),
	.w6(32'hbc2b8988),
	.w7(32'h3987ad34),
	.w8(32'hbb33c12b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20cc47),
	.w1(32'hbc9a917e),
	.w2(32'hbc2e1714),
	.w3(32'h3c5c1e4a),
	.w4(32'hbc5a8576),
	.w5(32'hbc7af3ef),
	.w6(32'h3cabaeca),
	.w7(32'hbc04821d),
	.w8(32'hbbafb07c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb24e98),
	.w1(32'h3acfc41c),
	.w2(32'hbbb6a681),
	.w3(32'h3cd6d901),
	.w4(32'h3b72512d),
	.w5(32'hbbebc40a),
	.w6(32'h3cb47723),
	.w7(32'h3c19cab5),
	.w8(32'h3c1d9458),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac08278),
	.w1(32'h3b93441c),
	.w2(32'h3b92f8cb),
	.w3(32'hbb88cf9e),
	.w4(32'h3bf2c1e7),
	.w5(32'h3c005b62),
	.w6(32'hbaf13217),
	.w7(32'h3b1e30ec),
	.w8(32'h3be2b56e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accab78),
	.w1(32'hbbd12fc1),
	.w2(32'hbbbc1f9d),
	.w3(32'hba484609),
	.w4(32'hbc1b919a),
	.w5(32'hbb9a4c12),
	.w6(32'h395db235),
	.w7(32'hbbe5f970),
	.w8(32'hbbcdae4a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb060b),
	.w1(32'h3bdd8337),
	.w2(32'h3b1b38c6),
	.w3(32'h3baf0a80),
	.w4(32'h3bf5d2ab),
	.w5(32'h3b93c610),
	.w6(32'h3bd6f695),
	.w7(32'h3b42bb88),
	.w8(32'h37aab0e1),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f6072),
	.w1(32'h3b2b090c),
	.w2(32'hbb879c0a),
	.w3(32'hb98e5d29),
	.w4(32'h3bd75983),
	.w5(32'h3af59108),
	.w6(32'hbb1822fa),
	.w7(32'h38afc7f9),
	.w8(32'hbbad6d27),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5dcbd0),
	.w1(32'h3ad0bfb6),
	.w2(32'hbb5d2c0b),
	.w3(32'hbc66cc55),
	.w4(32'h3ba6d5d6),
	.w5(32'hba5bd8fd),
	.w6(32'hbc6a4625),
	.w7(32'h3b8dfdd3),
	.w8(32'hbad284ec),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90c997),
	.w1(32'hbbd172ea),
	.w2(32'hbc140b74),
	.w3(32'hbca99c1a),
	.w4(32'hbba7917a),
	.w5(32'hbc3ca2ba),
	.w6(32'hbc449ba7),
	.w7(32'hba9f2e9e),
	.w8(32'hbbc94b59),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0b9f1),
	.w1(32'h39e2e43c),
	.w2(32'h3bc71933),
	.w3(32'h3bbda598),
	.w4(32'hbaa876e7),
	.w5(32'h3c17ef77),
	.w6(32'h3b9d2982),
	.w7(32'h3b118c57),
	.w8(32'h3bcac119),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f872c),
	.w1(32'hbbe3c183),
	.w2(32'hbc11824c),
	.w3(32'h3c175af8),
	.w4(32'hbb91a8c8),
	.w5(32'hbb8d9c76),
	.w6(32'h3bc9b6af),
	.w7(32'hbaa01de2),
	.w8(32'hbb96a55f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c02ee),
	.w1(32'h3a3d2aae),
	.w2(32'hbb6a220f),
	.w3(32'h3bbd2183),
	.w4(32'h3b73516d),
	.w5(32'hbc10c16c),
	.w6(32'hbae7b22c),
	.w7(32'h3b3369c5),
	.w8(32'hbb19eb0f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb984d6d),
	.w1(32'hbb911087),
	.w2(32'hbba85689),
	.w3(32'hbb8ae9fb),
	.w4(32'h3a2d185f),
	.w5(32'h39ad2b4f),
	.w6(32'h3b9d344a),
	.w7(32'hbb9d776a),
	.w8(32'hbaff1132),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6de3c),
	.w1(32'h3b7730be),
	.w2(32'hbad1bac1),
	.w3(32'h3ac6675b),
	.w4(32'h3befe0a1),
	.w5(32'h3a9bc104),
	.w6(32'hbc10685d),
	.w7(32'h3bb30c67),
	.w8(32'h3bddf988),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb414d54),
	.w1(32'h3bdd2c5b),
	.w2(32'h3c10cd36),
	.w3(32'hbbb116f1),
	.w4(32'h3c0336a3),
	.w5(32'h3c7709e6),
	.w6(32'h3ab3ee4e),
	.w7(32'h3b896ca9),
	.w8(32'h3bf85c2a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbeb640),
	.w1(32'hbb947bb6),
	.w2(32'h3c40c4b9),
	.w3(32'h3bd1bf63),
	.w4(32'h3b8f2603),
	.w5(32'h3c8b06c0),
	.w6(32'h3b3faf1b),
	.w7(32'h3bd49b91),
	.w8(32'h3bb4904b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb992d44),
	.w1(32'hbbcacb9c),
	.w2(32'hbba1bca2),
	.w3(32'h38e61402),
	.w4(32'hba1a8658),
	.w5(32'hbb2b3528),
	.w6(32'hbaeea86b),
	.w7(32'hbab4b99a),
	.w8(32'hbb4b2e25),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdf8cd),
	.w1(32'hbb71b193),
	.w2(32'h3bfa5408),
	.w3(32'hbb426242),
	.w4(32'hba47ceb5),
	.w5(32'h3b912dd3),
	.w6(32'h3b57f310),
	.w7(32'h3bcab001),
	.w8(32'h3b6157f6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba665d2),
	.w1(32'hbb528226),
	.w2(32'hbb37deab),
	.w3(32'hbbb987d8),
	.w4(32'hbbcdef53),
	.w5(32'hbb655592),
	.w6(32'hbbfbb60d),
	.w7(32'h3b6a78e5),
	.w8(32'h39957905),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3425ba),
	.w1(32'hbb6c132d),
	.w2(32'hbb2b0f4e),
	.w3(32'h3ca22f26),
	.w4(32'hbbcd3209),
	.w5(32'hbad13cc5),
	.w6(32'h3cc901e7),
	.w7(32'hbb1bcdc9),
	.w8(32'hbbce4ead),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b127adf),
	.w1(32'hbc32af08),
	.w2(32'h3a4ebd89),
	.w3(32'h3b9b1917),
	.w4(32'hbc2e83dc),
	.w5(32'hbb079aa4),
	.w6(32'hbbdcfceb),
	.w7(32'hbabab5b5),
	.w8(32'hb8e3a0fc),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72b1b8),
	.w1(32'hbab80706),
	.w2(32'h3b7a6a63),
	.w3(32'h3cb74b52),
	.w4(32'hbb587bae),
	.w5(32'hb8bf345c),
	.w6(32'h3c69012e),
	.w7(32'hbb67126a),
	.w8(32'hbbf4aa94),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addee94),
	.w1(32'hbaf1e22d),
	.w2(32'hbb993b53),
	.w3(32'h3ba5d7ad),
	.w4(32'h3ae390b1),
	.w5(32'hba21ffc9),
	.w6(32'hbb584152),
	.w7(32'hbad39388),
	.w8(32'hbbb8e662),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce7434),
	.w1(32'hbb36c21e),
	.w2(32'hbc0c4a37),
	.w3(32'h39b50526),
	.w4(32'hba9f586c),
	.w5(32'hbb84fdd7),
	.w6(32'hbbc25ead),
	.w7(32'h3bba1ebe),
	.w8(32'hbb1a1b5f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32e3cf),
	.w1(32'hbbdce28a),
	.w2(32'hbb3bd5da),
	.w3(32'hbb810a93),
	.w4(32'hbb950615),
	.w5(32'h3a43c6d1),
	.w6(32'hbc1fe500),
	.w7(32'hbb3b6de9),
	.w8(32'hbaac01e5),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6cb9c),
	.w1(32'hbc743de6),
	.w2(32'hbc290ba2),
	.w3(32'hbb47d725),
	.w4(32'hbc805efa),
	.w5(32'hbc331800),
	.w6(32'hbbbec70a),
	.w7(32'hbc1445bf),
	.w8(32'hbb294721),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc141728),
	.w1(32'hbc294e4a),
	.w2(32'hbbd10539),
	.w3(32'hbc700193),
	.w4(32'hbc1f1e23),
	.w5(32'hbbc309a0),
	.w6(32'hbc440287),
	.w7(32'hbbbd4262),
	.w8(32'hbb4e2ac7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b005b91),
	.w1(32'hbabc68a5),
	.w2(32'hbbc8b6e5),
	.w3(32'h3ca35593),
	.w4(32'h3b9bf53e),
	.w5(32'h3bb56afa),
	.w6(32'h3c614c95),
	.w7(32'h3a5ca2ec),
	.w8(32'h3be0877c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc379a70),
	.w1(32'h3bb8f9b1),
	.w2(32'h3bdc8c3c),
	.w3(32'hbc6ffd85),
	.w4(32'h3c0ff48e),
	.w5(32'h3be50110),
	.w6(32'hbc4d2df9),
	.w7(32'h3bfbf2a2),
	.w8(32'h3bcc693b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44f958),
	.w1(32'hbc1b1ff3),
	.w2(32'hbc6f5e80),
	.w3(32'h3ba9426c),
	.w4(32'hbb21c15f),
	.w5(32'hbc376f26),
	.w6(32'h3c14aaca),
	.w7(32'hba60c4d4),
	.w8(32'h3acfc5b7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeed38b),
	.w1(32'hbb70e36f),
	.w2(32'h3b9e492e),
	.w3(32'h3a471ca5),
	.w4(32'hba55cba9),
	.w5(32'h3c31732b),
	.w6(32'h3b9eecf6),
	.w7(32'h3b82cc37),
	.w8(32'h3be669e1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadd682),
	.w1(32'hbbebb7cf),
	.w2(32'h3b0a754e),
	.w3(32'hbac362a3),
	.w4(32'hba7aa221),
	.w5(32'h3b80ddcb),
	.w6(32'h3abc9351),
	.w7(32'h3bd9e500),
	.w8(32'h3c4fa3b5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5cd6a3),
	.w1(32'hbb89fb7c),
	.w2(32'hbb670600),
	.w3(32'h3cce089d),
	.w4(32'h3a835e1e),
	.w5(32'hba162fa5),
	.w6(32'h3c8e4df0),
	.w7(32'hbbc84696),
	.w8(32'hbba58dcb),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca15892),
	.w1(32'hbb3b7aa9),
	.w2(32'hbc5bfa5c),
	.w3(32'hbca65144),
	.w4(32'h3a9ce735),
	.w5(32'hbbd8a662),
	.w6(32'hbc65338a),
	.w7(32'h3af0ea8b),
	.w8(32'hbbea6221),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe296a8),
	.w1(32'hbbdd958d),
	.w2(32'hbc2133cc),
	.w3(32'hb9352a10),
	.w4(32'hbb886cab),
	.w5(32'hbbc7a3f6),
	.w6(32'h3b670745),
	.w7(32'hba157972),
	.w8(32'hba6103b6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6cb866),
	.w1(32'hbba7b2da),
	.w2(32'hbbc7b986),
	.w3(32'h3c52632a),
	.w4(32'hbae2d302),
	.w5(32'hbbd1b2c4),
	.w6(32'h3c4edc07),
	.w7(32'h3a8ce13c),
	.w8(32'h3c7bc11b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9737c),
	.w1(32'hbc2c3e03),
	.w2(32'hbb877c90),
	.w3(32'h3bc8f3f2),
	.w4(32'hbbe7b451),
	.w5(32'hba8f43db),
	.w6(32'h3c92513a),
	.w7(32'hbc469f38),
	.w8(32'h3aad0836),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912fdf4),
	.w1(32'h3c5b90dd),
	.w2(32'hbaf6609a),
	.w3(32'h3bcb31ab),
	.w4(32'h3c975280),
	.w5(32'h3c113ce4),
	.w6(32'h3bcb9435),
	.w7(32'h3ca58e43),
	.w8(32'h3c188c0b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc579571),
	.w1(32'hbb8f1cfc),
	.w2(32'h3b4abdf0),
	.w3(32'hbc90f052),
	.w4(32'hbbb66bfb),
	.w5(32'h3c117b85),
	.w6(32'hbc89bc94),
	.w7(32'h3be2838a),
	.w8(32'h3bbfeb59),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1f4c9),
	.w1(32'h39d5707f),
	.w2(32'hbb55acab),
	.w3(32'h3c0df6fd),
	.w4(32'hbb48edd9),
	.w5(32'hbbc46358),
	.w6(32'h3c3ccd73),
	.w7(32'hbbd5e6d8),
	.w8(32'hbb2cb863),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b5add),
	.w1(32'hbb33d97a),
	.w2(32'h3c375a5b),
	.w3(32'hbc46c4ff),
	.w4(32'hbb9f9df4),
	.w5(32'h3c545de8),
	.w6(32'hbc5c7aae),
	.w7(32'hbc39abeb),
	.w8(32'h3c5c21b6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67bded),
	.w1(32'h3b86cf94),
	.w2(32'hbb95bbef),
	.w3(32'h3bbc963a),
	.w4(32'h3ba74656),
	.w5(32'h3b7e477e),
	.w6(32'h3bd9ddbf),
	.w7(32'h3b4ca5b3),
	.w8(32'hbc304466),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9472050),
	.w1(32'hbaa99fa0),
	.w2(32'h3bb8c4a7),
	.w3(32'hbbad8c68),
	.w4(32'hbb662ae8),
	.w5(32'h3b93fdb0),
	.w6(32'hbc8e5073),
	.w7(32'hbb97c121),
	.w8(32'hbc00d969),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50c166),
	.w1(32'h3c1a07b3),
	.w2(32'h3915c321),
	.w3(32'h3ba91ebc),
	.w4(32'h3bf173e1),
	.w5(32'h3b21f00e),
	.w6(32'h3a17987b),
	.w7(32'h3c0e5e6a),
	.w8(32'h3bd3018a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc7fad),
	.w1(32'hbc025239),
	.w2(32'hbb9e432d),
	.w3(32'h3b4513d0),
	.w4(32'hbbb5d61c),
	.w5(32'hbc4d0c8b),
	.w6(32'hb95b2310),
	.w7(32'hbb434ed1),
	.w8(32'hbc1af242),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03d56b),
	.w1(32'hba3ebef8),
	.w2(32'hbba1f3e5),
	.w3(32'hba4ed768),
	.w4(32'hbad94fc3),
	.w5(32'hb9f6cf2a),
	.w6(32'hbba908d5),
	.w7(32'hbb781097),
	.w8(32'hbada4c60),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac6823),
	.w1(32'h3a9289c5),
	.w2(32'hba22053f),
	.w3(32'h3b5a73a5),
	.w4(32'h3b655174),
	.w5(32'hbbb46f29),
	.w6(32'h3b8eed6f),
	.w7(32'h3bfd9ae2),
	.w8(32'hbbbb4864),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92fa3f),
	.w1(32'hbb3554af),
	.w2(32'h3baf3479),
	.w3(32'hb76452da),
	.w4(32'hbbc972bc),
	.w5(32'h3be606fb),
	.w6(32'hbbc1fc5d),
	.w7(32'hbbd99910),
	.w8(32'h3b652890),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0cb51f),
	.w1(32'hbbfca6c1),
	.w2(32'hbcce9b68),
	.w3(32'hbcd6fb40),
	.w4(32'hbb7e4bf1),
	.w5(32'hbc6fbc76),
	.w6(32'hbc9cd18d),
	.w7(32'h3a9f1d93),
	.w8(32'h3a09b3ad),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ec17a),
	.w1(32'h3bebff14),
	.w2(32'hbabdfd23),
	.w3(32'hbc0a5ded),
	.w4(32'h3c85b308),
	.w5(32'h3b8358d3),
	.w6(32'h3a26588c),
	.w7(32'h3c8ae4ce),
	.w8(32'h3c6a53e1),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c030640),
	.w1(32'h3afb3e06),
	.w2(32'h3a1cd026),
	.w3(32'h3bdf2d7a),
	.w4(32'h3bb0511c),
	.w5(32'h3b871e88),
	.w6(32'h3c0c35fd),
	.w7(32'h3ac3b180),
	.w8(32'h3b672088),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a00a5),
	.w1(32'h3b0003b1),
	.w2(32'h3c521343),
	.w3(32'hbbe7d1f1),
	.w4(32'h3be30ac7),
	.w5(32'h3c4c9490),
	.w6(32'hbbc27024),
	.w7(32'h3b67160b),
	.w8(32'h3bcfbd1e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b56bd),
	.w1(32'h39962fae),
	.w2(32'h3b23282c),
	.w3(32'hbb3f409b),
	.w4(32'hbb33bf01),
	.w5(32'h3aa26a45),
	.w6(32'hbba54f03),
	.w7(32'hb9870b6f),
	.w8(32'h3b8342a6),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf44782),
	.w1(32'hbb2349b5),
	.w2(32'h3b0a6b9c),
	.w3(32'h3b8b98eb),
	.w4(32'h3a5d50f5),
	.w5(32'h3b07ce90),
	.w6(32'h3c2679bf),
	.w7(32'h3ae3d53c),
	.w8(32'h3ba7f132),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b996e04),
	.w1(32'h3c40accc),
	.w2(32'hba4746d3),
	.w3(32'h3c346abc),
	.w4(32'h3c55c217),
	.w5(32'h3c25cf80),
	.w6(32'h3c6f89f7),
	.w7(32'h3c7f78a8),
	.w8(32'hba9e0881),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b9a34),
	.w1(32'hbb54fb89),
	.w2(32'hbc30ecd8),
	.w3(32'hbcd407a2),
	.w4(32'hbb1a390e),
	.w5(32'hbc48ccde),
	.w6(32'hbcbc570b),
	.w7(32'hbb2f094e),
	.w8(32'hbb9ca2e9),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e2373),
	.w1(32'hbc81aa3a),
	.w2(32'hbc56f1ed),
	.w3(32'hbb9887ae),
	.w4(32'hba078090),
	.w5(32'hbc14096d),
	.w6(32'hbae2d0da),
	.w7(32'hb9667db0),
	.w8(32'hbb3e6e3a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaff530),
	.w1(32'hbaa521e2),
	.w2(32'h3c0e530d),
	.w3(32'hbb119371),
	.w4(32'hb9576e4e),
	.w5(32'h3c57edc7),
	.w6(32'hbb77d25d),
	.w7(32'hbbac45c4),
	.w8(32'h3c189d6f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf424ff),
	.w1(32'hbbe8276d),
	.w2(32'hbc1c11ae),
	.w3(32'hbb80f123),
	.w4(32'hbb5e3c1f),
	.w5(32'hbb9d19a4),
	.w6(32'hbc06aeb4),
	.w7(32'hbb28607b),
	.w8(32'hbb2dad5c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e040d),
	.w1(32'hbaa5f7a2),
	.w2(32'hbb1712fb),
	.w3(32'hba7b80cf),
	.w4(32'hba522ebf),
	.w5(32'hbac87e62),
	.w6(32'hbabaf178),
	.w7(32'hba330fc7),
	.w8(32'hbaafbaa3),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba32e2),
	.w1(32'h3829d5de),
	.w2(32'h389fcfb0),
	.w3(32'h38430e33),
	.w4(32'hb61275b5),
	.w5(32'h38182199),
	.w6(32'h3857fbe7),
	.w7(32'h35e43cb1),
	.w8(32'h38162364),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeefb70),
	.w1(32'hba9b61bc),
	.w2(32'hb9b75959),
	.w3(32'hbaa1f9ff),
	.w4(32'hba4f7f93),
	.w5(32'h3903e516),
	.w6(32'hbad0f920),
	.w7(32'hba76da9c),
	.w8(32'hb98f988d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396620ab),
	.w1(32'h38b828bd),
	.w2(32'h3926ca7e),
	.w3(32'h38ee805e),
	.w4(32'hb717ac19),
	.w5(32'h389726ab),
	.w6(32'h3904b98d),
	.w7(32'h35f2ec58),
	.w8(32'h38b66650),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba04f38),
	.w1(32'hba96b2e2),
	.w2(32'hbb146755),
	.w3(32'hbaeeb787),
	.w4(32'h3aec5b73),
	.w5(32'hba1445b5),
	.w6(32'hbac7653c),
	.w7(32'h3a9e27ef),
	.w8(32'hb95ba879),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb743cf),
	.w1(32'h3ab5af54),
	.w2(32'h3af81e66),
	.w3(32'hbb550b23),
	.w4(32'h3bb2ba3c),
	.w5(32'h3b937e0a),
	.w6(32'hbad3b61b),
	.w7(32'h3bdb3233),
	.w8(32'h3b6ae6f7),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f8c52),
	.w1(32'hbad7fda9),
	.w2(32'hbb935e6b),
	.w3(32'hba1c94b6),
	.w4(32'h3a9c85c2),
	.w5(32'hba90db89),
	.w6(32'h3a2de23d),
	.w7(32'h3b1732d7),
	.w8(32'h393be76e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1b38e),
	.w1(32'h39691518),
	.w2(32'h3a961fa6),
	.w3(32'hbabc91ff),
	.w4(32'hb7a51c1b),
	.w5(32'h3a10073e),
	.w6(32'hbabbda1a),
	.w7(32'hb90690c8),
	.w8(32'h39b3bf87),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b83eb),
	.w1(32'hbb40356f),
	.w2(32'hbbc7ae40),
	.w3(32'hbac088d4),
	.w4(32'h39c1cfa7),
	.w5(32'hbaf1c311),
	.w6(32'hba662373),
	.w7(32'h3aa2fb08),
	.w8(32'hbada21d4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b0ed7),
	.w1(32'hbb13d16c),
	.w2(32'hbb93520b),
	.w3(32'hba89ff13),
	.w4(32'hb9b82423),
	.w5(32'hbb179b84),
	.w6(32'hba6c2962),
	.w7(32'hb98a85a3),
	.w8(32'hbaae3c23),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5573eb),
	.w1(32'hbbf2de93),
	.w2(32'hbc242a5f),
	.w3(32'hbc389e15),
	.w4(32'hbb9e1f3d),
	.w5(32'hbbf9dff2),
	.w6(32'hbc12c641),
	.w7(32'hbb1bffa9),
	.w8(32'hbbec0efb),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386998d7),
	.w1(32'hb608a03a),
	.w2(32'h360a56dd),
	.w3(32'h3850ad00),
	.w4(32'hb5a1d84c),
	.w5(32'h3669d6f4),
	.w6(32'h38a47c8d),
	.w7(32'h3729325e),
	.w8(32'h3762689c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38203bb4),
	.w1(32'h382f6f2f),
	.w2(32'h3795fc95),
	.w3(32'h3824265b),
	.w4(32'h37ee1d72),
	.w5(32'hb7ce242c),
	.w6(32'hb797714a),
	.w7(32'h380eaeb4),
	.w8(32'hb72d29d7),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba186db),
	.w1(32'hba91eb2d),
	.w2(32'hbb8a2628),
	.w3(32'hb9dde36e),
	.w4(32'h3ae5c39b),
	.w5(32'hbb13456f),
	.w6(32'hb9a55c1d),
	.w7(32'h3b60b262),
	.w8(32'hba21584b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacccc5),
	.w1(32'hba9c0564),
	.w2(32'hbbe7cc05),
	.w3(32'h39d8e814),
	.w4(32'h3ae3d64b),
	.w5(32'hbb9faa46),
	.w6(32'h3a98d1a9),
	.w7(32'h3b83529f),
	.w8(32'h3a1e24e0),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc87290),
	.w1(32'hbb653ad3),
	.w2(32'hbbf9d14b),
	.w3(32'hbb14926b),
	.w4(32'h3a4f3a48),
	.w5(32'hbb476798),
	.w6(32'hbad0e7d2),
	.w7(32'h3b160a1b),
	.w8(32'hbab24d53),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f1961),
	.w1(32'hba722ca0),
	.w2(32'hba790572),
	.w3(32'h3b0bda3f),
	.w4(32'h3999dbb4),
	.w5(32'h3838dbcc),
	.w6(32'h3b108c18),
	.w7(32'hb712e522),
	.w8(32'hbafb191a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d06dd2),
	.w1(32'h375a20cb),
	.w2(32'h38c777cd),
	.w3(32'h396f54a3),
	.w4(32'hb89f73ef),
	.w5(32'h38dd7972),
	.w6(32'hb75bc4d7),
	.w7(32'hb8c0e937),
	.w8(32'h38c54266),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f73ae8),
	.w1(32'hb9ed2892),
	.w2(32'hb9644420),
	.w3(32'hba10d247),
	.w4(32'hb9eddd33),
	.w5(32'hb92d1189),
	.w6(32'hba1b10e9),
	.w7(32'hb9d3058b),
	.w8(32'hb966ff89),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a25fb6),
	.w1(32'h3aab1e0e),
	.w2(32'hbb0edba4),
	.w3(32'h3b9bac97),
	.w4(32'hba1348c1),
	.w5(32'hbb9505e8),
	.w6(32'h3b45acbd),
	.w7(32'h3a831b36),
	.w8(32'hbad4433b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc279213),
	.w1(32'hbc00b3d6),
	.w2(32'hbc389376),
	.w3(32'hbbd82110),
	.w4(32'hbbca6543),
	.w5(32'hbbc79954),
	.w6(32'hbc03a20e),
	.w7(32'hbb765b0d),
	.w8(32'hbb91e01a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91d5c1),
	.w1(32'hb99e9e27),
	.w2(32'hbb94488e),
	.w3(32'h3b383af4),
	.w4(32'h3b25b6d1),
	.w5(32'hba7920ab),
	.w6(32'h3b3f7f80),
	.w7(32'h3b12c0e5),
	.w8(32'hba8a360d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f5b21),
	.w1(32'h3b17c513),
	.w2(32'h3aac9d73),
	.w3(32'hbb401ccc),
	.w4(32'h3b72774c),
	.w5(32'h3b2469ef),
	.w6(32'hbad24138),
	.w7(32'h3b57f52b),
	.w8(32'h39f76a4a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09e9d8),
	.w1(32'hbbb045af),
	.w2(32'hbbd9fdc6),
	.w3(32'hbbec2e9a),
	.w4(32'hbb1b6b93),
	.w5(32'hbb6b187b),
	.w6(32'hbb667ac1),
	.w7(32'h3a3103f6),
	.w8(32'hba9631be),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38499d9b),
	.w1(32'h37e6978a),
	.w2(32'h3818fdb1),
	.w3(32'h37e73753),
	.w4(32'h37145e46),
	.w5(32'h3797e531),
	.w6(32'h37f6c063),
	.w7(32'h37529006),
	.w8(32'h379a7c7e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3844fbf8),
	.w1(32'h378498f2),
	.w2(32'h38272bec),
	.w3(32'h37be91c5),
	.w4(32'hb72303aa),
	.w5(32'h37335c15),
	.w6(32'h380af3eb),
	.w7(32'hb684d4a8),
	.w8(32'h377ed99a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ed1dd),
	.w1(32'h39d23272),
	.w2(32'h399a9b87),
	.w3(32'h3af571ee),
	.w4(32'h39f2b0f8),
	.w5(32'h39a374aa),
	.w6(32'h38b53ccf),
	.w7(32'hb915884a),
	.w8(32'h3981df63),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3897a992),
	.w1(32'hb62ede71),
	.w2(32'h37ab2bc1),
	.w3(32'h3835d64d),
	.w4(32'hb81d90e7),
	.w5(32'hb6e0555f),
	.w6(32'h38593be6),
	.w7(32'hb8169f7d),
	.w8(32'hb750ab15),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08fae2),
	.w1(32'hb9ae2ad2),
	.w2(32'hb9da2b20),
	.w3(32'h3a192dfc),
	.w4(32'h389db122),
	.w5(32'hba2b57bd),
	.w6(32'h38dd1a5d),
	.w7(32'hb840dbc5),
	.w8(32'hb9da3ca5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb602890),
	.w1(32'hbabc3b87),
	.w2(32'hbbae7782),
	.w3(32'h38cd5961),
	.w4(32'h3a885075),
	.w5(32'hbb3ef92a),
	.w6(32'h39eb2acd),
	.w7(32'h3b097ae0),
	.w8(32'hba18075f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26d24d),
	.w1(32'hbab1f3f1),
	.w2(32'hbb51d732),
	.w3(32'hbac0f995),
	.w4(32'h39d5317d),
	.w5(32'hbaa0b347),
	.w6(32'h3994bcaf),
	.w7(32'h3a8bcf38),
	.w8(32'hb980996b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38626566),
	.w1(32'h384061a5),
	.w2(32'h38354fba),
	.w3(32'h384c1260),
	.w4(32'h382b230a),
	.w5(32'h37d3f6fc),
	.w6(32'h38114f1d),
	.w7(32'h38248a93),
	.w8(32'h380f875e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c315a),
	.w1(32'hbabb273b),
	.w2(32'hbbda17ef),
	.w3(32'h3b08ebe4),
	.w4(32'h3a9b7c65),
	.w5(32'hbb744e7d),
	.w6(32'h3a7c4ae7),
	.w7(32'h3a6b177c),
	.w8(32'hbb95ead1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6629ba),
	.w1(32'hb95dba3b),
	.w2(32'hbb1a90cd),
	.w3(32'h3a8dce90),
	.w4(32'h397f5984),
	.w5(32'hbac40445),
	.w6(32'h39cf445c),
	.w7(32'h3a872d29),
	.w8(32'hba1815a4),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3818e881),
	.w1(32'hb7538d13),
	.w2(32'h380e89dd),
	.w3(32'hb756f6ab),
	.w4(32'hb9355aa3),
	.w5(32'h33baf5a4),
	.w6(32'hb63fbc67),
	.w7(32'hb84f153d),
	.w8(32'hb8288c6c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba650fe6),
	.w1(32'hba3d5b53),
	.w2(32'hbb14fa73),
	.w3(32'h3ac7b754),
	.w4(32'h398fa9e3),
	.w5(32'hbaa7a42b),
	.w6(32'h3a2f6465),
	.w7(32'h375f9427),
	.w8(32'hbaa18f03),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390200c0),
	.w1(32'h38c4617e),
	.w2(32'h38c6faaf),
	.w3(32'h38b43f1c),
	.w4(32'h382c1f47),
	.w5(32'h37e4bdd0),
	.w6(32'hb681630d),
	.w7(32'h35de1b5d),
	.w8(32'hb7389bb6),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa005b),
	.w1(32'h369a1ab2),
	.w2(32'hb7a56077),
	.w3(32'hb7d78ce9),
	.w4(32'h387807ae),
	.w5(32'hb78154ae),
	.w6(32'h379e54da),
	.w7(32'hb86940e3),
	.w8(32'hb8af6c4b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381c5439),
	.w1(32'h381cbdcb),
	.w2(32'h3828818c),
	.w3(32'h37cd3a1d),
	.w4(32'h37a72ecd),
	.w5(32'h37efc24e),
	.w6(32'h37e21d3e),
	.w7(32'h3803d797),
	.w8(32'h37fabd0e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3898d34c),
	.w1(32'h38571d67),
	.w2(32'h3821bb06),
	.w3(32'h38788ba8),
	.w4(32'h3810be46),
	.w5(32'h37f5d567),
	.w6(32'h3881ac96),
	.w7(32'h380c5a5a),
	.w8(32'h37af5d32),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4accc),
	.w1(32'hb648307e),
	.w2(32'h3a25c78a),
	.w3(32'hbace4809),
	.w4(32'hb7700642),
	.w5(32'h3a5bf676),
	.w6(32'hbad8f6cc),
	.w7(32'h38e792ed),
	.w8(32'h39df1625),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9da0b4),
	.w1(32'hbba012fc),
	.w2(32'hbc245811),
	.w3(32'h39dcdf8a),
	.w4(32'hba0715d6),
	.w5(32'hbb9328ea),
	.w6(32'h3ab2e5e8),
	.w7(32'h3a1018ca),
	.w8(32'hbaf25818),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23d39a),
	.w1(32'hbab29104),
	.w2(32'hbb98fdb8),
	.w3(32'h3aa2e9fe),
	.w4(32'h3ac2b58b),
	.w5(32'hbaf26531),
	.w6(32'h3af4fa3e),
	.w7(32'h3b1f7c78),
	.w8(32'hb8881575),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89f68c),
	.w1(32'hbb9638da),
	.w2(32'hbc062368),
	.w3(32'hb896029b),
	.w4(32'hbab6e15a),
	.w5(32'hbbb03b15),
	.w6(32'hb9cb2ba2),
	.w7(32'hba874868),
	.w8(32'hbb4d1784),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3863dd17),
	.w1(32'h38b9ca5b),
	.w2(32'h38902052),
	.w3(32'hb78c9bcf),
	.w4(32'h38937b83),
	.w5(32'h3857da8a),
	.w6(32'h3811785a),
	.w7(32'h38d74831),
	.w8(32'h3828125d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9411cc5),
	.w1(32'hb9834d6c),
	.w2(32'hb8ced41e),
	.w3(32'hb773e432),
	.w4(32'hb9426883),
	.w5(32'h37634981),
	.w6(32'hb8fb5c2a),
	.w7(32'hb980c293),
	.w8(32'hb7f52427),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d4b3f2),
	.w1(32'hb61b3acc),
	.w2(32'h377baed3),
	.w3(32'hb804c624),
	.w4(32'hb837322a),
	.w5(32'hb796fd8d),
	.w6(32'hb8485c48),
	.w7(32'hb8433a44),
	.w8(32'hb7ba86fe),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382bc213),
	.w1(32'h37e01f01),
	.w2(32'h3849d122),
	.w3(32'h3784d2a6),
	.w4(32'h36038932),
	.w5(32'h38182e64),
	.w6(32'h374824c6),
	.w7(32'hb780a33d),
	.w8(32'hb6dd35dc),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a60ed),
	.w1(32'hbb0ae10b),
	.w2(32'hbbb8aa23),
	.w3(32'h3a7f125c),
	.w4(32'h3ab0a5c5),
	.w5(32'hba9b2e2f),
	.w6(32'h3aa111ab),
	.w7(32'h3b02a3f6),
	.w8(32'hb9a4938d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ca925),
	.w1(32'hb91c0f01),
	.w2(32'hb905b08d),
	.w3(32'hb942542f),
	.w4(32'hb989c8ac),
	.w5(32'hb970691f),
	.w6(32'hb96a4036),
	.w7(32'hb9aa608f),
	.w8(32'hb9a9a933),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9264d7),
	.w1(32'h39335556),
	.w2(32'h3934d031),
	.w3(32'hba90ebd6),
	.w4(32'hb83f700c),
	.w5(32'hb998f269),
	.w6(32'hbab6bbea),
	.w7(32'h39208898),
	.w8(32'hba023a6f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1069b1),
	.w1(32'hba25a55b),
	.w2(32'hb9b31685),
	.w3(32'hbb0173ef),
	.w4(32'hb9d99814),
	.w5(32'h3960482e),
	.w6(32'hbac811d2),
	.w7(32'hb9a3700b),
	.w8(32'h39721a98),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ec387d),
	.w1(32'hb766159d),
	.w2(32'hb894166b),
	.w3(32'hb8009770),
	.w4(32'hb8e12c10),
	.w5(32'hb92615d3),
	.w6(32'hb7b106d0),
	.w7(32'hb8ea97ee),
	.w8(32'hb9365c0c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88e77e),
	.w1(32'hba80122f),
	.w2(32'hbb01c911),
	.w3(32'hba09f66e),
	.w4(32'hba123902),
	.w5(32'hbab55ed6),
	.w6(32'hb916310b),
	.w7(32'hba2c7159),
	.w8(32'hbab5a4ee),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e8eff),
	.w1(32'hb94de05c),
	.w2(32'hb8504a58),
	.w3(32'hb9228585),
	.w4(32'hb954716c),
	.w5(32'hb86cc938),
	.w6(32'hb939d11e),
	.w7(32'hb974b9e0),
	.w8(32'hb94dd697),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8497b),
	.w1(32'hbb6d0c20),
	.w2(32'hbc00eb5e),
	.w3(32'h3a8662e6),
	.w4(32'h39a7cb81),
	.w5(32'hbaefc090),
	.w6(32'h398c8781),
	.w7(32'h3a858139),
	.w8(32'hb90f29e0),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38974ec9),
	.w1(32'h36e6d5d3),
	.w2(32'h36e2a192),
	.w3(32'h391ec8bd),
	.w4(32'h35141678),
	.w5(32'h3749b32d),
	.w6(32'h38098ea0),
	.w7(32'hb85ad6b3),
	.w8(32'hb614fa7b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28b1d0),
	.w1(32'h3b175b01),
	.w2(32'h3a973a6c),
	.w3(32'hba5a0cb4),
	.w4(32'h3b91fcde),
	.w5(32'h3b4af314),
	.w6(32'hbb62aeaa),
	.w7(32'h3b733575),
	.w8(32'h3b6167fc),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule