module layer_6_featuremap_21(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2147f9),
	.w1(32'h3b3d6828),
	.w2(32'h3b1cb842),
	.w3(32'hbae65202),
	.w4(32'h3bc96399),
	.w5(32'h3bd12890),
	.w6(32'hba8dac9d),
	.w7(32'hbabf7364),
	.w8(32'hbacb923b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888124b),
	.w1(32'h3a2b7a6c),
	.w2(32'h3ae5a4e5),
	.w3(32'h3b99e59e),
	.w4(32'hb644b2f4),
	.w5(32'h3a4c7070),
	.w6(32'hb9ddb33c),
	.w7(32'hb80048bb),
	.w8(32'h39052a38),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8ece3),
	.w1(32'hbc13cb71),
	.w2(32'hbb9b53d1),
	.w3(32'hbc17bf8e),
	.w4(32'hbc0b7636),
	.w5(32'hbbb36c2e),
	.w6(32'hbc197b4e),
	.w7(32'hbba48d00),
	.w8(32'hbb65e8d3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd1336),
	.w1(32'hbb812b05),
	.w2(32'hbb8082df),
	.w3(32'hbbe7c5b5),
	.w4(32'hbb227227),
	.w5(32'hbbbc44c5),
	.w6(32'hbc1b5136),
	.w7(32'hbc18892a),
	.w8(32'hbc10a4c0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ac829),
	.w1(32'h3a83c4fc),
	.w2(32'hba281602),
	.w3(32'h3b33a5a1),
	.w4(32'h3a461f8b),
	.w5(32'hbab37698),
	.w6(32'h3b16f96f),
	.w7(32'h3912bb2d),
	.w8(32'hbb19cce6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f6aa9),
	.w1(32'h3a2d3400),
	.w2(32'h3a044770),
	.w3(32'hb8ac2d46),
	.w4(32'hb9869743),
	.w5(32'hb9fc4c8c),
	.w6(32'hbac71407),
	.w7(32'hbac5b826),
	.w8(32'hbaa802b0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71e0bc),
	.w1(32'hbb0d706b),
	.w2(32'hbb3199be),
	.w3(32'h3a87275d),
	.w4(32'hbb95aa02),
	.w5(32'hbb81e3ac),
	.w6(32'h3c2471ed),
	.w7(32'h3b968eb2),
	.w8(32'h3b9a35b0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9ed51),
	.w1(32'h3ae42994),
	.w2(32'h3aa0fd3a),
	.w3(32'hb7ed0d14),
	.w4(32'h3b20a7d9),
	.w5(32'h3ae932b3),
	.w6(32'h3b501c01),
	.w7(32'h3b260da9),
	.w8(32'h3b249489),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2a407),
	.w1(32'hbbc0fbad),
	.w2(32'hbaf65838),
	.w3(32'hbbc79fc9),
	.w4(32'hbbaee8e5),
	.w5(32'hbb864007),
	.w6(32'hbc13fb05),
	.w7(32'hbba1f948),
	.w8(32'hbb4b5af8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b76eb8),
	.w1(32'hba4275b3),
	.w2(32'h38e77dc6),
	.w3(32'hbb8b5412),
	.w4(32'hbb455a70),
	.w5(32'h39fb083b),
	.w6(32'h3a3f9a19),
	.w7(32'h38f4fa58),
	.w8(32'h3b70be88),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf22e02),
	.w1(32'h3b947e3a),
	.w2(32'h3b12cccb),
	.w3(32'h3beae55a),
	.w4(32'h3b32b51c),
	.w5(32'hbb08076f),
	.w6(32'h3bfafe3c),
	.w7(32'h3bb78940),
	.w8(32'h3b539ee0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b403d4),
	.w1(32'h3bb9c448),
	.w2(32'h3b98ea80),
	.w3(32'hbaf8f72a),
	.w4(32'h3b9ed8cd),
	.w5(32'h3b09d198),
	.w6(32'h3bd08dbc),
	.w7(32'h3bc3bdfe),
	.w8(32'h3b725177),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1be5a0),
	.w1(32'h3b42fe38),
	.w2(32'h3ac6e738),
	.w3(32'hbb46e378),
	.w4(32'h3b1708ab),
	.w5(32'h3ad45542),
	.w6(32'h3b2d4a04),
	.w7(32'h3b02cc83),
	.w8(32'h3a84f51b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85d7ff),
	.w1(32'h3b6c966c),
	.w2(32'h3b975b21),
	.w3(32'h3b3aa05a),
	.w4(32'h38aa2f2e),
	.w5(32'hba51dd6c),
	.w6(32'h3ba60d5e),
	.w7(32'hba3571bc),
	.w8(32'h37d169c0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39592560),
	.w1(32'hb986bb0c),
	.w2(32'h3acdb2bf),
	.w3(32'hba9cbe60),
	.w4(32'hb90c2f2d),
	.w5(32'h3a80eb0a),
	.w6(32'hbac254d9),
	.w7(32'hb9b49edf),
	.w8(32'h390d42e7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc747b),
	.w1(32'hbb0722eb),
	.w2(32'hbb30fb35),
	.w3(32'hbb1fa3f7),
	.w4(32'hbb4bfcdd),
	.w5(32'hbb419397),
	.w6(32'h390e1925),
	.w7(32'hba849524),
	.w8(32'hba927a8c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba58ea),
	.w1(32'h3ba83f2e),
	.w2(32'h3ba60d66),
	.w3(32'h3ab1825a),
	.w4(32'hbb697cf6),
	.w5(32'hbb4cd9c1),
	.w6(32'hbaab400c),
	.w7(32'h39ab2f4f),
	.w8(32'h3b560eb2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b254d85),
	.w1(32'h3b97cc8b),
	.w2(32'h3a74c873),
	.w3(32'h3b50c378),
	.w4(32'h3b89f8b9),
	.w5(32'h3a13ee99),
	.w6(32'h3ba15a89),
	.w7(32'h3ab34095),
	.w8(32'hbb82d575),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cdcb6),
	.w1(32'hb9783fee),
	.w2(32'h39f14576),
	.w3(32'hbb47e9f2),
	.w4(32'h389418a6),
	.w5(32'h3aa6b2d5),
	.w6(32'h3b54d8ff),
	.w7(32'h3b435558),
	.w8(32'h3b7db4e7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b30f3),
	.w1(32'h3aec6376),
	.w2(32'h3b3692bf),
	.w3(32'hbacfdee5),
	.w4(32'h3a055cab),
	.w5(32'h3aea5ab3),
	.w6(32'h3a67ac27),
	.w7(32'h3b93ec9d),
	.w8(32'h3b5eba8e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15662a),
	.w1(32'hba3db3c6),
	.w2(32'hb8aadbe2),
	.w3(32'hbacb6773),
	.w4(32'hbb22bce0),
	.w5(32'hba869bd2),
	.w6(32'h39838d7d),
	.w7(32'h3a9db5cb),
	.w8(32'h3ab42743),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b289dda),
	.w1(32'h3a195d29),
	.w2(32'h3ae1ff2f),
	.w3(32'h3b748c45),
	.w4(32'h3b1831ac),
	.w5(32'hbad3d23f),
	.w6(32'hbb7429ac),
	.w7(32'h3ab44593),
	.w8(32'hbb2f8766),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbefd73),
	.w1(32'hbacf0a5f),
	.w2(32'hbb25365f),
	.w3(32'hbb841a84),
	.w4(32'hb8d4fdf0),
	.w5(32'hbaae5d41),
	.w6(32'h3ad40e58),
	.w7(32'h39b7ae0f),
	.w8(32'hb97f9983),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba884fc),
	.w1(32'hbb0106a6),
	.w2(32'hbb07f5ad),
	.w3(32'h3bdece33),
	.w4(32'hbb974056),
	.w5(32'hbbbd7071),
	.w6(32'h3c15e501),
	.w7(32'hbb1b4984),
	.w8(32'hbb00adf9),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f02c7),
	.w1(32'hbb111930),
	.w2(32'hbbd0ea93),
	.w3(32'hbb9b0b92),
	.w4(32'hbb189dc6),
	.w5(32'hbc1c874e),
	.w6(32'hbbe4029d),
	.w7(32'hbb13fd24),
	.w8(32'hbb11638e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61133c),
	.w1(32'hbba6c550),
	.w2(32'hbb88c638),
	.w3(32'hbc90915d),
	.w4(32'hbba2bd25),
	.w5(32'hbbc88961),
	.w6(32'hbc8003a9),
	.w7(32'hbbeea18b),
	.w8(32'hbbeae8e1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b215bee),
	.w1(32'hbae55989),
	.w2(32'hba1aef02),
	.w3(32'h3b2fdaed),
	.w4(32'hbb21fa5f),
	.w5(32'hbadca4ca),
	.w6(32'h3abc9c28),
	.w7(32'h394ea17a),
	.w8(32'h3977c348),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba819b36),
	.w1(32'h3a11840e),
	.w2(32'h399c5476),
	.w3(32'hbaef3bf8),
	.w4(32'h3b2d3bf3),
	.w5(32'h3aeb3b3c),
	.w6(32'hbab668f0),
	.w7(32'hba0959cf),
	.w8(32'hba5c32bb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20daf9),
	.w1(32'h39089336),
	.w2(32'h3a3ea663),
	.w3(32'h3ad4573c),
	.w4(32'hba4383a9),
	.w5(32'hba6dd677),
	.w6(32'hb99907fe),
	.w7(32'h3994b2cd),
	.w8(32'hb96483cd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd390b6),
	.w1(32'hbc5980e2),
	.w2(32'hbc7bcb38),
	.w3(32'hbd225721),
	.w4(32'hbc7f075d),
	.w5(32'hbc981ad0),
	.w6(32'hbd0920d6),
	.w7(32'hbc9b5cb3),
	.w8(32'hbcb15897),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f44df),
	.w1(32'hbb9bfb85),
	.w2(32'hbbe3fbb9),
	.w3(32'h3a73042c),
	.w4(32'hbb72b7b5),
	.w5(32'hbc46df23),
	.w6(32'hbba04d47),
	.w7(32'hbc4903ea),
	.w8(32'hbba7458f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf72d97),
	.w1(32'hb9633303),
	.w2(32'h3c21c64f),
	.w3(32'hbb4cad52),
	.w4(32'hbc252eba),
	.w5(32'hbc043744),
	.w6(32'h3a69c9a0),
	.w7(32'h3981d9c6),
	.w8(32'h3ae6887c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d3007),
	.w1(32'hba86d560),
	.w2(32'h3cf7283c),
	.w3(32'hbbfc0dd3),
	.w4(32'hbc3b7d89),
	.w5(32'hbc197372),
	.w6(32'h3b8c4479),
	.w7(32'h3ce0ade9),
	.w8(32'h3c2c024b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96a60e),
	.w1(32'h3b6a435d),
	.w2(32'h3b981347),
	.w3(32'hbc84b731),
	.w4(32'hbb8ad5f7),
	.w5(32'h3b02e12a),
	.w6(32'hbb000103),
	.w7(32'h3b526ac1),
	.w8(32'h3b300893),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b916cc3),
	.w1(32'h3b8fd85b),
	.w2(32'hbb8ffae1),
	.w3(32'h3b60e532),
	.w4(32'h3a16d377),
	.w5(32'hbb85fb53),
	.w6(32'h3a12ad0a),
	.w7(32'hbc183afb),
	.w8(32'hbc1aad0a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c3645),
	.w1(32'hbad62949),
	.w2(32'hbbd384e0),
	.w3(32'hbc617ef2),
	.w4(32'hbc9b298b),
	.w5(32'hbb5754d5),
	.w6(32'hbccbd542),
	.w7(32'h3aa102d8),
	.w8(32'hbc1ae457),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a428747),
	.w1(32'h3ae8f2de),
	.w2(32'hbb5a7da7),
	.w3(32'hbc561f19),
	.w4(32'h3b90ffa1),
	.w5(32'h3adc221e),
	.w6(32'h3a8295c3),
	.w7(32'hbb150c9b),
	.w8(32'h3ae8a0ab),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdfda4),
	.w1(32'hbbc540f5),
	.w2(32'hbbc991a6),
	.w3(32'h3b79788e),
	.w4(32'hbbd90ec0),
	.w5(32'hbc105991),
	.w6(32'hb956f0ae),
	.w7(32'hbc5e48ca),
	.w8(32'hbc92f31e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2c951),
	.w1(32'h3b7ec681),
	.w2(32'h3ba39f0c),
	.w3(32'h3c5f6156),
	.w4(32'h3a8fe8f3),
	.w5(32'h3ae47315),
	.w6(32'h3a40520f),
	.w7(32'h3b768e26),
	.w8(32'h3c04437b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca554e2),
	.w1(32'h3b9a79dd),
	.w2(32'h39d9c89c),
	.w3(32'h3c84e5b5),
	.w4(32'hbbdabfa0),
	.w5(32'hbc26e2e3),
	.w6(32'hbbad01cc),
	.w7(32'h3b2e30ac),
	.w8(32'hbb68773c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29680a),
	.w1(32'h3c30efb9),
	.w2(32'h3c03101f),
	.w3(32'hba595520),
	.w4(32'h3be7e53a),
	.w5(32'h3c724a63),
	.w6(32'h3beb3c78),
	.w7(32'h3c6b4945),
	.w8(32'h3c57c5a2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddb436),
	.w1(32'h397dd43d),
	.w2(32'hbb2177bb),
	.w3(32'h3c045584),
	.w4(32'hbb4e377a),
	.w5(32'hbb987330),
	.w6(32'hba99a60e),
	.w7(32'hbb2c2116),
	.w8(32'hba597926),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab42994),
	.w1(32'hba1dded8),
	.w2(32'hbbc25012),
	.w3(32'hb8650130),
	.w4(32'h3b51c58c),
	.w5(32'h3c3ebc07),
	.w6(32'h3bc0daf0),
	.w7(32'hbaf10641),
	.w8(32'hba4b3d63),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38350baa),
	.w1(32'h3cd3f308),
	.w2(32'hba54b0d2),
	.w3(32'h3c5fc45b),
	.w4(32'h3ca72627),
	.w5(32'hbcaa494c),
	.w6(32'hbc288961),
	.w7(32'h3cad10b2),
	.w8(32'hbc9b8277),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1c5b5),
	.w1(32'h3a87b7cc),
	.w2(32'h3bdbadea),
	.w3(32'hbcf46a05),
	.w4(32'hbc27a363),
	.w5(32'hbbf01f4f),
	.w6(32'h38128aea),
	.w7(32'h3a439776),
	.w8(32'hbaef786e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cd286),
	.w1(32'hbc7a6a7b),
	.w2(32'h3a87e487),
	.w3(32'h3a8547d0),
	.w4(32'hbc997e46),
	.w5(32'hbc7cf051),
	.w6(32'hbc849112),
	.w7(32'hbc9af675),
	.w8(32'hbc68c446),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fd599),
	.w1(32'hbc1c42b0),
	.w2(32'hbbc6b134),
	.w3(32'hbc137b87),
	.w4(32'hbb4849fa),
	.w5(32'h3b3877b0),
	.w6(32'hbbb5c932),
	.w7(32'hbc2a8ddb),
	.w8(32'hbbfc664c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa002c4),
	.w1(32'hbb0e0d5b),
	.w2(32'hbbb45dcd),
	.w3(32'h3bb99c4a),
	.w4(32'hbbf7c9c5),
	.w5(32'hbb27a890),
	.w6(32'hbaf1ee3a),
	.w7(32'hbc80b0c5),
	.w8(32'hbc3af006),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5e00f),
	.w1(32'h3bf33bd1),
	.w2(32'h3cdfe08d),
	.w3(32'h3cd4514b),
	.w4(32'h3bb8b2b6),
	.w5(32'h3b00bd8b),
	.w6(32'h3c09823e),
	.w7(32'h3b860b28),
	.w8(32'hbb23bb1d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb48552),
	.w1(32'hbc9eb4cd),
	.w2(32'hbd30bb44),
	.w3(32'hbb457f00),
	.w4(32'hbc0149e1),
	.w5(32'hbce7c89d),
	.w6(32'hbc8bcd75),
	.w7(32'hbc9741d5),
	.w8(32'h3bd63118),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c503a64),
	.w1(32'h3b3d9df0),
	.w2(32'hbb4dfc9d),
	.w3(32'hbc0d0f1c),
	.w4(32'h3ab30b5d),
	.w5(32'h3a38c511),
	.w6(32'h3bc1c980),
	.w7(32'h3a8127db),
	.w8(32'h3ad6e3d4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c207ac9),
	.w1(32'h3bb0a4fd),
	.w2(32'h3b56ee09),
	.w3(32'h3bdb5a76),
	.w4(32'hbc7de07b),
	.w5(32'hbc841ef6),
	.w6(32'hbb0fbeaa),
	.w7(32'hbad29e99),
	.w8(32'hbb489a5f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80ad0a),
	.w1(32'hbc463b03),
	.w2(32'hbca22d05),
	.w3(32'hbc73f185),
	.w4(32'hbc1c3849),
	.w5(32'hbc495b92),
	.w6(32'h3b86df9a),
	.w7(32'hbc4b253f),
	.w8(32'hbbaa3f88),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cec8166),
	.w1(32'h3cb33f94),
	.w2(32'h3c30a7a4),
	.w3(32'h3cea533f),
	.w4(32'h3caa1a75),
	.w5(32'h3c28419f),
	.w6(32'h3ccfa5ce),
	.w7(32'h3c3e8172),
	.w8(32'h3c110e7e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca38712),
	.w1(32'h3c48ab70),
	.w2(32'h3bef0c71),
	.w3(32'h3cbc2deb),
	.w4(32'h3c1a1e61),
	.w5(32'h3beddbe2),
	.w6(32'h3c85f1f2),
	.w7(32'h3bfd3ca9),
	.w8(32'h3c6ab3dd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40be27),
	.w1(32'hbc0ee637),
	.w2(32'h39a3d0d7),
	.w3(32'hb8b06eff),
	.w4(32'hbc41ac9e),
	.w5(32'hbbdb479a),
	.w6(32'hbc427fd4),
	.w7(32'hbbb1a514),
	.w8(32'hbcd76fea),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cccfd69),
	.w1(32'h3c9537b6),
	.w2(32'h3cb6780a),
	.w3(32'h3cb104ce),
	.w4(32'h3bf277a1),
	.w5(32'h3c0f5a94),
	.w6(32'h3c8425c6),
	.w7(32'h3ce9d9c5),
	.w8(32'h3c3c317c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79015b),
	.w1(32'hbc1ff078),
	.w2(32'h3b98bfff),
	.w3(32'hbcf1f6bf),
	.w4(32'hbc7e71e7),
	.w5(32'hba3e24c9),
	.w6(32'hbbaa468e),
	.w7(32'hbb80e12d),
	.w8(32'h3c12834c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd75369),
	.w1(32'hbb059d01),
	.w2(32'h3cdb0edb),
	.w3(32'h3b57ebeb),
	.w4(32'hbc310bfa),
	.w5(32'h3b696923),
	.w6(32'hbc13d0f2),
	.w7(32'hbbd89712),
	.w8(32'hbc050732),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b18df),
	.w1(32'hbc6e8d3b),
	.w2(32'h3be1c9a7),
	.w3(32'hbb597533),
	.w4(32'hbc826205),
	.w5(32'hbc6f20f5),
	.w6(32'hbccc37e2),
	.w7(32'hbc7035fa),
	.w8(32'hbc762c7e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c89be),
	.w1(32'hbc985e6f),
	.w2(32'hbc4f37f2),
	.w3(32'hbc2dfa5b),
	.w4(32'hbcbbfbac),
	.w5(32'hbc9c8fed),
	.w6(32'hbcdf4c6a),
	.w7(32'hbcaf5730),
	.w8(32'hbcba6194),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc044d7),
	.w1(32'hbb35bd67),
	.w2(32'h3c418a8e),
	.w3(32'hbb07e3a6),
	.w4(32'hb9a19f26),
	.w5(32'h3c027d5a),
	.w6(32'hbccf3603),
	.w7(32'hbb47bce3),
	.w8(32'hbbad90dd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58c863),
	.w1(32'hbd044c0f),
	.w2(32'hbd26db6a),
	.w3(32'hbc3ced88),
	.w4(32'hbcac9d23),
	.w5(32'hbcf939a8),
	.w6(32'hbc2de2cb),
	.w7(32'hbc94fe81),
	.w8(32'hbce82c4b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abedd7e),
	.w1(32'hbb3a6743),
	.w2(32'hbb5a4e2e),
	.w3(32'h3b215550),
	.w4(32'h397c7e1b),
	.w5(32'h3a54a413),
	.w6(32'hbb9b1d4e),
	.w7(32'hbbae8b8e),
	.w8(32'hbbf75170),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule