module layer_10_featuremap_322(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa22e02),
	.w1(32'hba735f36),
	.w2(32'hbb050b00),
	.w3(32'hba2c9857),
	.w4(32'hbaa21060),
	.w5(32'h3a29d3c8),
	.w6(32'hbbf9a86f),
	.w7(32'hbb2f2606),
	.w8(32'hbac1bca7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b081aa4),
	.w1(32'h39629623),
	.w2(32'hbc013d91),
	.w3(32'hbb4a6e54),
	.w4(32'hbc2ebec6),
	.w5(32'hbc84c9d6),
	.w6(32'hbb911599),
	.w7(32'hbc60df44),
	.w8(32'hbbd146aa),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe85952),
	.w1(32'hbbcbd118),
	.w2(32'hbbce20e8),
	.w3(32'hbb5d7db4),
	.w4(32'hbb3d26b8),
	.w5(32'hbb662208),
	.w6(32'h3b3d6c0e),
	.w7(32'hba81a04e),
	.w8(32'hba48f8ab),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a11c44),
	.w1(32'h3b18576f),
	.w2(32'hbb602919),
	.w3(32'h39d27655),
	.w4(32'hbb13c2b1),
	.w5(32'hbbd75d42),
	.w6(32'h3b37083d),
	.w7(32'hbb8f38fe),
	.w8(32'hbb614709),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895e57),
	.w1(32'h3b830217),
	.w2(32'hbbcce697),
	.w3(32'hba9ef80f),
	.w4(32'h3ab51c53),
	.w5(32'hbb9a19c4),
	.w6(32'hba24a8b2),
	.w7(32'hbc778437),
	.w8(32'hbacf10fd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb9251),
	.w1(32'hba707c31),
	.w2(32'h3a96f0ad),
	.w3(32'h39b5810b),
	.w4(32'h3b6bdd49),
	.w5(32'hbb80c468),
	.w6(32'h39ba9a1f),
	.w7(32'h3a1766a1),
	.w8(32'hbb8f60e0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc047c6f),
	.w1(32'hbbceeb1c),
	.w2(32'h3c0a82f3),
	.w3(32'hbc310aad),
	.w4(32'h3b56dfbe),
	.w5(32'h3c30d190),
	.w6(32'hbc30a1f4),
	.w7(32'h3c1682c6),
	.w8(32'h3c5e959a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0d709),
	.w1(32'h3c5113c2),
	.w2(32'h3b80d28b),
	.w3(32'h3c930134),
	.w4(32'h3c9ee6ce),
	.w5(32'hbbd094d0),
	.w6(32'h3c220d7a),
	.w7(32'h3ce1a226),
	.w8(32'h3c8e4a42),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d1d48),
	.w1(32'hb9c67a70),
	.w2(32'h3b96cdf1),
	.w3(32'hba80d5bb),
	.w4(32'h3b98fb2c),
	.w5(32'hbb89f6ed),
	.w6(32'hbb651e38),
	.w7(32'h3b0fb9b6),
	.w8(32'hbaa7719b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08c10b),
	.w1(32'h3a840dd2),
	.w2(32'h3b28b4ab),
	.w3(32'hbb8cdaf4),
	.w4(32'hbb2f489a),
	.w5(32'hbb998257),
	.w6(32'h3b058f5c),
	.w7(32'h3af45824),
	.w8(32'h3bfc2892),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9133a5),
	.w1(32'hbb23aa6e),
	.w2(32'hbb2d29c7),
	.w3(32'h3b8b7cdf),
	.w4(32'h3ad5a856),
	.w5(32'hbac2993b),
	.w6(32'h3c45f379),
	.w7(32'hbb5e6918),
	.w8(32'hba1620c2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab84ada),
	.w1(32'hbb3104dd),
	.w2(32'h3bb6fa4f),
	.w3(32'hbc069e2d),
	.w4(32'hba4a66b2),
	.w5(32'h3c572f8e),
	.w6(32'hbc772b37),
	.w7(32'h3c2513ef),
	.w8(32'h3c453a88),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c8ca0),
	.w1(32'h3afeac55),
	.w2(32'hba5961df),
	.w3(32'hbb8fe4ed),
	.w4(32'hbb42bf96),
	.w5(32'hbbc2c71a),
	.w6(32'hbbcb0417),
	.w7(32'hbb55439d),
	.w8(32'hbb2fc082),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc140cf8),
	.w1(32'hbc32d2ce),
	.w2(32'h3c99b0ac),
	.w3(32'hbc328257),
	.w4(32'h3c2fe363),
	.w5(32'h3b391059),
	.w6(32'hbc29c24f),
	.w7(32'h3bae5613),
	.w8(32'h3b5ea11b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e5599),
	.w1(32'hba325c24),
	.w2(32'h3b888450),
	.w3(32'hbaf54854),
	.w4(32'hbbfe3f79),
	.w5(32'hbc1ccddb),
	.w6(32'hbb3a3fd5),
	.w7(32'hbb82f32e),
	.w8(32'hbc58d358),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb440bc1),
	.w1(32'hbbe52437),
	.w2(32'hbc02b128),
	.w3(32'hb927a49f),
	.w4(32'hbc143d24),
	.w5(32'hbc54ae8f),
	.w6(32'h3c5ce740),
	.w7(32'h3b2918d0),
	.w8(32'hb994b23a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3883e7c6),
	.w1(32'h3b982bca),
	.w2(32'h3bd518d4),
	.w3(32'h383d222e),
	.w4(32'h3c09fa26),
	.w5(32'hbb052273),
	.w6(32'hbba7034a),
	.w7(32'h3b8224cc),
	.w8(32'h3ae5833d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b800bae),
	.w1(32'h3b601509),
	.w2(32'h3c6a5d22),
	.w3(32'h3c17d92d),
	.w4(32'h3cfbb222),
	.w5(32'h3c006835),
	.w6(32'h3c945de6),
	.w7(32'h3d09a60f),
	.w8(32'h3cbe0046),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee6404),
	.w1(32'hb9a66027),
	.w2(32'h3c5c57dd),
	.w3(32'hbaaffc83),
	.w4(32'h3c4a3a22),
	.w5(32'h3c89d73a),
	.w6(32'h3b21d484),
	.w7(32'h3c8bfcd4),
	.w8(32'h3c7b39fd),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1aed6b),
	.w1(32'hbc4d86b2),
	.w2(32'hbb52c8e3),
	.w3(32'hbc45b827),
	.w4(32'h3b5f9ecd),
	.w5(32'hbbb28a27),
	.w6(32'hbc2e8a9c),
	.w7(32'hbb3d286d),
	.w8(32'hbbfe0f1f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a18f7),
	.w1(32'h3c0cb057),
	.w2(32'h3b78fe8a),
	.w3(32'h3c5065d1),
	.w4(32'h3bd1297d),
	.w5(32'h3a258009),
	.w6(32'h3c54875b),
	.w7(32'hb9f987cb),
	.w8(32'hbb14551f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b208e93),
	.w1(32'h3b9b1658),
	.w2(32'h3c0a7eed),
	.w3(32'hba71d1f1),
	.w4(32'h3b4ad344),
	.w5(32'hbb8b837b),
	.w6(32'hbbc21c32),
	.w7(32'h39edf50e),
	.w8(32'h3a838656),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7da4a),
	.w1(32'h3c210581),
	.w2(32'h3d43434f),
	.w3(32'h3c99208f),
	.w4(32'h3d37301c),
	.w5(32'h3cb771aa),
	.w6(32'h3d3fdad5),
	.w7(32'h3da30137),
	.w8(32'h3d123f7c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3bb29),
	.w1(32'hbb83521e),
	.w2(32'h3a93f3c9),
	.w3(32'hbb58568b),
	.w4(32'hbc599046),
	.w5(32'h3bb5bd05),
	.w6(32'h3c12ebc7),
	.w7(32'hbc52a180),
	.w8(32'h3c15e2aa),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2c228),
	.w1(32'hbc5468a0),
	.w2(32'hbc2f09a4),
	.w3(32'hbc3c97c6),
	.w4(32'hbcd3f61f),
	.w5(32'hbc48c5f6),
	.w6(32'hbc987147),
	.w7(32'hbcf4e330),
	.w8(32'hbc85a76a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabb1c0),
	.w1(32'hbafd5d44),
	.w2(32'h3b19288d),
	.w3(32'hbaf58de8),
	.w4(32'h39ad1607),
	.w5(32'hbb90ac43),
	.w6(32'hbb29d4a7),
	.w7(32'h3abf9d98),
	.w8(32'hbbcb3d89),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a4468),
	.w1(32'h3bd83010),
	.w2(32'h3b2c219a),
	.w3(32'h3bfbd761),
	.w4(32'hba7c1782),
	.w5(32'hbb15b2a8),
	.w6(32'h3a3cdda9),
	.w7(32'h3a4c633c),
	.w8(32'hbb72693f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1cc0f),
	.w1(32'h3c18e4a1),
	.w2(32'h3bebc69c),
	.w3(32'h3b404546),
	.w4(32'hbb15c669),
	.w5(32'hbc2f4b42),
	.w6(32'hbbe3df0f),
	.w7(32'hbc129afe),
	.w8(32'hbca75162),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98e51c),
	.w1(32'hbcb035c4),
	.w2(32'hbc8d5d3f),
	.w3(32'hbcd93f4c),
	.w4(32'hbc37bba1),
	.w5(32'hbb2d4168),
	.w6(32'hbc8dbc9a),
	.w7(32'hbce0bec8),
	.w8(32'h3b3fcfe9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f55c55),
	.w1(32'h3aa7f94e),
	.w2(32'hbb823f3c),
	.w3(32'hbb1c477c),
	.w4(32'hbc808228),
	.w5(32'hbc27cca0),
	.w6(32'h3bb09b3b),
	.w7(32'hbc8078df),
	.w8(32'hbc7d1e7a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b28f9d),
	.w1(32'hbc44f2a5),
	.w2(32'hbae9b271),
	.w3(32'hbb172ca6),
	.w4(32'h3b5c309f),
	.w5(32'hbc2c87c0),
	.w6(32'hba9ebd5c),
	.w7(32'h3b249d28),
	.w8(32'hbb933613),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ed4be),
	.w1(32'hbbf9e891),
	.w2(32'hbb040fb7),
	.w3(32'hbc260062),
	.w4(32'hbc2a40f6),
	.w5(32'hbb753c04),
	.w6(32'hbc0fa1e3),
	.w7(32'hbbc4c46e),
	.w8(32'h3a580300),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8af0b),
	.w1(32'hbc20e7bf),
	.w2(32'h38538b6e),
	.w3(32'hbc97b835),
	.w4(32'h3a4c0d2e),
	.w5(32'hbaea69a7),
	.w6(32'hbc6b5a7c),
	.w7(32'h3a470e6d),
	.w8(32'h3b419325),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b095ac9),
	.w1(32'hba5f86d8),
	.w2(32'hbc24608c),
	.w3(32'hba0e0ec4),
	.w4(32'hbc38c0ed),
	.w5(32'h3ca8717e),
	.w6(32'h3b976f20),
	.w7(32'hbca36b0c),
	.w8(32'h3ca57158),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13c847),
	.w1(32'h3b99f494),
	.w2(32'h3cab7b04),
	.w3(32'h3bb28303),
	.w4(32'hb7468b73),
	.w5(32'h3b6dcf12),
	.w6(32'h3d002363),
	.w7(32'h3c2ff99b),
	.w8(32'h3b923ffc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3999bc),
	.w1(32'hbbc0361c),
	.w2(32'h3aef885b),
	.w3(32'h393a1645),
	.w4(32'h3b187afe),
	.w5(32'hba2adb34),
	.w6(32'hbb950c1e),
	.w7(32'hb9d14420),
	.w8(32'h3bf2ed22),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c2ce80),
	.w1(32'hbd049c65),
	.w2(32'h3bf1a560),
	.w3(32'hbd03fad8),
	.w4(32'hbd0cfb0c),
	.w5(32'h3c230dd7),
	.w6(32'hbce7cfaa),
	.w7(32'hbb955868),
	.w8(32'h3cba4718),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91d99a),
	.w1(32'h3c54550e),
	.w2(32'hbc1edecf),
	.w3(32'h3c045157),
	.w4(32'hbc9d4f6a),
	.w5(32'hbcd01af5),
	.w6(32'h3b0b1bf7),
	.w7(32'hbcf263d2),
	.w8(32'hbcc443dc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19328e),
	.w1(32'h3cb6d611),
	.w2(32'h3c1b58d6),
	.w3(32'h3b93b132),
	.w4(32'h3ab29064),
	.w5(32'h3a82e364),
	.w6(32'hbc2a8ba2),
	.w7(32'hbc8bd9ae),
	.w8(32'hbc8aa708),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b100402),
	.w1(32'hba8d304d),
	.w2(32'h3b25e638),
	.w3(32'h390233a3),
	.w4(32'h3b0a51c5),
	.w5(32'hbb2a6760),
	.w6(32'hbbebf25e),
	.w7(32'hba907aac),
	.w8(32'hbb8bf774),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf248c),
	.w1(32'h3c0c55aa),
	.w2(32'hbba1dcb8),
	.w3(32'h3bd985af),
	.w4(32'hbae3b6ef),
	.w5(32'hbbb0bd8a),
	.w6(32'h3cde9a61),
	.w7(32'hbc2837c4),
	.w8(32'hbbd3576b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b8c3a),
	.w1(32'hbb1d664d),
	.w2(32'hbb53a281),
	.w3(32'hbbfeee2e),
	.w4(32'hbbc831b3),
	.w5(32'hbc113433),
	.w6(32'hbbfbdaea),
	.w7(32'hbbbd61b2),
	.w8(32'hbb551c21),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c3f59),
	.w1(32'hbbfc58eb),
	.w2(32'hbb04c5d1),
	.w3(32'hbb10a065),
	.w4(32'hbbd5245b),
	.w5(32'hbb9a0867),
	.w6(32'hbbacc362),
	.w7(32'hbc22c37a),
	.w8(32'h3ba71749),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d3f16),
	.w1(32'hbb46c362),
	.w2(32'hbad0a748),
	.w3(32'h3ca339b6),
	.w4(32'h3c93022b),
	.w5(32'h3b9adb56),
	.w6(32'h3ccb6193),
	.w7(32'h3c15492d),
	.w8(32'h3b9920d3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63e012),
	.w1(32'hba0658ff),
	.w2(32'hbbba3e3c),
	.w3(32'hba546a2f),
	.w4(32'hbc8eecff),
	.w5(32'hbba0629f),
	.w6(32'h392a98db),
	.w7(32'hbc7fa35f),
	.w8(32'hbb7ea5c4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0865be),
	.w1(32'hb89ca62d),
	.w2(32'hbb8c862d),
	.w3(32'hbb253836),
	.w4(32'hbb7aaec3),
	.w5(32'hbb003e51),
	.w6(32'hbb5c7012),
	.w7(32'hbc0a30f5),
	.w8(32'hbae6a166),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b0234),
	.w1(32'h3b16a403),
	.w2(32'hbc2d0710),
	.w3(32'hb9a815a2),
	.w4(32'hbc626b32),
	.w5(32'hbbffe860),
	.w6(32'h3c1b11fc),
	.w7(32'hbbb7bc7e),
	.w8(32'hbba23d1b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bbfe3),
	.w1(32'h3beba849),
	.w2(32'h3d06fec6),
	.w3(32'hba99e7df),
	.w4(32'h3d10eb3b),
	.w5(32'h3d0a6398),
	.w6(32'h3ba4e702),
	.w7(32'h3d2dfa00),
	.w8(32'h3d3dcec1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93a182),
	.w1(32'hbab1d4a1),
	.w2(32'hba8511e6),
	.w3(32'hbba86f30),
	.w4(32'hbbedb3d2),
	.w5(32'hbacb5b55),
	.w6(32'hbb86b3f2),
	.w7(32'hbbcc82c9),
	.w8(32'hbb75bc2f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e1640),
	.w1(32'h3baafe2f),
	.w2(32'h3ae6625d),
	.w3(32'hba092da2),
	.w4(32'h39b8ea4f),
	.w5(32'h3bb1c190),
	.w6(32'hbbb6746c),
	.w7(32'hba6c65ba),
	.w8(32'hbbdec9c9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0afc41),
	.w1(32'h3c78f608),
	.w2(32'h3ca4b50b),
	.w3(32'h3c607ac1),
	.w4(32'h3c2482b2),
	.w5(32'h3a9c65c2),
	.w6(32'h3cc4b4c5),
	.w7(32'h3aff3b23),
	.w8(32'h3a8d4c69),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9a35e),
	.w1(32'hb96705e7),
	.w2(32'h3b349e27),
	.w3(32'h3b97d754),
	.w4(32'h3bd67358),
	.w5(32'hbc26c306),
	.w6(32'h3a07cc9f),
	.w7(32'hba903311),
	.w8(32'hbc0c4b2f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21b0a6),
	.w1(32'hbcb2ecaa),
	.w2(32'hbc156beb),
	.w3(32'hbc8d2209),
	.w4(32'hbcb6f34a),
	.w5(32'hbbb0af88),
	.w6(32'hbb9b4f16),
	.w7(32'hbcd60a90),
	.w8(32'h39bc39a0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb906fb),
	.w1(32'h3c0cf66b),
	.w2(32'h3c9acaef),
	.w3(32'h3ba4f1df),
	.w4(32'h3c6fb4e7),
	.w5(32'h3b5f7ef0),
	.w6(32'h3c61729e),
	.w7(32'h3cf78643),
	.w8(32'h3c2927c5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd47aad),
	.w1(32'hbbf408f0),
	.w2(32'hbc282a0f),
	.w3(32'hbb974d99),
	.w4(32'hbc7e2db0),
	.w5(32'h3b2caf11),
	.w6(32'h3a94992e),
	.w7(32'hbc5fbc63),
	.w8(32'h3c753470),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfe8ab),
	.w1(32'h3c985aba),
	.w2(32'hbb0fab13),
	.w3(32'hbb89d2f9),
	.w4(32'hbc968dfe),
	.w5(32'h3cbd1fcc),
	.w6(32'h3cb35b1a),
	.w7(32'hbcc64110),
	.w8(32'h3c88f8da),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42fca9),
	.w1(32'h3c88bad1),
	.w2(32'h3c0e9ef9),
	.w3(32'h3c7f62e6),
	.w4(32'hbb47222d),
	.w5(32'hbb521bfb),
	.w6(32'h3cb30445),
	.w7(32'hbbbd2ae9),
	.w8(32'hbb3b771a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9a98c),
	.w1(32'h3a516d48),
	.w2(32'hbbb9c25e),
	.w3(32'h3b3002a2),
	.w4(32'hba616c1f),
	.w5(32'hbb92363e),
	.w6(32'h3ca59684),
	.w7(32'hbc4b3b60),
	.w8(32'hbbf61359),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20aabe),
	.w1(32'h3b079b25),
	.w2(32'hbafbc7ed),
	.w3(32'hba888d8b),
	.w4(32'hbbaf30e8),
	.w5(32'hbbebce86),
	.w6(32'hbbca8890),
	.w7(32'hbbaf8bf6),
	.w8(32'hbc0b3d31),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc024a36),
	.w1(32'hbbbbf99c),
	.w2(32'hba42186c),
	.w3(32'hbc3ca251),
	.w4(32'hbb357529),
	.w5(32'h3a389281),
	.w6(32'hbc2875e9),
	.w7(32'hba0b8856),
	.w8(32'h3a6a3c19),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e5702),
	.w1(32'h3ad4ac36),
	.w2(32'h3bba820d),
	.w3(32'hbb68892f),
	.w4(32'h3bbaa93f),
	.w5(32'h3be9a189),
	.w6(32'h3bb31861),
	.w7(32'h3c190893),
	.w8(32'h3bb047b5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e695e),
	.w1(32'hbabea8d4),
	.w2(32'hbb1b40ae),
	.w3(32'h3c5bc9d5),
	.w4(32'h3bb88380),
	.w5(32'h3ba9b6df),
	.w6(32'h3c3ec5ad),
	.w7(32'h3c074b39),
	.w8(32'h3bc6befd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ff804),
	.w1(32'hbc8bdc19),
	.w2(32'h3c62f0e6),
	.w3(32'hbbc1053c),
	.w4(32'hbb1ca2f3),
	.w5(32'h3c7489e8),
	.w6(32'h3b754d46),
	.w7(32'hbae35ca1),
	.w8(32'h3c198c4e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34efc),
	.w1(32'h3c969daa),
	.w2(32'h3c48ce70),
	.w3(32'h3c850f96),
	.w4(32'h3b2f7b33),
	.w5(32'h3bc44420),
	.w6(32'h3cd5da90),
	.w7(32'h3b6b46a3),
	.w8(32'h3b020820),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8af839),
	.w1(32'h3c787a5f),
	.w2(32'h3c45b777),
	.w3(32'h3c1837dd),
	.w4(32'hbc9b441d),
	.w5(32'hbc82b3f8),
	.w6(32'h3d0f0a60),
	.w7(32'hbc15901c),
	.w8(32'hbc404e97),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f30e3),
	.w1(32'hbcb90672),
	.w2(32'hbc804475),
	.w3(32'hbc342032),
	.w4(32'hbc8f1415),
	.w5(32'hba61c251),
	.w6(32'hbc1eceeb),
	.w7(32'hbcb544b4),
	.w8(32'hbabac8bd),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f15e1),
	.w1(32'hbc22a873),
	.w2(32'hbb3941a0),
	.w3(32'hbc06506c),
	.w4(32'hbbc00548),
	.w5(32'hbcb73db9),
	.w6(32'h3aa52056),
	.w7(32'h3c5a7480),
	.w8(32'hbc0b4866),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc90f8c),
	.w1(32'h3c4c49b7),
	.w2(32'h3c0aa679),
	.w3(32'hb9575c9f),
	.w4(32'h3ae9cd70),
	.w5(32'hba8a99c9),
	.w6(32'hbbb64ab2),
	.w7(32'hba978da1),
	.w8(32'h3c31fba4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27509d),
	.w1(32'h3c9e863a),
	.w2(32'hbc033ba5),
	.w3(32'h3cbcdaeb),
	.w4(32'hbb7c7586),
	.w5(32'h3c449d23),
	.w6(32'h3d313067),
	.w7(32'hbbad1de1),
	.w8(32'h3c0e4bef),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82e3f4),
	.w1(32'h3c1e29f1),
	.w2(32'hbb4049da),
	.w3(32'h3ba7fc6b),
	.w4(32'hbc7c8d89),
	.w5(32'hbcac36c8),
	.w6(32'hbbf794f0),
	.w7(32'hbcb60f57),
	.w8(32'hbc8f44ce),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1dca5),
	.w1(32'h3a374e20),
	.w2(32'h3b161cde),
	.w3(32'hbb6c5f5c),
	.w4(32'hbb022033),
	.w5(32'hba5a086d),
	.w6(32'hbbc927e1),
	.w7(32'h3ac83a27),
	.w8(32'hbc6002b5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22e233),
	.w1(32'hb7528eb1),
	.w2(32'h3ab2b8f7),
	.w3(32'hbbffcb7d),
	.w4(32'hba154e93),
	.w5(32'h39017704),
	.w6(32'hb9b98741),
	.w7(32'hbb2037a8),
	.w8(32'hbb5ce580),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67ce07),
	.w1(32'h37e49d72),
	.w2(32'hba7d0193),
	.w3(32'hbb1a953b),
	.w4(32'hbba5c687),
	.w5(32'h3ae30606),
	.w6(32'hbb4bf99e),
	.w7(32'h3ad68947),
	.w8(32'hbb00cd5c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d506e),
	.w1(32'hbaca7037),
	.w2(32'h3c21c2e7),
	.w3(32'hb8de9d0d),
	.w4(32'h3ba8acf3),
	.w5(32'h3b9963c6),
	.w6(32'h3c0d1693),
	.w7(32'h3c12fa93),
	.w8(32'h3be1ccbd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ba74c),
	.w1(32'hbb7789eb),
	.w2(32'hbadf7301),
	.w3(32'h3b835b53),
	.w4(32'h3a32e3e2),
	.w5(32'h38d75841),
	.w6(32'h3b95cc56),
	.w7(32'hba793af0),
	.w8(32'h3b4beaff),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b471c9d),
	.w1(32'h3bf7e91c),
	.w2(32'h3c3f2632),
	.w3(32'h3acbade2),
	.w4(32'h3c3c6e8a),
	.w5(32'h3bec7721),
	.w6(32'h3c1dffa2),
	.w7(32'h3c5fc04c),
	.w8(32'h3ceb6940),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c655001),
	.w1(32'h3b88cf7a),
	.w2(32'hbc183f37),
	.w3(32'h3c7cd54a),
	.w4(32'h3c926df6),
	.w5(32'h3c623ca4),
	.w6(32'h3cd87536),
	.w7(32'h3cd37d3c),
	.w8(32'h3cdbe7f9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc88905),
	.w1(32'hbb34ff59),
	.w2(32'hbba1e3bf),
	.w3(32'h3b5ad73b),
	.w4(32'hbb174f43),
	.w5(32'hbb291f52),
	.w6(32'h3ab08dca),
	.w7(32'hbbcd5819),
	.w8(32'hbbaceb47),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9eb17d),
	.w1(32'hbafb9b52),
	.w2(32'h3b586cd3),
	.w3(32'hbbd91707),
	.w4(32'h3b08f7f6),
	.w5(32'h3950457a),
	.w6(32'hbb820b24),
	.w7(32'h3c433424),
	.w8(32'h3b15704f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d89a6),
	.w1(32'h3b5fa53a),
	.w2(32'h3c22dfa0),
	.w3(32'hba85aab1),
	.w4(32'h3b949c4c),
	.w5(32'hbb9aa0a8),
	.w6(32'hbbd37ba1),
	.w7(32'h3bce087b),
	.w8(32'hbac8a2aa),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8220a),
	.w1(32'h3a89c996),
	.w2(32'h3b501366),
	.w3(32'hbb6f3934),
	.w4(32'hbbefb73b),
	.w5(32'h3b0be330),
	.w6(32'hbaf0e001),
	.w7(32'hbaf7ae38),
	.w8(32'hba79c47f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b568069),
	.w1(32'hb95223ab),
	.w2(32'h3c261acc),
	.w3(32'hbb4c14b2),
	.w4(32'h3bf8ef54),
	.w5(32'h3a67cb5f),
	.w6(32'h3b336587),
	.w7(32'h3c215525),
	.w8(32'h3cca8b2f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf04b2c),
	.w1(32'h3c306042),
	.w2(32'hbc852213),
	.w3(32'h3c038b1d),
	.w4(32'hbafdbfca),
	.w5(32'hba0f32f9),
	.w6(32'h3d1367a5),
	.w7(32'h3b4cc7ea),
	.w8(32'h3a945ed5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ee28a),
	.w1(32'hbb4b3eb6),
	.w2(32'hbc0f9941),
	.w3(32'h3afb288e),
	.w4(32'hbbe68108),
	.w5(32'hbc50281b),
	.w6(32'h3b373032),
	.w7(32'hbc36f4c9),
	.w8(32'hbbdf8ea4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb688093),
	.w1(32'h3c4e134a),
	.w2(32'h3c36ef58),
	.w3(32'hbbe0502b),
	.w4(32'h3c15019c),
	.w5(32'hbc375ebd),
	.w6(32'h3b650c2e),
	.w7(32'h3cdbc90d),
	.w8(32'h3aed485e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a82e39),
	.w1(32'hbb16e2b5),
	.w2(32'hbb0befa8),
	.w3(32'h3b281012),
	.w4(32'h3a572496),
	.w5(32'h3ac36538),
	.w6(32'h3bd1a0b3),
	.w7(32'hba501ea6),
	.w8(32'h3990a7c6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b3a92),
	.w1(32'hbc057235),
	.w2(32'hbc2e84a1),
	.w3(32'hbb169416),
	.w4(32'hbcafacb9),
	.w5(32'hbb8e7bdd),
	.w6(32'hbad696f2),
	.w7(32'hbc5173ca),
	.w8(32'h3bc56ba2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a7742),
	.w1(32'hbc0161de),
	.w2(32'hbbf19a66),
	.w3(32'hbb42c0e1),
	.w4(32'h3c176170),
	.w5(32'hba310743),
	.w6(32'hbc092aba),
	.w7(32'hbbcc6367),
	.w8(32'hbae5d5b5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04182e),
	.w1(32'hbaabe660),
	.w2(32'h3bd595c2),
	.w3(32'h39826f2a),
	.w4(32'h3b9b9a94),
	.w5(32'h3b5abde2),
	.w6(32'hbbee9d2f),
	.w7(32'hb96ef13d),
	.w8(32'h3c6e89b1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5abf5a),
	.w1(32'h3be7a419),
	.w2(32'h3c3326da),
	.w3(32'h3c14e4fd),
	.w4(32'h3cf125b9),
	.w5(32'h3c8ed0cb),
	.w6(32'h3cddea96),
	.w7(32'h3cf3488b),
	.w8(32'h3cfe84ca),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24c901),
	.w1(32'hb986df01),
	.w2(32'h3a2794af),
	.w3(32'h3b33563d),
	.w4(32'hbb894756),
	.w5(32'hbb5235fa),
	.w6(32'hbb5bb0f5),
	.w7(32'hbbdd5e35),
	.w8(32'h3bb6fbbc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac4fb6),
	.w1(32'hbcb4f312),
	.w2(32'hbaaf858b),
	.w3(32'hbce86002),
	.w4(32'hbc8ad26d),
	.w5(32'hbbcbf8ca),
	.w6(32'hbbcc3f68),
	.w7(32'h3b97bc0b),
	.w8(32'h3be044aa),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01b5e1),
	.w1(32'h3c2e597e),
	.w2(32'hbaa9a748),
	.w3(32'h3b7f65d2),
	.w4(32'h3c27b498),
	.w5(32'hbb3a763b),
	.w6(32'hba3cbb77),
	.w7(32'hbaaf0440),
	.w8(32'hbb2c92a1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b917d99),
	.w1(32'h3a9f1d0b),
	.w2(32'hbb15969d),
	.w3(32'hbb8582f5),
	.w4(32'hbbe8fdce),
	.w5(32'hbc10d4e0),
	.w6(32'h3c3d1062),
	.w7(32'h39b6b617),
	.w8(32'h3ac3ccf3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b815402),
	.w1(32'hbb840ec8),
	.w2(32'hbb87c15b),
	.w3(32'hbc25a438),
	.w4(32'hbc61bf20),
	.w5(32'hbc51419e),
	.w6(32'hbc0df9c8),
	.w7(32'hbc293118),
	.w8(32'hbc34653e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b231564),
	.w1(32'hbbc44caa),
	.w2(32'hbb341b21),
	.w3(32'hbc1ac088),
	.w4(32'hbc7f683a),
	.w5(32'h3a9fb0be),
	.w6(32'hbc76bb9e),
	.w7(32'hbc1f2ab0),
	.w8(32'hbc02d454),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f47cc),
	.w1(32'h3ae43553),
	.w2(32'h39d914e8),
	.w3(32'h3b87ec6c),
	.w4(32'h3a10b4df),
	.w5(32'h3b9f28c1),
	.w6(32'hbb1ec887),
	.w7(32'h3ba9359c),
	.w8(32'h3c27a4bc),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb20fe6),
	.w1(32'hbc034a8b),
	.w2(32'h3a6f2aa5),
	.w3(32'h3c0af55a),
	.w4(32'h3c162acb),
	.w5(32'h3b689880),
	.w6(32'h3c7349bd),
	.w7(32'h3a22c3fb),
	.w8(32'h3b846149),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaf649),
	.w1(32'hbabdfb00),
	.w2(32'h3b815574),
	.w3(32'hbb494b83),
	.w4(32'hbaa09baa),
	.w5(32'h3c785746),
	.w6(32'hbc5674a1),
	.w7(32'h3c092c43),
	.w8(32'h3cffb73e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac59157),
	.w1(32'hbc949b60),
	.w2(32'h3a5e1487),
	.w3(32'hbc90980f),
	.w4(32'hbc273d94),
	.w5(32'h3caed5be),
	.w6(32'hbc9ca3a3),
	.w7(32'hbca064a7),
	.w8(32'h3c960422),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb41364),
	.w1(32'hbb72ce4d),
	.w2(32'hbc57dca3),
	.w3(32'hbbc5f7a2),
	.w4(32'hbcbd4909),
	.w5(32'hbc7f7cf5),
	.w6(32'hbb6a6b5f),
	.w7(32'hbd027094),
	.w8(32'hbc63ad35),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71f774),
	.w1(32'hbbd71607),
	.w2(32'hbca82bf0),
	.w3(32'h3be56708),
	.w4(32'hbc0531c0),
	.w5(32'h3b02469d),
	.w6(32'hb92a7ce8),
	.w7(32'hbc9ff22d),
	.w8(32'h3b26b51c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b251ef2),
	.w1(32'hbc8aa9fe),
	.w2(32'h35d11d30),
	.w3(32'hbc1cc564),
	.w4(32'hbc5cc6d5),
	.w5(32'h3b4a29f9),
	.w6(32'hbc0f90bc),
	.w7(32'hbbd102fa),
	.w8(32'hbb379396),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b541c),
	.w1(32'hbbd42b52),
	.w2(32'h3c177311),
	.w3(32'hbc2b588a),
	.w4(32'hba40601c),
	.w5(32'hb9ae7a2a),
	.w6(32'h3c0c1413),
	.w7(32'h3c42086b),
	.w8(32'hbc229e03),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c264955),
	.w1(32'h3b4514f1),
	.w2(32'h3c90f119),
	.w3(32'h3bc2ca25),
	.w4(32'h3bd8c763),
	.w5(32'h3d38b7d6),
	.w6(32'h3b0aba1e),
	.w7(32'h3c54cb03),
	.w8(32'h3d86aac6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c895d5a),
	.w1(32'hbb103ddd),
	.w2(32'hbc3d1c00),
	.w3(32'hbc30cac9),
	.w4(32'hbcb7b3c0),
	.w5(32'h3d08719c),
	.w6(32'hbc965964),
	.w7(32'hbd28f559),
	.w8(32'h3ccd03e6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36db68),
	.w1(32'hbb907320),
	.w2(32'h39b92eaf),
	.w3(32'hbbb403b8),
	.w4(32'hbb4dec28),
	.w5(32'h398f50dd),
	.w6(32'hbc82b585),
	.w7(32'hbbe0b09d),
	.w8(32'hbac35fb2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5caa6f),
	.w1(32'hbbc39860),
	.w2(32'hbb3c5cd3),
	.w3(32'hbb1934fd),
	.w4(32'hbbda7ba0),
	.w5(32'hbb2733aa),
	.w6(32'h3b0c03f4),
	.w7(32'hbb0f9030),
	.w8(32'hbc3e617b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc813e0a),
	.w1(32'hbbf8a78c),
	.w2(32'hbbad5ab2),
	.w3(32'hbb906947),
	.w4(32'h3a63b2e0),
	.w5(32'hbaaa831b),
	.w6(32'hbbb5e667),
	.w7(32'h3b7b27e4),
	.w8(32'hbb154f78),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8146df),
	.w1(32'h3babbd4d),
	.w2(32'h3b97e24a),
	.w3(32'h3b94a52d),
	.w4(32'h3b83f36d),
	.w5(32'h3b4a5a33),
	.w6(32'hbb6f2236),
	.w7(32'hbaff4be9),
	.w8(32'hbb94bb37),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3c03e),
	.w1(32'h3c23f645),
	.w2(32'h3c07fd6b),
	.w3(32'h3c346452),
	.w4(32'h3b04b1bc),
	.w5(32'h3ccd97c9),
	.w6(32'h3c080bf3),
	.w7(32'h387995aa),
	.w8(32'h3c9d4ff1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd64647),
	.w1(32'hbc129850),
	.w2(32'hbc1a6577),
	.w3(32'h3b1b1b64),
	.w4(32'hbc214b6e),
	.w5(32'h3b07790b),
	.w6(32'h3b61e091),
	.w7(32'hbc405012),
	.w8(32'h3be06fee),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4dd35),
	.w1(32'hbc3e3330),
	.w2(32'hbbb0b89f),
	.w3(32'h3b1d6418),
	.w4(32'h3a316938),
	.w5(32'h3b109518),
	.w6(32'hbbf5414c),
	.w7(32'hbc019870),
	.w8(32'h3b4574f3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5140a8),
	.w1(32'hbad1b230),
	.w2(32'hbb107a7f),
	.w3(32'h3bb3fccc),
	.w4(32'hbbf8022c),
	.w5(32'hbc1b816e),
	.w6(32'h3bce7670),
	.w7(32'hb99adb42),
	.w8(32'h3c6506d9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d0969),
	.w1(32'hbbcf671d),
	.w2(32'hbc216ba3),
	.w3(32'hbbb8e548),
	.w4(32'hbb93af19),
	.w5(32'h3c33c7ac),
	.w6(32'hb96d97f4),
	.w7(32'hbc2717fa),
	.w8(32'h3c2c3d80),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b644b08),
	.w1(32'hbb924373),
	.w2(32'hbbf25fbc),
	.w3(32'h3be482ca),
	.w4(32'hbb66bf80),
	.w5(32'hbc415390),
	.w6(32'h3c3dec07),
	.w7(32'hbbdf9270),
	.w8(32'hbc7c0495),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b6ad5),
	.w1(32'hba412818),
	.w2(32'h3bfcb430),
	.w3(32'h3a5c9bf2),
	.w4(32'h3b518289),
	.w5(32'h3c0ad1f4),
	.w6(32'hbaaedde8),
	.w7(32'h3b8c2a74),
	.w8(32'h3c7fd944),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc101c9),
	.w1(32'h39d27f86),
	.w2(32'hbb825e66),
	.w3(32'hba9fa596),
	.w4(32'hb9edc399),
	.w5(32'hba4bf569),
	.w6(32'hbbde59ea),
	.w7(32'hbb8624b1),
	.w8(32'hbbd8e6f2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bdc27),
	.w1(32'hba0798a9),
	.w2(32'h3abf3b36),
	.w3(32'hbb215220),
	.w4(32'hbac62527),
	.w5(32'h3a6bd119),
	.w6(32'hbc1d56ff),
	.w7(32'hbbd8d475),
	.w8(32'hbc0d0388),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10bd02),
	.w1(32'hbc44658f),
	.w2(32'h393d4254),
	.w3(32'hbbbfe8e1),
	.w4(32'hbbecca92),
	.w5(32'h3afb0dd9),
	.w6(32'hbb829d35),
	.w7(32'h3a915755),
	.w8(32'hbbf32052),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15cb16),
	.w1(32'hbba6ffbe),
	.w2(32'hbc2be1ec),
	.w3(32'h3b588f58),
	.w4(32'hbb9ccd4d),
	.w5(32'h3bf7d805),
	.w6(32'h3c0fc769),
	.w7(32'hbc093587),
	.w8(32'h3c4482b4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9faf2),
	.w1(32'h3a9eefbd),
	.w2(32'h3b435d3a),
	.w3(32'hbc4fffc6),
	.w4(32'hb9baad54),
	.w5(32'h3bb9b870),
	.w6(32'hbb78bf49),
	.w7(32'h3b1b6e24),
	.w8(32'h3cc4fbab),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c825ccd),
	.w1(32'h39a2d068),
	.w2(32'hbc5aaa7c),
	.w3(32'hbaf0d4d2),
	.w4(32'hbc8e6c88),
	.w5(32'h3c31cf8d),
	.w6(32'hbb2e8f9e),
	.w7(32'hbc746deb),
	.w8(32'h3c2111a1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60c21e),
	.w1(32'hbb8df66b),
	.w2(32'hba3916cc),
	.w3(32'h3b66f38b),
	.w4(32'hbacbd4b3),
	.w5(32'hbac41272),
	.w6(32'hbb85f879),
	.w7(32'h3a5fd03f),
	.w8(32'h3bc69a8a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6c7ed),
	.w1(32'h3b5eb6c5),
	.w2(32'hbb50adfd),
	.w3(32'hb7c13433),
	.w4(32'hbb8e540c),
	.w5(32'h3a89e41d),
	.w6(32'h3b280399),
	.w7(32'hba433e57),
	.w8(32'h3b182388),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4f69d),
	.w1(32'hb7f4e6a1),
	.w2(32'hbbd294b8),
	.w3(32'hbb430375),
	.w4(32'h39d7e538),
	.w5(32'hbb703d0f),
	.w6(32'h3902e9d4),
	.w7(32'hbb9098e9),
	.w8(32'h3a3ec744),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3973c4f8),
	.w1(32'hbbbb0cf8),
	.w2(32'h3a005523),
	.w3(32'h3a98be78),
	.w4(32'h399e359c),
	.w5(32'hbae1ed61),
	.w6(32'h3b0993a9),
	.w7(32'h3ba12d3c),
	.w8(32'h3bb844f7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23967a),
	.w1(32'hbb968dc2),
	.w2(32'hb8b188e2),
	.w3(32'hbca2fc2a),
	.w4(32'hba033e26),
	.w5(32'h3bd0710f),
	.w6(32'hbc719e1f),
	.w7(32'hbba7cfd5),
	.w8(32'h3bac1e3a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc213352),
	.w1(32'hbb1afd62),
	.w2(32'h3c0298c0),
	.w3(32'h3b44f35f),
	.w4(32'h3c017497),
	.w5(32'h3b03c95d),
	.w6(32'h3c15c156),
	.w7(32'h3c92b5b3),
	.w8(32'h3c5a7226),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68a09f),
	.w1(32'hbaa13cc0),
	.w2(32'hba17ac07),
	.w3(32'hbb5bb4d6),
	.w4(32'hba9b5a3b),
	.w5(32'h3c762751),
	.w6(32'h3b190031),
	.w7(32'h393136b4),
	.w8(32'h3c7b402c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3316ed),
	.w1(32'h395a87fc),
	.w2(32'hbc76327e),
	.w3(32'h3c2c1c6d),
	.w4(32'hbb9faf62),
	.w5(32'h3b32161e),
	.w6(32'h3c11bb55),
	.w7(32'hbc100aae),
	.w8(32'h3bd0e6ab),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b421adf),
	.w1(32'h3b47c4bf),
	.w2(32'h3b74b13e),
	.w3(32'h3bbbda29),
	.w4(32'h3b30ce18),
	.w5(32'h3c3c973f),
	.w6(32'h3adfd584),
	.w7(32'h3b0edad2),
	.w8(32'h3cc02bcd),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7827e3),
	.w1(32'hbcb85dc2),
	.w2(32'hbbe402d2),
	.w3(32'hbc5fdf79),
	.w4(32'hbbd11647),
	.w5(32'hbc095fb3),
	.w6(32'hbc81a238),
	.w7(32'h395b6276),
	.w8(32'hbb9dd4a7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0edd2f),
	.w1(32'hbb0d76ad),
	.w2(32'hbaf2d630),
	.w3(32'h3af6a886),
	.w4(32'hbbee8156),
	.w5(32'hbc7fa3fb),
	.w6(32'h3b86bd19),
	.w7(32'hbb070f4f),
	.w8(32'hbbd9dab8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c2a06),
	.w1(32'hbb375ca2),
	.w2(32'h3c977825),
	.w3(32'h38a933be),
	.w4(32'h3c57a334),
	.w5(32'h3a6b5c71),
	.w6(32'h3b80be5c),
	.w7(32'h3cf3e431),
	.w8(32'h3c2a21d7),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb13143),
	.w1(32'h3b18ff15),
	.w2(32'h3b36c4b7),
	.w3(32'hbc0a5518),
	.w4(32'hbc38fc98),
	.w5(32'hbbd0fc27),
	.w6(32'hbbcb3579),
	.w7(32'hba5634b9),
	.w8(32'hbc34b21c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba125d96),
	.w1(32'hbb53cb7b),
	.w2(32'h3b8c057b),
	.w3(32'hbb30fa99),
	.w4(32'hbaf5decd),
	.w5(32'hbb071b24),
	.w6(32'hba1c467d),
	.w7(32'h3ba21699),
	.w8(32'h3aad3092),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf26bf0),
	.w1(32'hbb5263f4),
	.w2(32'h3c854e77),
	.w3(32'h39f86f6c),
	.w4(32'h3c912113),
	.w5(32'h3baeeac7),
	.w6(32'h3b997904),
	.w7(32'h3ca6a207),
	.w8(32'h3c878e16),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12703e),
	.w1(32'hbb1fc2e8),
	.w2(32'hbab1f45d),
	.w3(32'hbb157327),
	.w4(32'hbbcf1212),
	.w5(32'h3bf3801c),
	.w6(32'h3af0f1fc),
	.w7(32'hbbf3b9f4),
	.w8(32'h3b236442),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b966e12),
	.w1(32'h3b5ec4be),
	.w2(32'h3b679241),
	.w3(32'hbae8ce3e),
	.w4(32'hbc82a967),
	.w5(32'h3c501bc8),
	.w6(32'h3a0dad2b),
	.w7(32'hbb64fce7),
	.w8(32'h3c91ccc9),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d766f),
	.w1(32'hbb905195),
	.w2(32'hbba7d254),
	.w3(32'hbbb56c1c),
	.w4(32'hbc70a5c8),
	.w5(32'h3a8e280e),
	.w6(32'hbc172605),
	.w7(32'hbba836fc),
	.w8(32'h3cac5e60),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c343303),
	.w1(32'h39a2f8fd),
	.w2(32'hbb39c947),
	.w3(32'hbc91b23e),
	.w4(32'hbbbf76ca),
	.w5(32'h3ba1a6a1),
	.w6(32'hbc90f88c),
	.w7(32'hbca235fe),
	.w8(32'hb9289649),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378c7c84),
	.w1(32'h3ab56128),
	.w2(32'h3a03f845),
	.w3(32'h3a97732b),
	.w4(32'hbbb4d1ee),
	.w5(32'hb98b7901),
	.w6(32'h3b9299b0),
	.w7(32'h3acac56f),
	.w8(32'h3bbc660c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fed72),
	.w1(32'hbc1f779e),
	.w2(32'hba958c0d),
	.w3(32'hbc2daf44),
	.w4(32'hbb10ba0f),
	.w5(32'h3b8378c9),
	.w6(32'hbc2f82a5),
	.w7(32'hbb191d0e),
	.w8(32'h3b0059dc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d16d5f),
	.w1(32'hbbbde253),
	.w2(32'hbb2c83d3),
	.w3(32'hbb2a160b),
	.w4(32'hbba40fc7),
	.w5(32'h3c30af07),
	.w6(32'hba3d5136),
	.w7(32'hbb2168bb),
	.w8(32'h3ccd4e15),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9dabcc),
	.w1(32'hbb07bc63),
	.w2(32'hbc7ae61d),
	.w3(32'hbc0c2713),
	.w4(32'hbc5bd5e7),
	.w5(32'h3c7eb737),
	.w6(32'hbb9de2e8),
	.w7(32'hbc9b7083),
	.w8(32'h3c9468ec),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada11d1),
	.w1(32'hbb45ca39),
	.w2(32'h3b278979),
	.w3(32'hbc3ed085),
	.w4(32'hbcd32ddc),
	.w5(32'h3be590cd),
	.w6(32'h3b5bb9ce),
	.w7(32'hbcc9e983),
	.w8(32'h3cd1704a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce96931),
	.w1(32'h3bbb4ac5),
	.w2(32'hbc71f720),
	.w3(32'hbbe3167c),
	.w4(32'hbbc9f006),
	.w5(32'h3c07f7ef),
	.w6(32'hbb666b41),
	.w7(32'hbc5e2838),
	.w8(32'h3b41195d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89f5f0),
	.w1(32'h3a455f28),
	.w2(32'hb9ec7d3c),
	.w3(32'hbb0b7762),
	.w4(32'h3bac1aa5),
	.w5(32'hbc934d92),
	.w6(32'hba636914),
	.w7(32'h3a5d0536),
	.w8(32'hbcce5292),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0dfe3),
	.w1(32'hba6583fd),
	.w2(32'h3c8a4636),
	.w3(32'h39cd2673),
	.w4(32'h3c845790),
	.w5(32'h3b9f8d73),
	.w6(32'h3ba88ecf),
	.w7(32'h3cca06e6),
	.w8(32'h3c2a608a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba996a4),
	.w1(32'hbb11337c),
	.w2(32'hbb90eea5),
	.w3(32'h3be2ebdf),
	.w4(32'hbb9d3d53),
	.w5(32'hbb69421e),
	.w6(32'h3b97a9d1),
	.w7(32'hbc1a3991),
	.w8(32'h3b96c6ee),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ade9e3),
	.w1(32'hbbc22d70),
	.w2(32'h3c40f059),
	.w3(32'hbcab19b6),
	.w4(32'hbb3d5bb3),
	.w5(32'h3c2b730f),
	.w6(32'hbc998da8),
	.w7(32'h3c5de298),
	.w8(32'h3cc533d8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e8e18),
	.w1(32'h3c383208),
	.w2(32'h3a9593eb),
	.w3(32'h3bef1ae5),
	.w4(32'hbc04b0da),
	.w5(32'h3acf6b4e),
	.w6(32'h3b61a0a4),
	.w7(32'hbc45c6ba),
	.w8(32'h3b8e50e8),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc180b),
	.w1(32'hbb56cbfb),
	.w2(32'hbbd08098),
	.w3(32'hbb86d9af),
	.w4(32'hbc2586b0),
	.w5(32'hbba46dc6),
	.w6(32'hb972a0ca),
	.w7(32'hbc1e2d67),
	.w8(32'hbc099223),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9030e),
	.w1(32'hbb5b5f16),
	.w2(32'hba49eaf1),
	.w3(32'hbb6b252a),
	.w4(32'hbb241913),
	.w5(32'hbbc659c0),
	.w6(32'hbb7c4976),
	.w7(32'hbb94771f),
	.w8(32'hbc0c9949),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64d5a6),
	.w1(32'hbbb22865),
	.w2(32'hba90a851),
	.w3(32'h3aa853d7),
	.w4(32'h3a4cbe86),
	.w5(32'hba0c8211),
	.w6(32'hbbb5b650),
	.w7(32'hbba3a486),
	.w8(32'h3c65de3d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c613596),
	.w1(32'hbaf5eb45),
	.w2(32'hbc229175),
	.w3(32'hbc5996ff),
	.w4(32'hbc1d755d),
	.w5(32'h3a1d0b32),
	.w6(32'hbaec9691),
	.w7(32'hbc4cab38),
	.w8(32'h3c1df079),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c287c41),
	.w1(32'hbc27b3f8),
	.w2(32'hbbc59cfb),
	.w3(32'hbc41be89),
	.w4(32'hbbd53d52),
	.w5(32'h3c28b9b9),
	.w6(32'hbc7017ef),
	.w7(32'hbc1bf7f6),
	.w8(32'hba196b02),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada64ba),
	.w1(32'hbbae77b0),
	.w2(32'hbba96ac4),
	.w3(32'hb91f2dfa),
	.w4(32'hba3fa3c5),
	.w5(32'h3b3cc178),
	.w6(32'hbb885899),
	.w7(32'hbac290c3),
	.w8(32'h3be527c9),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b6bf5),
	.w1(32'h3b8322cd),
	.w2(32'hbb2d3d60),
	.w3(32'h3b736255),
	.w4(32'hbaa0b906),
	.w5(32'h3a8d9631),
	.w6(32'hb9d0d840),
	.w7(32'hba9cef58),
	.w8(32'h3b8efbc9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47fc89),
	.w1(32'hbc44ec8b),
	.w2(32'h3bf01bf6),
	.w3(32'hbc55acfd),
	.w4(32'hbb32db9f),
	.w5(32'h3c7716a6),
	.w6(32'hbb22a0b5),
	.w7(32'h3ac2786c),
	.w8(32'h3d1c5315),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb7a2da),
	.w1(32'hbb62bec3),
	.w2(32'hbc810f02),
	.w3(32'hbc760bd3),
	.w4(32'hbc8d679f),
	.w5(32'h3b704e17),
	.w6(32'hbc824f21),
	.w7(32'hbca2d532),
	.w8(32'h3b4fa477),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5a1c0),
	.w1(32'h3bd5763a),
	.w2(32'hb948967c),
	.w3(32'h3b6ce273),
	.w4(32'h3b2da198),
	.w5(32'h3c95eaf1),
	.w6(32'h3bf304bb),
	.w7(32'hbc1bf9af),
	.w8(32'h3cb58a17),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98fc85),
	.w1(32'hbadbf668),
	.w2(32'hbc22d6fd),
	.w3(32'hbc13185d),
	.w4(32'hbca64f50),
	.w5(32'h3c125087),
	.w6(32'hbb56af70),
	.w7(32'hbce0fa95),
	.w8(32'h3bf73a00),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4b71a),
	.w1(32'h399f328f),
	.w2(32'hba953da4),
	.w3(32'hbc43539f),
	.w4(32'hbb147cc5),
	.w5(32'hbc4338f1),
	.w6(32'hbb425763),
	.w7(32'h3a904afa),
	.w8(32'h3c2198ef),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfae6e1),
	.w1(32'hbaa05089),
	.w2(32'hba684944),
	.w3(32'hb9ea3efb),
	.w4(32'hba22b9dd),
	.w5(32'h3bec4264),
	.w6(32'h3c17eb82),
	.w7(32'hbb6b2d24),
	.w8(32'h3c4b6a36),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c188231),
	.w1(32'hb9b42787),
	.w2(32'hbadcfdf9),
	.w3(32'h3b2fcac0),
	.w4(32'hbb07b8a1),
	.w5(32'hbc98da87),
	.w6(32'h3b1a4559),
	.w7(32'hbaefd38d),
	.w8(32'hbce2df70),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3d6f0),
	.w1(32'hbb6db02b),
	.w2(32'h3c44ff1e),
	.w3(32'hbb3d1991),
	.w4(32'h3b84f1b3),
	.w5(32'h3c5e54ee),
	.w6(32'h399867cb),
	.w7(32'h3c4a13e8),
	.w8(32'h3c351d30),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7846f),
	.w1(32'hbb0da4bb),
	.w2(32'h3a80378a),
	.w3(32'hbb07970a),
	.w4(32'h3a6571ba),
	.w5(32'h3b42ca98),
	.w6(32'h3acc5fb4),
	.w7(32'h3a09929b),
	.w8(32'h3c458628),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb91bb0),
	.w1(32'hbbbe954f),
	.w2(32'hbadf1efe),
	.w3(32'hbb6a1b5c),
	.w4(32'hbb0636c5),
	.w5(32'h3c07de35),
	.w6(32'hbb5a8d22),
	.w7(32'hbaf7568e),
	.w8(32'h3c7436db),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c3b5a),
	.w1(32'h3bc64586),
	.w2(32'hbb0889fc),
	.w3(32'h3c6baaf5),
	.w4(32'h3825bb5c),
	.w5(32'h3c5a8b3f),
	.w6(32'h3bdb78b8),
	.w7(32'hbc5775da),
	.w8(32'h3cb326d2),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0cdde),
	.w1(32'hbc37075f),
	.w2(32'hbbe12806),
	.w3(32'hbb8a11a2),
	.w4(32'hbc84d764),
	.w5(32'h3af5c4c9),
	.w6(32'hbbab7f13),
	.w7(32'hbcba0695),
	.w8(32'hbc52c1dd),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1c6e3),
	.w1(32'hba387a7b),
	.w2(32'h3becd7e7),
	.w3(32'h3c1a49a5),
	.w4(32'h3c7ed106),
	.w5(32'h3c04aba0),
	.w6(32'h3c0710e9),
	.w7(32'h3ca697c2),
	.w8(32'h3bbaf2a7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cbebd),
	.w1(32'h3c11a337),
	.w2(32'h3bd562c1),
	.w3(32'hbacb310c),
	.w4(32'hbae23996),
	.w5(32'h3bada6d5),
	.w6(32'h3bb8c3d2),
	.w7(32'h3bd66ea6),
	.w8(32'hb96e25c6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03f6dc),
	.w1(32'hbbb5484e),
	.w2(32'h3bd1039f),
	.w3(32'hbc025504),
	.w4(32'hba3df65b),
	.w5(32'hbbdf4263),
	.w6(32'h3b6e0fc5),
	.w7(32'h3c42a79e),
	.w8(32'hbc0b5a2d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81f0af),
	.w1(32'hb5ecbfaf),
	.w2(32'h3c44ece5),
	.w3(32'h3babd266),
	.w4(32'h3c7ef1d9),
	.w5(32'h39db2137),
	.w6(32'hbabbd82d),
	.w7(32'h3c8a1dbf),
	.w8(32'h3b8f4517),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb26085),
	.w1(32'hbbb941a3),
	.w2(32'hbc5d7279),
	.w3(32'hbbc6294d),
	.w4(32'hbc927353),
	.w5(32'hbca3f2ac),
	.w6(32'hbc2830aa),
	.w7(32'hbc39496e),
	.w8(32'hbcbfc257),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94a1f7),
	.w1(32'hbb01fdfa),
	.w2(32'h3c4c18a4),
	.w3(32'hba0ce819),
	.w4(32'h3c5cdd93),
	.w5(32'h3c320e18),
	.w6(32'h3acf4d10),
	.w7(32'h3c70ec36),
	.w8(32'h3c30e3b9),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb66059),
	.w1(32'hbc254581),
	.w2(32'hbb680407),
	.w3(32'hbb565fd5),
	.w4(32'h3af8192c),
	.w5(32'h3a9e0b50),
	.w6(32'h398f375c),
	.w7(32'hbba944ce),
	.w8(32'h3c975596),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ffc81),
	.w1(32'hb9b00065),
	.w2(32'hbbe4e477),
	.w3(32'hbac66d0f),
	.w4(32'hbbc5e4e8),
	.w5(32'h3c415c9f),
	.w6(32'hbb19ddae),
	.w7(32'hbc84d12b),
	.w8(32'h3c29f8dc),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5501f),
	.w1(32'hbc0ade09),
	.w2(32'hbbdd5acc),
	.w3(32'h3bcaea73),
	.w4(32'hbc43d1b5),
	.w5(32'h3bf0b1e3),
	.w6(32'h3bf5d3b6),
	.w7(32'hbbb2bf89),
	.w8(32'h3c18dca2),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c083dc1),
	.w1(32'hbbc6651e),
	.w2(32'hbc294ab9),
	.w3(32'hbc389374),
	.w4(32'hbc6eb292),
	.w5(32'h3c42a896),
	.w6(32'hbc057686),
	.w7(32'hbc8b1895),
	.w8(32'h3c8f833c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a8f40),
	.w1(32'h3b40bfc2),
	.w2(32'hbc0d8510),
	.w3(32'h39bfa722),
	.w4(32'hbbccb744),
	.w5(32'hbb004f1f),
	.w6(32'hbb3967e4),
	.w7(32'hbc601fb0),
	.w8(32'h3c7cc11a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe7735),
	.w1(32'h3b3d175e),
	.w2(32'hbc0ffdf2),
	.w3(32'hbb58b048),
	.w4(32'h3b02047c),
	.w5(32'h3b11162a),
	.w6(32'h393d0b4a),
	.w7(32'hbc0d5dd5),
	.w8(32'h3ba9cda4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a055547),
	.w1(32'h3b8b53cd),
	.w2(32'h3b0040fc),
	.w3(32'h3b123556),
	.w4(32'hbbe32d0b),
	.w5(32'h3c3063ef),
	.w6(32'hbba5005c),
	.w7(32'hbb5f30d7),
	.w8(32'h3c9ed6e1),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c298f36),
	.w1(32'hbc23b877),
	.w2(32'hbb03efde),
	.w3(32'hbc114fbb),
	.w4(32'hbc19b505),
	.w5(32'hbbe7de6e),
	.w6(32'hbc1c2b5b),
	.w7(32'hbbe405b8),
	.w8(32'hbb8fd5ca),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44a140),
	.w1(32'hb9707f68),
	.w2(32'h3c031bbf),
	.w3(32'h3b05cea8),
	.w4(32'h3c20a22e),
	.w5(32'hbc96b562),
	.w6(32'hbafc0637),
	.w7(32'h3c00d0bf),
	.w8(32'hbc5001ee),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced8f90),
	.w1(32'h3c662e3e),
	.w2(32'h3cecc380),
	.w3(32'h3bc99f5b),
	.w4(32'h3cc6819b),
	.w5(32'h3c7dc1f1),
	.w6(32'h3cf66443),
	.w7(32'h3d28791f),
	.w8(32'h3ca3e43d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac0653),
	.w1(32'hbb507514),
	.w2(32'hbbfe6277),
	.w3(32'h3b0f9dbf),
	.w4(32'hbc981aaf),
	.w5(32'hbc167b28),
	.w6(32'h3bf3c960),
	.w7(32'hbc6bd0b4),
	.w8(32'h3b55783e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25f66c),
	.w1(32'hba3f5ddc),
	.w2(32'h3b70cccc),
	.w3(32'hbb3fedcb),
	.w4(32'h3a7b45cd),
	.w5(32'h3b96c312),
	.w6(32'h3ba25a1c),
	.w7(32'h3c023a8d),
	.w8(32'h3bb7c025),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a6136),
	.w1(32'h3b8ba231),
	.w2(32'h3c043492),
	.w3(32'hbbc0c215),
	.w4(32'hbaf77353),
	.w5(32'h3c70eb73),
	.w6(32'hbabe1bff),
	.w7(32'h3b1a27fa),
	.w8(32'h3cb74f69),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c762ccf),
	.w1(32'h3b8f3a98),
	.w2(32'hbbb965e7),
	.w3(32'hbb85ebde),
	.w4(32'hbba60cb9),
	.w5(32'h3c030843),
	.w6(32'hbb13bbfb),
	.w7(32'hbc6ae8ad),
	.w8(32'h3c9abd1e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f74f7),
	.w1(32'hbb8770c8),
	.w2(32'hbb00767a),
	.w3(32'hbbc396c5),
	.w4(32'hbb8aaa26),
	.w5(32'h3c0faf29),
	.w6(32'hbc0c8409),
	.w7(32'hbc329bc1),
	.w8(32'h3c21d586),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48c243),
	.w1(32'hbc115192),
	.w2(32'hbb991d2d),
	.w3(32'h3b05da2c),
	.w4(32'hbc3d7772),
	.w5(32'h3b0aee8f),
	.w6(32'hbb9dd816),
	.w7(32'hbc39cd92),
	.w8(32'h3bf06f08),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade0ce6),
	.w1(32'h3b7562b5),
	.w2(32'h3b9d9926),
	.w3(32'hbb640ecb),
	.w4(32'h3afb5088),
	.w5(32'h3b9fa26b),
	.w6(32'h3bc33fc7),
	.w7(32'h3c65d7ca),
	.w8(32'h3c03717e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20b616),
	.w1(32'h3bb06798),
	.w2(32'hbc03e943),
	.w3(32'h3c3858ed),
	.w4(32'hbc1846ba),
	.w5(32'hbbffa3df),
	.w6(32'hbb9989a9),
	.w7(32'hbc9fa8b7),
	.w8(32'h3aaf221e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a55e6),
	.w1(32'hbc233d27),
	.w2(32'hbc47d460),
	.w3(32'hbbf68601),
	.w4(32'hbbf690d3),
	.w5(32'h3c8ec8b4),
	.w6(32'hbb3c3952),
	.w7(32'hbc3fb8d5),
	.w8(32'h3cb44e02),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c085c43),
	.w1(32'hbbf50680),
	.w2(32'hbba90e8f),
	.w3(32'h3a9d856f),
	.w4(32'hbb4e7a1d),
	.w5(32'h3c5dcac8),
	.w6(32'hbb9f9e62),
	.w7(32'hbc6c5e27),
	.w8(32'h3c43b2cf),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b5018),
	.w1(32'h3b083d6a),
	.w2(32'hb98143cd),
	.w3(32'h3c2a2ddd),
	.w4(32'h3b6d7003),
	.w5(32'h3b7add4a),
	.w6(32'h3c165390),
	.w7(32'hbc23b46f),
	.w8(32'hbb8307cf),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab31f3f),
	.w1(32'hb6bd7cc0),
	.w2(32'h3a5a56a7),
	.w3(32'hba882f2d),
	.w4(32'hb7ddc6ea),
	.w5(32'h3a5a09d4),
	.w6(32'h3b9c285f),
	.w7(32'h3a802039),
	.w8(32'h3c4db26d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50dafc),
	.w1(32'h3be5bd8b),
	.w2(32'h3bbdbfc1),
	.w3(32'h3c22a50f),
	.w4(32'h3a9b8532),
	.w5(32'h3c461c8f),
	.w6(32'h3bc6c08b),
	.w7(32'hbbbd739a),
	.w8(32'h3c5acac0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c107967),
	.w1(32'hbbb69979),
	.w2(32'hbc4c71de),
	.w3(32'hbc6699dc),
	.w4(32'hbc5e74d8),
	.w5(32'h3987975f),
	.w6(32'hbc0424d5),
	.w7(32'hbc98b57e),
	.w8(32'h3c12ce65),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe309e),
	.w1(32'hbad97df6),
	.w2(32'h3c00705f),
	.w3(32'hbb0e280d),
	.w4(32'hba6f03f8),
	.w5(32'h3ca90577),
	.w6(32'h3b4a4611),
	.w7(32'h3c078aaa),
	.w8(32'h3cfc306a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb53ff8),
	.w1(32'hba6d7f63),
	.w2(32'hbc70c972),
	.w3(32'hbba8d9d1),
	.w4(32'hbcc44add),
	.w5(32'h3c1aecb7),
	.w6(32'hbb4d2414),
	.w7(32'hbcbdea4c),
	.w8(32'h3ba28654),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa44e0e),
	.w1(32'hbc23783c),
	.w2(32'hbba56e97),
	.w3(32'h3c0c8ea4),
	.w4(32'hbc6c4334),
	.w5(32'h3c6e1c98),
	.w6(32'hbb8f2e48),
	.w7(32'hbc7dc3d8),
	.w8(32'h3c41a7bb),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e6ea7),
	.w1(32'hbbf84cb7),
	.w2(32'hb9a2ce41),
	.w3(32'hbba3de78),
	.w4(32'hbb853cce),
	.w5(32'hbbf8ba0d),
	.w6(32'hbc1c113e),
	.w7(32'hbbaff9a1),
	.w8(32'hbc06d502),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f7c87),
	.w1(32'h3a15a6be),
	.w2(32'hbbc13af2),
	.w3(32'hbb502eab),
	.w4(32'hbc58d2c6),
	.w5(32'hbb576d1a),
	.w6(32'h3bc78c02),
	.w7(32'hbc18c212),
	.w8(32'hbb3514cd),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdeeab4),
	.w1(32'hbb942ec4),
	.w2(32'hbb837d42),
	.w3(32'h3a930d63),
	.w4(32'h3a1cdf01),
	.w5(32'hbc5baaa1),
	.w6(32'hb90e2d2d),
	.w7(32'h3bbf9790),
	.w8(32'hbd0ab6b1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9128d4),
	.w1(32'h3c299a0f),
	.w2(32'h3c7aab79),
	.w3(32'h3c2cf280),
	.w4(32'h3c72ec02),
	.w5(32'h3c90bbe5),
	.w6(32'h3aecfdbf),
	.w7(32'h3cb53c99),
	.w8(32'h3cf651f9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dba06),
	.w1(32'hbb8fa376),
	.w2(32'hbc2f49a4),
	.w3(32'hbb6b644e),
	.w4(32'hbc738ada),
	.w5(32'h3c0b5036),
	.w6(32'hb956c98d),
	.w7(32'hbc980341),
	.w8(32'h3c0fc118),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c1667),
	.w1(32'hbc4c083f),
	.w2(32'hbc0d3950),
	.w3(32'h3b8c35d7),
	.w4(32'h3940f284),
	.w5(32'hbbb38017),
	.w6(32'h3c3eaa25),
	.w7(32'hbbbf1b69),
	.w8(32'hbbcc289e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f0dc1),
	.w1(32'h3b447327),
	.w2(32'hbb346d23),
	.w3(32'hbb0bee50),
	.w4(32'h3aedfcee),
	.w5(32'h3ca7cda9),
	.w6(32'hbb9adc4d),
	.w7(32'h3b0c06b9),
	.w8(32'h3c65ddb6),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6d891),
	.w1(32'h3a95dd30),
	.w2(32'hb848bacb),
	.w3(32'h3c2dd714),
	.w4(32'h3c2ce092),
	.w5(32'h3c6d7502),
	.w6(32'h3ca1951c),
	.w7(32'h3b57f647),
	.w8(32'h3ceebc13),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf64aee),
	.w1(32'hbc05065f),
	.w2(32'hbc7acc2f),
	.w3(32'hbb4052ce),
	.w4(32'hbc9c50e7),
	.w5(32'h3b38a6dd),
	.w6(32'hbaf4a96f),
	.w7(32'hbc576ba8),
	.w8(32'h3b8b1fbd),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f6057),
	.w1(32'hbc307d5d),
	.w2(32'h3be42665),
	.w3(32'hbc6800b0),
	.w4(32'hbc330d80),
	.w5(32'h3b883494),
	.w6(32'hbcc7d091),
	.w7(32'hb91b50fc),
	.w8(32'h3bb2c8a1),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9adc36),
	.w1(32'hba2aaf54),
	.w2(32'hbbe3df84),
	.w3(32'h3aff2b9a),
	.w4(32'h39ff1a9c),
	.w5(32'hbb5834b6),
	.w6(32'h3abe5a24),
	.w7(32'hbb196aa9),
	.w8(32'hbb307e8e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb362809),
	.w1(32'hba0be9a9),
	.w2(32'h3bbad04c),
	.w3(32'h3a42b781),
	.w4(32'h3abe1355),
	.w5(32'h3b8b99ea),
	.w6(32'h399a011e),
	.w7(32'h3b2e7748),
	.w8(32'h3c2ca46a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b9d4a),
	.w1(32'hbc08ad11),
	.w2(32'h3c1ad627),
	.w3(32'hbbfe37ca),
	.w4(32'hba1c8df0),
	.w5(32'h3caa19cd),
	.w6(32'hbcc3b3c2),
	.w7(32'hbc0ec844),
	.w8(32'h3c79c35d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f21496),
	.w1(32'h3c232f9b),
	.w2(32'h3c2fc583),
	.w3(32'h3b9e1a90),
	.w4(32'h3c9e42af),
	.w5(32'h3c0299ab),
	.w6(32'h398546c4),
	.w7(32'h3cdc13eb),
	.w8(32'h3d09ca22),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac873a4),
	.w1(32'hbcb88947),
	.w2(32'h3a61e2bf),
	.w3(32'hbcb31525),
	.w4(32'hb9d59063),
	.w5(32'h3c2bcb44),
	.w6(32'hbbdfe4c1),
	.w7(32'h3be725bb),
	.w8(32'h3cb536a9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66293c),
	.w1(32'hbb94e801),
	.w2(32'hbc10f9dc),
	.w3(32'hbc09bfdc),
	.w4(32'hbc2c684a),
	.w5(32'hbc728e3d),
	.w6(32'hbc0819a8),
	.w7(32'hbcad383c),
	.w8(32'hbc8759e8),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1374a9),
	.w1(32'h3c05ee12),
	.w2(32'hbb27e66c),
	.w3(32'h3bba2baf),
	.w4(32'hbc1e1024),
	.w5(32'hbc78ab8a),
	.w6(32'h3aad6c0e),
	.w7(32'hbc42c850),
	.w8(32'hbc46ecfa),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ec1f5),
	.w1(32'h3b276666),
	.w2(32'h3ba5b08e),
	.w3(32'h3a2e8d67),
	.w4(32'h3bf74c64),
	.w5(32'hbbd76963),
	.w6(32'h3b727485),
	.w7(32'h3b896661),
	.w8(32'h3bfaadbe),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f6efa),
	.w1(32'h3c417f73),
	.w2(32'h3abf3eee),
	.w3(32'h3bcd9e7b),
	.w4(32'hba471a6a),
	.w5(32'hbcbbee21),
	.w6(32'h3c48f29c),
	.w7(32'hbbaea00e),
	.w8(32'hbcbc2160),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc783b47),
	.w1(32'h3b54652f),
	.w2(32'h3c39196b),
	.w3(32'hbb0bcbdf),
	.w4(32'h3c07be93),
	.w5(32'h3b1e92d3),
	.w6(32'h3c2d2ab4),
	.w7(32'h3cac3d10),
	.w8(32'h3b60f9cc),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a27b5),
	.w1(32'hbbeb9fac),
	.w2(32'hbb0aee5a),
	.w3(32'hbab52309),
	.w4(32'hbbae7903),
	.w5(32'h3b92b830),
	.w6(32'h3b484ae7),
	.w7(32'hbc133f11),
	.w8(32'h39ec0cdc),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39c29a),
	.w1(32'h3b653a53),
	.w2(32'h3b3642ec),
	.w3(32'hb9c1f3e1),
	.w4(32'hb937f83c),
	.w5(32'hbb1f755f),
	.w6(32'hbb9185a0),
	.w7(32'hbaf47716),
	.w8(32'hbbd7e011),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63bb03),
	.w1(32'h3bfee70b),
	.w2(32'h3bf8dedb),
	.w3(32'hbb4d5adc),
	.w4(32'hbacbd7cf),
	.w5(32'h3b5fcdef),
	.w6(32'h3c916719),
	.w7(32'h3b6cad40),
	.w8(32'hbb837d58),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf668c3),
	.w1(32'hbba22975),
	.w2(32'h3b4c1da4),
	.w3(32'hbbee948d),
	.w4(32'hba13e889),
	.w5(32'hb9b7d610),
	.w6(32'hbc4dbe55),
	.w7(32'h3b04146a),
	.w8(32'h3c91fda7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82bc83),
	.w1(32'h399f02a5),
	.w2(32'hbabb95aa),
	.w3(32'h3c072678),
	.w4(32'h3c28e999),
	.w5(32'hba44eead),
	.w6(32'h3ce5c5f7),
	.w7(32'hbb076fcb),
	.w8(32'hbbf666bc),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20153f),
	.w1(32'hbc245e72),
	.w2(32'h3c5f59f0),
	.w3(32'hbc6949fd),
	.w4(32'h3a6b55fa),
	.w5(32'h3b7e9be6),
	.w6(32'hbc421cbd),
	.w7(32'h3c655301),
	.w8(32'h3bf544ea),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05a09a),
	.w1(32'h3b0a7454),
	.w2(32'h3b59921d),
	.w3(32'h3999c28f),
	.w4(32'h3bb22966),
	.w5(32'hbb8eed69),
	.w6(32'h3bcd46ef),
	.w7(32'h3c8ce03d),
	.w8(32'h3b9ad1c6),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f70db),
	.w1(32'hbbde681f),
	.w2(32'hbb1cf886),
	.w3(32'hbbd38f60),
	.w4(32'h3b1790d2),
	.w5(32'hbba76e7d),
	.w6(32'hbc351d0c),
	.w7(32'hbb80e4b0),
	.w8(32'hbb823dec),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2561c6),
	.w1(32'h3b386616),
	.w2(32'h3c013d23),
	.w3(32'hbb9d1ee4),
	.w4(32'h3bbc8305),
	.w5(32'hba4f3d40),
	.w6(32'hbc328e08),
	.w7(32'h3bedfedd),
	.w8(32'h3c441b55),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e7b2d),
	.w1(32'hbb6bdf9e),
	.w2(32'h390aa75a),
	.w3(32'h3bd7a32f),
	.w4(32'hbb870c49),
	.w5(32'h3beeed44),
	.w6(32'h3c335a09),
	.w7(32'h3b2f4fa5),
	.w8(32'h3bfef972),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a106b),
	.w1(32'hbbda4e40),
	.w2(32'h3c2729ff),
	.w3(32'hbc30fedd),
	.w4(32'h3b9a0179),
	.w5(32'h3b689a17),
	.w6(32'hbc00e14b),
	.w7(32'h3bdd5c97),
	.w8(32'h3ab757bb),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a87b3),
	.w1(32'h3badabfb),
	.w2(32'hba6c6fda),
	.w3(32'h3bd5582d),
	.w4(32'hbabe3edf),
	.w5(32'h3aa84dbc),
	.w6(32'h3b03e4ff),
	.w7(32'hbb2c166e),
	.w8(32'hbaa52409),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcd86f),
	.w1(32'hb9c19762),
	.w2(32'hbaa72cbf),
	.w3(32'hbb925eee),
	.w4(32'hbb06c13e),
	.w5(32'h3bbf491a),
	.w6(32'hbae04b20),
	.w7(32'hbb2cec88),
	.w8(32'hbaba65d4),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bb095),
	.w1(32'h3b68fea3),
	.w2(32'hbafba9b8),
	.w3(32'h3b9eca98),
	.w4(32'hba67bd81),
	.w5(32'h3c11bd57),
	.w6(32'h3ab13ed2),
	.w7(32'h394dcfcc),
	.w8(32'h3c93e36d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ef3fb),
	.w1(32'h3c4caa5c),
	.w2(32'hbadf093d),
	.w3(32'h3c3d5381),
	.w4(32'hbbd926a0),
	.w5(32'hbadef0b4),
	.w6(32'h3c938a70),
	.w7(32'h3b3e73ae),
	.w8(32'h3b84358a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a47681),
	.w1(32'hbad83f4c),
	.w2(32'h3c153876),
	.w3(32'hbb221ff0),
	.w4(32'h3bfce8ef),
	.w5(32'h3c4f627d),
	.w6(32'hbbac3c67),
	.w7(32'h3bd677ec),
	.w8(32'h3c3bea21),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd64107),
	.w1(32'h3c1cfc03),
	.w2(32'h3c1024ee),
	.w3(32'h3c2b7002),
	.w4(32'h3b4b7fd7),
	.w5(32'h3ba1e63e),
	.w6(32'hba3bac42),
	.w7(32'h399fceaf),
	.w8(32'h3a518f2b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c4dc6),
	.w1(32'h3c014730),
	.w2(32'hb9d2c589),
	.w3(32'hbb1f081f),
	.w4(32'h3b8754e2),
	.w5(32'h3c0ce1ce),
	.w6(32'h389c6e8a),
	.w7(32'h3b50ed4a),
	.w8(32'h3cb1ae3c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cababd8),
	.w1(32'h3c9dfd7a),
	.w2(32'hbb9863b0),
	.w3(32'h3cb29284),
	.w4(32'h3bf1998b),
	.w5(32'h3aefb60e),
	.w6(32'h3cec5709),
	.w7(32'hbb57ca93),
	.w8(32'hbac155ef),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfc7a5),
	.w1(32'hbb8c113a),
	.w2(32'h3ac79023),
	.w3(32'hbb4f6ce6),
	.w4(32'h3b0c65c3),
	.w5(32'hbc1babba),
	.w6(32'hbb00eba0),
	.w7(32'h3abbec3f),
	.w8(32'hbb0f06d2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1be05b),
	.w1(32'hbb8c1e7d),
	.w2(32'hbc06c4ef),
	.w3(32'hbc19e526),
	.w4(32'hbb61cf00),
	.w5(32'h3c349f8a),
	.w6(32'hbc5b70a7),
	.w7(32'hbb185ac0),
	.w8(32'h3bfe57a8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be11e3f),
	.w1(32'hbb597881),
	.w2(32'h3bab9b68),
	.w3(32'hbb9c68dc),
	.w4(32'hbaa74a84),
	.w5(32'h3babe6e8),
	.w6(32'hbb861d94),
	.w7(32'h3a24f5ee),
	.w8(32'h3b39266f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d075e),
	.w1(32'h3b0fb7d8),
	.w2(32'hbb28966e),
	.w3(32'h3b264877),
	.w4(32'hbb786808),
	.w5(32'hbb7d7106),
	.w6(32'hbbc63ef3),
	.w7(32'hbbeecc67),
	.w8(32'h3a84c009),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacc8e8),
	.w1(32'h3b3b6255),
	.w2(32'h3bf41bb0),
	.w3(32'hbb87cf0e),
	.w4(32'hbba3587c),
	.w5(32'hbb19df85),
	.w6(32'h3c5ef945),
	.w7(32'h3c4b8afc),
	.w8(32'hbb898a62),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2a915),
	.w1(32'h3a301e3b),
	.w2(32'hbc0a4b84),
	.w3(32'h3b3cfff4),
	.w4(32'hbb7bca02),
	.w5(32'hbbbba83c),
	.w6(32'h3bdbad03),
	.w7(32'hbc14ab97),
	.w8(32'hbc387309),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57bdc7),
	.w1(32'hbbc7f442),
	.w2(32'hbada1388),
	.w3(32'hbb2d862e),
	.w4(32'hbc0db46f),
	.w5(32'hbbd9ca3c),
	.w6(32'hbb135ae8),
	.w7(32'hbc37c0bd),
	.w8(32'hbbed7334),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e3555),
	.w1(32'h3a1dd611),
	.w2(32'hbb42ec4b),
	.w3(32'hbb01e297),
	.w4(32'h3bcecb74),
	.w5(32'hbb7d5fab),
	.w6(32'hbb0311c2),
	.w7(32'h3a94119b),
	.w8(32'hbb9dbdd8),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b84dd),
	.w1(32'hbb2c139f),
	.w2(32'hbbbe278b),
	.w3(32'hbb96b1ed),
	.w4(32'hbc19c387),
	.w5(32'h3a368e90),
	.w6(32'hbb66da9c),
	.w7(32'hbb9ec082),
	.w8(32'hba61a201),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f1dbd),
	.w1(32'hbc87eef3),
	.w2(32'hbc3469f9),
	.w3(32'hbb5078b4),
	.w4(32'hbc26eaba),
	.w5(32'hbc46bc67),
	.w6(32'h3c1bb6a7),
	.w7(32'h3c65b88b),
	.w8(32'hbbbd3cfd),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58c2c5),
	.w1(32'hbb36f4f6),
	.w2(32'h3b0cf82d),
	.w3(32'hbb5a04e9),
	.w4(32'hb9a424e8),
	.w5(32'h3c97ed75),
	.w6(32'hbbe9bdcc),
	.w7(32'hbb79ecec),
	.w8(32'h3ca98f6a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58daae),
	.w1(32'h3c2b18c8),
	.w2(32'h3a2166ac),
	.w3(32'h3ab24896),
	.w4(32'hbb4d0585),
	.w5(32'h3b1be788),
	.w6(32'hbba165f8),
	.w7(32'hbc150e19),
	.w8(32'h3c67c89d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule