module layer_10_featuremap_68(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92937f),
	.w1(32'hbbbc84f6),
	.w2(32'hb8959f41),
	.w3(32'hbcd640b1),
	.w4(32'hbc3b6001),
	.w5(32'hbbf32a96),
	.w6(32'hbc107058),
	.w7(32'hbc4c5fec),
	.w8(32'hbb64b895),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b9e2c),
	.w1(32'hbbb3fead),
	.w2(32'hbae306f9),
	.w3(32'h3a9c3fea),
	.w4(32'hba41b667),
	.w5(32'hba8e1b84),
	.w6(32'h3bbea4c6),
	.w7(32'h3aec4861),
	.w8(32'hbb27f613),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a211f7a),
	.w1(32'hbb65637f),
	.w2(32'h3b5fcd4b),
	.w3(32'h3a6686e9),
	.w4(32'hba2491dd),
	.w5(32'h3bab07d5),
	.w6(32'h3bada56e),
	.w7(32'hb91f0904),
	.w8(32'h3bb5caf5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9640ef),
	.w1(32'hbb0c9ef5),
	.w2(32'hbc92257a),
	.w3(32'h3b24369b),
	.w4(32'h3b2617b1),
	.w5(32'hbc9f465d),
	.w6(32'h3bf309e7),
	.w7(32'hbb07a4dd),
	.w8(32'hbbc0b99c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70ef1a),
	.w1(32'hbc3f6c77),
	.w2(32'hbb7abc35),
	.w3(32'hbc337249),
	.w4(32'hbc821a15),
	.w5(32'hbb7b5776),
	.w6(32'hbbfca1af),
	.w7(32'hbc177fc6),
	.w8(32'hbbcacdf1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac5a20),
	.w1(32'h39735fd8),
	.w2(32'hbb49a30d),
	.w3(32'hbb561b84),
	.w4(32'hbb345a26),
	.w5(32'h3a14f641),
	.w6(32'hbc20c394),
	.w7(32'hbbe59dad),
	.w8(32'h39cac509),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0b09b),
	.w1(32'hbc21aae8),
	.w2(32'hbc237560),
	.w3(32'hba8d682e),
	.w4(32'hbbd594f9),
	.w5(32'hbce71e90),
	.w6(32'hbb0ce2e4),
	.w7(32'hbc08bb91),
	.w8(32'hbc397bde),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb981f2),
	.w1(32'hbc72d352),
	.w2(32'hbb371dcb),
	.w3(32'hbcc587a9),
	.w4(32'hbc83cc90),
	.w5(32'h3bbe181e),
	.w6(32'hbc172adf),
	.w7(32'hbbdbbf53),
	.w8(32'h3b5dc5f5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf43407),
	.w1(32'hbc01f2d5),
	.w2(32'hbc99e043),
	.w3(32'hbbf14b8c),
	.w4(32'hbc324ee4),
	.w5(32'hbc348b48),
	.w6(32'h3aba1e4f),
	.w7(32'h3ac16fe9),
	.w8(32'hbb3ec2af),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc251351),
	.w1(32'h3b39d299),
	.w2(32'hbb29b686),
	.w3(32'h3a5f4cfa),
	.w4(32'h3c208245),
	.w5(32'hb9952d0c),
	.w6(32'hbb419aba),
	.w7(32'h3a484275),
	.w8(32'hbb0317e0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2d73d),
	.w1(32'hbbae7e3d),
	.w2(32'h3b953d7b),
	.w3(32'hbacdee12),
	.w4(32'hbab28ab3),
	.w5(32'h3c2b8f52),
	.w6(32'hba02c0df),
	.w7(32'h39dca6be),
	.w8(32'h3b398a40),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9f7aa),
	.w1(32'h3c2c078d),
	.w2(32'h3c8398c7),
	.w3(32'h3c042a63),
	.w4(32'hbb7118d2),
	.w5(32'h3c4c8bc5),
	.w6(32'h3bc6c7a7),
	.w7(32'hbbf1c677),
	.w8(32'h3b015ecd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00a6fc),
	.w1(32'h3b67e2bc),
	.w2(32'hb9291628),
	.w3(32'h3b9e40a9),
	.w4(32'hba9889e7),
	.w5(32'h3b8288e6),
	.w6(32'hbb0c98c3),
	.w7(32'hbb82d54f),
	.w8(32'h395f39f0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87506f),
	.w1(32'hbb06c0b0),
	.w2(32'h3bcf84c7),
	.w3(32'h39fb288c),
	.w4(32'h3b85ce42),
	.w5(32'h3b9e2f75),
	.w6(32'h3bdda829),
	.w7(32'h3b96d91d),
	.w8(32'hbac83210),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2124a),
	.w1(32'hbc734123),
	.w2(32'h3a2c66ff),
	.w3(32'hbbdb769a),
	.w4(32'hbca3943b),
	.w5(32'hb954a892),
	.w6(32'hbc32ddd9),
	.w7(32'hbc485ef1),
	.w8(32'hbae7e3c6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab54cab),
	.w1(32'h3b640d18),
	.w2(32'h39958868),
	.w3(32'hbae709bb),
	.w4(32'h3b1f7a06),
	.w5(32'h3b51291d),
	.w6(32'hb9ece059),
	.w7(32'h3bd5df98),
	.w8(32'h3a72f98a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9fc8e),
	.w1(32'hbbd21e7a),
	.w2(32'h3c9f9a7b),
	.w3(32'hbb160798),
	.w4(32'hbb2b3898),
	.w5(32'h3cc0d148),
	.w6(32'h39756ce5),
	.w7(32'h3a9f955e),
	.w8(32'h3c5bcef3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95b0c4),
	.w1(32'h3ae1f80f),
	.w2(32'hbab7fa5c),
	.w3(32'h3cb28cf9),
	.w4(32'hbb28796f),
	.w5(32'hba29cd31),
	.w6(32'h3bd66883),
	.w7(32'hbc9004bf),
	.w8(32'h379fd152),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e0875),
	.w1(32'h3aa9eef4),
	.w2(32'h3a22a858),
	.w3(32'h3bb278b8),
	.w4(32'hbb9245e8),
	.w5(32'h3bda0609),
	.w6(32'hbb36d612),
	.w7(32'hbb96f41b),
	.w8(32'h3b986c8e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac32ad3),
	.w1(32'h3a53545e),
	.w2(32'h3bfb3f55),
	.w3(32'h3c1a2904),
	.w4(32'hbc1a0cf2),
	.w5(32'h3c056380),
	.w6(32'h3c063c7d),
	.w7(32'hbb095201),
	.w8(32'h3ad7cad8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01be7f),
	.w1(32'hbade95d7),
	.w2(32'hbad763b3),
	.w3(32'h3babd624),
	.w4(32'hbad77164),
	.w5(32'h3c1436ae),
	.w6(32'hb9837bde),
	.w7(32'hbb823113),
	.w8(32'h3b4af71b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde0547),
	.w1(32'h3c206652),
	.w2(32'h3a5225ff),
	.w3(32'h3c0e0f93),
	.w4(32'h3b787755),
	.w5(32'hbbe557cf),
	.w6(32'h3bb9a95e),
	.w7(32'hbbfdbf94),
	.w8(32'hbbeb79fe),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c2634),
	.w1(32'hbbce95bd),
	.w2(32'h3bc751e2),
	.w3(32'hbaf383ac),
	.w4(32'hbc27cb1d),
	.w5(32'h3bb765cf),
	.w6(32'hbbf6584e),
	.w7(32'hbc0fad97),
	.w8(32'hbb0c3f96),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53427e),
	.w1(32'h3b69d7a1),
	.w2(32'h3b0e17d7),
	.w3(32'hba9c98b0),
	.w4(32'hba119f91),
	.w5(32'hbb9932f5),
	.w6(32'hbb87bced),
	.w7(32'hbb99d34c),
	.w8(32'h3b8cd7a7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beff8cf),
	.w1(32'hb9e4010d),
	.w2(32'h3bf8744d),
	.w3(32'h3b143451),
	.w4(32'h3ba49993),
	.w5(32'h3b872fc1),
	.w6(32'h3b30f2ed),
	.w7(32'h3c2f92ba),
	.w8(32'hbabe9715),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d294e),
	.w1(32'hbbe55740),
	.w2(32'h3ae26048),
	.w3(32'hbbe69f69),
	.w4(32'hbbe1554f),
	.w5(32'hbb601ecc),
	.w6(32'hbbc30f91),
	.w7(32'hbc81ca1f),
	.w8(32'h39339a85),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13b8ed),
	.w1(32'hbb143a92),
	.w2(32'h3a3e253d),
	.w3(32'hbb23407e),
	.w4(32'hbc09bdeb),
	.w5(32'h3a10ee20),
	.w6(32'hbc0e9cc6),
	.w7(32'h3aa5deec),
	.w8(32'h3895023c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63a252),
	.w1(32'h3b10f55a),
	.w2(32'h3cd199c2),
	.w3(32'h3b6ed9af),
	.w4(32'hbb44b5e5),
	.w5(32'h3ce34c1b),
	.w6(32'h3b021a64),
	.w7(32'h397d13ae),
	.w8(32'h3c880292),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce06bff),
	.w1(32'h3c82c19a),
	.w2(32'h3c0ec6c5),
	.w3(32'h3cf5b83c),
	.w4(32'h3c64e4df),
	.w5(32'h3c18a94e),
	.w6(32'h3c3f054e),
	.w7(32'hbb4bbff7),
	.w8(32'hbb2a8d31),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17d61f),
	.w1(32'h3be76b06),
	.w2(32'hbc1030ee),
	.w3(32'h3bfc3dea),
	.w4(32'hbb9afd47),
	.w5(32'hbc0bb605),
	.w6(32'h3beb20a0),
	.w7(32'hbb184982),
	.w8(32'hbb2a3074),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fedeb),
	.w1(32'h3ba67a6c),
	.w2(32'hbbd7ed81),
	.w3(32'h3b947d9d),
	.w4(32'h3bffa4b4),
	.w5(32'h3b48f69b),
	.w6(32'h3b8cbd60),
	.w7(32'h3b47368b),
	.w8(32'hbb9d80d0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d4f1c),
	.w1(32'hbb9e5a7e),
	.w2(32'h3bf58f82),
	.w3(32'h3a45f4c5),
	.w4(32'hbbac28b6),
	.w5(32'hbb145234),
	.w6(32'hbac38e3a),
	.w7(32'hb9f27d26),
	.w8(32'hbbe53f19),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81e463),
	.w1(32'hba1a6daf),
	.w2(32'h3be2c318),
	.w3(32'hbbe36230),
	.w4(32'hbbb370db),
	.w5(32'h3c086a04),
	.w6(32'hbb675668),
	.w7(32'hbaa1c046),
	.w8(32'hbba71596),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c0bf2),
	.w1(32'h3b3d0bb1),
	.w2(32'h3b57f8d6),
	.w3(32'h3b9d5c2d),
	.w4(32'hbbc26259),
	.w5(32'h3ba54e5a),
	.w6(32'hbc5398bf),
	.w7(32'hbcab3efe),
	.w8(32'hbb9d1899),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0307f4),
	.w1(32'h3b63e181),
	.w2(32'h3bbd42b3),
	.w3(32'h3b90572c),
	.w4(32'hbb1d6b60),
	.w5(32'h3b9a1df3),
	.w6(32'hbbca2a82),
	.w7(32'hbc648260),
	.w8(32'hbb4a48ed),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2de94),
	.w1(32'hbb3e2f02),
	.w2(32'h3c46f8e5),
	.w3(32'hbb09d4d0),
	.w4(32'hbc163b03),
	.w5(32'h3b2357dd),
	.w6(32'hbbdf4877),
	.w7(32'hbc244ff6),
	.w8(32'hbc21c515),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b956ea9),
	.w1(32'hbc3a917e),
	.w2(32'h3cdaa7f3),
	.w3(32'hbbffe796),
	.w4(32'hbc285089),
	.w5(32'h3cd4ff9b),
	.w6(32'hbc493288),
	.w7(32'h3a56b5e0),
	.w8(32'hb9fd5c6b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d01da50),
	.w1(32'h3bd72c90),
	.w2(32'h3a7a94e1),
	.w3(32'h3c44e54d),
	.w4(32'hbc2db4e3),
	.w5(32'hb9f1b907),
	.w6(32'hbc86c997),
	.w7(32'hbd0e76b2),
	.w8(32'h3b9b273c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf79a64),
	.w1(32'h3c33e5be),
	.w2(32'hbab0e870),
	.w3(32'h3b1e02cf),
	.w4(32'h3b33f052),
	.w5(32'hbafac4c3),
	.w6(32'h3b9eb2e4),
	.w7(32'h3b0ed035),
	.w8(32'hbc7738b3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b962b27),
	.w1(32'h3a96277f),
	.w2(32'h3b0b1e18),
	.w3(32'h3c2eda9e),
	.w4(32'h3af18066),
	.w5(32'h3a57fbfb),
	.w6(32'hba0e4454),
	.w7(32'h3af7caa3),
	.w8(32'h37424321),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97bd7a),
	.w1(32'hba5b45e8),
	.w2(32'h3aa54ba1),
	.w3(32'hbb776f3a),
	.w4(32'h3b869f5f),
	.w5(32'h3bf72543),
	.w6(32'h3a04db43),
	.w7(32'h3c419b19),
	.w8(32'hb9ee0cdd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffdf5b),
	.w1(32'h3a170e52),
	.w2(32'hbaad0b03),
	.w3(32'h3c1756b3),
	.w4(32'h3a965a0e),
	.w5(32'h3b497f1d),
	.w6(32'h3a076665),
	.w7(32'h3b8a4d46),
	.w8(32'h3b29a1ba),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a982913),
	.w1(32'hba9e0b2c),
	.w2(32'h3c6ec13d),
	.w3(32'h3ba2ab7a),
	.w4(32'hba001b51),
	.w5(32'h3c2d7fed),
	.w6(32'hba367888),
	.w7(32'h3b4cfabf),
	.w8(32'h395c558c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11c0a4),
	.w1(32'hbae43cae),
	.w2(32'h3b119fdf),
	.w3(32'hb9c61896),
	.w4(32'hbc2bb09e),
	.w5(32'h3b722b67),
	.w6(32'hbc033d3c),
	.w7(32'hbc562fda),
	.w8(32'h3bebd090),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43716a),
	.w1(32'hbaa45fa2),
	.w2(32'hbb51efe7),
	.w3(32'h3b9cb3bc),
	.w4(32'h3b9c99c1),
	.w5(32'hbc022a03),
	.w6(32'h3c176389),
	.w7(32'hba921b15),
	.w8(32'hbba3e48d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3951ee66),
	.w1(32'hbb0f8b92),
	.w2(32'hbbb43923),
	.w3(32'hbc1c817f),
	.w4(32'hbc38756a),
	.w5(32'hba6d5219),
	.w6(32'hbc04e70c),
	.w7(32'hbb9db1fb),
	.w8(32'hbbfcbf06),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd186a7),
	.w1(32'hbc0e8dae),
	.w2(32'hbc364ae7),
	.w3(32'h3b96be73),
	.w4(32'h39aaadcf),
	.w5(32'hbc3f06df),
	.w6(32'hbbb0c6f0),
	.w7(32'hbb0cb473),
	.w8(32'hbb77412d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc07f9),
	.w1(32'h39909761),
	.w2(32'h3c63ec64),
	.w3(32'hbb8ecb0b),
	.w4(32'hbbf72888),
	.w5(32'h3c519a61),
	.w6(32'hbbdbbc56),
	.w7(32'hbc73bb66),
	.w8(32'h3baa4540),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c724ada),
	.w1(32'h3ba8943b),
	.w2(32'hbbcafe86),
	.w3(32'h3bf21a57),
	.w4(32'hbb0ff734),
	.w5(32'hba5ea285),
	.w6(32'h3ae173f8),
	.w7(32'hbbc06f78),
	.w8(32'h3bb67fd9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88f988),
	.w1(32'h3b8caf0c),
	.w2(32'h3bd8d1f6),
	.w3(32'h3b9d599b),
	.w4(32'h3bc43fc2),
	.w5(32'hbab7c156),
	.w6(32'h3bcf8ace),
	.w7(32'h3bedbb76),
	.w8(32'hbb8af79a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d8a95),
	.w1(32'hbb660be0),
	.w2(32'hbc57701b),
	.w3(32'hbc3f2731),
	.w4(32'hbbf24b8b),
	.w5(32'hbcdfe1e1),
	.w6(32'hbbc96595),
	.w7(32'hba197410),
	.w8(32'hbc8f8158),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccfccdf),
	.w1(32'hbc6ca3d7),
	.w2(32'h3b94470d),
	.w3(32'hbca8b09f),
	.w4(32'hba402589),
	.w5(32'hbb9a11aa),
	.w6(32'hbc883ffd),
	.w7(32'hbc0ef98e),
	.w8(32'h3b539104),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75d75e),
	.w1(32'h39bf4279),
	.w2(32'hbcb6eee5),
	.w3(32'hbbb75b90),
	.w4(32'hb8fa1214),
	.w5(32'hbd1391c3),
	.w6(32'h3a556b70),
	.w7(32'h3ba16a03),
	.w8(32'hbc8f4395),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfb6c33),
	.w1(32'hbcffddaa),
	.w2(32'hbb665083),
	.w3(32'hbd1bc4c1),
	.w4(32'hbce09807),
	.w5(32'h3bb87557),
	.w6(32'hbc9a8170),
	.w7(32'hbc849ada),
	.w8(32'h3ba1c01b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc179197),
	.w1(32'hbbbd1e06),
	.w2(32'h3b54e666),
	.w3(32'hbb30ab95),
	.w4(32'h3a236637),
	.w5(32'hbc0dd61c),
	.w6(32'hbba7174d),
	.w7(32'hbbbca9c3),
	.w8(32'hb93f3afc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93127b),
	.w1(32'hbb9855ff),
	.w2(32'hbbb74fec),
	.w3(32'hbc1e06b2),
	.w4(32'hbc155acd),
	.w5(32'h3b8b96ad),
	.w6(32'hbbee5a7f),
	.w7(32'hbc22efb2),
	.w8(32'h3c4a9c1a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d027a),
	.w1(32'h3c1f1423),
	.w2(32'hba25fa60),
	.w3(32'h3bbe5737),
	.w4(32'h3b9d4413),
	.w5(32'h3cdac644),
	.w6(32'h3c1598b6),
	.w7(32'h3c136634),
	.w8(32'h3d27eb95),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cde2a3e),
	.w1(32'h3d3ae4e2),
	.w2(32'h3b067a9f),
	.w3(32'h3d655961),
	.w4(32'h3d47b35e),
	.w5(32'h3bdc8cb9),
	.w6(32'h3d585bfa),
	.w7(32'h3d00d7fd),
	.w8(32'h3b9528cd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3869bb),
	.w1(32'h3c6031eb),
	.w2(32'hbba265f7),
	.w3(32'h3c296e33),
	.w4(32'h3c72e0e7),
	.w5(32'h3c44a119),
	.w6(32'h3bf19f32),
	.w7(32'h3c6d3c92),
	.w8(32'h3cd40acd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8552c7),
	.w1(32'h3ca363d7),
	.w2(32'hbc5884a9),
	.w3(32'h3d20e1fb),
	.w4(32'h3cb8c017),
	.w5(32'hbc80fe91),
	.w6(32'h3d00d02d),
	.w7(32'h3c0c1110),
	.w8(32'hbc2bdbff),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e7d09),
	.w1(32'hbc1aac5e),
	.w2(32'hbb96308d),
	.w3(32'hbb820900),
	.w4(32'hbad04fed),
	.w5(32'h3b87ca55),
	.w6(32'h3985a64b),
	.w7(32'hb93ff095),
	.w8(32'hbb9099fd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdb0da),
	.w1(32'h3a5bebf3),
	.w2(32'hbb4aff43),
	.w3(32'h3a49934a),
	.w4(32'hbb51f854),
	.w5(32'hbb98ebaf),
	.w6(32'hbb3055e1),
	.w7(32'hbc0f91e4),
	.w8(32'hbba2b8f0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e81ca),
	.w1(32'hbb935546),
	.w2(32'h3927e10d),
	.w3(32'h381881d4),
	.w4(32'hba3a8ace),
	.w5(32'h3ca077a0),
	.w6(32'hbbf22e74),
	.w7(32'hbb572a3f),
	.w8(32'hbb51e049),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c021fe4),
	.w1(32'h3b1f6c9d),
	.w2(32'hbb5a017c),
	.w3(32'h3cf4f965),
	.w4(32'h3c5b8012),
	.w5(32'hbb0e15e4),
	.w6(32'h3bcfed4d),
	.w7(32'h3c007c95),
	.w8(32'h3b860475),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981ae7a),
	.w1(32'h3a34d023),
	.w2(32'hbbe0c294),
	.w3(32'h3aeb13b1),
	.w4(32'h3b94ba62),
	.w5(32'hbbc29168),
	.w6(32'h3b41fde4),
	.w7(32'h3a7d64e9),
	.w8(32'hbba943cf),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fb34c),
	.w1(32'hbbcf6e5c),
	.w2(32'h3bb3c72b),
	.w3(32'hbc19e5c4),
	.w4(32'hbbaa9f8c),
	.w5(32'h3b5b72e8),
	.w6(32'hbc0bc486),
	.w7(32'hbb4b9691),
	.w8(32'hbc10b34f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9612a6),
	.w1(32'hbbd29fed),
	.w2(32'hbb252475),
	.w3(32'hba426890),
	.w4(32'hbc000f17),
	.w5(32'h3a4b6872),
	.w6(32'hbc3dedc5),
	.w7(32'hbc6290dd),
	.w8(32'h3a24df27),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2442a),
	.w1(32'h3ab1582d),
	.w2(32'h3c34a246),
	.w3(32'hbaadb459),
	.w4(32'hbbb1746a),
	.w5(32'h3aea5392),
	.w6(32'hbbdcd3b9),
	.w7(32'hbb961ac4),
	.w8(32'hba834197),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b984613),
	.w1(32'h3bb30b5d),
	.w2(32'h3b03f65e),
	.w3(32'hbb87d2ef),
	.w4(32'hbb53bb5f),
	.w5(32'h3b183a5a),
	.w6(32'hbc1da280),
	.w7(32'hb9d81230),
	.w8(32'h3b39ef3a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb8991),
	.w1(32'h3b9d07a9),
	.w2(32'hbc9a7dfa),
	.w3(32'hba53b215),
	.w4(32'h3b3e8c63),
	.w5(32'hbd082057),
	.w6(32'h3b81923f),
	.w7(32'h3b5ad706),
	.w8(32'hbce30e1a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd27daef),
	.w1(32'hbccb3549),
	.w2(32'hbb4fe000),
	.w3(32'hbd341111),
	.w4(32'hbcb84e68),
	.w5(32'h3b7d25c5),
	.w6(32'hbcf9bc51),
	.w7(32'hbc2c645b),
	.w8(32'h3a6dce18),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ce244),
	.w1(32'h3ba4166b),
	.w2(32'hbb8d401c),
	.w3(32'h3beaa62e),
	.w4(32'h3c02efcc),
	.w5(32'hbb2c248f),
	.w6(32'h3c08fa4b),
	.w7(32'h3a90c581),
	.w8(32'hbbe0b7c4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad36dcc),
	.w1(32'hbb7e988f),
	.w2(32'h3be6356e),
	.w3(32'hb98b78ea),
	.w4(32'h38fc44d8),
	.w5(32'h3c15bf0f),
	.w6(32'hbbcffc4d),
	.w7(32'hbb897c2a),
	.w8(32'h3bf42be3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac0993),
	.w1(32'h3b66181d),
	.w2(32'hb901c8ac),
	.w3(32'h3c363c30),
	.w4(32'h3b9167d1),
	.w5(32'h3b51756f),
	.w6(32'h3bf9d288),
	.w7(32'hbb30d60e),
	.w8(32'h3bdb56fb),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabee1c5),
	.w1(32'hb83861e1),
	.w2(32'hbc7ebb1f),
	.w3(32'h39303309),
	.w4(32'hbb5cbf31),
	.w5(32'hbc1cc8fb),
	.w6(32'h3b11e878),
	.w7(32'hbb1e9a66),
	.w8(32'hbc3937d3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c5e34),
	.w1(32'hbc4ce5ea),
	.w2(32'h3c078606),
	.w3(32'hbc0b1fa3),
	.w4(32'hbc82fb18),
	.w5(32'hba9a89cb),
	.w6(32'hbc22366d),
	.w7(32'hbc93db1c),
	.w8(32'h3ac242ee),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1da71),
	.w1(32'hb9843ae4),
	.w2(32'h3a73547e),
	.w3(32'hbb93a7ae),
	.w4(32'hbbd1bcb8),
	.w5(32'hbbec225c),
	.w6(32'h39d506bd),
	.w7(32'hbac12984),
	.w8(32'hbc09d69b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc195a2a),
	.w1(32'hbc29dded),
	.w2(32'hbc05ce63),
	.w3(32'hbc411bf7),
	.w4(32'hbbdba459),
	.w5(32'hbb19b11e),
	.w6(32'hbba6d5df),
	.w7(32'hbb2ad214),
	.w8(32'h3b6a0de1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b459b),
	.w1(32'h3bfc933f),
	.w2(32'h3b21c722),
	.w3(32'h3baa9c80),
	.w4(32'hba25731d),
	.w5(32'hbbd32d31),
	.w6(32'h3bb868be),
	.w7(32'h3b771a5a),
	.w8(32'h3a578912),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc663061),
	.w1(32'h3a684b15),
	.w2(32'hbc6eae3d),
	.w3(32'hbcb12d25),
	.w4(32'hbbf71f51),
	.w5(32'hbcd51ea3),
	.w6(32'hbc5d8726),
	.w7(32'hb9bccf3e),
	.w8(32'hbc74d457),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc60f2),
	.w1(32'hbc334916),
	.w2(32'h3c124eb9),
	.w3(32'hbcd952d5),
	.w4(32'hbc831004),
	.w5(32'h3c1be998),
	.w6(32'hbcb1f592),
	.w7(32'hbc8026a1),
	.w8(32'h3b0ad5dc),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39de54),
	.w1(32'h3c192f7e),
	.w2(32'h3c4641f1),
	.w3(32'h3c37b291),
	.w4(32'h3c02f585),
	.w5(32'h3c3b1468),
	.w6(32'h3a099b19),
	.w7(32'hbaf6e787),
	.w8(32'h3bcef759),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5837c),
	.w1(32'hbb216fcd),
	.w2(32'hb9e3b22b),
	.w3(32'hbb350da2),
	.w4(32'h39badfb1),
	.w5(32'h3bc3c99b),
	.w6(32'hbb946be1),
	.w7(32'hbb844975),
	.w8(32'h3b48a2ff),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc06a0),
	.w1(32'hbb100e96),
	.w2(32'hbb2da680),
	.w3(32'h3abb6d39),
	.w4(32'h3994f1e6),
	.w5(32'h3b689e8f),
	.w6(32'hbac63c98),
	.w7(32'hb97f5412),
	.w8(32'h3b870f29),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62dd46),
	.w1(32'hbb089c5c),
	.w2(32'h3b21f396),
	.w3(32'h3b38564a),
	.w4(32'hba9026a0),
	.w5(32'h3c8a6a02),
	.w6(32'h3ac80be6),
	.w7(32'hbbc972b8),
	.w8(32'h3b800e33),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be88110),
	.w1(32'h3b92fb0b),
	.w2(32'h3c858693),
	.w3(32'h3bda5e6c),
	.w4(32'hbb854579),
	.w5(32'h3cb5a89e),
	.w6(32'hbb7afa8d),
	.w7(32'hbc45b87c),
	.w8(32'h3c80d130),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d06f6c5),
	.w1(32'h3c6f7e97),
	.w2(32'h3aa108ae),
	.w3(32'h3d0f72cd),
	.w4(32'h3c9b3474),
	.w5(32'h3b654578),
	.w6(32'h3c8d454b),
	.w7(32'h3bcdf5de),
	.w8(32'h3b2b6a19),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1d1ae),
	.w1(32'h3b57c907),
	.w2(32'h3b06197b),
	.w3(32'h39edd12c),
	.w4(32'h3b2e8579),
	.w5(32'hbb7fda96),
	.w6(32'h3a6657c9),
	.w7(32'h3b6d59a2),
	.w8(32'hbb952faa),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcadd26),
	.w1(32'hbbb794f1),
	.w2(32'hbc15adf8),
	.w3(32'hbc258df9),
	.w4(32'hbb4b9a6f),
	.w5(32'hbc57063c),
	.w6(32'hbbc7d134),
	.w7(32'hbc0f3503),
	.w8(32'hbbbe5b74),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1385d8),
	.w1(32'hbb10063e),
	.w2(32'hbcb4604f),
	.w3(32'hbc85457e),
	.w4(32'hbc414a97),
	.w5(32'hbcee3f43),
	.w6(32'hbc2bb5da),
	.w7(32'hbc348b76),
	.w8(32'hbcf618d5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcedb254),
	.w1(32'hbcf0f448),
	.w2(32'hbcd2355b),
	.w3(32'hbd12ea89),
	.w4(32'hbca1ac07),
	.w5(32'hbcb97a55),
	.w6(32'hbcd19e74),
	.w7(32'hbc9202a4),
	.w8(32'hbc772bdb),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6992c4),
	.w1(32'hbb8c196e),
	.w2(32'h3bf1fced),
	.w3(32'h3b377fe6),
	.w4(32'h3c51d729),
	.w5(32'h3b90096a),
	.w6(32'h3c3ae992),
	.w7(32'h3c6f184f),
	.w8(32'h3a8e0232),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b949c16),
	.w1(32'h3a2c26ce),
	.w2(32'hbc351f0b),
	.w3(32'hbb731b48),
	.w4(32'hbb89c65d),
	.w5(32'hbc096725),
	.w6(32'hbbc6a157),
	.w7(32'hbba962ff),
	.w8(32'h3a84fa68),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc160eb0),
	.w1(32'h3b24b5fa),
	.w2(32'h3bd74266),
	.w3(32'hb99e6ccc),
	.w4(32'h3c215253),
	.w5(32'h3c33633e),
	.w6(32'h3c0c3091),
	.w7(32'h3c4388ca),
	.w8(32'h3c0a3500),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a2e32),
	.w1(32'h3a563005),
	.w2(32'h3c065f89),
	.w3(32'h3bad0790),
	.w4(32'hbaaca5d0),
	.w5(32'h3be91695),
	.w6(32'h3a136682),
	.w7(32'hba257c10),
	.w8(32'h3c0ebbe6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5421c1),
	.w1(32'h3c0fafa2),
	.w2(32'h3ae897ed),
	.w3(32'h3c02d7b3),
	.w4(32'h3b56d82c),
	.w5(32'h3a45a86e),
	.w6(32'h3c0a84ab),
	.w7(32'h3bc77393),
	.w8(32'hbb0ef29a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc15066),
	.w1(32'h3bdb83a4),
	.w2(32'h3baa33ac),
	.w3(32'h3b126b36),
	.w4(32'hbc02dc2f),
	.w5(32'h3a4e1fdd),
	.w6(32'hbbfdb5aa),
	.w7(32'hb9f7639a),
	.w8(32'h3ade73dc),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64cb6e),
	.w1(32'h3b53b409),
	.w2(32'hbb05a4ea),
	.w3(32'h3acb55dc),
	.w4(32'h3b735927),
	.w5(32'hbc12aa2b),
	.w6(32'h3b9c6bf4),
	.w7(32'h3aec0cb6),
	.w8(32'hbc66024b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd7b6f),
	.w1(32'hbb953767),
	.w2(32'h3bbde31d),
	.w3(32'hbc01f1cc),
	.w4(32'hbc93fe3e),
	.w5(32'hbc40a180),
	.w6(32'hbcc6eefa),
	.w7(32'hbcb1e54f),
	.w8(32'hbc6f024d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18dba0),
	.w1(32'hbc90cf90),
	.w2(32'hbbc3c721),
	.w3(32'hbcc79b28),
	.w4(32'hbc9d5ec4),
	.w5(32'hb98b4aa8),
	.w6(32'hbca0d422),
	.w7(32'hbc51d03c),
	.w8(32'hba59b6d0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c5738),
	.w1(32'hbc02e67f),
	.w2(32'h3b5b2d0c),
	.w3(32'hbbf616e5),
	.w4(32'hbc0a93ac),
	.w5(32'hbbcf1a28),
	.w6(32'hba4beb03),
	.w7(32'hbbea5eff),
	.w8(32'hbb9cccfb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadad150),
	.w1(32'hbb5e74ae),
	.w2(32'hbb0b8a71),
	.w3(32'hbba7744e),
	.w4(32'hbba74864),
	.w5(32'h3af11a73),
	.w6(32'hbbcf5ea0),
	.w7(32'hbbda9ce8),
	.w8(32'h3a0e6bea),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdaf5dd),
	.w1(32'h3b9aeaf8),
	.w2(32'hbcf66930),
	.w3(32'h3cf7ef5b),
	.w4(32'h3ac47dbe),
	.w5(32'hbd15bbc6),
	.w6(32'h3c34abea),
	.w7(32'hbc3327a0),
	.w8(32'hbcd954d3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2481c0),
	.w1(32'hbcd40669),
	.w2(32'h3b3b5569),
	.w3(32'hbd44f2fb),
	.w4(32'hbcdec038),
	.w5(32'h3b770ab0),
	.w6(32'hbd0b54b8),
	.w7(32'hbcdc52f0),
	.w8(32'hbb3faa6c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba416ffb),
	.w1(32'hbb4dc56b),
	.w2(32'h3b94233e),
	.w3(32'hbb06341b),
	.w4(32'hbae4f8cb),
	.w5(32'h3c54557e),
	.w6(32'hbc2b8184),
	.w7(32'hbbcb2639),
	.w8(32'h3c226288),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e64e2),
	.w1(32'h3c102848),
	.w2(32'h3c2ab1d0),
	.w3(32'h3c966458),
	.w4(32'h3c00674f),
	.w5(32'h3c6836bd),
	.w6(32'h3c100d04),
	.w7(32'hbb6ae7ba),
	.w8(32'h3c3ba414),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d13b9),
	.w1(32'h3c4e2d01),
	.w2(32'hbb2eb24c),
	.w3(32'h3c7338ce),
	.w4(32'h3c444189),
	.w5(32'hbc1f6a92),
	.w6(32'h3c0d48ee),
	.w7(32'h3adb0903),
	.w8(32'hbb306ecb),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba67618),
	.w1(32'hbb165a7b),
	.w2(32'hbb346903),
	.w3(32'hbc301ab6),
	.w4(32'hbc287d17),
	.w5(32'hbb3db344),
	.w6(32'hbc0bf9fe),
	.w7(32'hbc5ea3b4),
	.w8(32'hbc136a21),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaaf444),
	.w1(32'hbab1a7d6),
	.w2(32'hbb4d6e1a),
	.w3(32'h3ac910a4),
	.w4(32'h3b0f0d1d),
	.w5(32'h3b28073f),
	.w6(32'hbb2d5cc7),
	.w7(32'hbbc2b3f3),
	.w8(32'h3b588007),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04ff5e),
	.w1(32'hbc47eb95),
	.w2(32'h39ae0159),
	.w3(32'h3b85cb2f),
	.w4(32'hbb1c59fa),
	.w5(32'h3b03a754),
	.w6(32'h3a7ffd1b),
	.w7(32'hbb9c8e54),
	.w8(32'hba307144),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb322053),
	.w1(32'h3b900a07),
	.w2(32'hba73c820),
	.w3(32'h3c07c273),
	.w4(32'h3acfe3fe),
	.w5(32'h3b84dec0),
	.w6(32'h3bb62bc0),
	.w7(32'hbade783f),
	.w8(32'hba9b3668),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd2883),
	.w1(32'hbb83ba28),
	.w2(32'h3c449cc9),
	.w3(32'h3b8028be),
	.w4(32'hba52608d),
	.w5(32'h3b66fcd3),
	.w6(32'h3be0263e),
	.w7(32'hbbd8627c),
	.w8(32'hbb50c953),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb889851),
	.w1(32'hbc362651),
	.w2(32'h3ba17ad6),
	.w3(32'hbc3b6ddd),
	.w4(32'hbc59c99b),
	.w5(32'h3a2d8371),
	.w6(32'hbc8177bd),
	.w7(32'hbc1d0a69),
	.w8(32'h3a8c883d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b235980),
	.w1(32'h3b14696d),
	.w2(32'h3c4cd569),
	.w3(32'h3be91328),
	.w4(32'h3b28b6c4),
	.w5(32'h3bbc2aac),
	.w6(32'h3b42c81d),
	.w7(32'h3b70a9dd),
	.w8(32'hbb40491e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60407a),
	.w1(32'h3c3d960c),
	.w2(32'h3c389826),
	.w3(32'h3c10df43),
	.w4(32'h3bbcdbe2),
	.w5(32'h3c1ed7bf),
	.w6(32'h3aa31d74),
	.w7(32'h3a1be6da),
	.w8(32'h3be93c79),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc1754),
	.w1(32'h3cae13ad),
	.w2(32'hbcf7d598),
	.w3(32'h3ca49208),
	.w4(32'h3c80f3fe),
	.w5(32'hbd425fb7),
	.w6(32'h3c785565),
	.w7(32'h3c253ef4),
	.w8(32'hbd26b91f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd31671a),
	.w1(32'hbd16fa1b),
	.w2(32'h3c7e6302),
	.w3(32'hbd573c25),
	.w4(32'hbd134e08),
	.w5(32'h3cbdb9a8),
	.w6(32'hbd0140e8),
	.w7(32'hbc64eca6),
	.w8(32'h3c8c293f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce6f7f1),
	.w1(32'h3cb2ae0a),
	.w2(32'hbc98808d),
	.w3(32'h3d09e5ad),
	.w4(32'h3cb95853),
	.w5(32'hbc1b5476),
	.w6(32'h3ce041de),
	.w7(32'h3c761fd9),
	.w8(32'hbc2c03e1),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e1ea2),
	.w1(32'hbc501b72),
	.w2(32'hbbff164e),
	.w3(32'hbc5c1d6e),
	.w4(32'hbc895ffa),
	.w5(32'hbbae967c),
	.w6(32'hbc365188),
	.w7(32'hbc2da635),
	.w8(32'hba2638fb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb405788),
	.w1(32'hb934867b),
	.w2(32'hbc18f657),
	.w3(32'hbbad008b),
	.w4(32'hbb4a061e),
	.w5(32'h3aaf0dad),
	.w6(32'hbb7d000e),
	.w7(32'hbb38c8c9),
	.w8(32'hbb9073a4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4318c7),
	.w1(32'hbb14184f),
	.w2(32'hbae1e8ef),
	.w3(32'hbbb61649),
	.w4(32'hbb9d0a34),
	.w5(32'h3b447f9b),
	.w6(32'hbc45b33b),
	.w7(32'hbc0fe794),
	.w8(32'h3bc3ea93),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd9864),
	.w1(32'h3b2e2977),
	.w2(32'hbbd54472),
	.w3(32'h3bb84eb9),
	.w4(32'h3bb4169a),
	.w5(32'hbb58bea1),
	.w6(32'h3bba8c6f),
	.w7(32'h3b58671f),
	.w8(32'h3ae14edf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb863d77),
	.w1(32'h3b8c9a58),
	.w2(32'h3af30f2c),
	.w3(32'h3b8d14eb),
	.w4(32'h3be8186e),
	.w5(32'h3c31e871),
	.w6(32'h3bd7f9d1),
	.w7(32'h3bd908d8),
	.w8(32'hbad32c80),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44bf68),
	.w1(32'h3a3a7e97),
	.w2(32'h3cbecfc2),
	.w3(32'h3c7a50c1),
	.w4(32'h3ba6ae18),
	.w5(32'h3d0dc34f),
	.w6(32'h3b9d8663),
	.w7(32'hbbc052ac),
	.w8(32'h3cf64715),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd1dfe2),
	.w1(32'h3cbcb757),
	.w2(32'hbc782354),
	.w3(32'h3d0a14ac),
	.w4(32'h3cb78cae),
	.w5(32'hbcc29947),
	.w6(32'h3ccef2c1),
	.w7(32'h3c4521a0),
	.w8(32'hbc28b71a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7fc3ae),
	.w1(32'hbc03d39b),
	.w2(32'hbb595aad),
	.w3(32'hbc433b37),
	.w4(32'hbc92595a),
	.w5(32'h388faf3f),
	.w6(32'hbc8b68c4),
	.w7(32'hbc571812),
	.w8(32'hb8e2188a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc66e8e),
	.w1(32'hbc0e249d),
	.w2(32'hbb3014a3),
	.w3(32'hbba02da2),
	.w4(32'hbbe71131),
	.w5(32'hbb9ad484),
	.w6(32'hbb93568f),
	.w7(32'hbbf70a93),
	.w8(32'hbbaf5ae0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ebaf8),
	.w1(32'hbaf972af),
	.w2(32'hbb702548),
	.w3(32'hbaa90fad),
	.w4(32'hbb3b3866),
	.w5(32'h3b911925),
	.w6(32'hbbe33dd1),
	.w7(32'hbbbfb313),
	.w8(32'h3bc848aa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f5991),
	.w1(32'h3a29a07e),
	.w2(32'hbb4356f8),
	.w3(32'h3bdc1722),
	.w4(32'h3b0d2e16),
	.w5(32'hba9e9aeb),
	.w6(32'h3b2b0bc9),
	.w7(32'h3a956983),
	.w8(32'h3b162e10),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac45f23),
	.w1(32'hbab25fbf),
	.w2(32'h3c40ebe2),
	.w3(32'h3c271d19),
	.w4(32'h3a8260e1),
	.w5(32'h3b91a900),
	.w6(32'h3aaec267),
	.w7(32'h3a98c702),
	.w8(32'h3b7731fd),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff52b1),
	.w1(32'hbbaf0ee3),
	.w2(32'hbaf2c227),
	.w3(32'hbb0ba63f),
	.w4(32'hbbcf0474),
	.w5(32'hbaae743a),
	.w6(32'hbbdd0b2d),
	.w7(32'h3b885c6d),
	.w8(32'hbbb590a8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33fb22),
	.w1(32'hbb9454f7),
	.w2(32'hbb212047),
	.w3(32'h3b3fa0d2),
	.w4(32'h3965b628),
	.w5(32'h3b06d6d0),
	.w6(32'h3b21db34),
	.w7(32'hbafc8319),
	.w8(32'hbb18461d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9e28c),
	.w1(32'h3b2cc6f4),
	.w2(32'hbb967bec),
	.w3(32'hbc46977a),
	.w4(32'hbc4205a0),
	.w5(32'hbb3589c3),
	.w6(32'hbc4a57ad),
	.w7(32'hbbb83ea5),
	.w8(32'h3b655089),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6461e0),
	.w1(32'h3ad77110),
	.w2(32'h3a97c0a7),
	.w3(32'h3aaf98af),
	.w4(32'h3b3cd93d),
	.w5(32'h3ba58328),
	.w6(32'hbb50b76b),
	.w7(32'h3ab58a9f),
	.w8(32'h3bf88637),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fd94c),
	.w1(32'h3b3fc7e0),
	.w2(32'h3be7bafa),
	.w3(32'h3bef8871),
	.w4(32'h3b45a89f),
	.w5(32'h3c573472),
	.w6(32'h3c013085),
	.w7(32'h3bb8f042),
	.w8(32'h3b573078),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88d36e),
	.w1(32'h3c8acdb3),
	.w2(32'hbc6d6e23),
	.w3(32'h3c8d351b),
	.w4(32'h3c3be7f1),
	.w5(32'hbc68a01d),
	.w6(32'hba5fe06e),
	.w7(32'hbcb2d83c),
	.w8(32'hbc453100),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86fb41),
	.w1(32'hbc12c401),
	.w2(32'h3b54c4eb),
	.w3(32'hbc777ca5),
	.w4(32'hbc679dcf),
	.w5(32'hbaa0b028),
	.w6(32'hbcb65b8f),
	.w7(32'hbc73aef2),
	.w8(32'hbc08c98c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a23c69),
	.w1(32'hbb314f9b),
	.w2(32'hbc73f9f5),
	.w3(32'hbb01a69c),
	.w4(32'hbacbd4e1),
	.w5(32'hbc50252d),
	.w6(32'hbb1c3f5e),
	.w7(32'h398f1789),
	.w8(32'hbbcace55),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c7d21),
	.w1(32'hbb88401f),
	.w2(32'hbb4db883),
	.w3(32'hbb57e0fb),
	.w4(32'h3b9a3c89),
	.w5(32'hba0ee5d1),
	.w6(32'h39cc4143),
	.w7(32'h3bb40e68),
	.w8(32'h3a7ea65c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe63fd),
	.w1(32'hbb5576df),
	.w2(32'hbbbc3765),
	.w3(32'h3b026706),
	.w4(32'hbb367e55),
	.w5(32'hba9db414),
	.w6(32'h3b8f6fd9),
	.w7(32'hbc33af73),
	.w8(32'h3bd10538),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c5d8c),
	.w1(32'h3b8b436a),
	.w2(32'hbb294451),
	.w3(32'h3b1de26a),
	.w4(32'h3bade6e4),
	.w5(32'h3b63e288),
	.w6(32'h3c0a1da1),
	.w7(32'h3bbe478f),
	.w8(32'h3b843a43),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba583387),
	.w1(32'h38c4bc5c),
	.w2(32'hbc278883),
	.w3(32'h3b4897ed),
	.w4(32'hbba51e00),
	.w5(32'hbc215c60),
	.w6(32'h3b79dd49),
	.w7(32'h3b79571b),
	.w8(32'hbc94669e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99fb83),
	.w1(32'hbb8c78e7),
	.w2(32'h3c4c9ad7),
	.w3(32'hbc7434e5),
	.w4(32'hbc20be64),
	.w5(32'h3bb35c08),
	.w6(32'hbc8568b3),
	.w7(32'hbc35e256),
	.w8(32'h3c12414a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1f41b),
	.w1(32'h3bbc6728),
	.w2(32'hbc1d47a7),
	.w3(32'h3b59d95e),
	.w4(32'h3aedc626),
	.w5(32'hbc009582),
	.w6(32'h3ba3cec1),
	.w7(32'h3c2df4b2),
	.w8(32'h3a732767),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd93205),
	.w1(32'h3b78729e),
	.w2(32'hbc4774a9),
	.w3(32'h3b0540d0),
	.w4(32'h3c3c77a1),
	.w5(32'hbc5be127),
	.w6(32'h3c1f006e),
	.w7(32'h3c5a6b5b),
	.w8(32'h3bbfc147),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6dd18b),
	.w1(32'h3adcf2ed),
	.w2(32'hb922873b),
	.w3(32'hbc65afe2),
	.w4(32'hbbf27d59),
	.w5(32'hbb8b5970),
	.w6(32'hbc1825a1),
	.w7(32'hbc88e470),
	.w8(32'hbb75fc45),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22603a),
	.w1(32'hbb243efe),
	.w2(32'h3c0ffbea),
	.w3(32'hbad1ae9e),
	.w4(32'hbc0cef82),
	.w5(32'h3bcd62f8),
	.w6(32'hbb8132b3),
	.w7(32'hba0011eb),
	.w8(32'h3994e207),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2783ce),
	.w1(32'h3a438090),
	.w2(32'hbc13b694),
	.w3(32'h3b964434),
	.w4(32'hbb52eaaa),
	.w5(32'hbc9569e0),
	.w6(32'hbb67d45d),
	.w7(32'hbbd35821),
	.w8(32'hbc80251a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb0c28),
	.w1(32'hbc89781f),
	.w2(32'hbba3e5b4),
	.w3(32'hbd014a70),
	.w4(32'hbc9e91be),
	.w5(32'hbb608304),
	.w6(32'hbcced304),
	.w7(32'hbc41ce85),
	.w8(32'hbb66d157),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97678d),
	.w1(32'hba844218),
	.w2(32'h3ba02852),
	.w3(32'h3ba37142),
	.w4(32'h3bf88a81),
	.w5(32'h3b55f47f),
	.w6(32'hbb82bac4),
	.w7(32'h3b49ed3e),
	.w8(32'hbb19840d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2e951),
	.w1(32'hbaaf8a3d),
	.w2(32'h37f232f0),
	.w3(32'hbbea197b),
	.w4(32'hbc1178a8),
	.w5(32'h3b8c0818),
	.w6(32'hbc4caa28),
	.w7(32'hbb9d0941),
	.w8(32'h3b32cb54),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdafbeb),
	.w1(32'h3b9a1166),
	.w2(32'h3b5f2d96),
	.w3(32'h3c4a38c6),
	.w4(32'h3bab1558),
	.w5(32'h3be71760),
	.w6(32'h3bcfcc78),
	.w7(32'hbb6b8b68),
	.w8(32'h3b40df97),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc64f43),
	.w1(32'h3b9caaae),
	.w2(32'h3a53717a),
	.w3(32'h3c19f8f2),
	.w4(32'h3ae6629a),
	.w5(32'hb922da05),
	.w6(32'h3bdc49e1),
	.w7(32'h3af504bc),
	.w8(32'hba58d49f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab34d01),
	.w1(32'hbb556975),
	.w2(32'h39feb5d2),
	.w3(32'h3b533a71),
	.w4(32'hbab676f0),
	.w5(32'hbb683889),
	.w6(32'hbb9f0972),
	.w7(32'hbb64211a),
	.w8(32'hbb94798b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcba8f7),
	.w1(32'h3bc1b06e),
	.w2(32'h3a358577),
	.w3(32'hbbcb6da2),
	.w4(32'h3a8ef2cf),
	.w5(32'hba883ae6),
	.w6(32'hba9ef8a6),
	.w7(32'hbb5ab735),
	.w8(32'h3a8011b0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad26be7),
	.w1(32'h39e0b205),
	.w2(32'h3bb3b290),
	.w3(32'hbb432cc9),
	.w4(32'hbaced05d),
	.w5(32'h3b0e0455),
	.w6(32'hbae31b64),
	.w7(32'hba92f41f),
	.w8(32'hbc2c9375),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2eb0b4),
	.w1(32'h3b8de5e0),
	.w2(32'hb92344aa),
	.w3(32'h3bf56ee5),
	.w4(32'hba1487d6),
	.w5(32'hbc177121),
	.w6(32'hb9349bcd),
	.w7(32'hbc2a64c5),
	.w8(32'h3b81d947),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad324b1),
	.w1(32'hbc1516fb),
	.w2(32'h3aa6179b),
	.w3(32'hbcb3d837),
	.w4(32'hbb19475f),
	.w5(32'hbb647992),
	.w6(32'hbbcab06f),
	.w7(32'hbc228d58),
	.w8(32'hbb638fca),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98ce5e),
	.w1(32'h3b76ca91),
	.w2(32'h3b938d54),
	.w3(32'hba927a2a),
	.w4(32'h3ab648d8),
	.w5(32'h3ca07239),
	.w6(32'hbb7ddbe5),
	.w7(32'hbaf86437),
	.w8(32'h3c7955bb),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ec211),
	.w1(32'hbb847c8e),
	.w2(32'hb99cccb3),
	.w3(32'h3c67341e),
	.w4(32'hbaec0dfe),
	.w5(32'h3ba42470),
	.w6(32'h3c5d7977),
	.w7(32'hbb8768ee),
	.w8(32'h3afde842),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc030fda),
	.w1(32'hbc2bad9c),
	.w2(32'h3b2de60c),
	.w3(32'hbb3c5189),
	.w4(32'hbc580c59),
	.w5(32'hba0cdcbe),
	.w6(32'hbb87c643),
	.w7(32'hbca03b8d),
	.w8(32'hbb8a5f70),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66ca21),
	.w1(32'h3bc3ecb2),
	.w2(32'hbb8644cc),
	.w3(32'h3a70d519),
	.w4(32'h3bbcaac3),
	.w5(32'hbbf55d0d),
	.w6(32'hba255921),
	.w7(32'h3b428e44),
	.w8(32'hbbcff6c8),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b4247),
	.w1(32'hbb70766a),
	.w2(32'h3a3e638b),
	.w3(32'hbb28443a),
	.w4(32'hbb386d2d),
	.w5(32'h3b801628),
	.w6(32'hbcab3941),
	.w7(32'hbc2a18b2),
	.w8(32'hbaac7628),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b77be),
	.w1(32'h3957298d),
	.w2(32'hbc42809b),
	.w3(32'h3af232e3),
	.w4(32'hba0bd88e),
	.w5(32'hbcb59dcf),
	.w6(32'h39fc8a80),
	.w7(32'h3b01ef5c),
	.w8(32'hbc9a8565),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38f1f9),
	.w1(32'hbcab8fcc),
	.w2(32'h3ab28873),
	.w3(32'hbcf00900),
	.w4(32'hbcf87b46),
	.w5(32'hbbea6329),
	.w6(32'hbc95b3dc),
	.w7(32'hbc460eed),
	.w8(32'hbbdc266e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba153ba7),
	.w1(32'h3bdcb343),
	.w2(32'h3c4b7455),
	.w3(32'hbbb9a9e8),
	.w4(32'h3ada4c1e),
	.w5(32'h3b4fb9d6),
	.w6(32'hbbd225c4),
	.w7(32'hbafb25d3),
	.w8(32'h3c614ff3),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c94fb),
	.w1(32'hbab912c3),
	.w2(32'h3c01626e),
	.w3(32'h3b33b48b),
	.w4(32'hb8b7cc6c),
	.w5(32'hbbcae1fc),
	.w6(32'h3b715635),
	.w7(32'h3b2e7c31),
	.w8(32'hbcb2ca52),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda3dc4),
	.w1(32'h3bf6d268),
	.w2(32'hbc2e0b3c),
	.w3(32'h3c0b8851),
	.w4(32'h3bbab39f),
	.w5(32'hbbe96761),
	.w6(32'hbc25edaf),
	.w7(32'hbadbb755),
	.w8(32'h3bc5cbab),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f66d0),
	.w1(32'h39f7296f),
	.w2(32'h3c00146a),
	.w3(32'hbb6f9a66),
	.w4(32'h3c035d05),
	.w5(32'h3c089eec),
	.w6(32'h3b0d81d7),
	.w7(32'h3c5551e3),
	.w8(32'h3ca9a2f8),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b526683),
	.w1(32'hba821f62),
	.w2(32'h3c8e54d9),
	.w3(32'h3bde9aff),
	.w4(32'hbbd896ce),
	.w5(32'h3b91c59f),
	.w6(32'h3c4f385b),
	.w7(32'hba9b3529),
	.w8(32'hbc44fefd),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc01d5),
	.w1(32'h3be328cf),
	.w2(32'h3b727d34),
	.w3(32'hbc1c95bb),
	.w4(32'hbc1ec8c0),
	.w5(32'h3bc64207),
	.w6(32'hbccb1ef6),
	.w7(32'hbce35f90),
	.w8(32'h3ab12f43),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56786f),
	.w1(32'hba8fe3a1),
	.w2(32'hbb95b3a4),
	.w3(32'h3960e951),
	.w4(32'hbba57c3f),
	.w5(32'hbbe5db56),
	.w6(32'hb9e237f4),
	.w7(32'hbb2b7f2d),
	.w8(32'hbbaa1ed3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d5224),
	.w1(32'h3c85a246),
	.w2(32'hbb5bc198),
	.w3(32'h3c3a17b2),
	.w4(32'h3d04ff03),
	.w5(32'hbb9695a7),
	.w6(32'hb94b53af),
	.w7(32'h3c8fd51d),
	.w8(32'hbc264419),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996929a),
	.w1(32'hbbaf5215),
	.w2(32'hbbd3a71a),
	.w3(32'hbbdcfe21),
	.w4(32'h3c3cac48),
	.w5(32'hbcce0894),
	.w6(32'h3b0a30cb),
	.w7(32'h3bdb4f10),
	.w8(32'hbcab5998),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca2c29),
	.w1(32'h3ca1dd7c),
	.w2(32'h3beb4ccb),
	.w3(32'hbcde0bf6),
	.w4(32'hbaee227b),
	.w5(32'h3b448419),
	.w6(32'hbd335aca),
	.w7(32'hbc2b7bdb),
	.w8(32'hbbfd1827),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fa79b),
	.w1(32'h3c95bb32),
	.w2(32'hba749839),
	.w3(32'hbc8e3ec4),
	.w4(32'h3b27e4bc),
	.w5(32'h3adf327a),
	.w6(32'hbcfa98bc),
	.w7(32'hbc8213a6),
	.w8(32'h3b34ac55),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0eb1e2),
	.w1(32'hbb2c740d),
	.w2(32'hb92a34a5),
	.w3(32'hb968729f),
	.w4(32'hbb4bc18d),
	.w5(32'h3c71f5ac),
	.w6(32'hba9b602d),
	.w7(32'hba931cad),
	.w8(32'h3aa2b29c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81840f),
	.w1(32'hbbc2b684),
	.w2(32'h3c7280ea),
	.w3(32'h3c7d0d87),
	.w4(32'h3b4bbd61),
	.w5(32'h3bea09b8),
	.w6(32'hba684adf),
	.w7(32'hbb2eb635),
	.w8(32'hbcca1d73),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dd4a7),
	.w1(32'h3c15533f),
	.w2(32'h3c17fdf9),
	.w3(32'hb99ac012),
	.w4(32'h3b7c57ab),
	.w5(32'hbc6662bb),
	.w6(32'hbc863652),
	.w7(32'h3b56642e),
	.w8(32'hbc5e6ea9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb337424),
	.w1(32'h39419566),
	.w2(32'h3c76486c),
	.w3(32'hbc08c515),
	.w4(32'h3b8807ef),
	.w5(32'h3bbeebe3),
	.w6(32'h3b71ad1f),
	.w7(32'h3c8b9849),
	.w8(32'hbcd69d61),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ed617),
	.w1(32'h3bdc280e),
	.w2(32'hbbaa329e),
	.w3(32'h3bb40625),
	.w4(32'hbb1c447f),
	.w5(32'h3bc05765),
	.w6(32'hbc8a0e4c),
	.w7(32'hbafa9fa4),
	.w8(32'h3c780d4c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf19b02),
	.w1(32'hbc45ae3f),
	.w2(32'hbb87ac54),
	.w3(32'h3bc4b132),
	.w4(32'h3abd5ee5),
	.w5(32'hbbf6c4bf),
	.w6(32'h3c8f2a22),
	.w7(32'h3b69ce9b),
	.w8(32'h3bff4683),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5e358),
	.w1(32'hbc26b177),
	.w2(32'hbc774d14),
	.w3(32'hbc813a19),
	.w4(32'hbbd4e7b4),
	.w5(32'hbb525584),
	.w6(32'h3c9a3300),
	.w7(32'hbab86f60),
	.w8(32'h3c0e96cb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc617cc2),
	.w1(32'hbbb5a263),
	.w2(32'h3b274bb9),
	.w3(32'hbb102007),
	.w4(32'hbb20ea59),
	.w5(32'hbc6f121d),
	.w6(32'h3c995331),
	.w7(32'hbb04f133),
	.w8(32'hbd0ef390),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa298e5),
	.w1(32'hbb30678c),
	.w2(32'h3b5ed830),
	.w3(32'hbc39e8d4),
	.w4(32'h3b443397),
	.w5(32'hba69682c),
	.w6(32'hbccc4d74),
	.w7(32'hbaf39059),
	.w8(32'h39aafca8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb844fdb),
	.w1(32'h3b019821),
	.w2(32'hbabb72e8),
	.w3(32'hbbfa554e),
	.w4(32'h3c02d66b),
	.w5(32'hbb2f7265),
	.w6(32'hbc0df713),
	.w7(32'h3bebc6c4),
	.w8(32'h3ce130aa),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdad062),
	.w1(32'hbbfd0bbf),
	.w2(32'hbb1ca3ef),
	.w3(32'hbb964e5a),
	.w4(32'hbc0c842b),
	.w5(32'h3b88cf4b),
	.w6(32'h3ce2b244),
	.w7(32'h3cbc25fe),
	.w8(32'h3b0b65d6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5fef4),
	.w1(32'hbbc3705f),
	.w2(32'h3c08749c),
	.w3(32'h3af3cf72),
	.w4(32'hbbb728ef),
	.w5(32'h3c19daf7),
	.w6(32'h3b097633),
	.w7(32'hbbf84705),
	.w8(32'h3b093828),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b854e1b),
	.w1(32'hbb3bd917),
	.w2(32'h3bd2e170),
	.w3(32'h3bde5a08),
	.w4(32'hbb468ecb),
	.w5(32'hbbb1f1a7),
	.w6(32'h38e9904e),
	.w7(32'hbb9da370),
	.w8(32'hbc748991),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a93bb),
	.w1(32'h3be8956a),
	.w2(32'h3bc8b2dd),
	.w3(32'hbc024e31),
	.w4(32'h3aef994c),
	.w5(32'h3be0e5a1),
	.w6(32'hbcdbd1ad),
	.w7(32'hbc09a742),
	.w8(32'h3b1786be),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81c982),
	.w1(32'h3b40d987),
	.w2(32'h3ad96bfa),
	.w3(32'h3c0ae0a6),
	.w4(32'hb8f8c403),
	.w5(32'hb90c8acb),
	.w6(32'hbb07ac11),
	.w7(32'hba914184),
	.w8(32'hbb419bc3),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf9169),
	.w1(32'hbb14b6a1),
	.w2(32'hbbc0a693),
	.w3(32'h3ac156d2),
	.w4(32'h3b943a85),
	.w5(32'hbac2f305),
	.w6(32'h3baaad95),
	.w7(32'h3c0dddc3),
	.w8(32'h3c076aa3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d1c38),
	.w1(32'hbb22ef1b),
	.w2(32'hb925b22b),
	.w3(32'hbbda71e3),
	.w4(32'hba7e0cd3),
	.w5(32'h3b89456f),
	.w6(32'h3c033c1b),
	.w7(32'h3be711af),
	.w8(32'h3bec3acb),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397c9b3e),
	.w1(32'hbac7cc5e),
	.w2(32'h3b545e0c),
	.w3(32'h3bc6544b),
	.w4(32'h3b327355),
	.w5(32'h3a35280d),
	.w6(32'h3c1df1e7),
	.w7(32'h3bdbd9f7),
	.w8(32'hbb9fe872),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e51a7),
	.w1(32'h39416f9d),
	.w2(32'h3c25d5cd),
	.w3(32'hb9ffad3e),
	.w4(32'hbb6dbb9c),
	.w5(32'hbad0aa58),
	.w6(32'hbaf41f3e),
	.w7(32'hbb65b66c),
	.w8(32'hbc8e7f75),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a24b6),
	.w1(32'h3bdd40ea),
	.w2(32'h3be528ca),
	.w3(32'hbbcebe2b),
	.w4(32'h3b28306a),
	.w5(32'h3abbad4e),
	.w6(32'hbc912ea6),
	.w7(32'h3b2d0de4),
	.w8(32'hbbb1909d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa9519),
	.w1(32'hba57b4b3),
	.w2(32'hbc1389d6),
	.w3(32'h3c0311fd),
	.w4(32'h3b8cde47),
	.w5(32'hbc0559fd),
	.w6(32'hbbd21718),
	.w7(32'h3b4569ca),
	.w8(32'hbb59cc4d),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6c7db),
	.w1(32'hbc074af3),
	.w2(32'h3c120207),
	.w3(32'hbb7a3e0e),
	.w4(32'hbbcac318),
	.w5(32'hbb282801),
	.w6(32'h390f7b6b),
	.w7(32'hbb5cb523),
	.w8(32'hbc514fea),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c620d63),
	.w1(32'h3c1b0370),
	.w2(32'h3b9952bd),
	.w3(32'h3b795b8d),
	.w4(32'h3b17c25d),
	.w5(32'h3b707727),
	.w6(32'hbb3cf765),
	.w7(32'hbb0cabc8),
	.w8(32'hbb47320f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f6087),
	.w1(32'h3c03daf9),
	.w2(32'hbbc4a265),
	.w3(32'h3baa8508),
	.w4(32'h3bbb2091),
	.w5(32'hbc7d78a3),
	.w6(32'h399009a6),
	.w7(32'h3b991616),
	.w8(32'hbc91319f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0433f3),
	.w1(32'h3b6c4ca2),
	.w2(32'h3b6d8c02),
	.w3(32'hbca3e3ce),
	.w4(32'hbc0f33d5),
	.w5(32'hbb642649),
	.w6(32'hbccc0038),
	.w7(32'hbc4fae6c),
	.w8(32'hbabf86c6),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba68a49),
	.w1(32'hbc0f9dad),
	.w2(32'h3ae35504),
	.w3(32'hb9ba61fc),
	.w4(32'hbc16407c),
	.w5(32'h3b9591b2),
	.w6(32'h3b6d2f3e),
	.w7(32'hbba7c62b),
	.w8(32'h3ac91690),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a4145a),
	.w1(32'hba8c4dd7),
	.w2(32'h3986b777),
	.w3(32'h39d3e065),
	.w4(32'hbbab252b),
	.w5(32'hbbbcf508),
	.w6(32'hbb5b7199),
	.w7(32'hbbae03f4),
	.w8(32'hbbe857f4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb909ca2),
	.w1(32'hbbc5f6a2),
	.w2(32'h3b3aba2a),
	.w3(32'hbc285f53),
	.w4(32'hbc208958),
	.w5(32'hba0ad0f0),
	.w6(32'hbc72cee4),
	.w7(32'hbc2aee0a),
	.w8(32'hbbd15d92),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad295f8),
	.w1(32'hbb5fe6bb),
	.w2(32'h3b27655a),
	.w3(32'h3b025d80),
	.w4(32'h3b387a5d),
	.w5(32'hbb2c8362),
	.w6(32'h3bf55c43),
	.w7(32'h3b69e0a9),
	.w8(32'h3bf29490),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd05ad2),
	.w1(32'hbb86ce31),
	.w2(32'h3b60a9bb),
	.w3(32'h3c1692f9),
	.w4(32'hbb0feea2),
	.w5(32'hbbba8d80),
	.w6(32'h3c706330),
	.w7(32'h3bb665f5),
	.w8(32'hbb8dd212),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb706aa8),
	.w1(32'h3c50a1e3),
	.w2(32'hbb2809cd),
	.w3(32'hbcde5672),
	.w4(32'hbbe80536),
	.w5(32'hbb045c4e),
	.w6(32'hbcd2ece3),
	.w7(32'hbc9f3fbb),
	.w8(32'hb815f8e9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a3ff9),
	.w1(32'h3709a0ab),
	.w2(32'h3ba6c41e),
	.w3(32'hbb2fdddd),
	.w4(32'hba7f2335),
	.w5(32'hb9e9a74a),
	.w6(32'h39974a30),
	.w7(32'hb9207719),
	.w8(32'hbad0a118),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8843e2),
	.w1(32'h3b02331d),
	.w2(32'h3bfae8ec),
	.w3(32'hbb8c6d07),
	.w4(32'hb9dbb0ad),
	.w5(32'h3b6b77fa),
	.w6(32'hbba307a0),
	.w7(32'hb9f5680a),
	.w8(32'h3a1a49e4),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb76ae1),
	.w1(32'h3ae0213a),
	.w2(32'hbb27e9b9),
	.w3(32'h3b22452e),
	.w4(32'hbb3fb34e),
	.w5(32'hbcab8e63),
	.w6(32'h3ad87d27),
	.w7(32'hbaa4784e),
	.w8(32'hbc4be57a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffc1dc),
	.w1(32'hbbb7c27e),
	.w2(32'h3b2eacbb),
	.w3(32'hbca46140),
	.w4(32'hbca1c2db),
	.w5(32'hbc204ea4),
	.w6(32'hbcc82d23),
	.w7(32'hbbe77bbe),
	.w8(32'hbc1a0283),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13fded),
	.w1(32'h3cd5c9fd),
	.w2(32'hbbf6318c),
	.w3(32'hbcaa8109),
	.w4(32'h3b808087),
	.w5(32'hbc4b4bef),
	.w6(32'hbd0baedf),
	.w7(32'hbcfbb45a),
	.w8(32'hbc068d36),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac46838),
	.w1(32'h3b6da870),
	.w2(32'hbaa11ee5),
	.w3(32'hbc795353),
	.w4(32'hbbb27e9c),
	.w5(32'hbc8f3447),
	.w6(32'hbcaeae8f),
	.w7(32'hbca8d566),
	.w8(32'hbd0c7d04),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8152be),
	.w1(32'h3c1df935),
	.w2(32'h3b8736e3),
	.w3(32'hbca42132),
	.w4(32'h3c4524c0),
	.w5(32'h3bd3984e),
	.w6(32'hbbfc428c),
	.w7(32'h3c680dd7),
	.w8(32'h3b3cf196),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b51a1),
	.w1(32'h3bdd1c19),
	.w2(32'h3b874bd9),
	.w3(32'h39cacabc),
	.w4(32'h3bea91bf),
	.w5(32'h3ae12fe6),
	.w6(32'hb86dad30),
	.w7(32'h3b909e68),
	.w8(32'h3a421d50),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cb4f2),
	.w1(32'h39c307aa),
	.w2(32'h3c51f1e2),
	.w3(32'h3ae9a066),
	.w4(32'h3b85b515),
	.w5(32'h3be858bf),
	.w6(32'h3b1183a8),
	.w7(32'h381ae1d1),
	.w8(32'hbc9c9dd3),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82c40c),
	.w1(32'h3c2b41d4),
	.w2(32'h3a38a049),
	.w3(32'h3bd47f30),
	.w4(32'hba971b10),
	.w5(32'h3c33d50c),
	.w6(32'hbca63733),
	.w7(32'h3b89a7cc),
	.w8(32'h3c03b2cf),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fdeac),
	.w1(32'hbb08f6bf),
	.w2(32'h3aee6c47),
	.w3(32'h3bea2a7e),
	.w4(32'h3ba047e7),
	.w5(32'hbb9685ba),
	.w6(32'h3c72593e),
	.w7(32'h3b8eaace),
	.w8(32'hbab83216),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb964e18),
	.w1(32'hb903376e),
	.w2(32'h3af0daeb),
	.w3(32'hbb1bd5c6),
	.w4(32'hbbab1d10),
	.w5(32'h3b8db23b),
	.w6(32'h3ad97a53),
	.w7(32'hbbc88fa2),
	.w8(32'h3c605292),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1b225),
	.w1(32'hbbbfea22),
	.w2(32'hbc0060e3),
	.w3(32'h3b63683c),
	.w4(32'hbbada08b),
	.w5(32'hbc3f48f5),
	.w6(32'h3c4bef58),
	.w7(32'hbb322ad3),
	.w8(32'hbc0ee5d5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb883be9),
	.w1(32'h39b71523),
	.w2(32'hbac2cb21),
	.w3(32'hbc1d215d),
	.w4(32'hbb307ddb),
	.w5(32'hbb935736),
	.w6(32'hbbe8dc69),
	.w7(32'h389eba0b),
	.w8(32'hbbf4341b),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60db33),
	.w1(32'hbbc81a8b),
	.w2(32'h3c24b7f9),
	.w3(32'hbbe0ffd6),
	.w4(32'hbc253f83),
	.w5(32'h3b5b0263),
	.w6(32'hbc19f11e),
	.w7(32'hbc45d98e),
	.w8(32'hbb3cb222),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18adca),
	.w1(32'h3c0544c4),
	.w2(32'hbac4be9d),
	.w3(32'h3bd7a8e1),
	.w4(32'h3bd26613),
	.w5(32'h3c74312f),
	.w6(32'hbb5f04ab),
	.w7(32'h39433b58),
	.w8(32'h3ba4f95a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f7cec),
	.w1(32'hbc6d170b),
	.w2(32'hbbc1bbe6),
	.w3(32'h3c51db07),
	.w4(32'h3c1a5cce),
	.w5(32'hbb98543c),
	.w6(32'h3b180548),
	.w7(32'h3b9d3fcf),
	.w8(32'hbc0d5e0a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14c4c7),
	.w1(32'hbc0cf280),
	.w2(32'h3c4d1c30),
	.w3(32'hbbcbf48d),
	.w4(32'hbb39f336),
	.w5(32'hbb4c5b6c),
	.w6(32'hbc50067e),
	.w7(32'hbc1c1e26),
	.w8(32'h3b419ebc),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4dfa2c),
	.w1(32'h3c10e99d),
	.w2(32'hbb933f9e),
	.w3(32'hbc468366),
	.w4(32'hbb013e0a),
	.w5(32'h3beec1f7),
	.w6(32'hbcb46174),
	.w7(32'hbccd1de3),
	.w8(32'h3c2d0dbb),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9182df),
	.w1(32'hbc69188b),
	.w2(32'hba875f22),
	.w3(32'h3c79bd3c),
	.w4(32'hbaf91c46),
	.w5(32'hbb7b3a6f),
	.w6(32'h3c0f5027),
	.w7(32'h3ba3e382),
	.w8(32'hbb1dccd6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7e055),
	.w1(32'h3c131da9),
	.w2(32'h3a43f2be),
	.w3(32'hbba1637a),
	.w4(32'h3bf0f2a1),
	.w5(32'h3c7c7e4a),
	.w6(32'hbbaf9c41),
	.w7(32'h3ada71cd),
	.w8(32'h3c1d945c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafa8f3),
	.w1(32'hbbad7e96),
	.w2(32'hbbd357bf),
	.w3(32'h3c16b4ab),
	.w4(32'hbb62f684),
	.w5(32'h3c193533),
	.w6(32'h3aca5d60),
	.w7(32'hbb753dc3),
	.w8(32'h3ca9d0bf),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac883ca),
	.w1(32'hb9712111),
	.w2(32'h3ba7fe8a),
	.w3(32'h3c876821),
	.w4(32'hb955d127),
	.w5(32'h3c67fb19),
	.w6(32'h3cb23087),
	.w7(32'h3c1cd44f),
	.w8(32'h3a93b840),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0140dd),
	.w1(32'h3b584ee4),
	.w2(32'hbb84e747),
	.w3(32'h3c9ac968),
	.w4(32'h3c3944bc),
	.w5(32'h3a570163),
	.w6(32'h3b920d9f),
	.w7(32'hbb048760),
	.w8(32'hbb97a76f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fb87f),
	.w1(32'h3c06bf48),
	.w2(32'hb9ae3901),
	.w3(32'h3b589837),
	.w4(32'h3c6bbdd3),
	.w5(32'hbc802b24),
	.w6(32'h3b7fd1b6),
	.w7(32'h3c377474),
	.w8(32'hbd11aff7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b92fb),
	.w1(32'h3cc94c82),
	.w2(32'hba97768b),
	.w3(32'hbcdcf6f7),
	.w4(32'h3b8ca755),
	.w5(32'hba098da2),
	.w6(32'hbd3338a6),
	.w7(32'h3b68978d),
	.w8(32'hbaf1adac),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d4e6d),
	.w1(32'h3c19b901),
	.w2(32'h3b6eca84),
	.w3(32'h3b1d5a1d),
	.w4(32'h3c3e91c5),
	.w5(32'hbb65b9a6),
	.w6(32'h3b683e45),
	.w7(32'h3be4ff17),
	.w8(32'hbc1895c9),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d705b),
	.w1(32'h3c32d207),
	.w2(32'hba8bab21),
	.w3(32'h3adaa6c9),
	.w4(32'h3c06ba3d),
	.w5(32'h3baf969c),
	.w6(32'hbb08dc87),
	.w7(32'h3a97df93),
	.w8(32'h3ab3e3b4),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384c6f85),
	.w1(32'h3ba96e38),
	.w2(32'hbc254174),
	.w3(32'hbafa9af7),
	.w4(32'h3b932e87),
	.w5(32'hbc8e9ff2),
	.w6(32'hbb7984cd),
	.w7(32'hbbd9036b),
	.w8(32'hbc6e5189),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5e81e),
	.w1(32'h3b4246a8),
	.w2(32'h396ca71c),
	.w3(32'hbc809393),
	.w4(32'hba9f06ab),
	.w5(32'h3c7a9385),
	.w6(32'hbca567aa),
	.w7(32'hbbb9daf4),
	.w8(32'h3c1895ba),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b294d76),
	.w1(32'hbb1b36c3),
	.w2(32'h3c9c4355),
	.w3(32'h3bc915fd),
	.w4(32'hbc0de29f),
	.w5(32'h3a667e5c),
	.w6(32'h3be45716),
	.w7(32'hbc011487),
	.w8(32'hbbb4afab),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c51f9),
	.w1(32'h3c1ba829),
	.w2(32'h398f4df5),
	.w3(32'hbc1ff9b3),
	.w4(32'h3b1529f1),
	.w5(32'hbbaf1d40),
	.w6(32'hbcaaf121),
	.w7(32'hbcc01e85),
	.w8(32'hbc686864),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8d478),
	.w1(32'h3c62b3b4),
	.w2(32'hbb89e8a7),
	.w3(32'hbb8956ec),
	.w4(32'h3aefad95),
	.w5(32'hbc4e93b3),
	.w6(32'hbc7ea05c),
	.w7(32'hbbc02bbc),
	.w8(32'hbc8858c9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7576c),
	.w1(32'h3bb98381),
	.w2(32'h3c09c94b),
	.w3(32'hbb48255d),
	.w4(32'h3c19ea35),
	.w5(32'h3c933bbb),
	.w6(32'hbca863f3),
	.w7(32'hb9e4f6d7),
	.w8(32'h3af8f843),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39ca72),
	.w1(32'h3aa38204),
	.w2(32'hbbc61c55),
	.w3(32'h3c48f2bc),
	.w4(32'h3b00e1ff),
	.w5(32'hbbc59f48),
	.w6(32'hbc310f40),
	.w7(32'hbc8d9215),
	.w8(32'h3a9e0df5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0fb09),
	.w1(32'hbb0556b7),
	.w2(32'h3acf9401),
	.w3(32'h3be57418),
	.w4(32'hba111073),
	.w5(32'hbb988985),
	.w6(32'hb8c0cdce),
	.w7(32'hba22cf97),
	.w8(32'hbc0db3ea),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9517bd),
	.w1(32'h3a970ba2),
	.w2(32'h3a905b2b),
	.w3(32'hbad786ac),
	.w4(32'hbb3d1185),
	.w5(32'h3b90782d),
	.w6(32'hbbe6735b),
	.w7(32'hbbc5b2db),
	.w8(32'h3b97c235),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89d5e6),
	.w1(32'h3acf908a),
	.w2(32'h38ab9e7d),
	.w3(32'h3b0e744a),
	.w4(32'h3b9ce9e6),
	.w5(32'h3b79bd24),
	.w6(32'h3afbe9a7),
	.w7(32'hbbc33a58),
	.w8(32'h3c117ff1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b055b),
	.w1(32'hbb10c206),
	.w2(32'hbbbb0dee),
	.w3(32'h3a852c11),
	.w4(32'h3adc8bce),
	.w5(32'h3bcbe8fe),
	.w6(32'h3c342f52),
	.w7(32'h3c22bf76),
	.w8(32'h3c3cd6f1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe01ae4),
	.w1(32'hbac576bc),
	.w2(32'h3aaa2d7e),
	.w3(32'h3c0c75d9),
	.w4(32'hbc3dd3d0),
	.w5(32'h3c9ca1a2),
	.w6(32'h3cae2477),
	.w7(32'h3b2c6cb9),
	.w8(32'h3ca3c60b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cff21),
	.w1(32'h3b0ffaf2),
	.w2(32'h3c0dd916),
	.w3(32'h3b5b4ccd),
	.w4(32'hbb3f573d),
	.w5(32'h3c0d9c01),
	.w6(32'h3c82393b),
	.w7(32'h3babe975),
	.w8(32'hba2cc209),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be88b1a),
	.w1(32'h3bbb4c3f),
	.w2(32'hbb4a4c8c),
	.w3(32'hbb22785f),
	.w4(32'h3ba99e7d),
	.w5(32'hbb1ee050),
	.w6(32'hbb97a6b5),
	.w7(32'hbc14c61b),
	.w8(32'h39f0db08),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2a64a),
	.w1(32'h3ad88aa8),
	.w2(32'h39db3e17),
	.w3(32'h3b184058),
	.w4(32'h3b63bc23),
	.w5(32'hbba2f57a),
	.w6(32'h3b00db9e),
	.w7(32'h3bd10fae),
	.w8(32'hbb631d21),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31ba02),
	.w1(32'h3aec8cf7),
	.w2(32'h3b0d7843),
	.w3(32'hbb300720),
	.w4(32'h3a7cac09),
	.w5(32'h3bc1c008),
	.w6(32'hbba29d5a),
	.w7(32'hb9e54f0b),
	.w8(32'h3a3f5a8a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96526a),
	.w1(32'h3c694cde),
	.w2(32'h3b2c135c),
	.w3(32'hbbc5ec11),
	.w4(32'h3c8fdd85),
	.w5(32'h3b873d84),
	.w6(32'hbcaeb4b6),
	.w7(32'hbabf127e),
	.w8(32'h3be9c6dc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a5bf8),
	.w1(32'h3be4990f),
	.w2(32'h3b4ea92d),
	.w3(32'h3b8c0a13),
	.w4(32'h3bce8494),
	.w5(32'hbc11a520),
	.w6(32'h3bebc61b),
	.w7(32'h3b2e1f65),
	.w8(32'hbcccd329),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6e1bd),
	.w1(32'h3c21a70c),
	.w2(32'h3a8fa59e),
	.w3(32'hbc254fdd),
	.w4(32'h3c202138),
	.w5(32'hbbb7dd47),
	.w6(32'hbca74992),
	.w7(32'h3bc44927),
	.w8(32'hbcc545d8),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8190b),
	.w1(32'h3c3cc186),
	.w2(32'hbb29c8fd),
	.w3(32'hbc654d7d),
	.w4(32'hb9f8f4e7),
	.w5(32'hbc6a6692),
	.w6(32'hbd03abd6),
	.w7(32'h3aa10829),
	.w8(32'hbc99ac82),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a8730),
	.w1(32'h3ca18975),
	.w2(32'h3c5688b6),
	.w3(32'hbc9292a4),
	.w4(32'h3b12c532),
	.w5(32'h3c348886),
	.w6(32'hbcd3dd9d),
	.w7(32'h3931a7fc),
	.w8(32'hbbca1dd6),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule