module layer_6_featuremap_120(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11c4ea),
	.w1(32'h39607906),
	.w2(32'h3bc3b6e0),
	.w3(32'hbbf74f73),
	.w4(32'hbb858b7b),
	.w5(32'hbaa27e87),
	.w6(32'h3a59da94),
	.w7(32'h3c3be1b5),
	.w8(32'h3c0305dd),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fa12c),
	.w1(32'hbc21d2ac),
	.w2(32'hbbb5228f),
	.w3(32'h3b0fe971),
	.w4(32'h3b970ab4),
	.w5(32'h3af32aa8),
	.w6(32'h3ca37b48),
	.w7(32'h3c8c3510),
	.w8(32'h3c92a4ae),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d56b8),
	.w1(32'h3ac27cb8),
	.w2(32'h3bc646c0),
	.w3(32'h3bc9cd7f),
	.w4(32'hbcdc8212),
	.w5(32'hbc95a9fe),
	.w6(32'hbc78ae88),
	.w7(32'hbc971c3b),
	.w8(32'hbc00a128),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f6adb),
	.w1(32'hbb967bc1),
	.w2(32'hbbb11513),
	.w3(32'hbacb7594),
	.w4(32'h3adcd550),
	.w5(32'hbae9eb35),
	.w6(32'hb8c57da7),
	.w7(32'hbb0dd818),
	.w8(32'hbba24e9b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb0281),
	.w1(32'h3cda7e83),
	.w2(32'h3d452437),
	.w3(32'hbce0e60e),
	.w4(32'hbd2ef238),
	.w5(32'hbca538b1),
	.w6(32'h3c919d0a),
	.w7(32'h3d34aebc),
	.w8(32'h3d475368),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce87d26),
	.w1(32'hbb2bf6a6),
	.w2(32'h3a6133bd),
	.w3(32'hbc64361b),
	.w4(32'hbc6d3d0c),
	.w5(32'hbc14b2a5),
	.w6(32'hbc0554bf),
	.w7(32'hba4947c4),
	.w8(32'h3b44f5d2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c355746),
	.w1(32'hbb03ee5e),
	.w2(32'hbacdcc52),
	.w3(32'h3c992e93),
	.w4(32'h3c59faf7),
	.w5(32'h3b9edc23),
	.w6(32'h3c0494f2),
	.w7(32'hbad1248f),
	.w8(32'h3895c93f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03238c),
	.w1(32'hbc68464b),
	.w2(32'hbcc8652b),
	.w3(32'hbc50d8f9),
	.w4(32'h3c5bf222),
	.w5(32'h3cacee66),
	.w6(32'hbbfa7fb9),
	.w7(32'hba4089ec),
	.w8(32'h3c15cf06),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ef0a1),
	.w1(32'hbc1e566c),
	.w2(32'hbd337b2d),
	.w3(32'hbc289a70),
	.w4(32'h3c0590e5),
	.w5(32'h3c7d76fb),
	.w6(32'h3cc89d5d),
	.w7(32'h3d0b9220),
	.w8(32'h3caaaba4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcedfebf),
	.w1(32'hbb11e6b3),
	.w2(32'hbb2e0319),
	.w3(32'hbb8fbc5e),
	.w4(32'hb9f4e9a1),
	.w5(32'h397ff16c),
	.w6(32'h3b5ef9b3),
	.w7(32'h3c277a15),
	.w8(32'h3ba0751e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ca352),
	.w1(32'hbbd4f2fd),
	.w2(32'h3a7b2a6d),
	.w3(32'hbc64a830),
	.w4(32'hbc8d4262),
	.w5(32'hbc02aba4),
	.w6(32'hbcd258bd),
	.w7(32'hbc9d0d47),
	.w8(32'hbc6c2b64),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42430d),
	.w1(32'hbc0d274c),
	.w2(32'hbc1491d9),
	.w3(32'hbbf53ea6),
	.w4(32'hbba962aa),
	.w5(32'hba920acb),
	.w6(32'h3c450d94),
	.w7(32'h3c88ef77),
	.w8(32'h3c87c773),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67022c),
	.w1(32'hbb8a7c71),
	.w2(32'hbb087437),
	.w3(32'h3b362075),
	.w4(32'h39e848e5),
	.w5(32'hbb52aedf),
	.w6(32'hb83565ac),
	.w7(32'h3a070453),
	.w8(32'hbb945025),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe28893),
	.w1(32'hbc03c5f5),
	.w2(32'h3b373602),
	.w3(32'hbca62afa),
	.w4(32'hbcfe2374),
	.w5(32'hbc8a3450),
	.w6(32'h39508291),
	.w7(32'hbc52da6d),
	.w8(32'hbbb9bdf2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a908c),
	.w1(32'h3b453969),
	.w2(32'h3c830350),
	.w3(32'hbbcb7556),
	.w4(32'h3b500d04),
	.w5(32'hbb12e27b),
	.w6(32'h3bbd2f6a),
	.w7(32'h3c702a83),
	.w8(32'h3a74922e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00f960),
	.w1(32'hbac0d51d),
	.w2(32'h3ab53cc0),
	.w3(32'hbbab3a99),
	.w4(32'hbbddb7dc),
	.w5(32'hbbe5a92c),
	.w6(32'hba9d0180),
	.w7(32'hbb7e0ddc),
	.w8(32'h3ab070f9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99baa0d),
	.w1(32'h3bb1286b),
	.w2(32'hbb6b4fff),
	.w3(32'h3c329439),
	.w4(32'h3a31d3cf),
	.w5(32'hbc6bfa7f),
	.w6(32'h3ce2beb0),
	.w7(32'h3bec338b),
	.w8(32'hbc3abbdc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2769fd),
	.w1(32'hbb6b87d5),
	.w2(32'hba69ca62),
	.w3(32'hbb3f2be3),
	.w4(32'h3bd91ab1),
	.w5(32'h3bbc09f3),
	.w6(32'h3a8d5f3d),
	.w7(32'h3bcb5381),
	.w8(32'h3bdd2731),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b304145),
	.w1(32'hba3698a9),
	.w2(32'hb9d0cabb),
	.w3(32'h3bde9d12),
	.w4(32'h3b7023c8),
	.w5(32'h3bb714d6),
	.w6(32'h39a4ee81),
	.w7(32'h39779ddb),
	.w8(32'h3b3be76d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40f095),
	.w1(32'hbb989775),
	.w2(32'h3b409ccf),
	.w3(32'hbbba7d23),
	.w4(32'hbca73085),
	.w5(32'hbca42f43),
	.w6(32'hbc8faed8),
	.w7(32'hbc815cc5),
	.w8(32'hbc5a078b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9aeee),
	.w1(32'hbb4e9e8f),
	.w2(32'hbb917813),
	.w3(32'h3a43c398),
	.w4(32'h3a7196ef),
	.w5(32'h3ac70e47),
	.w6(32'h3a9abb23),
	.w7(32'hba4ad21e),
	.w8(32'h392f5f42),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc281ed6),
	.w1(32'hbbd9e480),
	.w2(32'h3aea4f70),
	.w3(32'hbc705be6),
	.w4(32'hbc6678a9),
	.w5(32'h38321c10),
	.w6(32'hbb6d867b),
	.w7(32'hbc030816),
	.w8(32'hbc28d8ad),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c1f4c),
	.w1(32'hbc7e5076),
	.w2(32'hbc036c78),
	.w3(32'hbbda8c7c),
	.w4(32'h3a52cd3f),
	.w5(32'h3bc5bcf1),
	.w6(32'h3cb26503),
	.w7(32'h3d2a7c32),
	.w8(32'h3d0298be),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0f9436),
	.w1(32'hbc380b84),
	.w2(32'hbc9beca6),
	.w3(32'hbac2aff3),
	.w4(32'h3c4bf4c6),
	.w5(32'h3c4ed216),
	.w6(32'h3bab3667),
	.w7(32'hbc8e73e6),
	.w8(32'hbd24109c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6755ed),
	.w1(32'h3b062e43),
	.w2(32'h3c4205e8),
	.w3(32'h3bde5338),
	.w4(32'h3c34c6c4),
	.w5(32'h3c898ed0),
	.w6(32'h3c55fcb4),
	.w7(32'h3c638884),
	.w8(32'h3cd5caea),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f5ca8),
	.w1(32'hbbaf95dc),
	.w2(32'h3c24e29b),
	.w3(32'h3c4158e3),
	.w4(32'h3b8813d8),
	.w5(32'h3c83fd15),
	.w6(32'h3c1e4154),
	.w7(32'h3bca08aa),
	.w8(32'h3b88c7e0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc688ff8),
	.w1(32'h3b614664),
	.w2(32'h3c8af471),
	.w3(32'hbb2daa5c),
	.w4(32'hbc09b6b7),
	.w5(32'hbb2271dc),
	.w6(32'h3befa90b),
	.w7(32'h3baaa3bd),
	.w8(32'h3c54ecea),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48f348),
	.w1(32'hbb6d4932),
	.w2(32'hbbdf9a76),
	.w3(32'h3c168e41),
	.w4(32'h3baa0d16),
	.w5(32'h3bafb53c),
	.w6(32'hbb2f6c4b),
	.w7(32'hbc4d479f),
	.w8(32'hbbf4a27f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a765e4e),
	.w1(32'h3ade2c69),
	.w2(32'hbb0f924c),
	.w3(32'hbb0ff7da),
	.w4(32'hbb7561e4),
	.w5(32'hbb23b955),
	.w6(32'h3a4441f3),
	.w7(32'hbb2c1e90),
	.w8(32'hbb22a42d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7192a7),
	.w1(32'hbd21262b),
	.w2(32'hbc73563b),
	.w3(32'h3c48d135),
	.w4(32'h3b26e338),
	.w5(32'hbbc5948d),
	.w6(32'hbc17e390),
	.w7(32'h3cb1e271),
	.w8(32'h3c6d1e6d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ccbc3),
	.w1(32'hbc3681aa),
	.w2(32'h3c23a464),
	.w3(32'h3aeffe8f),
	.w4(32'hbd02cd3c),
	.w5(32'hbcd6246e),
	.w6(32'hbd817ffe),
	.w7(32'hbdb473ae),
	.w8(32'hbd62df18),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf3ec20),
	.w1(32'h3c3f4c04),
	.w2(32'h3d09809f),
	.w3(32'hbd00f88c),
	.w4(32'hbd06cb16),
	.w5(32'hbd04810f),
	.w6(32'hbc278b48),
	.w7(32'hbaa5dffc),
	.w8(32'hbb5b514d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d17f796),
	.w1(32'hbb380931),
	.w2(32'hbc8a8320),
	.w3(32'hbc7432a6),
	.w4(32'hbcfa0ea3),
	.w5(32'hbcb9fb9a),
	.w6(32'hbba457d6),
	.w7(32'hbc2d41ea),
	.w8(32'hbc3761f6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0563b3),
	.w1(32'h3c0bbadc),
	.w2(32'h3c21a25d),
	.w3(32'hbb924266),
	.w4(32'h3b3bfb72),
	.w5(32'hb9f7aa2d),
	.w6(32'h3c84d429),
	.w7(32'h3cae1800),
	.w8(32'h3c2ab681),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfe2c4),
	.w1(32'hbb344235),
	.w2(32'hbbcdb973),
	.w3(32'hbc41f24b),
	.w4(32'hbc078354),
	.w5(32'hba9ce041),
	.w6(32'h3b7d4d6e),
	.w7(32'h3b9863ec),
	.w8(32'h3b89ec84),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe2f4c),
	.w1(32'h3b24d214),
	.w2(32'h3ba0f61d),
	.w3(32'hbb982088),
	.w4(32'h3a78ae93),
	.w5(32'hbbc85242),
	.w6(32'h3b92947e),
	.w7(32'h3bff0ca7),
	.w8(32'h3c57ddd1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac0240),
	.w1(32'h3a6350db),
	.w2(32'h3c52f72a),
	.w3(32'hbc141f29),
	.w4(32'hbc1a8172),
	.w5(32'hbbdbf764),
	.w6(32'hbbd17b94),
	.w7(32'h3bb08939),
	.w8(32'h3ada6dba),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76b7bb),
	.w1(32'hbad8d087),
	.w2(32'hba3ec08e),
	.w3(32'h3c292a71),
	.w4(32'h3bf1fff2),
	.w5(32'h3c003787),
	.w6(32'h3b82b519),
	.w7(32'h39bcfd2e),
	.w8(32'h3ba5786d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d27603),
	.w1(32'h3b1b72c7),
	.w2(32'h3c58226a),
	.w3(32'h3b60d5dc),
	.w4(32'h39a5247c),
	.w5(32'h3bce3f58),
	.w6(32'hbc437f78),
	.w7(32'hbc06df19),
	.w8(32'hbbc43c3f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e844f),
	.w1(32'h3bfd8fcd),
	.w2(32'h3cb0382a),
	.w3(32'hbd6715b5),
	.w4(32'hbd930e9d),
	.w5(32'hbceca0df),
	.w6(32'hbc027b53),
	.w7(32'hbcf48047),
	.w8(32'hbd0a5b56),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cde7bba),
	.w1(32'hbca6b6db),
	.w2(32'hbd11a23b),
	.w3(32'h3b1647ce),
	.w4(32'h3c7546ac),
	.w5(32'h3c571e37),
	.w6(32'hbcdb9f25),
	.w7(32'hbce82e80),
	.w8(32'hbd232a48),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdb18f6),
	.w1(32'hbb747266),
	.w2(32'hbb408a7c),
	.w3(32'h3b2364eb),
	.w4(32'h3ac35383),
	.w5(32'h3a1f2a83),
	.w6(32'hb88a2eb2),
	.w7(32'hba93f724),
	.w8(32'h3a0f437f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c00ef),
	.w1(32'h3a9f2726),
	.w2(32'h3b3cfc5f),
	.w3(32'hba5a0adb),
	.w4(32'h3b6d5a99),
	.w5(32'h3c287f37),
	.w6(32'h3b7a528a),
	.w7(32'h3c27f592),
	.w8(32'h3c1db65d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b7987),
	.w1(32'hbce2a8e0),
	.w2(32'hbc8742d9),
	.w3(32'h3ceb1aaf),
	.w4(32'h3babd50b),
	.w5(32'hbb22f92d),
	.w6(32'h3bcc9d07),
	.w7(32'h3cc3f975),
	.w8(32'h3cd5d495),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00ebc7),
	.w1(32'h3b0ee7ec),
	.w2(32'h3b97dbcc),
	.w3(32'hbbf69f6d),
	.w4(32'hbbf7daa8),
	.w5(32'h3b585fd6),
	.w6(32'h3af412ea),
	.w7(32'hbc0104dc),
	.w8(32'hbc1adf9d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35676c),
	.w1(32'h37fe1a2b),
	.w2(32'hbb5046c7),
	.w3(32'hbcac9550),
	.w4(32'hbccabd0f),
	.w5(32'hbca26b46),
	.w6(32'hbc553215),
	.w7(32'h3c19718e),
	.w8(32'h3c02b6f1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2acbd),
	.w1(32'hbaa955c7),
	.w2(32'hbb729697),
	.w3(32'h3bae4710),
	.w4(32'h3c719652),
	.w5(32'h3c868335),
	.w6(32'h3bcb62ef),
	.w7(32'hbb71cd47),
	.w8(32'hbc364145),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39e0fd),
	.w1(32'hbcbcde58),
	.w2(32'hbb6ad9a9),
	.w3(32'hbcaf5ec0),
	.w4(32'hbcd3a4d6),
	.w5(32'hbca2f1ee),
	.w6(32'h3c340f24),
	.w7(32'h3c31730a),
	.w8(32'h3c108682),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6838e),
	.w1(32'hba8b922d),
	.w2(32'hba108ef6),
	.w3(32'hbafbad28),
	.w4(32'hbb926527),
	.w5(32'hbb293bb8),
	.w6(32'hbab97e7e),
	.w7(32'hbb97836c),
	.w8(32'hbb9563c9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ecffb),
	.w1(32'h3b28fca1),
	.w2(32'h3c770dfe),
	.w3(32'hbd23c7c2),
	.w4(32'hbd595cb7),
	.w5(32'hbd076c66),
	.w6(32'hbcbc5ca6),
	.w7(32'hbc9ac3e3),
	.w8(32'hbc1133bd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2a6f25),
	.w1(32'h3b5fd31d),
	.w2(32'h3a9975c5),
	.w3(32'h3c0bd315),
	.w4(32'h3c3c4c67),
	.w5(32'h3bb2b3ba),
	.w6(32'h3c3d3f57),
	.w7(32'h3c1cbf49),
	.w8(32'h3bcc6d6f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05e657),
	.w1(32'hbbacaef7),
	.w2(32'hbbf760c9),
	.w3(32'h3c0c958b),
	.w4(32'h38c110ac),
	.w5(32'h3c1b0cee),
	.w6(32'h3b0198bf),
	.w7(32'hbb811837),
	.w8(32'h3c00c6d9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3af8fb),
	.w1(32'h3bb18489),
	.w2(32'h3a6a6646),
	.w3(32'h3c017e18),
	.w4(32'h3be2c18a),
	.w5(32'h3c53ec72),
	.w6(32'h3bd45550),
	.w7(32'hbc31e332),
	.w8(32'hbb92c5bb),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58b759),
	.w1(32'hbc494bb0),
	.w2(32'hbc281a21),
	.w3(32'h3b144a32),
	.w4(32'h3b966cb7),
	.w5(32'h3acaf82c),
	.w6(32'h3b962724),
	.w7(32'h3ae4fee4),
	.w8(32'hbb7444fe),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb228ef1),
	.w1(32'hbc3b201f),
	.w2(32'hbc7ac73c),
	.w3(32'hbba09916),
	.w4(32'h3ae3eaca),
	.w5(32'hbb62ff55),
	.w6(32'hb981e66d),
	.w7(32'h3b0e4990),
	.w8(32'hbb72050b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a5f66),
	.w1(32'h3c88a0ed),
	.w2(32'h3cc3a19f),
	.w3(32'h3ca99d3f),
	.w4(32'h3cb54e89),
	.w5(32'h3c4870f1),
	.w6(32'hbc56b70c),
	.w7(32'h3bcb89db),
	.w8(32'h3bb7e801),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f5cdf),
	.w1(32'hbbd3d008),
	.w2(32'hbbdd7ab1),
	.w3(32'hbb50ccd0),
	.w4(32'hbbb3853c),
	.w5(32'hbb04fa2f),
	.w6(32'h39fc67d8),
	.w7(32'h3941d635),
	.w8(32'h3a4d199b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacda6ef),
	.w1(32'h3c098193),
	.w2(32'h3bfc8d63),
	.w3(32'h3c17cae7),
	.w4(32'h3c8acb8b),
	.w5(32'h3bbb58f1),
	.w6(32'hbbed0266),
	.w7(32'hbcb70720),
	.w8(32'hbcae7d47),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32d493),
	.w1(32'hbb8b6bb7),
	.w2(32'hbb3cceed),
	.w3(32'hbb556e00),
	.w4(32'hbba0f1b0),
	.w5(32'hbb97ab40),
	.w6(32'hbb79eef1),
	.w7(32'hbb3262c6),
	.w8(32'hbb85b0ae),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d168c),
	.w1(32'hbb4b3e74),
	.w2(32'hb9da38f4),
	.w3(32'h3ae53d3a),
	.w4(32'h3b250a45),
	.w5(32'h3bf2f309),
	.w6(32'h3c90684c),
	.w7(32'hbba328c6),
	.w8(32'hbc4f942b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce6775),
	.w1(32'hbb64b896),
	.w2(32'hba859c19),
	.w3(32'h3c1ab552),
	.w4(32'h3bd394e1),
	.w5(32'h383d1afd),
	.w6(32'h3b76b1af),
	.w7(32'h3af18d05),
	.w8(32'h39b6fbe6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8282a),
	.w1(32'hbc24113b),
	.w2(32'h3bbd3680),
	.w3(32'h3bbf6b39),
	.w4(32'h3c3c08d4),
	.w5(32'h3c9e833b),
	.w6(32'h3c9160e6),
	.w7(32'h3bfec786),
	.w8(32'h3c1e4147),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc623c97),
	.w1(32'hbd1c65ec),
	.w2(32'hbce3e1b6),
	.w3(32'hbaa2619d),
	.w4(32'hbd67decf),
	.w5(32'hbd32722d),
	.w6(32'h3d000941),
	.w7(32'h3d3e3457),
	.w8(32'h3d2fb1e5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6b5d8),
	.w1(32'h3a49f8b4),
	.w2(32'hbb25d83c),
	.w3(32'h3bd73ba2),
	.w4(32'h3c14397a),
	.w5(32'h3bb69abf),
	.w6(32'hbc254b20),
	.w7(32'hbc419baa),
	.w8(32'hbc289276),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule