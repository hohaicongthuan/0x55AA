module layer_8_featuremap_25(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad59a57),
	.w1(32'hb998a8a2),
	.w2(32'hbac27b88),
	.w3(32'h3aa7a691),
	.w4(32'h3a00e704),
	.w5(32'hbabec5ab),
	.w6(32'h365cf612),
	.w7(32'h3a2f9f48),
	.w8(32'hbafec993),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3790e261),
	.w1(32'h3785b11b),
	.w2(32'hba47f546),
	.w3(32'hb8ccc26a),
	.w4(32'hb84b534b),
	.w5(32'hbaad8555),
	.w6(32'hb9a7a16b),
	.w7(32'hb82c1e19),
	.w8(32'hb9e60d19),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f7d89),
	.w1(32'hbab386a5),
	.w2(32'hba97bf5a),
	.w3(32'hb89a0f2a),
	.w4(32'h3a3bf1c8),
	.w5(32'hba7cc0e2),
	.w6(32'h38e2ff1d),
	.w7(32'h39ab8ad1),
	.w8(32'hbb83c78a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb320c4a),
	.w1(32'hbaaface2),
	.w2(32'h39be10a7),
	.w3(32'hbb23b06e),
	.w4(32'hbb26557f),
	.w5(32'hbab8ec08),
	.w6(32'hbb68541f),
	.w7(32'hbaab88e1),
	.w8(32'h399d788b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f9a8f),
	.w1(32'h3a487872),
	.w2(32'h3a1ca028),
	.w3(32'h3a91da53),
	.w4(32'h3b00ed00),
	.w5(32'h3a77d5ac),
	.w6(32'h3a548b13),
	.w7(32'h3ab1f4a7),
	.w8(32'h37a41ff3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f5247),
	.w1(32'hba4f87c5),
	.w2(32'h3b29cb32),
	.w3(32'h3a1ac9b4),
	.w4(32'hb8c07dd0),
	.w5(32'h3b19b388),
	.w6(32'hb998a653),
	.w7(32'h3ab9a78d),
	.w8(32'h39a98a45),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f9cb5),
	.w1(32'hb9c9aabd),
	.w2(32'h389dc4c5),
	.w3(32'h3ab84183),
	.w4(32'h3a05630e),
	.w5(32'hb82137c2),
	.w6(32'h37326269),
	.w7(32'h39e00a39),
	.w8(32'hb9170f71),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f6fc4),
	.w1(32'hba99a0e5),
	.w2(32'hbb3d7420),
	.w3(32'h3af7005d),
	.w4(32'h3b2d1af5),
	.w5(32'hbaa6b180),
	.w6(32'hbaacff0c),
	.w7(32'hba11ac6a),
	.w8(32'hbb7895c4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b345aa6),
	.w1(32'h3b883251),
	.w2(32'hba59967e),
	.w3(32'h3ba73f37),
	.w4(32'h3bbd6a7d),
	.w5(32'hba797575),
	.w6(32'h3af1ba13),
	.w7(32'h3b025bcd),
	.w8(32'hbbbbee83),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2abb2a),
	.w1(32'h3a197766),
	.w2(32'h38f8b2e0),
	.w3(32'hbb888e97),
	.w4(32'hbbb2c24b),
	.w5(32'hbb858b6b),
	.w6(32'hba8c88ba),
	.w7(32'hba009dcf),
	.w8(32'hba73c247),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7849b),
	.w1(32'h3a78af1c),
	.w2(32'hbb007cb7),
	.w3(32'h3b080f0e),
	.w4(32'h3b394b74),
	.w5(32'hbafd8eb3),
	.w6(32'h3ab6ab68),
	.w7(32'h3a926418),
	.w8(32'hba98bcb8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0b076),
	.w1(32'h39025d56),
	.w2(32'hba8d2b43),
	.w3(32'h3a9a3293),
	.w4(32'h3abbcbfd),
	.w5(32'hba223692),
	.w6(32'h3a0b21a1),
	.w7(32'h3a871c3c),
	.w8(32'hba39fa21),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e334b),
	.w1(32'hba97d7a8),
	.w2(32'hbb45754e),
	.w3(32'h3aa343b1),
	.w4(32'h3a6e3450),
	.w5(32'hbb38046b),
	.w6(32'hbad8e029),
	.w7(32'hbad66e26),
	.w8(32'hbb315e41),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab37b78),
	.w1(32'hba168415),
	.w2(32'h3b2166cd),
	.w3(32'h3a8f83fd),
	.w4(32'h39b80592),
	.w5(32'h3b0d8a33),
	.w6(32'hb91f1d00),
	.w7(32'h3af21e7b),
	.w8(32'hba5eee31),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2241b4),
	.w1(32'h39211efe),
	.w2(32'h3ac5b2fa),
	.w3(32'h3a5d4839),
	.w4(32'h3a2110b6),
	.w5(32'h3b0241f2),
	.w6(32'h39e741a2),
	.w7(32'h3acadf4f),
	.w8(32'h3a2bd014),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86771a),
	.w1(32'h3917dd40),
	.w2(32'h399c1ee1),
	.w3(32'h38bcdedc),
	.w4(32'hb99aadfa),
	.w5(32'hba603d5d),
	.w6(32'h384a2ac5),
	.w7(32'hb91521ec),
	.w8(32'hbab52a47),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57328f),
	.w1(32'h3a356ef7),
	.w2(32'h3b82f171),
	.w3(32'h3b15a39b),
	.w4(32'h3b6d80e7),
	.w5(32'h37e6a2aa),
	.w6(32'h3a8c11c7),
	.w7(32'h3b8e6fe7),
	.w8(32'hb9b962bb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8eeb2),
	.w1(32'hbb1792cd),
	.w2(32'hbb3276a5),
	.w3(32'hbad13d97),
	.w4(32'hbb0768de),
	.w5(32'hbb4fff0c),
	.w6(32'hbb132889),
	.w7(32'hbb05f93d),
	.w8(32'hbb49b09d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f4729),
	.w1(32'h3b5d927d),
	.w2(32'hbb9fe375),
	.w3(32'h3b74ad6a),
	.w4(32'h3b48c963),
	.w5(32'hbbaec8b7),
	.w6(32'h3aca3ee1),
	.w7(32'hbaa479d3),
	.w8(32'hbbd75fec),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6b1c7),
	.w1(32'h3af910a6),
	.w2(32'hbb86b56e),
	.w3(32'hbabb342a),
	.w4(32'hbb1a82e0),
	.w5(32'hbbdf44f0),
	.w6(32'h3a484c64),
	.w7(32'hbbb661d7),
	.w8(32'h3b49f43e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b000006),
	.w1(32'h3ad6ed2f),
	.w2(32'h3a496fa3),
	.w3(32'h3b4ab676),
	.w4(32'h3b133435),
	.w5(32'h3abd7cd6),
	.w6(32'h3b2abe37),
	.w7(32'h3ac05a44),
	.w8(32'h3aa0b5a0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cb1eb),
	.w1(32'hbaf5d3a2),
	.w2(32'h3a0cecfd),
	.w3(32'h3a84502b),
	.w4(32'hb9b138e9),
	.w5(32'h39bb4779),
	.w6(32'hbae66581),
	.w7(32'hba140f95),
	.w8(32'h3a03546d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12b22d),
	.w1(32'h3a93b1fc),
	.w2(32'hbaaef2c7),
	.w3(32'h3b02cfe0),
	.w4(32'h3b8adcb1),
	.w5(32'hba88749c),
	.w6(32'h3a155a49),
	.w7(32'h3b78da9c),
	.w8(32'hbb88287a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba425f71),
	.w1(32'hb994888a),
	.w2(32'hba4ce59f),
	.w3(32'hb9a21c26),
	.w4(32'h39ce81da),
	.w5(32'hba1459ee),
	.w6(32'hbac04517),
	.w7(32'hb8bf4c17),
	.w8(32'hbab65e78),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e2572),
	.w1(32'h3ad5d2e6),
	.w2(32'hbb9fef6e),
	.w3(32'hbb563e91),
	.w4(32'hbb1d54db),
	.w5(32'hbbd0977f),
	.w6(32'hbac96e0b),
	.w7(32'hbbcfd3cb),
	.w8(32'h3b34ae9d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accd788),
	.w1(32'h39ce65fe),
	.w2(32'hba40f299),
	.w3(32'h3a1af265),
	.w4(32'h3ab5e7ab),
	.w5(32'h3a2706a3),
	.w6(32'hbac3a6b2),
	.w7(32'h3ab0a7d7),
	.w8(32'h3a3e4268),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9d0b5),
	.w1(32'hb999eb75),
	.w2(32'h3a67b3dd),
	.w3(32'h3afba41e),
	.w4(32'h398d234a),
	.w5(32'h3a5c51dc),
	.w6(32'h3977f960),
	.w7(32'h3a341417),
	.w8(32'h3a80e20d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31a026),
	.w1(32'h3b8852b6),
	.w2(32'h3b5ad38f),
	.w3(32'h3b8f7497),
	.w4(32'h3b53486f),
	.w5(32'h3bd5c151),
	.w6(32'h3ba7db99),
	.w7(32'h3b894175),
	.w8(32'h3bade72f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab04f90),
	.w1(32'hbb899809),
	.w2(32'h3aa0ba21),
	.w3(32'hbb913c13),
	.w4(32'hbbc392ec),
	.w5(32'hbaf15a41),
	.w6(32'hba047d35),
	.w7(32'hbadade60),
	.w8(32'hba9675c2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f87ab),
	.w1(32'hba1fd4b1),
	.w2(32'hb9c79576),
	.w3(32'h39c358f1),
	.w4(32'hb83255c3),
	.w5(32'hb9db26ca),
	.w6(32'hb8b74a79),
	.w7(32'hb9082004),
	.w8(32'hbb723651),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb953edc),
	.w1(32'hbb6aeca0),
	.w2(32'hbb05dd0c),
	.w3(32'hbc13282d),
	.w4(32'hbad49ac8),
	.w5(32'h3953a442),
	.w6(32'hbbd9fdda),
	.w7(32'hbbeb84c3),
	.w8(32'h3b6778a9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2057ef),
	.w1(32'h38a48ce3),
	.w2(32'hbb39dc53),
	.w3(32'h3b253c83),
	.w4(32'h3a6d5983),
	.w5(32'hbb0c8039),
	.w6(32'h3affd4d0),
	.w7(32'h3718b528),
	.w8(32'hbb1bd8f4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60f1f2),
	.w1(32'h3904e2f0),
	.w2(32'h3b1d306d),
	.w3(32'hbb65f4f3),
	.w4(32'h3b31a6f2),
	.w5(32'h3b961b56),
	.w6(32'hba5bf9b5),
	.w7(32'hbab209d2),
	.w8(32'h3a73f3b2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13d755),
	.w1(32'h38397e54),
	.w2(32'hb9d5f976),
	.w3(32'hbbb5d962),
	.w4(32'hbb62dd8a),
	.w5(32'h3a8a9e2e),
	.w6(32'h3a13373c),
	.w7(32'hbb4ba33a),
	.w8(32'h39cd9dec),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab36cda),
	.w1(32'h3937f47a),
	.w2(32'h3b89de76),
	.w3(32'h3a9e586d),
	.w4(32'h3a9007c6),
	.w5(32'h3b836a60),
	.w6(32'h3a0d2f74),
	.w7(32'h3b373d4d),
	.w8(32'h392c0c2a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d2dd5),
	.w1(32'h3b117d93),
	.w2(32'h3a73045a),
	.w3(32'h3a363f90),
	.w4(32'h3b0273a8),
	.w5(32'h39fc4848),
	.w6(32'h39b056af),
	.w7(32'h3a918bc8),
	.w8(32'h391dd937),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0a41c),
	.w1(32'h3af2c4e9),
	.w2(32'hbb2a763d),
	.w3(32'h396240c1),
	.w4(32'h38f74141),
	.w5(32'hbb4b0961),
	.w6(32'hb9a9f917),
	.w7(32'hbb19467b),
	.w8(32'h39249b93),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba355bea),
	.w1(32'hba9f3bf1),
	.w2(32'hba976914),
	.w3(32'h39c7169f),
	.w4(32'h38cbe663),
	.w5(32'hba7c48a7),
	.w6(32'hba850bb2),
	.w7(32'hb9bbbab6),
	.w8(32'hbb164bfa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a923b29),
	.w1(32'h3a3c1de3),
	.w2(32'h3b203f76),
	.w3(32'h3aef2006),
	.w4(32'h3af0209a),
	.w5(32'h3b95ee98),
	.w6(32'h3a210aef),
	.w7(32'h3b4840bb),
	.w8(32'hb92ca477),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb846fb43),
	.w1(32'hba3161ab),
	.w2(32'hbb4bf65f),
	.w3(32'hba39f35a),
	.w4(32'hbae84092),
	.w5(32'hbb354c2c),
	.w6(32'hba181588),
	.w7(32'hbb0e6666),
	.w8(32'h3a66b746),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f863df),
	.w1(32'h3a75c4e4),
	.w2(32'h3aa170be),
	.w3(32'h3a0c7b89),
	.w4(32'h3a9b1e17),
	.w5(32'h3a96b701),
	.w6(32'hb96c3307),
	.w7(32'h39a5d145),
	.w8(32'h3a7341f3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5ed97),
	.w1(32'h3adf4479),
	.w2(32'h3a842f18),
	.w3(32'h3a127375),
	.w4(32'h3a7c6c1f),
	.w5(32'h3a0771cf),
	.w6(32'h3acbfa61),
	.w7(32'h3ab0e603),
	.w8(32'h3aa09e91),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af887e1),
	.w1(32'hbafbe4fd),
	.w2(32'hbad7cedf),
	.w3(32'h3b1362a1),
	.w4(32'hba1718fe),
	.w5(32'hba0e4684),
	.w6(32'hbaa3e060),
	.w7(32'hba641514),
	.w8(32'h3a255791),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0631f4),
	.w1(32'h3b11f90c),
	.w2(32'h3a45728b),
	.w3(32'h3a762d24),
	.w4(32'h3aecb129),
	.w5(32'h3a0ea201),
	.w6(32'h3aea7c0a),
	.w7(32'h3ab252a5),
	.w8(32'h3a925426),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c338c),
	.w1(32'h3b125255),
	.w2(32'hba88d626),
	.w3(32'h3b1c728c),
	.w4(32'h3b50779d),
	.w5(32'h350de5d5),
	.w6(32'h3b19a0d0),
	.w7(32'h3b62be7a),
	.w8(32'hb9ebea13),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6876e),
	.w1(32'h3aba8c32),
	.w2(32'h3aaf94e3),
	.w3(32'h3ad6367e),
	.w4(32'h3a222484),
	.w5(32'h390b9f21),
	.w6(32'h3ab75c4a),
	.w7(32'h3b005a82),
	.w8(32'h39aebda1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902397e),
	.w1(32'h3abee3fa),
	.w2(32'h39907487),
	.w3(32'hb895ed27),
	.w4(32'hba617ce5),
	.w5(32'hbadee9e3),
	.w6(32'h3a86eb90),
	.w7(32'h3ae1352f),
	.w8(32'h3afb4d72),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c0e45),
	.w1(32'h3b8bb523),
	.w2(32'hba2e36f4),
	.w3(32'h3b406c18),
	.w4(32'h3b9ae6ee),
	.w5(32'hb9ba16f6),
	.w6(32'h3b39f7b0),
	.w7(32'h3b298361),
	.w8(32'hbbac99fb),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb098ec3),
	.w1(32'hbaf762e3),
	.w2(32'hbb2d1d63),
	.w3(32'hbb0a25aa),
	.w4(32'hbb13d497),
	.w5(32'hbb2e172a),
	.w6(32'hbb28d090),
	.w7(32'hbb1c7e37),
	.w8(32'hb8c899fd),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad03517),
	.w1(32'h3a823acb),
	.w2(32'hba828a45),
	.w3(32'h3a4e8c4b),
	.w4(32'h3965f2dc),
	.w5(32'hba986334),
	.w6(32'h3aad641f),
	.w7(32'h3a8a508b),
	.w8(32'hba26d015),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13d00d),
	.w1(32'h389a4ef9),
	.w2(32'h3b0db5ab),
	.w3(32'h3aa97cb5),
	.w4(32'h39c51ef5),
	.w5(32'h3ac94e58),
	.w6(32'h3a423550),
	.w7(32'hba1d2826),
	.w8(32'h3ae43847),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9752e9),
	.w1(32'h3b645e3a),
	.w2(32'hb8fdc474),
	.w3(32'h3ba9bc57),
	.w4(32'h3b97c4e9),
	.w5(32'hb94588d1),
	.w6(32'h3b7d8292),
	.w7(32'h3b4ca2d6),
	.w8(32'hbaf9cc27),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b480e2e),
	.w1(32'h3a78d8e0),
	.w2(32'hb8d6a639),
	.w3(32'h3b0b38c0),
	.w4(32'h3ac85a36),
	.w5(32'hba2ecfe0),
	.w6(32'h3a62a78f),
	.w7(32'h3b74e1cd),
	.w8(32'hbb9b5107),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab29742),
	.w1(32'h39d85de5),
	.w2(32'hba5dfd4f),
	.w3(32'hbad5b629),
	.w4(32'hba1ac23d),
	.w5(32'hbab3c712),
	.w6(32'hba4227ae),
	.w7(32'hb9dc6767),
	.w8(32'hba9ee159),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2829b3),
	.w1(32'hb8ad0208),
	.w2(32'hbadbc2a3),
	.w3(32'hba5f3e67),
	.w4(32'h3a558212),
	.w5(32'hbaa168ae),
	.w6(32'h3a525593),
	.w7(32'hba83cb3f),
	.w8(32'hba206e52),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efddff),
	.w1(32'h3b78d47b),
	.w2(32'hb9b2b8bf),
	.w3(32'h3b2b2c09),
	.w4(32'h3bae1a03),
	.w5(32'h3a64e407),
	.w6(32'h3b366431),
	.w7(32'h3b6d7013),
	.w8(32'hbb074296),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d3b53),
	.w1(32'hb77d96dd),
	.w2(32'hb996f409),
	.w3(32'hb9828641),
	.w4(32'h39c717de),
	.w5(32'hba85b659),
	.w6(32'h39104f8f),
	.w7(32'h3a7464f1),
	.w8(32'h3a7e525a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6c989),
	.w1(32'h3abaeb4c),
	.w2(32'h399d6010),
	.w3(32'h3ab83753),
	.w4(32'h3af505f0),
	.w5(32'h39f13daf),
	.w6(32'hb985cbf1),
	.w7(32'hbad07725),
	.w8(32'h3aec35e2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d5d6b),
	.w1(32'h3a10699d),
	.w2(32'h3744e097),
	.w3(32'h3a8642ad),
	.w4(32'h3a27c571),
	.w5(32'hb9466e9d),
	.w6(32'h3a6e79c1),
	.w7(32'h3a78d407),
	.w8(32'hba31dfb3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba854ba7),
	.w1(32'hbb23c27a),
	.w2(32'hb9ec2f7f),
	.w3(32'hb9bb6750),
	.w4(32'hbaaf71a4),
	.w5(32'h3968c17a),
	.w6(32'hbabeea86),
	.w7(32'h3a1fbb75),
	.w8(32'h3b3734cb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc2bb7),
	.w1(32'h3a4aead3),
	.w2(32'h3a1197c3),
	.w3(32'h3abcc8ce),
	.w4(32'h3a2544ac),
	.w5(32'hbb64334c),
	.w6(32'h3b344ade),
	.w7(32'h3b5c85d1),
	.w8(32'hb98ded57),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14e1e4),
	.w1(32'h3a9ad583),
	.w2(32'h3b047c75),
	.w3(32'h3aee8574),
	.w4(32'h3ad998ae),
	.w5(32'h3ac1583b),
	.w6(32'h3a14cd7a),
	.w7(32'h3accf8f2),
	.w8(32'h3b43e079),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b678b),
	.w1(32'h3b120499),
	.w2(32'h3accd985),
	.w3(32'h3b66649b),
	.w4(32'h3b4290bb),
	.w5(32'h3ae884d9),
	.w6(32'h3b143e54),
	.w7(32'h3b8ae9d5),
	.w8(32'h3a172e9f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4967e),
	.w1(32'h393dcb84),
	.w2(32'hbae0d99b),
	.w3(32'h3b376e02),
	.w4(32'h3b3de40c),
	.w5(32'h3aa30535),
	.w6(32'h3a360b2b),
	.w7(32'h38ac800b),
	.w8(32'hba87e558),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37e78f),
	.w1(32'h3a8d54fb),
	.w2(32'hb8ca60ac),
	.w3(32'hb96544d9),
	.w4(32'h3a8ba38b),
	.w5(32'hb9acc6c3),
	.w6(32'h3a7c9fac),
	.w7(32'h393bdab3),
	.w8(32'hb9529eb8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3ebae),
	.w1(32'h3af56208),
	.w2(32'h3a819585),
	.w3(32'h3ac1c387),
	.w4(32'h3b285fde),
	.w5(32'h3a86a529),
	.w6(32'h3b040fe6),
	.w7(32'h3b308e75),
	.w8(32'h3a00575f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83621d),
	.w1(32'hb9993a76),
	.w2(32'hb88113b2),
	.w3(32'hb9cc9b8b),
	.w4(32'h3a9cdb5a),
	.w5(32'h3a5959e7),
	.w6(32'h3a093a25),
	.w7(32'h3ae9a071),
	.w8(32'hb9e6fe96),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b279e89),
	.w1(32'h3afa5ae2),
	.w2(32'h3b4ad148),
	.w3(32'h3ac129d5),
	.w4(32'h3abf768e),
	.w5(32'h3a95d93c),
	.w6(32'h391dfed4),
	.w7(32'h3a9f2fb2),
	.w8(32'h3a5c80c9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4aa59),
	.w1(32'h3a846d7e),
	.w2(32'h3a63d799),
	.w3(32'h3a8035a0),
	.w4(32'h3a57c745),
	.w5(32'h3a60ad87),
	.w6(32'h3ab10b09),
	.w7(32'h3a946cb2),
	.w8(32'h3ba2ca00),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd65557),
	.w1(32'h3bc74637),
	.w2(32'h3b722b24),
	.w3(32'h3ba20916),
	.w4(32'h3be0fc0f),
	.w5(32'h3bb19377),
	.w6(32'h3bafdb06),
	.w7(32'h3be3a49e),
	.w8(32'h3b0ff317),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5115dd),
	.w1(32'h3aa29394),
	.w2(32'h3a8e967c),
	.w3(32'h38d6c855),
	.w4(32'h3a4aa474),
	.w5(32'h3a67332a),
	.w6(32'h3a91b5f4),
	.w7(32'h3a3b5907),
	.w8(32'h39dfeaa0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb00e7),
	.w1(32'h3b0b7d53),
	.w2(32'hb9a7871c),
	.w3(32'h3a2a0f7f),
	.w4(32'h3b04b23c),
	.w5(32'hb9c59ffe),
	.w6(32'h3a7d8ce2),
	.w7(32'h3af36938),
	.w8(32'h3a32ffbe),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeefea3),
	.w1(32'h3aef0552),
	.w2(32'h3a9d80bb),
	.w3(32'h3a91dc04),
	.w4(32'h3a8d7ad6),
	.w5(32'h3a860978),
	.w6(32'h3b0f298e),
	.w7(32'h3aa79b70),
	.w8(32'h3a5cd2c9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb259df6),
	.w1(32'h39985c49),
	.w2(32'hbac304d3),
	.w3(32'hbaa6d7a2),
	.w4(32'hba5deda7),
	.w5(32'h38961498),
	.w6(32'hb89b33d4),
	.w7(32'hba9bc054),
	.w8(32'h3a0d65e6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84bb68),
	.w1(32'h3a48d97d),
	.w2(32'h3a90c3fb),
	.w3(32'h39fd8c41),
	.w4(32'h39941569),
	.w5(32'h3a29b134),
	.w6(32'h3a87606f),
	.w7(32'h3a94a907),
	.w8(32'h3a52c7ee),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2064e),
	.w1(32'h3a7289cb),
	.w2(32'h3a22923a),
	.w3(32'h3a907e56),
	.w4(32'h3a961f34),
	.w5(32'h3a94c73d),
	.w6(32'h3a9d9e21),
	.w7(32'h3aedebc0),
	.w8(32'h3ab857f3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a909716),
	.w1(32'h3a58c10b),
	.w2(32'h3a6367cb),
	.w3(32'h3a0e0fc1),
	.w4(32'h39f392fc),
	.w5(32'h3a24e35a),
	.w6(32'h3a90fc72),
	.w7(32'h3a5d2ba7),
	.w8(32'h3bb64b18),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2437e),
	.w1(32'h3b8d7103),
	.w2(32'h3ae53123),
	.w3(32'h3b98c82b),
	.w4(32'h3b982506),
	.w5(32'h3ad30aa5),
	.w6(32'h3b9cb7bc),
	.w7(32'h3bbfbe57),
	.w8(32'h3acab891),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48e243),
	.w1(32'h3b2631f1),
	.w2(32'h3b5a72b3),
	.w3(32'h3b276e16),
	.w4(32'h3b3ed173),
	.w5(32'h3b3ad8bc),
	.w6(32'h3b581a13),
	.w7(32'h3b73a080),
	.w8(32'h3a0a41ff),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0d073),
	.w1(32'h3a07bb7a),
	.w2(32'hb742b909),
	.w3(32'h38b58cbd),
	.w4(32'h398e3de9),
	.w5(32'hb8b99fe1),
	.w6(32'h39b41611),
	.w7(32'hb9cb9e7e),
	.w8(32'h3aab3485),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f9d37),
	.w1(32'hb95ea5c8),
	.w2(32'h3a5f5ec2),
	.w3(32'h3a8d6720),
	.w4(32'h3a5b9b57),
	.w5(32'h3a9bc280),
	.w6(32'h3b2736bc),
	.w7(32'h3acaaaee),
	.w8(32'h3a6fd730),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1cf8b),
	.w1(32'h3accc349),
	.w2(32'h3afbbcfc),
	.w3(32'h3aae7958),
	.w4(32'h3b0a00a6),
	.w5(32'h3ab43cda),
	.w6(32'h3ad32043),
	.w7(32'h3b10d1ba),
	.w8(32'h39a5b2b3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13921c),
	.w1(32'h3b1289d4),
	.w2(32'hbab2b082),
	.w3(32'h3aa980ed),
	.w4(32'h3b3bde09),
	.w5(32'hba973d5c),
	.w6(32'h3a4c87c9),
	.w7(32'h3ad79b07),
	.w8(32'hbb2ca4b7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4aece8),
	.w1(32'h39fb67bd),
	.w2(32'h39cb38fa),
	.w3(32'h3a440450),
	.w4(32'h38912cf7),
	.w5(32'h38ca60dc),
	.w6(32'hbacf13da),
	.w7(32'hb9105a24),
	.w8(32'h3a51b251),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d1caf),
	.w1(32'h3b911fb4),
	.w2(32'hbae8bf16),
	.w3(32'h3b632788),
	.w4(32'h3bdc11db),
	.w5(32'hba2ecd97),
	.w6(32'h3b34493d),
	.w7(32'h3bafbf2c),
	.w8(32'hba3da0a2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1e54e),
	.w1(32'h3b70b6bc),
	.w2(32'h3a4bc3d2),
	.w3(32'h3b81e4ff),
	.w4(32'h3b7c9bfd),
	.w5(32'h3adc3281),
	.w6(32'h3b5b080f),
	.w7(32'h3b767715),
	.w8(32'hbb856447),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb482ce0),
	.w1(32'hbb1f4154),
	.w2(32'hbb1f63e9),
	.w3(32'hbb1ca796),
	.w4(32'hbb28825f),
	.w5(32'hbb147d6d),
	.w6(32'hbb31662a),
	.w7(32'hbb3574da),
	.w8(32'h3a4a76ef),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13092a),
	.w1(32'h3960be44),
	.w2(32'hb708171d),
	.w3(32'h3a083e9c),
	.w4(32'h3a43da9a),
	.w5(32'h38faf145),
	.w6(32'h3a886a36),
	.w7(32'h39a4ae59),
	.w8(32'h38a81b84),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96fbe04),
	.w1(32'hbaff8280),
	.w2(32'hba85614e),
	.w3(32'hb9b2b1ba),
	.w4(32'hbab1472f),
	.w5(32'hba30160e),
	.w6(32'hbabc674e),
	.w7(32'hba52a675),
	.w8(32'hbb1e84d0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb633797),
	.w1(32'hbadb3877),
	.w2(32'hbb53eb85),
	.w3(32'hbb2ef127),
	.w4(32'hbadacbe2),
	.w5(32'hbb485d70),
	.w6(32'hbb3357c2),
	.w7(32'hbb01dfd0),
	.w8(32'hbb40b9aa),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d9466),
	.w1(32'hbae0ebc6),
	.w2(32'hbaec11b7),
	.w3(32'hbb01860e),
	.w4(32'hbae987e2),
	.w5(32'hbb059fa6),
	.w6(32'hbb060585),
	.w7(32'hbafd5777),
	.w8(32'h39955c21),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d82d8),
	.w1(32'h3b13845f),
	.w2(32'h3ac8d99f),
	.w3(32'h39f83517),
	.w4(32'h3aa5a04e),
	.w5(32'h3a937440),
	.w6(32'h3ab52dc9),
	.w7(32'h3ac7284d),
	.w8(32'hba024e76),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca0e1f),
	.w1(32'h3a82103c),
	.w2(32'hbae1132f),
	.w3(32'h3941fa41),
	.w4(32'h3b4dae1e),
	.w5(32'h3a04e286),
	.w6(32'h3ae2d58c),
	.w7(32'hba298119),
	.w8(32'hb9315249),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabf38c),
	.w1(32'h3a1f3d67),
	.w2(32'hbad07f7c),
	.w3(32'h3a6ba2a4),
	.w4(32'h3a3cd4d3),
	.w5(32'hbab1e0ee),
	.w6(32'h3a9ba5d4),
	.w7(32'h3a98ca81),
	.w8(32'hbaef5f47),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2077c8),
	.w1(32'hba971dd8),
	.w2(32'h3991fe99),
	.w3(32'hba0b1a6c),
	.w4(32'hbacfcd77),
	.w5(32'hbabd4e58),
	.w6(32'hba82ef15),
	.w7(32'h39938126),
	.w8(32'h3acdf547),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af71daa),
	.w1(32'h3ae69eba),
	.w2(32'h3a5c10a0),
	.w3(32'h3b89451e),
	.w4(32'h3b747a5f),
	.w5(32'h3b073072),
	.w6(32'h3b29420f),
	.w7(32'h3b607cff),
	.w8(32'hbafd8b8b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81f10c),
	.w1(32'h3b3b3b29),
	.w2(32'hba4e619d),
	.w3(32'hb8829002),
	.w4(32'h3b5889e9),
	.w5(32'hbb1d433c),
	.w6(32'h3a94dfcc),
	.w7(32'h3b53e55a),
	.w8(32'hbb1b8a43),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba862eab),
	.w1(32'hb9c8f327),
	.w2(32'hb8a5f07f),
	.w3(32'h3a19e670),
	.w4(32'h3aa752a9),
	.w5(32'h3a7d5567),
	.w6(32'h3a52c0c0),
	.w7(32'h3b002ea5),
	.w8(32'h3b9f7a63),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b651571),
	.w1(32'h3b0f9fb3),
	.w2(32'h3b25651c),
	.w3(32'h3b51bd0c),
	.w4(32'h3b22cbc1),
	.w5(32'h3b1d8ee0),
	.w6(32'h3b7bf0c5),
	.w7(32'h3b8103a2),
	.w8(32'h3a0c96b2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a277496),
	.w1(32'h3a458216),
	.w2(32'hb68970a1),
	.w3(32'h399d8cb2),
	.w4(32'h3a520637),
	.w5(32'h3624fadb),
	.w6(32'h3abc85f6),
	.w7(32'h3a0e2cdd),
	.w8(32'h39ae7131),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac5cc8),
	.w1(32'h3a3efb90),
	.w2(32'h3a74ab11),
	.w3(32'h38d9c069),
	.w4(32'h39171223),
	.w5(32'h393028af),
	.w6(32'h39971e09),
	.w7(32'h3a29e2bd),
	.w8(32'h3a7b73d8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44fec3),
	.w1(32'h3a8685f0),
	.w2(32'h3a0f54f9),
	.w3(32'h3ac05912),
	.w4(32'h3acfd04f),
	.w5(32'h3a2cc299),
	.w6(32'h3ac8bf8b),
	.w7(32'h3ad3cc40),
	.w8(32'h3ba08f46),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb5771),
	.w1(32'h3b7400ac),
	.w2(32'h3b7202f5),
	.w3(32'h3b922335),
	.w4(32'h3b56d602),
	.w5(32'h3b2c1749),
	.w6(32'h3baaf7ed),
	.w7(32'h3baa3f47),
	.w8(32'hb9e3e2f5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af64cb3),
	.w1(32'h3b74e98d),
	.w2(32'h39203118),
	.w3(32'h3a5953b6),
	.w4(32'h3b3d5ab8),
	.w5(32'h399310a2),
	.w6(32'h3b23e35d),
	.w7(32'h3b2f8db1),
	.w8(32'hba9f4298),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf2265),
	.w1(32'hba8065db),
	.w2(32'hba514385),
	.w3(32'hba898743),
	.w4(32'hba99fccf),
	.w5(32'hba42328b),
	.w6(32'hba9f1182),
	.w7(32'hbaa08358),
	.w8(32'h3a41b010),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9c179),
	.w1(32'hb9e6f422),
	.w2(32'hbb67e131),
	.w3(32'h3a3cc05a),
	.w4(32'hb89de071),
	.w5(32'hbb682db8),
	.w6(32'h3ad75ab7),
	.w7(32'h3aac16ef),
	.w8(32'hbba7446e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77a947),
	.w1(32'hbad0e578),
	.w2(32'h3b8b9317),
	.w3(32'h3b182def),
	.w4(32'h3c13bcb7),
	.w5(32'h3bd6571e),
	.w6(32'hbbceb628),
	.w7(32'h3b9fb863),
	.w8(32'hbb05556c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0498b7),
	.w1(32'hba99406c),
	.w2(32'hbb0a3a52),
	.w3(32'hba4ef393),
	.w4(32'hbafb4a31),
	.w5(32'hbb2c9fe4),
	.w6(32'h3805313d),
	.w7(32'hba29f5fc),
	.w8(32'hba0207a1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb854676a),
	.w1(32'hb9ec6cad),
	.w2(32'h3abf1065),
	.w3(32'hba31a524),
	.w4(32'hba817b6d),
	.w5(32'h3a8fcea9),
	.w6(32'h38e03119),
	.w7(32'h37d00294),
	.w8(32'h3b7653e8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9473eb6),
	.w1(32'hba8359d3),
	.w2(32'hbafe0b78),
	.w3(32'h39b29716),
	.w4(32'h3b2f5f29),
	.w5(32'hbaec2f8d),
	.w6(32'h3b55c4de),
	.w7(32'h3b0057b5),
	.w8(32'hbbad9a0a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15ba19),
	.w1(32'hbb200bbd),
	.w2(32'hbb5cbc31),
	.w3(32'hbbdeb40a),
	.w4(32'hbbb128ba),
	.w5(32'hba7687b1),
	.w6(32'hbb8a5cda),
	.w7(32'hbbb6ec69),
	.w8(32'hba820e7b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef1657),
	.w1(32'hbad8f812),
	.w2(32'h3b49bc8b),
	.w3(32'hbaabaf74),
	.w4(32'hbae3a866),
	.w5(32'hbb04fe76),
	.w6(32'hbb2c5bb6),
	.w7(32'hba95e4da),
	.w8(32'h3b53677d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a777357),
	.w1(32'hb97f2c99),
	.w2(32'h39ed5225),
	.w3(32'h3a7e6084),
	.w4(32'h3a4d515e),
	.w5(32'h3b227f36),
	.w6(32'h3ad4df9c),
	.w7(32'h3b1299ae),
	.w8(32'h3b03e22d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3af5b5),
	.w1(32'hb9f62492),
	.w2(32'h39439efc),
	.w3(32'h398da916),
	.w4(32'hb9208533),
	.w5(32'hb95b726d),
	.w6(32'h39ae7fbe),
	.w7(32'hb8ea87d7),
	.w8(32'h392bedb2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b1458),
	.w1(32'hb9ca436f),
	.w2(32'hb9965c42),
	.w3(32'hb979633c),
	.w4(32'hba47f103),
	.w5(32'hba8304ff),
	.w6(32'hb3674684),
	.w7(32'h39105d41),
	.w8(32'h38966936),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb927e180),
	.w1(32'hbb0bec2d),
	.w2(32'hbaf3c9e0),
	.w3(32'hba95d62d),
	.w4(32'hbb34866f),
	.w5(32'hbb40df68),
	.w6(32'h39d6b284),
	.w7(32'hb9f6c9cd),
	.w8(32'hbb831725),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75dc01),
	.w1(32'hba268c2d),
	.w2(32'h3aa575c7),
	.w3(32'h3b2be49b),
	.w4(32'h3bf8aa87),
	.w5(32'h3bd84d67),
	.w6(32'hbbd8f1d7),
	.w7(32'hbb6ebe9b),
	.w8(32'h3b58f1ba),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f90e2),
	.w1(32'h392af823),
	.w2(32'hbb19b14d),
	.w3(32'h3a69d4af),
	.w4(32'hb9cafd68),
	.w5(32'hbb0d9c59),
	.w6(32'h3af14eb1),
	.w7(32'hb70181ff),
	.w8(32'hbba50938),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16832d),
	.w1(32'hba9e4f24),
	.w2(32'hbb2f723f),
	.w3(32'hb84931e9),
	.w4(32'h3b127e4a),
	.w5(32'hbb5b0ada),
	.w6(32'hbc0d992c),
	.w7(32'hbb6da8b1),
	.w8(32'h3bb40ac1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75a469),
	.w1(32'hbb9e3c14),
	.w2(32'hbbab1b60),
	.w3(32'hb8587254),
	.w4(32'hbae9851b),
	.w5(32'hba1fbea7),
	.w6(32'h3abe6801),
	.w7(32'hba41018b),
	.w8(32'hbad6d42c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04e17d),
	.w1(32'hb9d68cc2),
	.w2(32'hbb33fb8f),
	.w3(32'hb9f6839c),
	.w4(32'hbb6c49b8),
	.w5(32'hba05bdcc),
	.w6(32'h3b06b110),
	.w7(32'hbb015e38),
	.w8(32'hbb4d5420),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9821d8),
	.w1(32'hbae1b448),
	.w2(32'h3b0a28cf),
	.w3(32'hb88cc146),
	.w4(32'h3aca1df6),
	.w5(32'h3b1703fe),
	.w6(32'hbb77be88),
	.w7(32'h3bc02804),
	.w8(32'h3a77774b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a393af0),
	.w1(32'h39e7f6d0),
	.w2(32'h3af1046b),
	.w3(32'h3ad44329),
	.w4(32'h3a8b1793),
	.w5(32'h3b2528cd),
	.w6(32'h3aa6c841),
	.w7(32'h3b27bf7f),
	.w8(32'hb94c0401),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c95a2),
	.w1(32'h3b1d86f0),
	.w2(32'h3ac153c6),
	.w3(32'hbb27d494),
	.w4(32'hb98a588e),
	.w5(32'h3b3c0945),
	.w6(32'hbadadb42),
	.w7(32'hb9d66fb4),
	.w8(32'h3bed37f7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba87d15),
	.w1(32'h39430b30),
	.w2(32'hbaa8de4f),
	.w3(32'hbb20623d),
	.w4(32'hbb279df3),
	.w5(32'h3c17404f),
	.w6(32'h3b1d19a5),
	.w7(32'hbb12610a),
	.w8(32'h38a1fbca),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5228f2),
	.w1(32'hb76ebb0f),
	.w2(32'h3a08a592),
	.w3(32'h3a45d62c),
	.w4(32'hbafe051d),
	.w5(32'hbb2faf89),
	.w6(32'h39d6f7f0),
	.w7(32'hba98ca23),
	.w8(32'h3a627109),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fbd72),
	.w1(32'h3a11c1cf),
	.w2(32'h396f1613),
	.w3(32'h3ad0d50c),
	.w4(32'hb988afb3),
	.w5(32'hb9a7f673),
	.w6(32'h3b65ae64),
	.w7(32'h3adfb158),
	.w8(32'hbb7877f0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcf2a7),
	.w1(32'hbbc813d2),
	.w2(32'h3b0d4f08),
	.w3(32'hbb18f328),
	.w4(32'h3a8767f6),
	.w5(32'h3aaf996c),
	.w6(32'hbbc08066),
	.w7(32'h3a2ce5fa),
	.w8(32'hb6d8e960),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule