module layer_10_featuremap_299(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f3bad),
	.w1(32'h3c05f8fa),
	.w2(32'h3c0d37df),
	.w3(32'h3baf919a),
	.w4(32'h3bc0e006),
	.w5(32'h3a95b53b),
	.w6(32'hba0a665a),
	.w7(32'h3bad4163),
	.w8(32'h3a814902),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72c8c1),
	.w1(32'h3b7981de),
	.w2(32'hbb09a9c1),
	.w3(32'hb84c2294),
	.w4(32'h3b44434d),
	.w5(32'hbb0e78ec),
	.w6(32'h3b1e202d),
	.w7(32'hbafc8666),
	.w8(32'h3b606137),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c751e),
	.w1(32'h3b6f85f1),
	.w2(32'h3c2d91fc),
	.w3(32'hb894cc76),
	.w4(32'hbbc404cf),
	.w5(32'h39b731c8),
	.w6(32'hbab1ff23),
	.w7(32'h3b1bc0f6),
	.w8(32'hbad58e90),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b8cb2),
	.w1(32'h3acc42dd),
	.w2(32'h3a6d1a57),
	.w3(32'hbbaa7ab0),
	.w4(32'hbb049a85),
	.w5(32'h3c0cbca5),
	.w6(32'hbb5f0bef),
	.w7(32'hbb013b92),
	.w8(32'h3c0bca77),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82cb77),
	.w1(32'hbc0abbe4),
	.w2(32'h3b8e3fb4),
	.w3(32'hbc3c88d6),
	.w4(32'h3b362a84),
	.w5(32'hba08d443),
	.w6(32'hbc211cd0),
	.w7(32'hba97e4ee),
	.w8(32'h3b3a4a95),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0694c7),
	.w1(32'h3a56c30d),
	.w2(32'h3b6359e7),
	.w3(32'hbb2d5714),
	.w4(32'h3a8f63ae),
	.w5(32'h3ad037ee),
	.w6(32'hba7a506e),
	.w7(32'h3b82471c),
	.w8(32'hb9c1aefa),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb682bd),
	.w1(32'hbaf69662),
	.w2(32'hbb5c5370),
	.w3(32'hbb851dcb),
	.w4(32'hbb102b6b),
	.w5(32'hbaf3fd75),
	.w6(32'hbbe2b587),
	.w7(32'hbbe0cbee),
	.w8(32'hbc0cfd86),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb96577),
	.w1(32'hbc07c3e7),
	.w2(32'hbbf8bcb2),
	.w3(32'hbbc0d12b),
	.w4(32'hbb900f96),
	.w5(32'hbb6a4088),
	.w6(32'hbc885c02),
	.w7(32'hbbfa9801),
	.w8(32'h3a291d69),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b109fad),
	.w1(32'h3a85af0f),
	.w2(32'h3a9c2fc6),
	.w3(32'h399e1296),
	.w4(32'h3a65f2e0),
	.w5(32'hbb01e0b6),
	.w6(32'hb91e77b2),
	.w7(32'h3a718b6f),
	.w8(32'hbb1b9f69),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb714f7b4),
	.w1(32'hbac85aac),
	.w2(32'h3b4d77c4),
	.w3(32'hbba2d6bb),
	.w4(32'h3b36bf93),
	.w5(32'hbb57bf6f),
	.w6(32'hbb81b9a6),
	.w7(32'h3bc3263c),
	.w8(32'hbb2d9a3e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10560c),
	.w1(32'hbbdfbb62),
	.w2(32'h3ba6c683),
	.w3(32'hbc7e4490),
	.w4(32'hbbc63d2e),
	.w5(32'h39f9c2b0),
	.w6(32'hbc5b2451),
	.w7(32'hbb8cb417),
	.w8(32'h3bdd9723),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7d74a),
	.w1(32'hbabfb196),
	.w2(32'h388ccbb9),
	.w3(32'h3b59232b),
	.w4(32'hbb35ed1f),
	.w5(32'h3a1b12ad),
	.w6(32'h3bd0dbe3),
	.w7(32'h3ae508c7),
	.w8(32'hbbae2821),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e557a0),
	.w1(32'hbabf86d1),
	.w2(32'h3aaff91a),
	.w3(32'h3aab32d1),
	.w4(32'h3c026efa),
	.w5(32'hb88f5954),
	.w6(32'h3a87d8b1),
	.w7(32'h3b3d1956),
	.w8(32'hb897e1f1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ed509),
	.w1(32'h3b96fff8),
	.w2(32'hb9212b88),
	.w3(32'h3aba16e4),
	.w4(32'h3a084c09),
	.w5(32'hb9d3b3db),
	.w6(32'h3aa578ad),
	.w7(32'h3b0a76d5),
	.w8(32'hbb1889e1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd98163),
	.w1(32'h39c8bec1),
	.w2(32'h3b02e5c0),
	.w3(32'hbb14c7e0),
	.w4(32'h3ae3c3fa),
	.w5(32'h3b3ffbde),
	.w6(32'hbae64bc0),
	.w7(32'hba30bfff),
	.w8(32'h3ae1bcfc),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada89be),
	.w1(32'h3b301807),
	.w2(32'h3b08325d),
	.w3(32'h3b0e2bf9),
	.w4(32'h3b6c7551),
	.w5(32'hbae4b887),
	.w6(32'hba87d51e),
	.w7(32'hba8f7a7f),
	.w8(32'hbb12b404),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86256d),
	.w1(32'h3a808301),
	.w2(32'hbb52ef63),
	.w3(32'h3a1e40d1),
	.w4(32'hbb7b6d4b),
	.w5(32'hba04509b),
	.w6(32'h3af3ea73),
	.w7(32'hbb3496af),
	.w8(32'h3b7be4ec),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec23ba),
	.w1(32'hbba7ff32),
	.w2(32'hbca8f71f),
	.w3(32'hba0f783e),
	.w4(32'hbc8441fd),
	.w5(32'hbc5a41a8),
	.w6(32'hba8391d5),
	.w7(32'hbc37991e),
	.w8(32'hbbdb3d77),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7b1cf),
	.w1(32'hbb9f7770),
	.w2(32'hbc2b5823),
	.w3(32'hbb53b113),
	.w4(32'hbc0f099f),
	.w5(32'hbb5e5a8c),
	.w6(32'h3b9564e3),
	.w7(32'h3a5b20a0),
	.w8(32'hbb66816b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4d660),
	.w1(32'hbb8fb168),
	.w2(32'hbb2d01d7),
	.w3(32'h3735c254),
	.w4(32'hbb1f1bb6),
	.w5(32'h38d0a536),
	.w6(32'hb90e586c),
	.w7(32'hba871bf5),
	.w8(32'h396a6a3e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab15978),
	.w1(32'hbb71b0e9),
	.w2(32'hbb516d4b),
	.w3(32'hbb0678b5),
	.w4(32'hb9e6835b),
	.w5(32'hbaf0f995),
	.w6(32'hbb40cc0b),
	.w7(32'hbae5c5b5),
	.w8(32'hba53e890),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb2933),
	.w1(32'h3bbb33eb),
	.w2(32'h3bb89bff),
	.w3(32'h39b6e254),
	.w4(32'h3a4a8b62),
	.w5(32'h3ac7ac59),
	.w6(32'h3b1a28bc),
	.w7(32'h3a691d86),
	.w8(32'h3a1c66ab),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39399955),
	.w1(32'hbc0398a1),
	.w2(32'hbc856d21),
	.w3(32'hbb3a6090),
	.w4(32'hbc1e7e8b),
	.w5(32'hbc22239a),
	.w6(32'hbc8cecd5),
	.w7(32'hbc5db297),
	.w8(32'hbc75297e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1b4d1),
	.w1(32'hbad2520b),
	.w2(32'hb96f50c9),
	.w3(32'h3bb0e61b),
	.w4(32'h3c14655c),
	.w5(32'h3af8ceb1),
	.w6(32'h3a896e0e),
	.w7(32'h3b538bad),
	.w8(32'h3b3f4d84),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c041dc7),
	.w1(32'h3c1902ce),
	.w2(32'h3b0e3bd8),
	.w3(32'h3b8cf66d),
	.w4(32'h3ad1158e),
	.w5(32'h3b8d8396),
	.w6(32'h3bfbed77),
	.w7(32'hb9f422aa),
	.w8(32'hbba0df83),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57e371),
	.w1(32'hba77d8bc),
	.w2(32'h3ad5b1ca),
	.w3(32'hbb37c689),
	.w4(32'h3af56f07),
	.w5(32'h3b04c7a9),
	.w6(32'hbb9824fd),
	.w7(32'h390a3b5b),
	.w8(32'h3b8f26c8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398532ad),
	.w1(32'hbb9c040f),
	.w2(32'hbb512675),
	.w3(32'hbacd9e14),
	.w4(32'hb9634f94),
	.w5(32'h3b225ce4),
	.w6(32'h3aa0d1d2),
	.w7(32'hbaffacde),
	.w8(32'h3b17b0f9),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ab236),
	.w1(32'h3c1d8e57),
	.w2(32'h3bfd65ec),
	.w3(32'h3c442c7c),
	.w4(32'h3c0d15d0),
	.w5(32'h3a23b3ea),
	.w6(32'h3c3c3f4d),
	.w7(32'h3be48afa),
	.w8(32'h3b559851),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b756faf),
	.w1(32'h3b49cb3e),
	.w2(32'hbb5d2381),
	.w3(32'h3b37e179),
	.w4(32'h3a96ece1),
	.w5(32'hbb1b81af),
	.w6(32'hba439fbf),
	.w7(32'hbb0382aa),
	.w8(32'hbb362cbb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8d42f),
	.w1(32'hbaac5b6a),
	.w2(32'h3bf0fb1f),
	.w3(32'hba636f38),
	.w4(32'h3b8167b8),
	.w5(32'h3a10e299),
	.w6(32'h3a1993a8),
	.w7(32'h3bb94375),
	.w8(32'h3b9213d2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6feacd),
	.w1(32'hb8100c57),
	.w2(32'h3b191f9c),
	.w3(32'hbb92293f),
	.w4(32'hbb014e9d),
	.w5(32'hbb932292),
	.w6(32'h3b10ad84),
	.w7(32'h3a85cad7),
	.w8(32'h3b62ee02),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd6d33),
	.w1(32'hb8e06b50),
	.w2(32'hbb9c3cd0),
	.w3(32'hbb551193),
	.w4(32'hbc2563c5),
	.w5(32'hbba78d78),
	.w6(32'h3b8551a8),
	.w7(32'h3b2d3a6b),
	.w8(32'h3a0c8d9d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e8ff3),
	.w1(32'h3b1cbbf9),
	.w2(32'hbb380cf8),
	.w3(32'h3a38e0d3),
	.w4(32'hbc003622),
	.w5(32'hba3b2fc0),
	.w6(32'h3b9bc743),
	.w7(32'hbb127671),
	.w8(32'h3b39a53d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1448ec),
	.w1(32'h3b59925b),
	.w2(32'hbb9f869b),
	.w3(32'h3bede488),
	.w4(32'hbaa5f3bc),
	.w5(32'hb915af41),
	.w6(32'h3c097ed2),
	.w7(32'h39042b3b),
	.w8(32'h3afc4fdb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b3b345),
	.w1(32'h3a082e36),
	.w2(32'h3a8228aa),
	.w3(32'h3a9ad069),
	.w4(32'h3ba01f68),
	.w5(32'hbb31b752),
	.w6(32'h3a787fa9),
	.w7(32'h3a958614),
	.w8(32'h3b2c544d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fadf8),
	.w1(32'hba6dba0c),
	.w2(32'hbbb73aa2),
	.w3(32'hba9b32f9),
	.w4(32'hbba3073c),
	.w5(32'h3acaf84c),
	.w6(32'h3bdc51ea),
	.w7(32'h3b19f1a7),
	.w8(32'hba5e73c6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5056d),
	.w1(32'h39bb730b),
	.w2(32'hbc648526),
	.w3(32'hbb9a8c68),
	.w4(32'hbb5b3392),
	.w5(32'h3999e67a),
	.w6(32'hbc176963),
	.w7(32'hbb5526a2),
	.w8(32'h3bd6c8cb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae47b37),
	.w1(32'h3aa1b63e),
	.w2(32'h3c5b6ab2),
	.w3(32'hbba2839a),
	.w4(32'h3bd70d18),
	.w5(32'h3bc24f5a),
	.w6(32'h3bd738fd),
	.w7(32'h3c2415b3),
	.w8(32'h3c1c4121),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33b600),
	.w1(32'h3c397e77),
	.w2(32'h3c1afb30),
	.w3(32'h3c01afe5),
	.w4(32'h3bbc8523),
	.w5(32'h3bbbd0cf),
	.w6(32'h3c8e9efb),
	.w7(32'h3b3a05f4),
	.w8(32'h3be22564),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83e889),
	.w1(32'h3bd2c164),
	.w2(32'h3bff8bc8),
	.w3(32'h3ba3a23f),
	.w4(32'h3b785ffd),
	.w5(32'hba4e27d6),
	.w6(32'h3bcd5ab9),
	.w7(32'h3ba51c86),
	.w8(32'hba1a0a17),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb276932),
	.w1(32'hbb892449),
	.w2(32'hbb28011c),
	.w3(32'hbb4e3800),
	.w4(32'hbb76e398),
	.w5(32'hbade3207),
	.w6(32'hbaccb4d6),
	.w7(32'hb8ec3037),
	.w8(32'hbb967d86),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6749d),
	.w1(32'hbb54de2b),
	.w2(32'hb8801acd),
	.w3(32'hbb507d30),
	.w4(32'h3b4a0d2c),
	.w5(32'hbba27709),
	.w6(32'hbb9c492b),
	.w7(32'hbacf5302),
	.w8(32'h3af7d660),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba091de8),
	.w1(32'h398f1ea3),
	.w2(32'h3b083092),
	.w3(32'hbc0145a5),
	.w4(32'hbb99f726),
	.w5(32'hbb49e5bc),
	.w6(32'h3ba2f38e),
	.w7(32'h3b713fdf),
	.w8(32'h3c003d1c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c4d05),
	.w1(32'h3b67869d),
	.w2(32'hbb3fc85e),
	.w3(32'hbc0264c4),
	.w4(32'hbb7a64b9),
	.w5(32'hbb75601e),
	.w6(32'h3baed5c8),
	.w7(32'h3c2c3e2e),
	.w8(32'hbb430f3a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9ac48),
	.w1(32'h3bd784d6),
	.w2(32'hba4155ff),
	.w3(32'h3b78dc46),
	.w4(32'h3b121e7c),
	.w5(32'h3b8ed5b9),
	.w6(32'h3bdca0a5),
	.w7(32'h3ac69aed),
	.w8(32'hba47f51e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccc5ca),
	.w1(32'h3b9c2f51),
	.w2(32'h3abd3002),
	.w3(32'h3bf467f2),
	.w4(32'h3c2dbf12),
	.w5(32'h3ba844b4),
	.w6(32'h3c275739),
	.w7(32'h3c0d40ff),
	.w8(32'h3af3e4e8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d3ac6),
	.w1(32'h3934d53b),
	.w2(32'h393eca4d),
	.w3(32'h3bb14347),
	.w4(32'h39c957ab),
	.w5(32'h390fb079),
	.w6(32'h3be2504b),
	.w7(32'h3937723a),
	.w8(32'hbb961604),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b740ab2),
	.w1(32'hbc1e7d76),
	.w2(32'hbc81b0a6),
	.w3(32'hbbdc11a4),
	.w4(32'hbbf67051),
	.w5(32'hbc1c50f4),
	.w6(32'hbc6fa59a),
	.w7(32'hbc560c10),
	.w8(32'hbc203610),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7882c42),
	.w1(32'hba0d3c28),
	.w2(32'h3b1ef645),
	.w3(32'h3b3acd4c),
	.w4(32'h3be9111e),
	.w5(32'hbb36b408),
	.w6(32'h3ad013cc),
	.w7(32'h3bbf0cd5),
	.w8(32'hbb2c333a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c0b8d),
	.w1(32'hb75bfec5),
	.w2(32'h3b7fdc8a),
	.w3(32'hbbae9996),
	.w4(32'h3b3a1cb6),
	.w5(32'h3b362577),
	.w6(32'hbb78c832),
	.w7(32'h3aea4cc7),
	.w8(32'h3b85f8db),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba446feb),
	.w1(32'hbbccd586),
	.w2(32'hbb66dbe8),
	.w3(32'h3be12ff2),
	.w4(32'h3b70b6d6),
	.w5(32'h39c5d405),
	.w6(32'h3b347cbd),
	.w7(32'hbb68bdad),
	.w8(32'h3c33f90a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46e562),
	.w1(32'hbb1a75a1),
	.w2(32'hbbf4745f),
	.w3(32'hbb76eda4),
	.w4(32'hbbacf843),
	.w5(32'h3b774358),
	.w6(32'h3bea294b),
	.w7(32'hb890f9c5),
	.w8(32'h3b22ba94),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f6cf66),
	.w1(32'hbb12187b),
	.w2(32'h3a3dedbc),
	.w3(32'hbaa56ac7),
	.w4(32'hbc04e8ea),
	.w5(32'hba41d3d2),
	.w6(32'hbb716f75),
	.w7(32'hba6a40a5),
	.w8(32'hbb72993b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02a464),
	.w1(32'hbc153e05),
	.w2(32'hbc28abf8),
	.w3(32'hb9aff2ab),
	.w4(32'hb9169807),
	.w5(32'hbb8f7132),
	.w6(32'hbbbbbe32),
	.w7(32'hbabd37fa),
	.w8(32'hbb1139cf),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba34997),
	.w1(32'hbb89dfc9),
	.w2(32'hbc06c609),
	.w3(32'hba8ee97f),
	.w4(32'hbbca5e15),
	.w5(32'hb93d3c6c),
	.w6(32'h39b3e323),
	.w7(32'hbbb2c460),
	.w8(32'h3b3e0b70),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ae515),
	.w1(32'hbb8ef9d1),
	.w2(32'hbb935fc2),
	.w3(32'hbb512bc2),
	.w4(32'h39eb9d98),
	.w5(32'hbac18bf1),
	.w6(32'hbbc52d42),
	.w7(32'hbb4a627f),
	.w8(32'hba624275),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e4656),
	.w1(32'hbb029882),
	.w2(32'hbaf657ea),
	.w3(32'hba66713d),
	.w4(32'h39d96a83),
	.w5(32'h3acf4689),
	.w6(32'hba4df490),
	.w7(32'h3a980b31),
	.w8(32'hbb542549),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ed03e),
	.w1(32'h3aec8aa3),
	.w2(32'h3b88c3ab),
	.w3(32'hb9631d36),
	.w4(32'hbbc3dd31),
	.w5(32'hbb06b192),
	.w6(32'hbac2ccb8),
	.w7(32'hba7ce730),
	.w8(32'hbb353ecd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66163b),
	.w1(32'hba872f7a),
	.w2(32'h3bc1ad11),
	.w3(32'hbbacd5e1),
	.w4(32'h3a0f8813),
	.w5(32'h3a336782),
	.w6(32'hbbbd20ba),
	.w7(32'h3a3d37b5),
	.w8(32'h3b749a54),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ce0ee),
	.w1(32'hba994a01),
	.w2(32'hbb0c5314),
	.w3(32'hb9507b2c),
	.w4(32'h3ad68233),
	.w5(32'h3b13ab2f),
	.w6(32'h3b256933),
	.w7(32'h3b2ed3be),
	.w8(32'h394125bc),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba831ac6),
	.w1(32'hbb0de480),
	.w2(32'hbb78a45d),
	.w3(32'hbac2bd7c),
	.w4(32'hbb4ffd15),
	.w5(32'hbb27486f),
	.w6(32'hbae121a4),
	.w7(32'hbb2fad86),
	.w8(32'hbbf4b118),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd6a63),
	.w1(32'hbb25ef4a),
	.w2(32'h3a4169c0),
	.w3(32'hbbafa48a),
	.w4(32'h39d8c019),
	.w5(32'h3b8b2cec),
	.w6(32'hbc0410b0),
	.w7(32'hbb2bb644),
	.w8(32'h3b75739d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a840aa0),
	.w1(32'h3ac845dd),
	.w2(32'hb9d9a09f),
	.w3(32'h3b517b53),
	.w4(32'h3b8fc6f2),
	.w5(32'hb9dd0cd8),
	.w6(32'h3b66bcea),
	.w7(32'h3aa08bcc),
	.w8(32'h3a845677),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace3b65),
	.w1(32'hbb59ab21),
	.w2(32'hbb161332),
	.w3(32'hbb7b94bd),
	.w4(32'hbb3bb7ba),
	.w5(32'hbaf79642),
	.w6(32'hbb8d9722),
	.w7(32'hba8fe64a),
	.w8(32'hbaa83858),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fa0ef),
	.w1(32'hbaf4dbaa),
	.w2(32'h3ab3fa50),
	.w3(32'hba989640),
	.w4(32'h3b96a72b),
	.w5(32'h3a8544f3),
	.w6(32'hbb8951d1),
	.w7(32'hb8c6614a),
	.w8(32'h3b9ecd07),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25b8d7),
	.w1(32'h3b168a31),
	.w2(32'hbb8d361a),
	.w3(32'hbb24c134),
	.w4(32'hbbd0c17a),
	.w5(32'h3bac5141),
	.w6(32'h3b8b11c3),
	.w7(32'h3ab389e0),
	.w8(32'hbb1e4cfb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31e3ad),
	.w1(32'hbadcac79),
	.w2(32'h3b0eb011),
	.w3(32'h3bb63f5d),
	.w4(32'hba48cb1e),
	.w5(32'hb7da3d8b),
	.w6(32'hbba51782),
	.w7(32'hbb96dd22),
	.w8(32'hbb4c3c30),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7df9bf),
	.w1(32'h3c00818c),
	.w2(32'h3c0dac75),
	.w3(32'h3c3188f8),
	.w4(32'h3c2b2488),
	.w5(32'h3a6449bc),
	.w6(32'h3bbf25e1),
	.w7(32'h3b8c06d5),
	.w8(32'hbb9fee40),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb38322),
	.w1(32'hbbde4c77),
	.w2(32'hbc4a06af),
	.w3(32'hbb3e12df),
	.w4(32'hbc419a88),
	.w5(32'hbc4145fa),
	.w6(32'hbbbfe7d2),
	.w7(32'hbc58cc1a),
	.w8(32'hbbf6e580),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf77e37),
	.w1(32'h3b982754),
	.w2(32'h3b38e808),
	.w3(32'h3931a293),
	.w4(32'h3aa5ada2),
	.w5(32'h3aa0d5a6),
	.w6(32'h3c3bd03b),
	.w7(32'h3c041759),
	.w8(32'h3b58de06),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeca1b2),
	.w1(32'hbb202b11),
	.w2(32'hba206b2c),
	.w3(32'hbbb0e97c),
	.w4(32'hbb4e878a),
	.w5(32'h3a3c5511),
	.w6(32'h39c4f537),
	.w7(32'h3b4cdd3a),
	.w8(32'hbaf1884f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83da39),
	.w1(32'hbaaaf6e8),
	.w2(32'hbb43c8fb),
	.w3(32'hb8b75cdf),
	.w4(32'hbb5744ef),
	.w5(32'h3a88682d),
	.w6(32'hba2d602d),
	.w7(32'hbb56254e),
	.w8(32'hb9000ab7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76c9a2),
	.w1(32'h3bc8b1fc),
	.w2(32'h3baceba6),
	.w3(32'h380201c3),
	.w4(32'h3a4170c8),
	.w5(32'hb9784d26),
	.w6(32'hb85d8f42),
	.w7(32'hbb062b24),
	.w8(32'h3af380f0),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b261ae3),
	.w1(32'hbae0fc08),
	.w2(32'hbb799ae9),
	.w3(32'h3b091e4e),
	.w4(32'h3a5a86f9),
	.w5(32'hbb92b8f7),
	.w6(32'h3acfcd1c),
	.w7(32'hbb1af0fb),
	.w8(32'h3ae768e1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2ce18),
	.w1(32'h3bfbf9fb),
	.w2(32'h3c874149),
	.w3(32'h3a8cd56d),
	.w4(32'h3b669315),
	.w5(32'h3a3d7f9c),
	.w6(32'h3b7d6436),
	.w7(32'h3c4bf542),
	.w8(32'h3b5af499),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7929f59),
	.w1(32'hbc09eba0),
	.w2(32'hbc5dea0e),
	.w3(32'hb93d0c4d),
	.w4(32'hbc101a99),
	.w5(32'hbba14ec5),
	.w6(32'hbb2c6546),
	.w7(32'hbc0e193c),
	.w8(32'hbb08bd0a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6bb1f),
	.w1(32'hbc162657),
	.w2(32'hbbe78c79),
	.w3(32'hbb9bb329),
	.w4(32'hbc0bfa83),
	.w5(32'hbc2b6afd),
	.w6(32'hbc3237a2),
	.w7(32'hbb9a82c7),
	.w8(32'hbb752442),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa850b),
	.w1(32'h3b4e29ea),
	.w2(32'h3ac4064c),
	.w3(32'h3a35362a),
	.w4(32'hba902b46),
	.w5(32'h3bcb103f),
	.w6(32'h3c2f3032),
	.w7(32'h3bf2021a),
	.w8(32'h3b22376d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c07de),
	.w1(32'hbae056cf),
	.w2(32'hbab22b36),
	.w3(32'h3b4f7482),
	.w4(32'h3b0ed5db),
	.w5(32'h3ac948b2),
	.w6(32'hbacd5bd4),
	.w7(32'hbb15b742),
	.w8(32'hbafabad6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f897e),
	.w1(32'hba845691),
	.w2(32'hbabbff8d),
	.w3(32'h3b697305),
	.w4(32'h3b7abada),
	.w5(32'hb94068b2),
	.w6(32'hbb33ee31),
	.w7(32'hba03536c),
	.w8(32'hbb050a0c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a669111),
	.w1(32'h3a27c481),
	.w2(32'h3bb056a2),
	.w3(32'h3b4df2bc),
	.w4(32'h3bd667be),
	.w5(32'hba3225d2),
	.w6(32'h3ba50c89),
	.w7(32'h3c04cdb4),
	.w8(32'h3ab3da51),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8dff3),
	.w1(32'hbb2319d4),
	.w2(32'hbbaec9f2),
	.w3(32'h3a2e64ca),
	.w4(32'hba71588f),
	.w5(32'hbb9b657e),
	.w6(32'h3b89f8b5),
	.w7(32'h3a421095),
	.w8(32'hbb847644),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91bdde),
	.w1(32'hbb5f2941),
	.w2(32'h3b936d74),
	.w3(32'hbb09c9b4),
	.w4(32'hba7886d5),
	.w5(32'hbad43074),
	.w6(32'hbbdba008),
	.w7(32'hba39b810),
	.w8(32'hbb18f020),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d7696),
	.w1(32'h3b8c6f54),
	.w2(32'h3a599445),
	.w3(32'h3b3e982c),
	.w4(32'hbb69772e),
	.w5(32'h3b3eb213),
	.w6(32'h3b130f42),
	.w7(32'hbbbd703a),
	.w8(32'h3b1703f7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c5029),
	.w1(32'h3b359293),
	.w2(32'h3b520669),
	.w3(32'h3b041a51),
	.w4(32'hbaef4682),
	.w5(32'hbb6a2547),
	.w6(32'hbaab5a8c),
	.w7(32'hbaa45018),
	.w8(32'h3a1f18e3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3739c84a),
	.w1(32'h3a75526a),
	.w2(32'h3bc681be),
	.w3(32'hbb8fb391),
	.w4(32'h3ad046f7),
	.w5(32'h38bae534),
	.w6(32'hbb4af23a),
	.w7(32'h3bc9cc05),
	.w8(32'hbb286283),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1be3dc),
	.w1(32'hbacc42e0),
	.w2(32'h3c96571d),
	.w3(32'h3925a2c0),
	.w4(32'h3bf5d450),
	.w5(32'h3ba6584d),
	.w6(32'h3a14903a),
	.w7(32'h3c14fba3),
	.w8(32'h3c01e138),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10d46f),
	.w1(32'h3b3a97ec),
	.w2(32'hb9d993ac),
	.w3(32'h3b6e6478),
	.w4(32'h3a982616),
	.w5(32'h3b6f77cf),
	.w6(32'h3c106cbe),
	.w7(32'h3b8a61e6),
	.w8(32'h3b712093),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92480a),
	.w1(32'hba194675),
	.w2(32'hba836136),
	.w3(32'h3a861183),
	.w4(32'h3b44b325),
	.w5(32'hbc03a998),
	.w6(32'h3a918bb9),
	.w7(32'h3ac8f61d),
	.w8(32'hbc1140ae),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8ce55),
	.w1(32'hbc032af0),
	.w2(32'hbbed0b5d),
	.w3(32'hbc0ca4f2),
	.w4(32'hbc82a43f),
	.w5(32'hbb4fe450),
	.w6(32'hbcb029c9),
	.w7(32'hbc4aa573),
	.w8(32'hbbd11b5f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62fc0f),
	.w1(32'hb9e77a8e),
	.w2(32'hbaa20e3e),
	.w3(32'h3bd10c89),
	.w4(32'h3bc3ee4b),
	.w5(32'hba6148f2),
	.w6(32'h3b830c4d),
	.w7(32'h3af6adc7),
	.w8(32'h3a636eb9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6302a),
	.w1(32'h3c831cf8),
	.w2(32'hbb74f92f),
	.w3(32'h3b6fa957),
	.w4(32'hbc41fc99),
	.w5(32'hbb29e62b),
	.w6(32'h3c059527),
	.w7(32'hb999cc6e),
	.w8(32'hbb9ea549),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba970816),
	.w1(32'h3b87aa83),
	.w2(32'h3b8386af),
	.w3(32'h3bf76d7a),
	.w4(32'h3b0f59af),
	.w5(32'h3c57f42d),
	.w6(32'h3b71ee8e),
	.w7(32'h3b8c6fb5),
	.w8(32'h3c9b3853),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc329c7a),
	.w1(32'h3d0cd627),
	.w2(32'h3a98e3e5),
	.w3(32'h3cd9ddf5),
	.w4(32'hbb5077c6),
	.w5(32'hbb7ef4f1),
	.w6(32'h3d08b3d8),
	.w7(32'h3cc0f7a1),
	.w8(32'hbba10192),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae77db9),
	.w1(32'h3c0116aa),
	.w2(32'h3b51a2f2),
	.w3(32'h3b1a7699),
	.w4(32'hbb0452c5),
	.w5(32'h390c2d6c),
	.w6(32'h3ba379f7),
	.w7(32'h3a994bad),
	.w8(32'h3ba0cf3f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0b3a9),
	.w1(32'hbba1e5b8),
	.w2(32'hbb4ded83),
	.w3(32'hbb73a567),
	.w4(32'hbb36bb4f),
	.w5(32'h3b3a2660),
	.w6(32'h3bcea2e2),
	.w7(32'h3bee923b),
	.w8(32'h3b9fdd52),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be33533),
	.w1(32'h3b7839d9),
	.w2(32'h3a90f5d7),
	.w3(32'h3bb3afe6),
	.w4(32'h3c000437),
	.w5(32'hbbacb404),
	.w6(32'h3b8eb1b8),
	.w7(32'h3a92ebbe),
	.w8(32'hbb1adcae),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10161d),
	.w1(32'h3b9d688d),
	.w2(32'hbbd25e78),
	.w3(32'h3c229d2f),
	.w4(32'h3c18cf98),
	.w5(32'hbb7328e8),
	.w6(32'h3bb13349),
	.w7(32'h3c047c58),
	.w8(32'hbc007ce2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae51c27),
	.w1(32'hbb82c561),
	.w2(32'hbb9224d1),
	.w3(32'hbbc69992),
	.w4(32'h3a634305),
	.w5(32'h3bc634b0),
	.w6(32'hbc371a10),
	.w7(32'hbb94b1b4),
	.w8(32'hbb917fd1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0284f5),
	.w1(32'hbc3b1cda),
	.w2(32'hbc22c839),
	.w3(32'hbb4047f1),
	.w4(32'hbbfdf19f),
	.w5(32'hbb9809cd),
	.w6(32'hbc837fea),
	.w7(32'hbc27844a),
	.w8(32'h3bdb0668),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb69975),
	.w1(32'h3c25f1d9),
	.w2(32'h3c425b34),
	.w3(32'h3b98e2d6),
	.w4(32'h3c8d83c7),
	.w5(32'h3c740250),
	.w6(32'h3becda74),
	.w7(32'h3c7d1766),
	.w8(32'h3b080f1e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedd993),
	.w1(32'h3b9a0d85),
	.w2(32'h3b1cfa04),
	.w3(32'h3c1a5a56),
	.w4(32'h3c585d14),
	.w5(32'h3ba9fe88),
	.w6(32'h3b311c67),
	.w7(32'h3be98b09),
	.w8(32'h3b7851c7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4bd9f),
	.w1(32'hbb332839),
	.w2(32'hbc120dbb),
	.w3(32'hbb6157d8),
	.w4(32'h3b365cf9),
	.w5(32'h3b1aa39b),
	.w6(32'hbba8d5e6),
	.w7(32'h3b41aa1a),
	.w8(32'hb923a191),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b090b26),
	.w1(32'h3b769554),
	.w2(32'h3b45c618),
	.w3(32'h3bba5fb8),
	.w4(32'h3bfa212c),
	.w5(32'h3bb0d6f4),
	.w6(32'h3bc9ae49),
	.w7(32'h3c0a913b),
	.w8(32'hbb2b0b01),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae148f1),
	.w1(32'hbc865cea),
	.w2(32'hbcd313a9),
	.w3(32'hbb1b85a0),
	.w4(32'hbc585546),
	.w5(32'hbc82726b),
	.w6(32'hbce2a09d),
	.w7(32'hbc890af1),
	.w8(32'hbc2e79c8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c53ec),
	.w1(32'h39ebc7f0),
	.w2(32'hbb4027b8),
	.w3(32'hba400f4f),
	.w4(32'hbb3b72af),
	.w5(32'h3c17c2c4),
	.w6(32'h3b19568f),
	.w7(32'hbb195e9e),
	.w8(32'hb9c7a5a8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e71ded),
	.w1(32'hbbee8b96),
	.w2(32'hbb1136b8),
	.w3(32'h3b90de8f),
	.w4(32'h3c1fbd3c),
	.w5(32'hbb3744b8),
	.w6(32'hbb9a889a),
	.w7(32'hbb9ef297),
	.w8(32'h3ac065e3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6437e8),
	.w1(32'hba10721f),
	.w2(32'hb9dda788),
	.w3(32'hbb12f1fa),
	.w4(32'hbb11d7c6),
	.w5(32'h3be0c39d),
	.w6(32'hbb285d83),
	.w7(32'hbb7a8ef8),
	.w8(32'h3b1992d4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b349000),
	.w1(32'h399166a9),
	.w2(32'hbadf98e2),
	.w3(32'hbb22a988),
	.w4(32'h3bac63f1),
	.w5(32'hbb4aefe7),
	.w6(32'hbc043ad6),
	.w7(32'hbb884903),
	.w8(32'hbb04f4d4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3ef7d),
	.w1(32'h3b63bfb2),
	.w2(32'hbaaae21e),
	.w3(32'hbb1d98dd),
	.w4(32'h3b176faf),
	.w5(32'h398df164),
	.w6(32'h39badbe0),
	.w7(32'h3b438bc9),
	.w8(32'hbc2256c2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc336796),
	.w1(32'hbc04a100),
	.w2(32'h3b8c05eb),
	.w3(32'h3c0b102e),
	.w4(32'h3c917da4),
	.w5(32'hbb60845c),
	.w6(32'hbbcb30a9),
	.w7(32'h3be016ba),
	.w8(32'hbb6699e5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2f385),
	.w1(32'hbb558ee2),
	.w2(32'hbb0ace00),
	.w3(32'hbb80c5f7),
	.w4(32'hbb85abb8),
	.w5(32'hbb9eed78),
	.w6(32'hbb80a20c),
	.w7(32'hbb2ad795),
	.w8(32'hba140a61),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8246b3),
	.w1(32'hbba09277),
	.w2(32'hbad3ec88),
	.w3(32'hbba7865a),
	.w4(32'hbaeea904),
	.w5(32'hbb25f34a),
	.w6(32'hbba1812a),
	.w7(32'h3b14ef43),
	.w8(32'h3b479252),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9181a9),
	.w1(32'hbb42cf12),
	.w2(32'hbb398228),
	.w3(32'hbc221347),
	.w4(32'hbbc7c750),
	.w5(32'h3adbc19e),
	.w6(32'hb9ca213c),
	.w7(32'hbb8586ad),
	.w8(32'hbba40642),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3e1c9),
	.w1(32'h3adcec38),
	.w2(32'h3ac92be3),
	.w3(32'hbb91e18b),
	.w4(32'hbb8b6cee),
	.w5(32'h3b13194b),
	.w6(32'h3c44033a),
	.w7(32'hbbd210b4),
	.w8(32'hbb8f2045),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b0938),
	.w1(32'hbb6e9a78),
	.w2(32'h39c17fc8),
	.w3(32'hbb42f30e),
	.w4(32'hbad5d846),
	.w5(32'hbabaf024),
	.w6(32'hbbd45097),
	.w7(32'hbb0c5090),
	.w8(32'h3bbc97f2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc152cb),
	.w1(32'h3bea0a1c),
	.w2(32'hbb4451c9),
	.w3(32'hbbb77d18),
	.w4(32'hbb7ad18b),
	.w5(32'h3bd3dff6),
	.w6(32'h3b20a64b),
	.w7(32'hbb67b0df),
	.w8(32'h3acc5932),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf609a5),
	.w1(32'hba546a00),
	.w2(32'hba021aba),
	.w3(32'h3b5182b8),
	.w4(32'h3b8b67da),
	.w5(32'h3b8ef616),
	.w6(32'hbb1756e5),
	.w7(32'h3ae1da2d),
	.w8(32'h3b346477),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bbe14),
	.w1(32'h3a99070b),
	.w2(32'h3b87b652),
	.w3(32'hb81671f8),
	.w4(32'h3bf11c29),
	.w5(32'hbc541f1f),
	.w6(32'hba2c99f5),
	.w7(32'h3b3684e3),
	.w8(32'hbc822522),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33af36),
	.w1(32'hbc5bab75),
	.w2(32'hbbcc220b),
	.w3(32'hbc712f17),
	.w4(32'hbb53fccf),
	.w5(32'h3a831a58),
	.w6(32'hbc8eae84),
	.w7(32'hbc3aefc2),
	.w8(32'hbb12bd31),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c28f5),
	.w1(32'hbb5f0ea1),
	.w2(32'hbb58677d),
	.w3(32'hbb7b4c27),
	.w4(32'hbb8b6056),
	.w5(32'h3b078c67),
	.w6(32'hbb9e9e9f),
	.w7(32'hba982ec3),
	.w8(32'h3b8535a3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b797cdd),
	.w1(32'hbb7d7e50),
	.w2(32'h3a0df250),
	.w3(32'h3acff63e),
	.w4(32'hba24667e),
	.w5(32'hbb85cd14),
	.w6(32'hbb947699),
	.w7(32'hb9f5b639),
	.w8(32'hbb42b3d4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cef59),
	.w1(32'h3ab858a8),
	.w2(32'h3b507ab3),
	.w3(32'h3b395099),
	.w4(32'h3bd6c70b),
	.w5(32'h3b71a591),
	.w6(32'h3bcee118),
	.w7(32'h3b0fd929),
	.w8(32'h3af28492),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd4f99),
	.w1(32'h3a842e42),
	.w2(32'h3b82d14f),
	.w3(32'hbb1e07dc),
	.w4(32'hbb98397d),
	.w5(32'h3b0ed861),
	.w6(32'hbac413d4),
	.w7(32'hbb0ae507),
	.w8(32'hbbbd88eb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8876c2),
	.w1(32'hbb1750d4),
	.w2(32'hba87b506),
	.w3(32'h3baf4507),
	.w4(32'h3afb9e25),
	.w5(32'hbb14f8a1),
	.w6(32'hbb1718f4),
	.w7(32'h3a73e32f),
	.w8(32'hba8a4257),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c6cd9),
	.w1(32'hba9392f1),
	.w2(32'h3950ba6e),
	.w3(32'h38fbff3a),
	.w4(32'h3a8de066),
	.w5(32'hbb3403b5),
	.w6(32'h3b8a8597),
	.w7(32'h38861764),
	.w8(32'h3b478325),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e0e46),
	.w1(32'h3a9dc3b5),
	.w2(32'hba9d1e01),
	.w3(32'hbb00f375),
	.w4(32'h3b954352),
	.w5(32'h3b900a6f),
	.w6(32'hbc00ff55),
	.w7(32'hb9f203c4),
	.w8(32'h3b95b01b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b038cfb),
	.w1(32'h3bc122e9),
	.w2(32'hba954f77),
	.w3(32'h3900457f),
	.w4(32'hb9da796e),
	.w5(32'hbc28ab2f),
	.w6(32'h3be1ee8c),
	.w7(32'hbabadc72),
	.w8(32'hbba81e29),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbede0d4),
	.w1(32'hbc43e84e),
	.w2(32'hbc7b7590),
	.w3(32'hbc7128f9),
	.w4(32'hbc760ec7),
	.w5(32'h3b6d47af),
	.w6(32'hbbecc70d),
	.w7(32'hbc1c0bd9),
	.w8(32'h39519540),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ff789),
	.w1(32'hbb92413d),
	.w2(32'hbb8376e8),
	.w3(32'h3a8b7038),
	.w4(32'hbc0057a0),
	.w5(32'hba868ba8),
	.w6(32'h3b37e40f),
	.w7(32'hbbff003f),
	.w8(32'hbb8ab3e9),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19e037),
	.w1(32'hbbe2e290),
	.w2(32'hbb5b9bf3),
	.w3(32'hba9226e3),
	.w4(32'h3b48df28),
	.w5(32'hbbddcc08),
	.w6(32'hbbc7134d),
	.w7(32'h3a25fa0e),
	.w8(32'hbb368f53),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19e9bd),
	.w1(32'hbb214f27),
	.w2(32'h3afbcb22),
	.w3(32'hbaebeb37),
	.w4(32'h3bdc9cca),
	.w5(32'h3b932300),
	.w6(32'hbbe2b8c8),
	.w7(32'h3b1cc35b),
	.w8(32'h3ba74195),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80593f),
	.w1(32'hbb90d9e4),
	.w2(32'hbb57bab6),
	.w3(32'h3bd90a99),
	.w4(32'h3c510e95),
	.w5(32'hbba5f678),
	.w6(32'hba6315bd),
	.w7(32'h3bec9642),
	.w8(32'hbaf7c292),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983dbda),
	.w1(32'h39bda130),
	.w2(32'h3b4b5282),
	.w3(32'hbbd28294),
	.w4(32'h3a9d6b80),
	.w5(32'h3bd54666),
	.w6(32'hbc3208ff),
	.w7(32'hba6b8d53),
	.w8(32'h3c44a210),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c081c82),
	.w1(32'h3b68f5cf),
	.w2(32'hbbfc3540),
	.w3(32'hbb31e864),
	.w4(32'hbb4d043f),
	.w5(32'hbc196bf1),
	.w6(32'hbc0f8195),
	.w7(32'hbbe00cde),
	.w8(32'hbc138625),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3821ceb5),
	.w1(32'hbb18f845),
	.w2(32'hbbc0f4d1),
	.w3(32'hbbe4d1b8),
	.w4(32'h3a1d0a89),
	.w5(32'hb57c7cee),
	.w6(32'hbbd6fe18),
	.w7(32'hbb8bcf19),
	.w8(32'h3b9b7ca8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba853606),
	.w1(32'hba40988b),
	.w2(32'hbbb82405),
	.w3(32'hbbdb341c),
	.w4(32'hba9c1958),
	.w5(32'hbbb4064d),
	.w6(32'hbb914c80),
	.w7(32'hbb0371e9),
	.w8(32'hbba2c45f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c866fe),
	.w1(32'hbbc0485d),
	.w2(32'hbbfd60f9),
	.w3(32'hbc0d8bad),
	.w4(32'hbb4e4ce1),
	.w5(32'hbc01e65f),
	.w6(32'hbc86320b),
	.w7(32'hbbc9b087),
	.w8(32'hbb44c402),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ea4faa),
	.w1(32'hba702f27),
	.w2(32'h3b004fe6),
	.w3(32'hbbcbdfe9),
	.w4(32'h3a54b624),
	.w5(32'h3a9f6225),
	.w6(32'hbc3ede1d),
	.w7(32'hbb44698a),
	.w8(32'h395a3030),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde0ffc),
	.w1(32'hbbc3453b),
	.w2(32'hbbc8a1a5),
	.w3(32'hbb05d9bc),
	.w4(32'h3b9115d8),
	.w5(32'hbbc64e17),
	.w6(32'hba495ebc),
	.w7(32'h3b8bdd01),
	.w8(32'hbbc5182e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc525ce),
	.w1(32'hbbecb6fd),
	.w2(32'hbbf16b3f),
	.w3(32'hbbd83fcb),
	.w4(32'hbbdf2da1),
	.w5(32'h3a9efc25),
	.w6(32'hbb920679),
	.w7(32'hbb98fe41),
	.w8(32'h3ae577cb),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06b571),
	.w1(32'h3b2ee387),
	.w2(32'h3b81bf25),
	.w3(32'h3afa5e92),
	.w4(32'h3ba744bf),
	.w5(32'h3b50b338),
	.w6(32'h3c07e3c9),
	.w7(32'h3baf87bb),
	.w8(32'hbaf06bcb),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93805c),
	.w1(32'h3afc5b46),
	.w2(32'h3c430af5),
	.w3(32'h3be643d7),
	.w4(32'h3c98e020),
	.w5(32'hbb2581ee),
	.w6(32'hbc0ab695),
	.w7(32'h3c4deb6d),
	.w8(32'hbaa2babb),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea3163),
	.w1(32'hbb181875),
	.w2(32'hbb19ca44),
	.w3(32'hbb02417e),
	.w4(32'h3bd4c74e),
	.w5(32'hba9a64c5),
	.w6(32'hbbd95cc3),
	.w7(32'h3b819099),
	.w8(32'h3b9bb1dd),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61505e),
	.w1(32'h3add39b3),
	.w2(32'h3a318675),
	.w3(32'hbb7ade9e),
	.w4(32'hbac88e71),
	.w5(32'h3ad7e608),
	.w6(32'hbb1aaa6e),
	.w7(32'hbaf4d266),
	.w8(32'hb9894f41),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7c532),
	.w1(32'hb8caefc8),
	.w2(32'h3aa129a6),
	.w3(32'hba8b23b1),
	.w4(32'hba4c2630),
	.w5(32'hbabd1288),
	.w6(32'hbaf299a7),
	.w7(32'hba9ea69b),
	.w8(32'hbc07e4fb),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70344d),
	.w1(32'hba2e902f),
	.w2(32'h3b85b51a),
	.w3(32'h3b5a221d),
	.w4(32'h3c25452d),
	.w5(32'hbb9c667a),
	.w6(32'hbb9d127f),
	.w7(32'h3b352c5d),
	.w8(32'h3979dade),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e23a01),
	.w1(32'hbb7bd609),
	.w2(32'hbb3b72a1),
	.w3(32'hbb910d45),
	.w4(32'hbbd6ae89),
	.w5(32'hbb9f419a),
	.w6(32'h3ab6cb18),
	.w7(32'hbb7f76d0),
	.w8(32'h3a6a847b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c4842),
	.w1(32'hb9870d69),
	.w2(32'hbb786a60),
	.w3(32'hbbc97862),
	.w4(32'h3ac8d834),
	.w5(32'hbb40c6fe),
	.w6(32'hbb9f8e52),
	.w7(32'hbafab720),
	.w8(32'h3b933a23),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40bbf1),
	.w1(32'h3bf36374),
	.w2(32'h3b364a89),
	.w3(32'h3ac2f067),
	.w4(32'h3b94037f),
	.w5(32'hbb8b3a3e),
	.w6(32'h3bb19ba9),
	.w7(32'h3bdbe760),
	.w8(32'h370d05f5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3931e47b),
	.w1(32'h3a786ec2),
	.w2(32'hba90d3e6),
	.w3(32'h3aa2f8c8),
	.w4(32'h3884349e),
	.w5(32'hbbe681e7),
	.w6(32'h3b91f162),
	.w7(32'hbaa7838a),
	.w8(32'hbc0ce80e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc294002),
	.w1(32'hbbe42224),
	.w2(32'hbc75fb0b),
	.w3(32'hbc2ebf4e),
	.w4(32'h393caa26),
	.w5(32'hbbb47fd2),
	.w6(32'hbc48ea71),
	.w7(32'hbae4cf01),
	.w8(32'hbc6ef3b7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0a772),
	.w1(32'hbb579f52),
	.w2(32'hba537e71),
	.w3(32'hbafb1c6a),
	.w4(32'h3b05c12e),
	.w5(32'hbb479d0d),
	.w6(32'hb910c685),
	.w7(32'hba5d0c11),
	.w8(32'h3a6af476),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1ea0a),
	.w1(32'h3b8a7db6),
	.w2(32'h3c0415b5),
	.w3(32'h3b1d5a6d),
	.w4(32'h3c38af3b),
	.w5(32'h3bbed226),
	.w6(32'hbc0df9a4),
	.w7(32'h3b6163c9),
	.w8(32'h3be140ec),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99cd6f),
	.w1(32'h37ff4cb7),
	.w2(32'hbb2ebdf0),
	.w3(32'h3b415a43),
	.w4(32'h3b800397),
	.w5(32'hbb80da87),
	.w6(32'h3a6baaa4),
	.w7(32'h3b34d9aa),
	.w8(32'hbb05b49e),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ecea7),
	.w1(32'hbbc05caa),
	.w2(32'hbc107d84),
	.w3(32'hbc494891),
	.w4(32'hbc253b11),
	.w5(32'hbb4edd84),
	.w6(32'hbb8e3544),
	.w7(32'hbb7044c5),
	.w8(32'hbadaec80),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf996c1),
	.w1(32'h3a6d8336),
	.w2(32'h3a98cf77),
	.w3(32'hbba99612),
	.w4(32'h39140a43),
	.w5(32'h3b8d0a4c),
	.w6(32'hbae5bbce),
	.w7(32'hbb8e092f),
	.w8(32'h3bad9eff),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e60ae),
	.w1(32'hbbad4edb),
	.w2(32'h3ad5ee3b),
	.w3(32'hbb34000f),
	.w4(32'hbba51fc3),
	.w5(32'hbacbb849),
	.w6(32'hbb8dfcce),
	.w7(32'hbb5120c4),
	.w8(32'hbc00c51d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc170ab0),
	.w1(32'hbbf6188d),
	.w2(32'hbb0be43f),
	.w3(32'hbb7cd997),
	.w4(32'hbb94a44b),
	.w5(32'hbac4fb22),
	.w6(32'hbb4970d7),
	.w7(32'hbbceda7b),
	.w8(32'h3b5bf598),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb795689),
	.w1(32'h3b1a623b),
	.w2(32'hbac06fd9),
	.w3(32'hbc3a0dda),
	.w4(32'hbbc46000),
	.w5(32'hbb2ddfa2),
	.w6(32'h3bd2195c),
	.w7(32'hbb230c69),
	.w8(32'hbb56fd0a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d9159),
	.w1(32'h3baef6e0),
	.w2(32'h3c002469),
	.w3(32'h3b460d5c),
	.w4(32'h3bdb85ae),
	.w5(32'hba901f28),
	.w6(32'h3abdcd58),
	.w7(32'h3a57820c),
	.w8(32'hbb3a68c2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaebf88),
	.w1(32'hba7a3ce7),
	.w2(32'h3a2f2de5),
	.w3(32'hb9d036bf),
	.w4(32'hbb129159),
	.w5(32'h3ae30944),
	.w6(32'hbb651e3a),
	.w7(32'hbb64a2b9),
	.w8(32'hbb90aeea),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b1580),
	.w1(32'h3a88c95a),
	.w2(32'h3a8804ab),
	.w3(32'h3adc93f7),
	.w4(32'h3b5f9e5b),
	.w5(32'hbae9d908),
	.w6(32'h3a5cb0be),
	.w7(32'hba962e1c),
	.w8(32'hbbb8de7c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74521e),
	.w1(32'hba81fdf0),
	.w2(32'hb9d05b81),
	.w3(32'hbbd2aef6),
	.w4(32'hbbb9730f),
	.w5(32'h3af3c3e1),
	.w6(32'hbb17feca),
	.w7(32'hbb242e3a),
	.w8(32'hbaf9a36a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06e484),
	.w1(32'h3b5baa99),
	.w2(32'h3b00e03d),
	.w3(32'h3c2f8f57),
	.w4(32'h3b0d3ffb),
	.w5(32'hba4125b9),
	.w6(32'h3becc0b6),
	.w7(32'h3ac0f782),
	.w8(32'h39197f3b),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baca345),
	.w1(32'hbaaee6d9),
	.w2(32'hbbbe006b),
	.w3(32'hbab0ae2e),
	.w4(32'h3bc33248),
	.w5(32'h3ad99e25),
	.w6(32'hbc3b2b70),
	.w7(32'hbad4bccc),
	.w8(32'hbb2cf83d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e8d71),
	.w1(32'h3b90015c),
	.w2(32'h3b8d7571),
	.w3(32'hba3b4dc0),
	.w4(32'hbb2dcaa9),
	.w5(32'hbb807a45),
	.w6(32'h3a739a00),
	.w7(32'h39a0bd85),
	.w8(32'h3c1bf7f3),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be327fe),
	.w1(32'h3af228c0),
	.w2(32'hbaf525e3),
	.w3(32'h3b2dcaac),
	.w4(32'hbabf4631),
	.w5(32'h3b556937),
	.w6(32'h3abdbbf9),
	.w7(32'h3bcf8a49),
	.w8(32'h3a352f4b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08f50b),
	.w1(32'hbbbd055c),
	.w2(32'hbb9b2748),
	.w3(32'hbb03dbad),
	.w4(32'hbb4fa07d),
	.w5(32'hba5b78c8),
	.w6(32'hbbc7a764),
	.w7(32'hbb8bdb10),
	.w8(32'h3bd5a876),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43177f),
	.w1(32'h3c0f5a5f),
	.w2(32'h3bbdf80c),
	.w3(32'h3ba55524),
	.w4(32'h3c34c587),
	.w5(32'hbb2e991e),
	.w6(32'hbb589be8),
	.w7(32'h3ba2c9bf),
	.w8(32'hbc19f00b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d2baf),
	.w1(32'hbbfcaf18),
	.w2(32'hbb6e3b1a),
	.w3(32'hbbaca7d0),
	.w4(32'h3a404e3c),
	.w5(32'h3be6f6d9),
	.w6(32'hbaeb52ee),
	.w7(32'h3b076cdb),
	.w8(32'hbb67516e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42672b),
	.w1(32'hbbc29148),
	.w2(32'h38cdd11c),
	.w3(32'hbb35e510),
	.w4(32'h3b847d6b),
	.w5(32'hbb976085),
	.w6(32'hbc2423cc),
	.w7(32'hbb992d4f),
	.w8(32'h3b123f7b),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03c6df),
	.w1(32'h3b467858),
	.w2(32'h3a3c5bae),
	.w3(32'hbb998aa3),
	.w4(32'hbb4ffcca),
	.w5(32'hbb92dc2c),
	.w6(32'hbba7b191),
	.w7(32'hbb9a4f62),
	.w8(32'h3b312890),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba827586),
	.w1(32'hbadc4bdd),
	.w2(32'hba82b7a4),
	.w3(32'hbb95d472),
	.w4(32'hbbb41ba2),
	.w5(32'hba674cb5),
	.w6(32'hbb26e29b),
	.w7(32'hba9d4519),
	.w8(32'hbb783e13),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeeb195),
	.w1(32'hbc2acaf1),
	.w2(32'hbb8b8501),
	.w3(32'hb996f441),
	.w4(32'h3b9f5146),
	.w5(32'hbb619d50),
	.w6(32'hbc637c25),
	.w7(32'hba1688e4),
	.w8(32'h393f3a9c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01c36b),
	.w1(32'h3b5bb2ce),
	.w2(32'h39c9a05d),
	.w3(32'h3b1fa48d),
	.w4(32'h3b252300),
	.w5(32'hbabab367),
	.w6(32'h3bfe7884),
	.w7(32'h3c0c3244),
	.w8(32'hb68a4180),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f18a0),
	.w1(32'hba3ecd84),
	.w2(32'hbba7ac35),
	.w3(32'hbaebb116),
	.w4(32'hbbbd7fc9),
	.w5(32'h3aa661d8),
	.w6(32'h3a369675),
	.w7(32'hbb9bac07),
	.w8(32'h3c2df526),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00dc6d),
	.w1(32'h3be848e8),
	.w2(32'h3b994498),
	.w3(32'h3b652812),
	.w4(32'h3c261509),
	.w5(32'h3c2bf4b5),
	.w6(32'h3b019bfa),
	.w7(32'h3bfd8b62),
	.w8(32'h3b32c8b3),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5e3f7),
	.w1(32'hbbec2712),
	.w2(32'hbb124d9a),
	.w3(32'hbb695cc4),
	.w4(32'hbbd6faac),
	.w5(32'h3ba5238e),
	.w6(32'hbc047648),
	.w7(32'hbbdc89ca),
	.w8(32'h3ab9b19b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b805af2),
	.w1(32'hbb53a2db),
	.w2(32'hba801f80),
	.w3(32'hbba78229),
	.w4(32'hbb215224),
	.w5(32'hbb8a7992),
	.w6(32'h3ab637d7),
	.w7(32'hbb6581c4),
	.w8(32'hbb901d7a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76aec6),
	.w1(32'hbb15f42c),
	.w2(32'h3b707cd6),
	.w3(32'h39d1a0a0),
	.w4(32'h3ac14850),
	.w5(32'h3a554582),
	.w6(32'h3a0a0a43),
	.w7(32'h3bb610bb),
	.w8(32'h3bc65ff4),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dbba4),
	.w1(32'hbb5e3207),
	.w2(32'h3737b296),
	.w3(32'h3bf093e9),
	.w4(32'h3a1cada1),
	.w5(32'hbbe98530),
	.w6(32'hbab564fd),
	.w7(32'h3aa442e1),
	.w8(32'hbabf0f1d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9e80e),
	.w1(32'hbb44279e),
	.w2(32'hbbb7c3f7),
	.w3(32'hbb697889),
	.w4(32'hbb770f3b),
	.w5(32'h3ba5d8c7),
	.w6(32'h394855ec),
	.w7(32'hbb6b8f5a),
	.w8(32'hbaffa99d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb473434),
	.w1(32'hbb71d084),
	.w2(32'hbb69fe52),
	.w3(32'hbabf1076),
	.w4(32'hba4b2c21),
	.w5(32'hbab0045e),
	.w6(32'hbb9d87aa),
	.w7(32'hbc02e552),
	.w8(32'hbb46787c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f9664),
	.w1(32'hb929ac41),
	.w2(32'hbb47d8da),
	.w3(32'hba6f8d50),
	.w4(32'hbbb050b6),
	.w5(32'h3a5a1eba),
	.w6(32'h3bdbd08b),
	.w7(32'hbbac67ae),
	.w8(32'h3a31ad42),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada6ae8),
	.w1(32'hbba892ac),
	.w2(32'hba6c126c),
	.w3(32'hbab7bdce),
	.w4(32'h39a9d7e6),
	.w5(32'h3b899e88),
	.w6(32'hbb954d07),
	.w7(32'h3ad69e04),
	.w8(32'h3c74a8c0),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c019398),
	.w1(32'h3bdd6669),
	.w2(32'h3b079672),
	.w3(32'h3a645379),
	.w4(32'h3be68090),
	.w5(32'hbc188173),
	.w6(32'h3a609fb2),
	.w7(32'h3b993892),
	.w8(32'hbaec694c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba8c11),
	.w1(32'hbbc61875),
	.w2(32'hbc7a28ec),
	.w3(32'hbb9ec8de),
	.w4(32'h3ba98431),
	.w5(32'hbc09a532),
	.w6(32'h3b133f80),
	.w7(32'h3b86bc61),
	.w8(32'hbc3f2455),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe182b3),
	.w1(32'hba910ce8),
	.w2(32'h3bfdc8e2),
	.w3(32'h3b432cfb),
	.w4(32'h3c4204e3),
	.w5(32'hbadbfcea),
	.w6(32'hbace8e58),
	.w7(32'h3bf2fce6),
	.w8(32'hba99e769),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e4600),
	.w1(32'hbc004ef4),
	.w2(32'hbb59696c),
	.w3(32'hbb45042f),
	.w4(32'h3b81cc1a),
	.w5(32'hb88512e7),
	.w6(32'hbc3ab61a),
	.w7(32'hb9d329d8),
	.w8(32'hbb91b972),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05c492),
	.w1(32'h3b3863db),
	.w2(32'h3a22df02),
	.w3(32'h3ab0c4a3),
	.w4(32'h3b33e93a),
	.w5(32'h3b9eaa3c),
	.w6(32'hba13be62),
	.w7(32'hbaaebe2d),
	.w8(32'h3b4f0aa4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28f88e),
	.w1(32'h3a2fd993),
	.w2(32'hba47a251),
	.w3(32'h3adca4c3),
	.w4(32'h3a7e5c76),
	.w5(32'h3999771d),
	.w6(32'h3add03a4),
	.w7(32'hbb670c67),
	.w8(32'h3aae453a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b398d78),
	.w1(32'hbbd71fd1),
	.w2(32'hbbf47a6f),
	.w3(32'hbbd3977e),
	.w4(32'hbbd57c0b),
	.w5(32'hba32941b),
	.w6(32'hbbf29acd),
	.w7(32'hbc2016c3),
	.w8(32'hbb2e0f23),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba571950),
	.w1(32'hba333cb9),
	.w2(32'hbb4ccc94),
	.w3(32'hbb3069f3),
	.w4(32'h3b1db1b5),
	.w5(32'hbc00c14f),
	.w6(32'hbaceec36),
	.w7(32'h3b0f8e4e),
	.w8(32'hbb8d9548),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28c7d7),
	.w1(32'hbbb6177a),
	.w2(32'h396ce01d),
	.w3(32'h3b1603fd),
	.w4(32'h3ba98629),
	.w5(32'h3bef68dc),
	.w6(32'hbbe32260),
	.w7(32'h3b9a5b9e),
	.w8(32'h3b967ad0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c1463),
	.w1(32'h3c600cf7),
	.w2(32'h3c6f4c9a),
	.w3(32'h3c42e376),
	.w4(32'h3c319c03),
	.w5(32'h3b1715e2),
	.w6(32'h3c765f6b),
	.w7(32'h3c37ee20),
	.w8(32'h3bca2b67),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a7cbc),
	.w1(32'hbb7c2100),
	.w2(32'hbb51033f),
	.w3(32'hbb670b4c),
	.w4(32'hba97d633),
	.w5(32'h3b36329c),
	.w6(32'hb952de34),
	.w7(32'hbbb51a5d),
	.w8(32'hbba698a2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61aa52),
	.w1(32'hbb1cb0de),
	.w2(32'hbb5cce09),
	.w3(32'hbb569053),
	.w4(32'h3b091be6),
	.w5(32'hbb77cfd2),
	.w6(32'hbb9558c8),
	.w7(32'hbab12826),
	.w8(32'hbbd95982),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb290241),
	.w1(32'hbb98eff1),
	.w2(32'hba5513ff),
	.w3(32'hb8802ac7),
	.w4(32'h3b2f62a9),
	.w5(32'h3aa5db8f),
	.w6(32'hbbe6f232),
	.w7(32'h399e48d1),
	.w8(32'hba18f305),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12933e),
	.w1(32'h3b004085),
	.w2(32'h39227648),
	.w3(32'h3ab43e83),
	.w4(32'hbb06b036),
	.w5(32'hbbafd741),
	.w6(32'h3aea479f),
	.w7(32'h3ad1867c),
	.w8(32'hbb231091),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba05cdc),
	.w1(32'hbbb34a00),
	.w2(32'hbbb5e607),
	.w3(32'hbbd18867),
	.w4(32'hbbe63865),
	.w5(32'hb6b98a5e),
	.w6(32'h3b90919f),
	.w7(32'hba22e29d),
	.w8(32'h3ac6e1c9),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0599df),
	.w1(32'h39c151a2),
	.w2(32'h3a930b72),
	.w3(32'hb9f6644a),
	.w4(32'hbbaa8db3),
	.w5(32'hbb97bd6a),
	.w6(32'hba365b63),
	.w7(32'hbb4c2f93),
	.w8(32'h3aceeb8d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e11e10),
	.w1(32'hbaaaab5d),
	.w2(32'h3b96703a),
	.w3(32'h3b2795a7),
	.w4(32'h3b1c6283),
	.w5(32'hbbc2b9b4),
	.w6(32'hbb22d7b4),
	.w7(32'h3be7e3af),
	.w8(32'hbc03adb5),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfddcf0),
	.w1(32'hbbfa62ea),
	.w2(32'hbbc31548),
	.w3(32'hbbd34800),
	.w4(32'hbc0e52b2),
	.w5(32'h3ade5c33),
	.w6(32'h3ad3fd0f),
	.w7(32'hbbd7e705),
	.w8(32'hbb4f6aa4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc92447),
	.w1(32'hbb849185),
	.w2(32'hba068098),
	.w3(32'h3b36bd53),
	.w4(32'h3bae2f66),
	.w5(32'h3b633d60),
	.w6(32'h3a1e0e7b),
	.w7(32'h3b8c7e22),
	.w8(32'h39a0b55b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae339b9),
	.w1(32'hbb88c853),
	.w2(32'h3a81d118),
	.w3(32'hba939e9e),
	.w4(32'h3b26c9bd),
	.w5(32'hbbe2898b),
	.w6(32'hbbb3a1ac),
	.w7(32'hb9e81c68),
	.w8(32'hbb0dc8b8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f4cf4),
	.w1(32'h3ae16be7),
	.w2(32'h3b1748a2),
	.w3(32'h3b6b3642),
	.w4(32'h3bb43f54),
	.w5(32'hb860e4d0),
	.w6(32'h3b615cf8),
	.w7(32'h3b816654),
	.w8(32'h3aac9833),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63ac01),
	.w1(32'hba59180c),
	.w2(32'h3aa87489),
	.w3(32'hbacc5892),
	.w4(32'h3ae0fbfc),
	.w5(32'hbc3b1fba),
	.w6(32'hbbe0ebea),
	.w7(32'h3b2cdba2),
	.w8(32'hbb179e21),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9974ec),
	.w1(32'hba214806),
	.w2(32'hbb074594),
	.w3(32'hbc02b5a9),
	.w4(32'hba86e051),
	.w5(32'hba419122),
	.w6(32'h3b950e36),
	.w7(32'hbab38025),
	.w8(32'hbaed0a0a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2d198),
	.w1(32'h39e6bd96),
	.w2(32'h3ab929d4),
	.w3(32'hba4d37b6),
	.w4(32'hbb168d47),
	.w5(32'h38d8f631),
	.w6(32'h3ad5ddf9),
	.w7(32'hb961a681),
	.w8(32'hba87cb78),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15c454),
	.w1(32'hbbbb7642),
	.w2(32'hbbb7b75e),
	.w3(32'hbb88e61a),
	.w4(32'hbb8cc6e0),
	.w5(32'h3ac266e7),
	.w6(32'hbb83b432),
	.w7(32'hbba727c4),
	.w8(32'h3c09912c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02d722),
	.w1(32'h3c01d43f),
	.w2(32'h3b9410fb),
	.w3(32'h3c217d77),
	.w4(32'h3c16ce4f),
	.w5(32'hbb515763),
	.w6(32'h3c1ebcfd),
	.w7(32'h3c3b4d62),
	.w8(32'hbb041227),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9d57c),
	.w1(32'hbb4ad337),
	.w2(32'hbc026757),
	.w3(32'hbba1cab5),
	.w4(32'hbbc73270),
	.w5(32'hbbb7da35),
	.w6(32'hbbe02358),
	.w7(32'hbc12cd4f),
	.w8(32'hbc04287e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd99559),
	.w1(32'hbb4e597d),
	.w2(32'hbb19b7d6),
	.w3(32'hbb0e2107),
	.w4(32'hba8f2e20),
	.w5(32'h3bd16904),
	.w6(32'hb931eec2),
	.w7(32'hbb48156b),
	.w8(32'h3bd5e2e0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81d8c2),
	.w1(32'hbbc2acab),
	.w2(32'hbbadcab1),
	.w3(32'h3bd2426e),
	.w4(32'h3bb30f11),
	.w5(32'h3aeee00f),
	.w6(32'hbba9e054),
	.w7(32'h3b6a0989),
	.w8(32'hbb17d608),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab9bc9),
	.w1(32'hbb634f9b),
	.w2(32'hbb5c5b21),
	.w3(32'h39f772d4),
	.w4(32'h3a21ef55),
	.w5(32'hba036613),
	.w6(32'h3aaf726e),
	.w7(32'hbad9f238),
	.w8(32'h3acf05dc),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b168e5d),
	.w1(32'h3adc87c5),
	.w2(32'h380159b4),
	.w3(32'hbb42826a),
	.w4(32'h3b222bee),
	.w5(32'h3aabcb9d),
	.w6(32'hbc1c910e),
	.w7(32'hba285bd4),
	.w8(32'h3abab8ae),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a165d),
	.w1(32'h3b91a151),
	.w2(32'hbb56a93d),
	.w3(32'hbbd4d5e7),
	.w4(32'hbabaa4ef),
	.w5(32'hbc054f9a),
	.w6(32'hbb5da22a),
	.w7(32'hbad7b1e2),
	.w8(32'h3ac45bc9),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2bdc4),
	.w1(32'hbb861b58),
	.w2(32'hbc241cbd),
	.w3(32'hbb394bf6),
	.w4(32'hbc0509f8),
	.w5(32'hbba1834d),
	.w6(32'hbbdb0d9d),
	.w7(32'hbbbfbbca),
	.w8(32'hbbf05f7d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a111f),
	.w1(32'hbbedfed7),
	.w2(32'hbc12a740),
	.w3(32'hbb59798c),
	.w4(32'hbb89fafd),
	.w5(32'hbb4be64e),
	.w6(32'hbc607632),
	.w7(32'hbc1b3798),
	.w8(32'hbb1909fd),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd2caa),
	.w1(32'h3b273e11),
	.w2(32'h3a8b25e4),
	.w3(32'hbad57c2d),
	.w4(32'h3b71f03a),
	.w5(32'h3b7dd7a0),
	.w6(32'h3a97f7a0),
	.w7(32'hbae5645e),
	.w8(32'h3b76e997),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e605d),
	.w1(32'h3b731a1f),
	.w2(32'h3b5345f9),
	.w3(32'h3a21c3d1),
	.w4(32'h3bae833d),
	.w5(32'hbb01a267),
	.w6(32'h3b9a3c3b),
	.w7(32'h3b937358),
	.w8(32'hb9c71be0),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03acb3),
	.w1(32'hbb0b45ee),
	.w2(32'hbbf0dc57),
	.w3(32'hbb8284a2),
	.w4(32'hb9b573f7),
	.w5(32'hba9187c0),
	.w6(32'hbbaf7ebf),
	.w7(32'hbb97b117),
	.w8(32'hbba488cf),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd987b5),
	.w1(32'hbb96bc71),
	.w2(32'hbb344622),
	.w3(32'hbbbf5df3),
	.w4(32'h3add171c),
	.w5(32'hbac29106),
	.w6(32'hbaacbb40),
	.w7(32'h3b0c4f29),
	.w8(32'h3a4f0752),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafafc7d),
	.w1(32'h3a104c6c),
	.w2(32'hbaf1c808),
	.w3(32'hbb1e3322),
	.w4(32'hbbd9dab9),
	.w5(32'hbabdf7b8),
	.w6(32'h3bd99ce9),
	.w7(32'hbacbc206),
	.w8(32'hbab3642e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2aa085),
	.w1(32'h39aeef8c),
	.w2(32'hbb91b37e),
	.w3(32'hbba19f6b),
	.w4(32'h3b5d658a),
	.w5(32'h3b8e2bb1),
	.w6(32'h39bc0f0b),
	.w7(32'hbb2b020c),
	.w8(32'h3b40b4ec),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e38d3),
	.w1(32'h3b8f91ad),
	.w2(32'h3b34a657),
	.w3(32'h3bbf953f),
	.w4(32'h3bab99d3),
	.w5(32'hbb97c1e1),
	.w6(32'h3b4e98f0),
	.w7(32'h3b599d39),
	.w8(32'hbb2352fe),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee12e8),
	.w1(32'hbbb5ee97),
	.w2(32'hba823fa4),
	.w3(32'hbb2bea13),
	.w4(32'h3b14195e),
	.w5(32'hbb4df767),
	.w6(32'hbb7b8287),
	.w7(32'h3a949413),
	.w8(32'hbb665e2e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfb381),
	.w1(32'h3ab265ce),
	.w2(32'hbb2ad7ae),
	.w3(32'h3af22fd5),
	.w4(32'h3b689245),
	.w5(32'h3bd1d604),
	.w6(32'h3bbe7f7b),
	.w7(32'h3aff2dde),
	.w8(32'hbaca21de),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989eaf0),
	.w1(32'hba0673c1),
	.w2(32'h3afd8f1f),
	.w3(32'h3b69c15d),
	.w4(32'h3b1c12cb),
	.w5(32'h3afa8ff4),
	.w6(32'hbb7b6ef6),
	.w7(32'hbacd5e69),
	.w8(32'h3995143b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b9d67),
	.w1(32'hbb37361f),
	.w2(32'hbc31957a),
	.w3(32'hbb0c48bf),
	.w4(32'hba8cb7c1),
	.w5(32'hbbe89754),
	.w6(32'hbc0045ae),
	.w7(32'hbb8335d5),
	.w8(32'hbbc92b9c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b1dfe),
	.w1(32'hbb5f1491),
	.w2(32'hbb8b8849),
	.w3(32'hbb4ad1d1),
	.w4(32'hbb2c0e61),
	.w5(32'hbac44f2e),
	.w6(32'hbb3723e9),
	.w7(32'hbb5a0e86),
	.w8(32'hbba12f52),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6fa8e),
	.w1(32'h3a60c651),
	.w2(32'h3a96c332),
	.w3(32'h3a866b00),
	.w4(32'h3abfd55f),
	.w5(32'hbb7722c8),
	.w6(32'hbb53cd2b),
	.w7(32'hbb98a4fb),
	.w8(32'hbb29efd3),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb819ba2),
	.w1(32'hbbb12274),
	.w2(32'hbbe108aa),
	.w3(32'hbba4dbb6),
	.w4(32'hbbaca448),
	.w5(32'hbc0e08aa),
	.w6(32'hbbc3f7b8),
	.w7(32'hbbc23deb),
	.w8(32'hbbbdc45e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29a195),
	.w1(32'hba371b96),
	.w2(32'hba2c2c15),
	.w3(32'hbaeb022a),
	.w4(32'h3ae3a815),
	.w5(32'hb948cfff),
	.w6(32'hb989b40a),
	.w7(32'h3a2bac01),
	.w8(32'h3a5e4ade),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c37013),
	.w1(32'hbb5ddd1b),
	.w2(32'hba80efe4),
	.w3(32'hbb5fde99),
	.w4(32'hb9840cd1),
	.w5(32'h3ba54b26),
	.w6(32'hbb338e20),
	.w7(32'hb9646434),
	.w8(32'h3afa796a),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15b693),
	.w1(32'h3a8f9c38),
	.w2(32'h3a96deb5),
	.w3(32'h3b97757a),
	.w4(32'h3ba4bd23),
	.w5(32'h3bc6797d),
	.w6(32'hb8817b4e),
	.w7(32'h3b1e7657),
	.w8(32'h36864632),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37fcea),
	.w1(32'h39b02518),
	.w2(32'h3b7dac74),
	.w3(32'h3b7ea120),
	.w4(32'h3b6a53aa),
	.w5(32'hbb6926fa),
	.w6(32'hbb50be84),
	.w7(32'hba8df2f5),
	.w8(32'hbab2689a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb845a6c4),
	.w1(32'hb8b00339),
	.w2(32'hbaed5f94),
	.w3(32'hbb3b7f9e),
	.w4(32'hba9392fe),
	.w5(32'h3b32f5fa),
	.w6(32'hbb022fa7),
	.w7(32'hbb27c4e7),
	.w8(32'h3adf514d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ba46c),
	.w1(32'h3a90d5ce),
	.w2(32'h3b5ba0fb),
	.w3(32'h3a24be6b),
	.w4(32'h3bbcc6a6),
	.w5(32'h3b91d006),
	.w6(32'h3a84c392),
	.w7(32'h3b90bb26),
	.w8(32'h3acdbc0b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8302ec),
	.w1(32'hb8fbb450),
	.w2(32'hb82dc91e),
	.w3(32'h3b2de3de),
	.w4(32'h3b48be12),
	.w5(32'hbb1707f4),
	.w6(32'h39e898ec),
	.w7(32'h3adfb89f),
	.w8(32'hbabe89b0),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bf842),
	.w1(32'hbb347010),
	.w2(32'hbb84b1ff),
	.w3(32'hbb1f1f07),
	.w4(32'hbb1a0035),
	.w5(32'hbadd5bbb),
	.w6(32'hbb21d7aa),
	.w7(32'hbb068ea3),
	.w8(32'hba89619a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacff207),
	.w1(32'h390f7856),
	.w2(32'h3b738853),
	.w3(32'hbb0904f9),
	.w4(32'hb8575a17),
	.w5(32'h3a9ace4b),
	.w6(32'hbb00e37c),
	.w7(32'h3b78e75d),
	.w8(32'hb70f96e6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4aa1e),
	.w1(32'hba8481be),
	.w2(32'h3b0948ac),
	.w3(32'hba8d4560),
	.w4(32'h3b501436),
	.w5(32'hba5361c5),
	.w6(32'hbadc8846),
	.w7(32'h3ac6f4de),
	.w8(32'hb9baa5f3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393252a4),
	.w1(32'h3b2421ad),
	.w2(32'h3a0dd85a),
	.w3(32'hbacd3517),
	.w4(32'hbae661e0),
	.w5(32'hbadb1813),
	.w6(32'h3a9812c0),
	.w7(32'h3a1cabb2),
	.w8(32'hbb33fc23),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed7d83),
	.w1(32'hbada123a),
	.w2(32'h3a861efc),
	.w3(32'hb5b2caf6),
	.w4(32'hb9ffaf84),
	.w5(32'h3bd0a0c5),
	.w6(32'hbab5ba72),
	.w7(32'hba5fb288),
	.w8(32'h3ab669a1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b830e67),
	.w1(32'h3b06996b),
	.w2(32'h3b8d4b6c),
	.w3(32'h3bfffc5d),
	.w4(32'h3bc066d7),
	.w5(32'h3b476f60),
	.w6(32'h39fe372c),
	.w7(32'h3ae8ca15),
	.w8(32'h3b0b497e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59b00c),
	.w1(32'h3bc3864d),
	.w2(32'h3b7c44ce),
	.w3(32'h3bcd49f7),
	.w4(32'h3bd01266),
	.w5(32'h3b3c9fbf),
	.w6(32'h3baa2c51),
	.w7(32'h3b9bea4c),
	.w8(32'h3b004930),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac060c),
	.w1(32'h3b803983),
	.w2(32'h3b814d3d),
	.w3(32'h3b8f6e39),
	.w4(32'h3b8ffc2c),
	.w5(32'h38ae30ef),
	.w6(32'h3bab09ff),
	.w7(32'h3bc1ef3c),
	.w8(32'hba8274d7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01e354),
	.w1(32'hbb5d2af3),
	.w2(32'hbb4edf93),
	.w3(32'hba70b645),
	.w4(32'hbaaa6857),
	.w5(32'hba8b81c0),
	.w6(32'hba8f5486),
	.w7(32'hbb3915e2),
	.w8(32'hbaa669ad),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ca22f),
	.w1(32'hbb6a2063),
	.w2(32'hbab1ffff),
	.w3(32'hbaf32c46),
	.w4(32'hbb5af9e0),
	.w5(32'h3a86fffd),
	.w6(32'hbb7d4f72),
	.w7(32'hbb0f0a9b),
	.w8(32'h3a358f0a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b5008),
	.w1(32'hba974071),
	.w2(32'hba831a50),
	.w3(32'hb7b5fcea),
	.w4(32'h38693a8b),
	.w5(32'h3832a7c2),
	.w6(32'h3a31c2d1),
	.w7(32'hb9b29615),
	.w8(32'hbb477ee1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01024b),
	.w1(32'hbb2808fc),
	.w2(32'hbae4b83f),
	.w3(32'hba6b2bda),
	.w4(32'hbb5932a7),
	.w5(32'h3b7a9d4c),
	.w6(32'hbb6014c8),
	.w7(32'hbb4c8a94),
	.w8(32'h3a79f6a5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95cf3e1),
	.w1(32'hbbc65db7),
	.w2(32'hbbe75095),
	.w3(32'h3a8677c9),
	.w4(32'hbb27afe8),
	.w5(32'hbb52bd53),
	.w6(32'hbb184073),
	.w7(32'hbbc5a7bb),
	.w8(32'hbb796a25),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3323a6),
	.w1(32'h3a9612b6),
	.w2(32'h39ead9ab),
	.w3(32'h3a9608ed),
	.w4(32'hb907d906),
	.w5(32'hb9421ec5),
	.w6(32'hba2611d2),
	.w7(32'hb9a42f6c),
	.w8(32'h375dcc5c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb597141),
	.w1(32'hbb374230),
	.w2(32'h3b271db2),
	.w3(32'hbb9be7b7),
	.w4(32'hba4833e7),
	.w5(32'h3bbb5af7),
	.w6(32'hbb46ecef),
	.w7(32'hb9b8645c),
	.w8(32'h3ae73990),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule