module layer_10_featuremap_110(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61f631b),
	.w1(32'hb5d02575),
	.w2(32'hb5fce73d),
	.w3(32'hb64ba547),
	.w4(32'hb5ca28ed),
	.w5(32'hb65f9a7b),
	.w6(32'hb6711330),
	.w7(32'hb64721ac),
	.w8(32'hb6462b33),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb907cee1),
	.w1(32'hb8000b0d),
	.w2(32'hb8ef57b0),
	.w3(32'hb92f3eb3),
	.w4(32'hb8851732),
	.w5(32'hb8c2b51d),
	.w6(32'hb8cdb9c1),
	.w7(32'h384679a3),
	.w8(32'hb7a1623c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3353fa66),
	.w1(32'hb4c9adc7),
	.w2(32'hb52ed785),
	.w3(32'hb2f1ffee),
	.w4(32'h33a0b108),
	.w5(32'hb50d7c20),
	.w6(32'hb49a8e75),
	.w7(32'hb4feb5b7),
	.w8(32'hb55302d9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3866dac7),
	.w1(32'hb86619df),
	.w2(32'hb83b827a),
	.w3(32'h389c1ccd),
	.w4(32'hb683784d),
	.w5(32'hb81db42b),
	.w6(32'h3867c87d),
	.w7(32'h382fe851),
	.w8(32'hb81ebeda),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fd3c2e),
	.w1(32'hb8383f64),
	.w2(32'hb79dfa4a),
	.w3(32'hb828df2c),
	.w4(32'hb849f7cb),
	.w5(32'hb808ae26),
	.w6(32'hb81592f1),
	.w7(32'hb811cdcb),
	.w8(32'hb800312e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36831c9d),
	.w1(32'h35ed1f75),
	.w2(32'h353a9421),
	.w3(32'hb48c7f7d),
	.w4(32'hb6c73be8),
	.w5(32'hb701dee1),
	.w6(32'h3581cd4c),
	.w7(32'hb5995105),
	.w8(32'hb6a8a63e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb835159d),
	.w1(32'hb858e7e9),
	.w2(32'h389f38c8),
	.w3(32'hb8941ebc),
	.w4(32'hb58b2035),
	.w5(32'h38c70331),
	.w6(32'hb8112314),
	.w7(32'h380d70cf),
	.w8(32'h38f45826),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb875a9f4),
	.w1(32'hb8725c00),
	.w2(32'h393b8498),
	.w3(32'hb7d6ee1d),
	.w4(32'h39069b64),
	.w5(32'h3938db02),
	.w6(32'h38e2e844),
	.w7(32'hb7f28194),
	.w8(32'h395831f1),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a3198),
	.w1(32'hb8f0cd9b),
	.w2(32'hb88a05e9),
	.w3(32'hb90b8cc0),
	.w4(32'hb85d52f7),
	.w5(32'h38083afe),
	.w6(32'hb9074d54),
	.w7(32'hb85ee7f5),
	.w8(32'h38afb536),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38df0366),
	.w1(32'h38a1d90a),
	.w2(32'h39b53d6c),
	.w3(32'h3923a15c),
	.w4(32'h36fae79f),
	.w5(32'h3998a094),
	.w6(32'h35d8d0f9),
	.w7(32'hb90a861d),
	.w8(32'h3960fb8e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3773dc56),
	.w1(32'h378e9835),
	.w2(32'h38d1c1db),
	.w3(32'hb7846638),
	.w4(32'h37a228a5),
	.w5(32'h38b229b5),
	.w6(32'h37a4b7b9),
	.w7(32'h387281ff),
	.w8(32'h38b352a2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b89cd5),
	.w1(32'hb9b964a4),
	.w2(32'hb8c5778b),
	.w3(32'hb82403b2),
	.w4(32'hb94481f1),
	.w5(32'hb802c046),
	.w6(32'h3873ece1),
	.w7(32'hb858766f),
	.w8(32'h35a713e9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3956e9b8),
	.w1(32'hb8d680f4),
	.w2(32'h39a23987),
	.w3(32'h3931367c),
	.w4(32'h3725e576),
	.w5(32'h399e93da),
	.w6(32'hb8ac0cd4),
	.w7(32'hb94a4dc6),
	.w8(32'h385bcf40),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb827fe30),
	.w1(32'hb93eaa0a),
	.w2(32'h389776cc),
	.w3(32'h38618b06),
	.w4(32'hb682c9ee),
	.w5(32'h38cd6375),
	.w6(32'hb8e83286),
	.w7(32'hb7c4b8c5),
	.w8(32'h38af3c48),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bf0cf0),
	.w1(32'hb8bcff54),
	.w2(32'hb89a529b),
	.w3(32'hb815ae1b),
	.w4(32'hb80ff9d5),
	.w5(32'hb8ab750b),
	.w6(32'hb89b1539),
	.w7(32'hb906162a),
	.w8(32'hb8611fef),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b50c5c),
	.w1(32'hb92ca734),
	.w2(32'h380def0c),
	.w3(32'h375e8993),
	.w4(32'hb8725bcf),
	.w5(32'h388e958d),
	.w6(32'hb84c2806),
	.w7(32'hb86c0367),
	.w8(32'h3910395b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dc317f),
	.w1(32'hb6c6d8b3),
	.w2(32'h348931d5),
	.w3(32'h36d8d488),
	.w4(32'h37c9174d),
	.w5(32'h37f9eae4),
	.w6(32'h35a2a8a1),
	.w7(32'h37b647e1),
	.w8(32'h37ce30b1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f84e2),
	.w1(32'hb93db5a1),
	.w2(32'h39d8a50f),
	.w3(32'h397495b7),
	.w4(32'h3861b930),
	.w5(32'h39ee83fc),
	.w6(32'h3940dd73),
	.w7(32'hb8ea4e1c),
	.w8(32'h39ffd229),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98720d4),
	.w1(32'hb8b59104),
	.w2(32'h38d689a0),
	.w3(32'h38963020),
	.w4(32'h3712a4b3),
	.w5(32'h3922c548),
	.w6(32'h388696b8),
	.w7(32'hb870f7a0),
	.w8(32'h38ebda8b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62fcac2),
	.w1(32'hb5fce158),
	.w2(32'hb588bb48),
	.w3(32'hb62a7d9a),
	.w4(32'hb5a66779),
	.w5(32'hb5056b0e),
	.w6(32'hb663d4fc),
	.w7(32'h355fae9a),
	.w8(32'h33bbbb34),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a7e2db),
	.w1(32'h36459ed2),
	.w2(32'h36896377),
	.w3(32'hb50c5e6f),
	.w4(32'h35979622),
	.w5(32'h366558e6),
	.w6(32'hb69274d2),
	.w7(32'hb65444ac),
	.w8(32'hb60dce7a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e14b7),
	.w1(32'hb868e9a5),
	.w2(32'hb8e292bc),
	.w3(32'hb9130cfc),
	.w4(32'hb8ae21bf),
	.w5(32'hb90f558f),
	.w6(32'hb893620f),
	.w7(32'hb789600d),
	.w8(32'hb8dda2dc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972ab53),
	.w1(32'hba3c6871),
	.w2(32'hb8810baf),
	.w3(32'h380fc821),
	.w4(32'hb9d74900),
	.w5(32'h391f4280),
	.w6(32'h3a1bbd27),
	.w7(32'h39662c71),
	.w8(32'h39a61578),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392fd95d),
	.w1(32'h362d9493),
	.w2(32'h385f62e3),
	.w3(32'h38a90fb5),
	.w4(32'hb7d99d58),
	.w5(32'h38e83e8e),
	.w6(32'hb6aab306),
	.w7(32'hb948466d),
	.w8(32'h38234e59),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dbf368),
	.w1(32'hb8c4106c),
	.w2(32'hb95dfb02),
	.w3(32'hb8ddd768),
	.w4(32'hb92c1383),
	.w5(32'hb9572b94),
	.w6(32'hb8f2b0e2),
	.w7(32'hb9055c1e),
	.w8(32'hb90b3a75),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb789d7cc),
	.w1(32'hb8c696f5),
	.w2(32'h3716216a),
	.w3(32'h38b77c6a),
	.w4(32'h35f26973),
	.w5(32'h38a9bf67),
	.w6(32'h383eda91),
	.w7(32'hb7157e6c),
	.w8(32'h37fb1cd6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3541562d),
	.w1(32'h3668abec),
	.w2(32'hb695cbeb),
	.w3(32'hb6ad1102),
	.w4(32'hb6efb19d),
	.w5(32'hb76763b7),
	.w6(32'hb685a9fb),
	.w7(32'hb6707672),
	.w8(32'hb739354c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cbeda3),
	.w1(32'hb7ddca24),
	.w2(32'hb8f2e56f),
	.w3(32'hb85de19d),
	.w4(32'hb714b758),
	.w5(32'hb82ddd97),
	.w6(32'hb7e5629a),
	.w7(32'hb6afa23f),
	.w8(32'hb832e528),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d16af2),
	.w1(32'h37ae1fea),
	.w2(32'hb8c87d50),
	.w3(32'hb7d8eb97),
	.w4(32'h3881c300),
	.w5(32'hb7dc8319),
	.w6(32'h3847015a),
	.w7(32'h38325463),
	.w8(32'hb81921c7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38adc4d4),
	.w1(32'hb88b6994),
	.w2(32'h38ca2683),
	.w3(32'h38d92ca2),
	.w4(32'hb5aa2c2a),
	.w5(32'h3976fd06),
	.w6(32'h372b7893),
	.w7(32'hb896702a),
	.w8(32'h395935d4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a92d9b),
	.w1(32'h35daa791),
	.w2(32'h361c8f57),
	.w3(32'h36a84713),
	.w4(32'h36a7a8db),
	.w5(32'h369c0212),
	.w6(32'h36646fae),
	.w7(32'h368c7502),
	.w8(32'h36811389),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76d8609),
	.w1(32'h367c9d56),
	.w2(32'h369dd985),
	.w3(32'hb6239804),
	.w4(32'h37462590),
	.w5(32'h37451b14),
	.w6(32'h32cb8dd6),
	.w7(32'h3707b985),
	.w8(32'h372205f9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b86cb5),
	.w1(32'hb85946bb),
	.w2(32'h38d2ecac),
	.w3(32'h37ec3506),
	.w4(32'hb8ae9c31),
	.w5(32'h38215666),
	.w6(32'hb83b2717),
	.w7(32'hb906e841),
	.w8(32'h379c9958),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37acf438),
	.w1(32'hb780b140),
	.w2(32'hb8627c32),
	.w3(32'h378f56d1),
	.w4(32'h373fd4a2),
	.w5(32'h37976a4a),
	.w6(32'h380a4172),
	.w7(32'h3858578a),
	.w8(32'h37d866de),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36de3b3d),
	.w1(32'h37e34140),
	.w2(32'h373704a1),
	.w3(32'h370154f0),
	.w4(32'h37d04e2e),
	.w5(32'h37f76b83),
	.w6(32'h37bdeec3),
	.w7(32'h382e80bd),
	.w8(32'h37c84dee),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f09b71),
	.w1(32'hb89dde34),
	.w2(32'h38818c09),
	.w3(32'hb6e8e5d2),
	.w4(32'h3863b65a),
	.w5(32'h390d75c3),
	.w6(32'hb745924e),
	.w7(32'hb7c70962),
	.w8(32'h388a7245),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952a514),
	.w1(32'hba0c51a2),
	.w2(32'h386b433d),
	.w3(32'h38abf09b),
	.w4(32'hb9b229c4),
	.w5(32'h392fe33d),
	.w6(32'h396a498f),
	.w7(32'hb81cef27),
	.w8(32'h38a89068),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b2ab1),
	.w1(32'hb8bbb342),
	.w2(32'hba25720a),
	.w3(32'h391eecf7),
	.w4(32'hb8bcbc82),
	.w5(32'hba0be71c),
	.w6(32'h39cd727b),
	.w7(32'h391f04a4),
	.w8(32'hb9bbc992),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9817473),
	.w1(32'hb94cdc1e),
	.w2(32'hba1c70b8),
	.w3(32'hb93f84d5),
	.w4(32'hb926e4ca),
	.w5(32'hb9e6bf72),
	.w6(32'h37197605),
	.w7(32'h3940838a),
	.w8(32'hb8fc5998),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3814d2a2),
	.w1(32'hb8b8c9ba),
	.w2(32'hb9027d75),
	.w3(32'h37dbd82d),
	.w4(32'hb90b40de),
	.w5(32'hb92c1b52),
	.w6(32'h3887a5e8),
	.w7(32'hb82d0da0),
	.w8(32'hb88fa4bf),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7879816),
	.w1(32'hb7bd8dc9),
	.w2(32'hb7664166),
	.w3(32'hb6693053),
	.w4(32'hb75dfdeb),
	.w5(32'h36844bb9),
	.w6(32'hb6a039b0),
	.w7(32'h36f49b53),
	.w8(32'h3801fca2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7264817),
	.w1(32'hb72f83e3),
	.w2(32'hb81d93e3),
	.w3(32'h356a8d45),
	.w4(32'hb58f186d),
	.w5(32'hb7db4327),
	.w6(32'hb5a8da9c),
	.w7(32'hb65a1741),
	.w8(32'hb7373ad1),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bf614b),
	.w1(32'hb8efecbe),
	.w2(32'hb98ebc3e),
	.w3(32'hb72c77d3),
	.w4(32'hb7d9d8ce),
	.w5(32'hb90ae0f0),
	.w6(32'h389836d2),
	.w7(32'hb86874bd),
	.w8(32'hb9172770),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb829bd3f),
	.w1(32'h38466019),
	.w2(32'h39aa51ce),
	.w3(32'h38e5d867),
	.w4(32'h379721f1),
	.w5(32'h39b0300f),
	.w6(32'hb89ddecc),
	.w7(32'hb8a1abbd),
	.w8(32'h39a93b90),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ef0ddd),
	.w1(32'h37f577b5),
	.w2(32'h38ef6576),
	.w3(32'h3908bb8e),
	.w4(32'hb5014f96),
	.w5(32'h391e9614),
	.w6(32'h3828cd2d),
	.w7(32'hb87f68de),
	.w8(32'h390a020b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a91680),
	.w1(32'hb8f3c05d),
	.w2(32'h3745a5d6),
	.w3(32'h3885eb2a),
	.w4(32'hb8beef1b),
	.w5(32'h382f6629),
	.w6(32'h37ce8b93),
	.w7(32'hb901d01c),
	.w8(32'h387a00a8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9147d66),
	.w1(32'hb9570dd0),
	.w2(32'hb8ede64c),
	.w3(32'hb77517e6),
	.w4(32'hb8001a2a),
	.w5(32'h38809eb9),
	.w6(32'h38fb5c5a),
	.w7(32'h389e7219),
	.w8(32'h3935c6d1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afff7c),
	.w1(32'hba0bb68a),
	.w2(32'h39b77bec),
	.w3(32'h39c184c8),
	.w4(32'hb7882dbe),
	.w5(32'h3a117992),
	.w6(32'h39f48168),
	.w7(32'hb882e84c),
	.w8(32'h39663e73),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83ba65e),
	.w1(32'hb816bfc4),
	.w2(32'hb83244ab),
	.w3(32'hb7d5f4c7),
	.w4(32'hb5ba62c2),
	.w5(32'hb664ef64),
	.w6(32'hb71d3dc8),
	.w7(32'h37a4608c),
	.w8(32'h382797df),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a8cc79),
	.w1(32'hb90770d2),
	.w2(32'hb912e6b5),
	.w3(32'h35aebe25),
	.w4(32'h3878a0e0),
	.w5(32'h380a7635),
	.w6(32'h3897cc07),
	.w7(32'h39353a22),
	.w8(32'h3917dc04),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb805bbb7),
	.w1(32'hb7dcd7bb),
	.w2(32'hb7ef4fcf),
	.w3(32'hb78a4ff7),
	.w4(32'h35d6808c),
	.w5(32'hb7650afc),
	.w6(32'hb6d80b6a),
	.w7(32'h37c351b0),
	.w8(32'hb79c4f0a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3916c53c),
	.w1(32'hb7b7ddc1),
	.w2(32'h38600637),
	.w3(32'h392049f3),
	.w4(32'hb85ef608),
	.w5(32'hb84b8a7d),
	.w6(32'h37cb44e9),
	.w7(32'hb894c724),
	.w8(32'hb78f6d5c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78d67a5),
	.w1(32'hb712aeea),
	.w2(32'h38197e9f),
	.w3(32'h3609f9e5),
	.w4(32'h37317754),
	.w5(32'h380f1855),
	.w6(32'h37b7b8e3),
	.w7(32'h38070851),
	.w8(32'h3864d0de),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b8caec),
	.w1(32'hb958d741),
	.w2(32'h3990d95c),
	.w3(32'h392f3d72),
	.w4(32'hb94e4df1),
	.w5(32'h378483a4),
	.w6(32'h3966cf6c),
	.w7(32'hb92c1c65),
	.w8(32'h3922740d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bfbdf2),
	.w1(32'hb7a48264),
	.w2(32'hb80c69f6),
	.w3(32'h379add95),
	.w4(32'hb74196f2),
	.w5(32'hb7e7dc66),
	.w6(32'h386b281f),
	.w7(32'h37aed596),
	.w8(32'h3603f571),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f234fa),
	.w1(32'hb792b0db),
	.w2(32'h378dec11),
	.w3(32'h36dd6061),
	.w4(32'hb708a604),
	.w5(32'h37b4c82b),
	.w6(32'h36406b4a),
	.w7(32'hb74113a3),
	.w8(32'h37456e58),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb625ddbb),
	.w1(32'h3640c2d9),
	.w2(32'hb31bf82e),
	.w3(32'hb690a1fb),
	.w4(32'h34a48bb1),
	.w5(32'hb5221a29),
	.w6(32'hb6ae5b90),
	.w7(32'hb5cdb30f),
	.w8(32'hb5671cf3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36abfdc5),
	.w1(32'h3767fd55),
	.w2(32'hb6a08736),
	.w3(32'h36118560),
	.w4(32'h370aac16),
	.w5(32'h36123bd8),
	.w6(32'h3638adb8),
	.w7(32'hb73b2fc8),
	.w8(32'hb637af1e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8311dc0),
	.w1(32'hb81a9b4d),
	.w2(32'hb8e3f902),
	.w3(32'hb8353d28),
	.w4(32'hb7d6d0a8),
	.w5(32'hb89bb5f8),
	.w6(32'hb6b6e8af),
	.w7(32'hb750be76),
	.w8(32'hb888b799),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ddeac4),
	.w1(32'h37c41cc5),
	.w2(32'hb7bf69b7),
	.w3(32'h381af219),
	.w4(32'h380677d9),
	.w5(32'hb7c6601c),
	.w6(32'h3654d0d0),
	.w7(32'h37260d6c),
	.w8(32'hb7adba6e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb803b5fe),
	.w1(32'h3839b720),
	.w2(32'h38d58427),
	.w3(32'hb6d77fe2),
	.w4(32'h38361072),
	.w5(32'h394a9f23),
	.w6(32'hb8327111),
	.w7(32'h37025d1d),
	.w8(32'h386e12c2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b4d77),
	.w1(32'h38988ddb),
	.w2(32'h38042fcf),
	.w3(32'h392b077a),
	.w4(32'h38cc5232),
	.w5(32'h38a51b4b),
	.w6(32'h39443894),
	.w7(32'h39341105),
	.w8(32'h38c9ba3e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a421f7),
	.w1(32'hb6c8db41),
	.w2(32'hb69b4069),
	.w3(32'hb5a49cd8),
	.w4(32'h36e1be60),
	.w5(32'h3741e3a8),
	.w6(32'h37029361),
	.w7(32'h379890ce),
	.w8(32'h37bf11ae),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h352c2509),
	.w1(32'h365f2040),
	.w2(32'h369aa536),
	.w3(32'h35cedbd3),
	.w4(32'h369604d8),
	.w5(32'h368c4bf1),
	.w6(32'h336db0a2),
	.w7(32'h360d4786),
	.w8(32'h35e6bd07),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70f1f54),
	.w1(32'h36d84271),
	.w2(32'h35ef415d),
	.w3(32'hb52a3eb8),
	.w4(32'h36da4d02),
	.w5(32'h36b13966),
	.w6(32'hb4a0b22b),
	.w7(32'h367f8018),
	.w8(32'h36a25ad9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b10415),
	.w1(32'h364b732a),
	.w2(32'hb589cc22),
	.w3(32'hb62f0806),
	.w4(32'hb65841ce),
	.w5(32'hb6b9ef77),
	.w6(32'hb6be7b9d),
	.w7(32'hb664ac7e),
	.w8(32'hb6dfbf52),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d5666),
	.w1(32'h3732bad3),
	.w2(32'hb8196361),
	.w3(32'hb78a8c2e),
	.w4(32'hb898dfa4),
	.w5(32'hb8c3485a),
	.w6(32'h38b44c01),
	.w7(32'h3948deb0),
	.w8(32'h38181847),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb850f1d0),
	.w1(32'hb7df8e00),
	.w2(32'hb7b261b2),
	.w3(32'hb939e969),
	.w4(32'hb8d042ee),
	.w5(32'hb890419a),
	.w6(32'hb8818ea3),
	.w7(32'hb7cd4a48),
	.w8(32'h37a6a7b9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81d8648),
	.w1(32'hb8b100e8),
	.w2(32'hb920328e),
	.w3(32'hb9284de5),
	.w4(32'hb830f50b),
	.w5(32'hb89130c3),
	.w6(32'h38a721aa),
	.w7(32'h38f4cb81),
	.w8(32'hb6997606),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7aac907),
	.w1(32'hb97217bd),
	.w2(32'hb904998f),
	.w3(32'hb992d82f),
	.w4(32'hb9583c7a),
	.w5(32'hb88fd452),
	.w6(32'hb951e52a),
	.w7(32'hb965ae56),
	.w8(32'hb87ef839),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35bb8d53),
	.w1(32'h3507fa2d),
	.w2(32'hb59bf738),
	.w3(32'h36757369),
	.w4(32'h3657edd3),
	.w5(32'hb4a60708),
	.w6(32'hb4ff6d29),
	.w7(32'h35bbf480),
	.w8(32'hb5937883),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb583c801),
	.w1(32'h353ead13),
	.w2(32'h35b83d8d),
	.w3(32'hb6073de6),
	.w4(32'h358c6cca),
	.w5(32'h35efc477),
	.w6(32'hb6bd18ef),
	.w7(32'hb5d1b859),
	.w8(32'hb5a7e79e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362e43f8),
	.w1(32'h36e63eb1),
	.w2(32'h372f7ed0),
	.w3(32'h35405ef9),
	.w4(32'h3678cfd7),
	.w5(32'h36e6362e),
	.w6(32'hb6b004ad),
	.w7(32'hb6c78e4d),
	.w8(32'h3549ad2d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7aa2ce5),
	.w1(32'h3815a553),
	.w2(32'h3818d7e6),
	.w3(32'h37586e4c),
	.w4(32'h35414468),
	.w5(32'hb72a89b8),
	.w6(32'h369db666),
	.w7(32'h3832c4c8),
	.w8(32'h3860ae99),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3531ccbe),
	.w1(32'hb6c08f83),
	.w2(32'hb7833211),
	.w3(32'h37354413),
	.w4(32'h371af6f4),
	.w5(32'h361448f5),
	.w6(32'h3708d502),
	.w7(32'h37686842),
	.w8(32'h37b3238e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c87b23),
	.w1(32'hb8e72de8),
	.w2(32'h393a0db0),
	.w3(32'h38b9782c),
	.w4(32'hb7df0d73),
	.w5(32'h38bb5721),
	.w6(32'h390b674e),
	.w7(32'h38e282bb),
	.w8(32'h3940637b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d7509),
	.w1(32'hb90b1e6b),
	.w2(32'h3980034a),
	.w3(32'hb7ca8983),
	.w4(32'h39491e82),
	.w5(32'h39e13d99),
	.w6(32'hb8e58cec),
	.w7(32'hb85662b6),
	.w8(32'h39b45cd5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900e9d4),
	.w1(32'hb8ba2aa8),
	.w2(32'h37b0a9df),
	.w3(32'h38bde653),
	.w4(32'hb8fd9a2e),
	.w5(32'hb72b8446),
	.w6(32'hb838d7dd),
	.w7(32'hb937d958),
	.w8(32'hb8c9edeb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cefbc9),
	.w1(32'h3908dde7),
	.w2(32'h391eb3e8),
	.w3(32'h378415d9),
	.w4(32'hb8580e66),
	.w5(32'hb6fb1f43),
	.w6(32'hb8b088c7),
	.w7(32'hb85a4530),
	.w8(32'h37e90b73),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb780f759),
	.w1(32'hb866aa7f),
	.w2(32'h37c0b31e),
	.w3(32'h378863c0),
	.w4(32'hb8343cd4),
	.w5(32'hb8101c5c),
	.w6(32'h38136720),
	.w7(32'h389b2c6f),
	.w8(32'h38d73632),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389bf33f),
	.w1(32'h3851015b),
	.w2(32'h38cb6827),
	.w3(32'h38e79977),
	.w4(32'h381c7057),
	.w5(32'h38f443eb),
	.w6(32'h384564d1),
	.w7(32'h37925951),
	.w8(32'h38c6b7c6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89085d7),
	.w1(32'hb8bfda25),
	.w2(32'h393c5619),
	.w3(32'h382eea2f),
	.w4(32'hb89ba692),
	.w5(32'h39292a1a),
	.w6(32'h381de5e9),
	.w7(32'hb77e78e7),
	.w8(32'h391d430c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35145904),
	.w1(32'hb412140a),
	.w2(32'hb5b50d30),
	.w3(32'hb55cf25d),
	.w4(32'hb5c1e456),
	.w5(32'hb618f71e),
	.w6(32'hb5b107e5),
	.w7(32'hb5f53f97),
	.w8(32'hb61ec977),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6935acc),
	.w1(32'hb684fc31),
	.w2(32'hb6be3151),
	.w3(32'hb649c8b7),
	.w4(32'hb57c642a),
	.w5(32'hb5d3d38c),
	.w6(32'hb53c96da),
	.w7(32'hb4b578d2),
	.w8(32'hb61428f9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360bd8fd),
	.w1(32'h3654af7f),
	.w2(32'hb60391d5),
	.w3(32'hb6933327),
	.w4(32'h360807ee),
	.w5(32'hb5fa7c00),
	.w6(32'hb6f44299),
	.w7(32'hb66c10eb),
	.w8(32'hb7040f1c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ec4714),
	.w1(32'hb4f65ca4),
	.w2(32'hb41eca30),
	.w3(32'h35db4417),
	.w4(32'hb62f45fc),
	.w5(32'hb4db4efb),
	.w6(32'h363ed1e5),
	.w7(32'hb6cc2ae9),
	.w8(32'hb6244cff),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385e72a7),
	.w1(32'h3776f1d2),
	.w2(32'hb99b1373),
	.w3(32'hb7d14ed2),
	.w4(32'hb9426f01),
	.w5(32'hb9870b6f),
	.w6(32'h3961d91e),
	.w7(32'h388e0c7b),
	.w8(32'hb8e8d520),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7940ffe),
	.w1(32'hb84b26d0),
	.w2(32'hb900bdbb),
	.w3(32'h3740f63d),
	.w4(32'hb57d82c3),
	.w5(32'hb8b17c0e),
	.w6(32'hb7a20341),
	.w7(32'hb81a7873),
	.w8(32'hb8c41b85),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382f44c7),
	.w1(32'hb8248e02),
	.w2(32'hb70e52dc),
	.w3(32'h350b9301),
	.w4(32'hb92a34ef),
	.w5(32'hb8900f0d),
	.w6(32'h37c5ed61),
	.w7(32'hb8b914d0),
	.w8(32'h3880b39a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900f838),
	.w1(32'h391bd7e6),
	.w2(32'h39aa3930),
	.w3(32'h3998a45d),
	.w4(32'h399eeb02),
	.w5(32'h39971803),
	.w6(32'h39fe67d1),
	.w7(32'h39bacb08),
	.w8(32'h3994c578),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb778810f),
	.w1(32'hb96bd17a),
	.w2(32'hb99c49df),
	.w3(32'h383a4b8b),
	.w4(32'hb89b467e),
	.w5(32'hb9726cd8),
	.w6(32'h390cca28),
	.w7(32'h391c37d8),
	.w8(32'hb8b21944),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397979ff),
	.w1(32'hb91322b0),
	.w2(32'h38a9b887),
	.w3(32'hb7575d06),
	.w4(32'hb92c556f),
	.w5(32'h3775ed7f),
	.w6(32'h38035ce6),
	.w7(32'h397b271a),
	.w8(32'h374bfb33),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903b878),
	.w1(32'hb7d60f7d),
	.w2(32'hb906f412),
	.w3(32'h38a3d242),
	.w4(32'hb8543327),
	.w5(32'hb83627d6),
	.w6(32'hb8835df3),
	.w7(32'hb9275ff5),
	.w8(32'hb90a5c7b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387bc5e1),
	.w1(32'hb87155d6),
	.w2(32'hb86bc45d),
	.w3(32'hb871c56c),
	.w4(32'hb9ac794d),
	.w5(32'hb9a6513a),
	.w6(32'hb902394b),
	.w7(32'hb8e2d58e),
	.w8(32'h37b56d35),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8288b40),
	.w1(32'hb8dee0e7),
	.w2(32'hb915f2d1),
	.w3(32'hb8315103),
	.w4(32'hb94b7e56),
	.w5(32'hb9110d49),
	.w6(32'hb7330c7f),
	.w7(32'h37b8ef5b),
	.w8(32'h3807a08b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f30af),
	.w1(32'hb898873b),
	.w2(32'hb92f0000),
	.w3(32'h38af9360),
	.w4(32'hb949060b),
	.w5(32'hb9a897fe),
	.w6(32'h390d7011),
	.w7(32'hb8575211),
	.w8(32'hb7f544b8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb710e3f5),
	.w1(32'hb80fd74f),
	.w2(32'hb88dbd04),
	.w3(32'hb6c333e0),
	.w4(32'hb7b4495d),
	.w5(32'hb81c6884),
	.w6(32'hb70ca87d),
	.w7(32'h37904778),
	.w8(32'h36827363),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972f834),
	.w1(32'hb986bee1),
	.w2(32'hb88b1f28),
	.w3(32'h38bd5c83),
	.w4(32'hb8200c47),
	.w5(32'hb6061472),
	.w6(32'h38930eec),
	.w7(32'hb9017c68),
	.w8(32'h38b4438a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3841de53),
	.w1(32'h36c6932f),
	.w2(32'hb9be7b8c),
	.w3(32'hb7c0222e),
	.w4(32'hb925a7f4),
	.w5(32'hb9909489),
	.w6(32'h38c7ecec),
	.w7(32'h39237cc7),
	.w8(32'hb90792f6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1c2bb),
	.w1(32'hb9bf2a02),
	.w2(32'h3939d0cd),
	.w3(32'h391c5883),
	.w4(32'h38663948),
	.w5(32'h39a8dbe3),
	.w6(32'h38bd0a34),
	.w7(32'h3970c82d),
	.w8(32'h3946939e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f6ebc),
	.w1(32'hba24f38f),
	.w2(32'hba86dbee),
	.w3(32'hb823409c),
	.w4(32'hb973008e),
	.w5(32'hba008daf),
	.w6(32'h399e31aa),
	.w7(32'h392bab39),
	.w8(32'hb9a1ac19),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389c2de9),
	.w1(32'hb94af322),
	.w2(32'hb735438a),
	.w3(32'h38a42428),
	.w4(32'hb819a601),
	.w5(32'h398ff2d5),
	.w6(32'h38340c21),
	.w7(32'hb95bda8f),
	.w8(32'h39888975),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8b0ec),
	.w1(32'hb9c9e5d8),
	.w2(32'h38c65637),
	.w3(32'hb8dccf59),
	.w4(32'hb98fbea2),
	.w5(32'h399aba07),
	.w6(32'h3920c655),
	.w7(32'h38dc0b7e),
	.w8(32'h396fc5b0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b63542),
	.w1(32'hb88acc40),
	.w2(32'hb8ebdb2e),
	.w3(32'hb7804c46),
	.w4(32'hb68449a1),
	.w5(32'hb8a8e7a0),
	.w6(32'hb7625dc9),
	.w7(32'hb828cd9b),
	.w8(32'hb886ca83),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e7728),
	.w1(32'hb892894a),
	.w2(32'h3862e91e),
	.w3(32'h39fae219),
	.w4(32'hb93105e4),
	.w5(32'hb84b3e0d),
	.w6(32'h394846b8),
	.w7(32'h3a062c22),
	.w8(32'h39b44df5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394581d5),
	.w1(32'hb85dca3c),
	.w2(32'h378896d1),
	.w3(32'h38c09d9d),
	.w4(32'hb900fb74),
	.w5(32'h39151cdb),
	.w6(32'hb806fe45),
	.w7(32'hb88439b0),
	.w8(32'hb8c0ce94),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb778a1f2),
	.w1(32'hb7a9d26f),
	.w2(32'hb7bb1772),
	.w3(32'hb73e49fd),
	.w4(32'hb795a979),
	.w5(32'hb7b7a613),
	.w6(32'hb797c093),
	.w7(32'hb767d873),
	.w8(32'hb7ab045f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7edcd38),
	.w1(32'h381d43f4),
	.w2(32'hb81025f7),
	.w3(32'hb5f86e46),
	.w4(32'h371592a1),
	.w5(32'h37a25825),
	.w6(32'h3835d0c7),
	.w7(32'h3917ca60),
	.w8(32'h380c20a3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8177498),
	.w1(32'hb9081602),
	.w2(32'h38caed2e),
	.w3(32'h38df3481),
	.w4(32'hb8eca379),
	.w5(32'h38f0934c),
	.w6(32'hb89f51b3),
	.w7(32'hb9a110d7),
	.w8(32'hb89f9cd1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e43471),
	.w1(32'hb8790036),
	.w2(32'h37e08118),
	.w3(32'h3717eba8),
	.w4(32'hb781b0c7),
	.w5(32'h395586a7),
	.w6(32'hb85522b7),
	.w7(32'hb8b660fc),
	.w8(32'h39430002),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8479162),
	.w1(32'hb722ef83),
	.w2(32'hb925eea3),
	.w3(32'h390fb22d),
	.w4(32'h389cc00d),
	.w5(32'hb942d4a2),
	.w6(32'h38ad2e3a),
	.w7(32'h38c63ee2),
	.w8(32'h3703483a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38691e8a),
	.w1(32'hb6496bd9),
	.w2(32'hb8770de9),
	.w3(32'h383b38b0),
	.w4(32'hb6bb2b78),
	.w5(32'hb8777143),
	.w6(32'h38941c81),
	.w7(32'h390acf17),
	.w8(32'h3913f727),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b52d03),
	.w1(32'hb956c58b),
	.w2(32'hb91118a2),
	.w3(32'h37fe6a1e),
	.w4(32'hb88fb9fe),
	.w5(32'hb8422280),
	.w6(32'h39513a32),
	.w7(32'h3859653d),
	.w8(32'hb832b404),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d328dc),
	.w1(32'hb8d73c18),
	.w2(32'h37aa3cbb),
	.w3(32'hb83b51b2),
	.w4(32'hb8b68b64),
	.w5(32'h38c792c5),
	.w6(32'h3808f441),
	.w7(32'h38be9f85),
	.w8(32'h39178426),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388915cf),
	.w1(32'hb80ad1bd),
	.w2(32'h38a86fa1),
	.w3(32'h3885aea4),
	.w4(32'hb7b27896),
	.w5(32'h38e338ff),
	.w6(32'hb7a2b638),
	.w7(32'hb91596c9),
	.w8(32'h37d8e001),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb601df7a),
	.w1(32'hb5ca64de),
	.w2(32'hb66f8108),
	.w3(32'hb6681c69),
	.w4(32'hb6081fba),
	.w5(32'hb52c979f),
	.w6(32'hb591947d),
	.w7(32'h316f773c),
	.w8(32'h355dbcc2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fc2b86),
	.w1(32'hb6d90312),
	.w2(32'hb762f93e),
	.w3(32'hb5a5cb08),
	.w4(32'hb6b9e1e3),
	.w5(32'hb73e3235),
	.w6(32'h366e9e49),
	.w7(32'h36e61030),
	.w8(32'hb5e1a69d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h31b0abf6),
	.w1(32'h368accda),
	.w2(32'h35b637dc),
	.w3(32'h35a61785),
	.w4(32'h36abfc00),
	.w5(32'hb59d28d1),
	.w6(32'hb5f269f0),
	.w7(32'h35c4e824),
	.w8(32'h35e7073b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cd8a05),
	.w1(32'hb85d702b),
	.w2(32'hb8926b1f),
	.w3(32'hb7a8887f),
	.w4(32'hb840f08d),
	.w5(32'hb84c7f73),
	.w6(32'h373821a1),
	.w7(32'h37bd9111),
	.w8(32'h371c1965),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bad37f),
	.w1(32'hb7bf524c),
	.w2(32'h3735de5e),
	.w3(32'h38c49834),
	.w4(32'hb77e3236),
	.w5(32'h3903ea34),
	.w6(32'hb6755304),
	.w7(32'hb8678489),
	.w8(32'h3905ff43),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385768d8),
	.w1(32'h3825dee1),
	.w2(32'hb75e2c74),
	.w3(32'h3730417f),
	.w4(32'hb7b13725),
	.w5(32'hb85d6700),
	.w6(32'hb7a2746d),
	.w7(32'h37a0fea5),
	.w8(32'h37b6c260),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83f2e47),
	.w1(32'hb91eaa1a),
	.w2(32'h37e8dd06),
	.w3(32'h38a99f82),
	.w4(32'h369988dc),
	.w5(32'h38975381),
	.w6(32'h391c1605),
	.w7(32'hb802afa1),
	.w8(32'h388b3819),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e5a4d),
	.w1(32'h3751f580),
	.w2(32'hb91d28d2),
	.w3(32'h37aa7439),
	.w4(32'h37d284b2),
	.w5(32'hb92b6814),
	.w6(32'h38cb4d17),
	.w7(32'h3797ed05),
	.w8(32'hb82cf2b9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c7bc8d),
	.w1(32'hb6a64578),
	.w2(32'hb62938c4),
	.w3(32'hb721a6e0),
	.w4(32'hb6ff0213),
	.w5(32'hb4ead398),
	.w6(32'hb726a6ef),
	.w7(32'hb71505a5),
	.w8(32'hb6b3e5ad),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d209cd),
	.w1(32'hb7bfe791),
	.w2(32'hb8166a78),
	.w3(32'hb7f81002),
	.w4(32'hb7a9c2dd),
	.w5(32'hb7c8c9e1),
	.w6(32'hb70075f1),
	.w7(32'hb4c505b8),
	.w8(32'h35dcbd09),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4dea5ce),
	.w1(32'h362c3199),
	.w2(32'hb61d6301),
	.w3(32'h3475f884),
	.w4(32'h3493f8b5),
	.w5(32'hb67f85f1),
	.w6(32'h34a9ad5f),
	.w7(32'hb52f2b3f),
	.w8(32'hb6b6c1f7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3758e06f),
	.w1(32'h3a02e8ff),
	.w2(32'h38f326b8),
	.w3(32'hb7debc08),
	.w4(32'h399b20c7),
	.w5(32'h39c0e394),
	.w6(32'h3a38bf7d),
	.w7(32'h3a2cb553),
	.w8(32'h3a17c0a5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9db21),
	.w1(32'h39e0ee06),
	.w2(32'h3a0d72ae),
	.w3(32'h3a0a5dd7),
	.w4(32'h39a6f816),
	.w5(32'h3938f806),
	.w6(32'h3a42b4b9),
	.w7(32'h3a0afdad),
	.w8(32'h39cd5b63),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3818c49a),
	.w1(32'h38c48595),
	.w2(32'h37812842),
	.w3(32'h393a313f),
	.w4(32'h3b0265e0),
	.w5(32'h3a908c2c),
	.w6(32'h39973727),
	.w7(32'h3949ff4b),
	.w8(32'hba1c1224),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9792c57),
	.w1(32'h3a686062),
	.w2(32'h3a8a9563),
	.w3(32'h385e5caa),
	.w4(32'h3a1e11b8),
	.w5(32'h39e7f33e),
	.w6(32'h3a17a56d),
	.w7(32'h3a4b86c8),
	.w8(32'h3a58103f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86e8ab),
	.w1(32'h39e9e85f),
	.w2(32'h3a1ce225),
	.w3(32'h39c0b88f),
	.w4(32'hb8ca5287),
	.w5(32'hb9cb630c),
	.w6(32'hb9b42f7c),
	.w7(32'h384326bf),
	.w8(32'h3a0a71e2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b966a),
	.w1(32'hba3e4fab),
	.w2(32'hb94087f4),
	.w3(32'hb7e7a310),
	.w4(32'hbafac11c),
	.w5(32'hbb226f3b),
	.w6(32'hbaaa151b),
	.w7(32'hbae0c7ff),
	.w8(32'hbafc4de8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3fd6b),
	.w1(32'hb9b7fb5a),
	.w2(32'hbaf8682b),
	.w3(32'hbabfc3ea),
	.w4(32'hba147b72),
	.w5(32'hba922703),
	.w6(32'hba5c5088),
	.w7(32'hbad01045),
	.w8(32'hba15ceb5),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d294bc),
	.w1(32'h3ab842f4),
	.w2(32'h3aa38265),
	.w3(32'hba5d7921),
	.w4(32'h3ac492dc),
	.w5(32'h3aad9c79),
	.w6(32'h3ad7e276),
	.w7(32'h3ae0f3fb),
	.w8(32'h3af4c5f3),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1d318),
	.w1(32'h3937a853),
	.w2(32'h3a8dfab3),
	.w3(32'h3ad24028),
	.w4(32'h39ead7e3),
	.w5(32'h3a42c386),
	.w6(32'hb8b80ddd),
	.w7(32'h3930a730),
	.w8(32'h3a0c5b71),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e90c4),
	.w1(32'h3a849bf3),
	.w2(32'h3a5415b6),
	.w3(32'h3a6dfe5d),
	.w4(32'h3a821f82),
	.w5(32'h3a313c52),
	.w6(32'h3a6c29ad),
	.w7(32'h3a532de5),
	.w8(32'h3a0b9517),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0bd92),
	.w1(32'h39f13fc2),
	.w2(32'h3a6298bf),
	.w3(32'h3a206094),
	.w4(32'hb896f48f),
	.w5(32'h39a2768c),
	.w6(32'h3a7d5451),
	.w7(32'h3a90f9df),
	.w8(32'h3a1b52b2),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27f9e5),
	.w1(32'hba982e7c),
	.w2(32'hb93e9e8c),
	.w3(32'h3a3a5bc7),
	.w4(32'hba39465a),
	.w5(32'hb905fd1a),
	.w6(32'hba1a4ce3),
	.w7(32'hba2d8319),
	.w8(32'h398fe53b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399519d3),
	.w1(32'hba829e9a),
	.w2(32'hba6e075a),
	.w3(32'h38044083),
	.w4(32'hba0922c5),
	.w5(32'hb886586d),
	.w6(32'hb9dcf2bb),
	.w7(32'hba9023de),
	.w8(32'hba9a0ebb),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7442e),
	.w1(32'hb9a41325),
	.w2(32'h3a79532c),
	.w3(32'hb78a9d27),
	.w4(32'hba0743ab),
	.w5(32'h39831df8),
	.w6(32'hba81f2de),
	.w7(32'hba9d7b30),
	.w8(32'hba80b379),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83ac4ef),
	.w1(32'h39a6889d),
	.w2(32'h399ca0f7),
	.w3(32'h36480e9e),
	.w4(32'h3a082f65),
	.w5(32'h3a306660),
	.w6(32'h3a05abb7),
	.w7(32'h39f10878),
	.w8(32'h3a092bd3),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984de3c),
	.w1(32'h3aa08157),
	.w2(32'h3a6e4ac5),
	.w3(32'h3a2b9270),
	.w4(32'h3af05281),
	.w5(32'h3aaaa342),
	.w6(32'h3a076fe9),
	.w7(32'h39bbb0ca),
	.w8(32'hb9730a70),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb783c935),
	.w1(32'hb98e22c9),
	.w2(32'hb9a5a731),
	.w3(32'h3a444583),
	.w4(32'hb933ac8d),
	.w5(32'hba436825),
	.w6(32'hbad09bb2),
	.w7(32'hbadd5674),
	.w8(32'hbaa15d16),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd597b),
	.w1(32'h3a4189be),
	.w2(32'h3a5fe729),
	.w3(32'hbab9df32),
	.w4(32'hb794267c),
	.w5(32'hb8d9ae88),
	.w6(32'h3a41935e),
	.w7(32'h3a78d0c2),
	.w8(32'h3a511b93),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf6b2b),
	.w1(32'h39fd4f48),
	.w2(32'h3a4c289f),
	.w3(32'h38b90c84),
	.w4(32'h3a177308),
	.w5(32'h3a18efa5),
	.w6(32'h394cb5a9),
	.w7(32'h3a3f78a4),
	.w8(32'hb8aa1b63),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ddbcaa),
	.w1(32'hb910daa2),
	.w2(32'h39d33f17),
	.w3(32'h3a7d0a6d),
	.w4(32'hb9c83129),
	.w5(32'hb9953459),
	.w6(32'hb866fbf6),
	.w7(32'h3965a615),
	.w8(32'h3a31e84f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398feac3),
	.w1(32'hb97a7d5b),
	.w2(32'h390fae37),
	.w3(32'h390e3ea0),
	.w4(32'hb8eb3ea2),
	.w5(32'hb6fba9ba),
	.w6(32'hb9983907),
	.w7(32'h39006562),
	.w8(32'h398d5322),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11ab61),
	.w1(32'h39cc7336),
	.w2(32'h3a35b0ba),
	.w3(32'h3912ea83),
	.w4(32'h395ce8c6),
	.w5(32'h3a1548e1),
	.w6(32'h39baa49b),
	.w7(32'h3a1aa29a),
	.w8(32'h38d1bfa7),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fef80b),
	.w1(32'h3a187c3b),
	.w2(32'h3a1ce7c4),
	.w3(32'h38fbe530),
	.w4(32'h3a92de64),
	.w5(32'h3aad5846),
	.w6(32'h3aaaaeee),
	.w7(32'h3ab3d4ff),
	.w8(32'h3a3cf148),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394075bb),
	.w1(32'h39a29677),
	.w2(32'h3ae13ff3),
	.w3(32'h3abcac69),
	.w4(32'h3abcc3b7),
	.w5(32'h3ab0452b),
	.w6(32'hba849737),
	.w7(32'hba2a6e94),
	.w8(32'hb7b0a374),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14306a),
	.w1(32'h39122f56),
	.w2(32'hba517160),
	.w3(32'h3a420ffe),
	.w4(32'hba5a0146),
	.w5(32'hba865813),
	.w6(32'h3a2211d0),
	.w7(32'hb9906ca5),
	.w8(32'hba077b21),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803a7e),
	.w1(32'h3a559b1a),
	.w2(32'h3a8ea673),
	.w3(32'hbaa3c5b9),
	.w4(32'h3a8076e0),
	.w5(32'h3a89a16b),
	.w6(32'h3aa388a2),
	.w7(32'h3a9014ad),
	.w8(32'h3a47da7b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccf289),
	.w1(32'h3998f2fe),
	.w2(32'h39fa74ba),
	.w3(32'h3a307539),
	.w4(32'hb9c5a026),
	.w5(32'hba5e405b),
	.w6(32'hb80747b4),
	.w7(32'h38ead283),
	.w8(32'h38abf992),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ac511),
	.w1(32'hb9c5340d),
	.w2(32'hba36d3b3),
	.w3(32'hb96c3190),
	.w4(32'h3959fc7f),
	.w5(32'hb7ff3e5a),
	.w6(32'hba4eaafe),
	.w7(32'hba8efcf8),
	.w8(32'hba9a7178),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21b9a5),
	.w1(32'h39a7afac),
	.w2(32'h388ba877),
	.w3(32'h38da3bbf),
	.w4(32'h3932e0b8),
	.w5(32'h39e1e7fa),
	.w6(32'h3a48eb5f),
	.w7(32'h3a1e7b58),
	.w8(32'h37b11240),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ef1db8),
	.w1(32'hba849aea),
	.w2(32'hba29fb11),
	.w3(32'h39ed701e),
	.w4(32'hbac8db06),
	.w5(32'hbada7a99),
	.w6(32'hba7e02e5),
	.w7(32'hba684da5),
	.w8(32'hb9cd172d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba783e03),
	.w1(32'hb9820a59),
	.w2(32'hba49cd1e),
	.w3(32'hbac9d7ac),
	.w4(32'hba1a50bc),
	.w5(32'hba4e6cd8),
	.w6(32'h36e728be),
	.w7(32'h395bd975),
	.w8(32'h376259ff),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6884b4),
	.w1(32'h3a3c45d5),
	.w2(32'h39ec9073),
	.w3(32'hba19603e),
	.w4(32'h3a234185),
	.w5(32'h396f4a2f),
	.w6(32'h3a3e9659),
	.w7(32'h3a6e5dd3),
	.w8(32'h3921b805),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b7382),
	.w1(32'h3a6a4e3c),
	.w2(32'h3a07fdbe),
	.w3(32'h397ae423),
	.w4(32'h3a8b75a3),
	.w5(32'h3a8640e8),
	.w6(32'h3aae981d),
	.w7(32'h3a976c58),
	.w8(32'h3a32f990),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947287d),
	.w1(32'h3a2eeb39),
	.w2(32'h39f9a01e),
	.w3(32'h3a732bef),
	.w4(32'h3a4c0e0b),
	.w5(32'h3a491996),
	.w6(32'h3a93294a),
	.w7(32'h3a810776),
	.w8(32'h3a385ef3),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cecf89),
	.w1(32'h3a09c310),
	.w2(32'h39335b7b),
	.w3(32'h3a6453aa),
	.w4(32'h3945f9ff),
	.w5(32'h3a70c817),
	.w6(32'h3916d320),
	.w7(32'hb9f7450c),
	.w8(32'hbad62a65),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99cdeb3),
	.w1(32'hba4cc4e9),
	.w2(32'hb99f3395),
	.w3(32'hb9964d3c),
	.w4(32'hba7764d1),
	.w5(32'h39702545),
	.w6(32'hb9ba585e),
	.w7(32'hba054630),
	.w8(32'hba06b616),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f9148),
	.w1(32'hb9a0506d),
	.w2(32'h394896fd),
	.w3(32'hb97f9891),
	.w4(32'hb9a98029),
	.w5(32'h39ccbb3c),
	.w6(32'hb9f35e97),
	.w7(32'hb99ab6ce),
	.w8(32'h39f04378),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a844aa0),
	.w1(32'hb970945f),
	.w2(32'hba205e0e),
	.w3(32'h3a235658),
	.w4(32'hb89aad81),
	.w5(32'hb95610ca),
	.w6(32'h38370c7b),
	.w7(32'hb9124c32),
	.w8(32'hb9d0bdab),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71419d),
	.w1(32'h3a4b258b),
	.w2(32'h3a77b65b),
	.w3(32'hb98190bd),
	.w4(32'h39fa4ac1),
	.w5(32'h3a255410),
	.w6(32'hb88f69e4),
	.w7(32'h39f2515e),
	.w8(32'h3a2ef768),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cb5eb),
	.w1(32'h3a127b9c),
	.w2(32'h3a45984b),
	.w3(32'h39545585),
	.w4(32'h3a06a46f),
	.w5(32'h39d2c348),
	.w6(32'h39aeb286),
	.w7(32'h3a321cf3),
	.w8(32'h3a2802ff),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12af35),
	.w1(32'h3a4735ba),
	.w2(32'h3a3398f9),
	.w3(32'h3a0c4a7d),
	.w4(32'h3a2595f5),
	.w5(32'h39a475da),
	.w6(32'h3a7b52ff),
	.w7(32'h3a80a864),
	.w8(32'h3a1add15),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39200c0f),
	.w1(32'h399c59ec),
	.w2(32'h3a2b429d),
	.w3(32'h39c24da9),
	.w4(32'h38cb1cbd),
	.w5(32'h397ca6a3),
	.w6(32'hb94cb83e),
	.w7(32'hb840c24f),
	.w8(32'h394cd782),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f17d31),
	.w1(32'h38d83fe4),
	.w2(32'hb9850c25),
	.w3(32'h396be5cc),
	.w4(32'h39a79e51),
	.w5(32'h38f76c49),
	.w6(32'h3a375db0),
	.w7(32'h3a3c12fb),
	.w8(32'h392aac45),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba940925),
	.w1(32'h39da530a),
	.w2(32'h39a7bc4b),
	.w3(32'hb9b8e4e3),
	.w4(32'h372f40be),
	.w5(32'hb955095a),
	.w6(32'hb86a98d6),
	.w7(32'hb981abd6),
	.w8(32'hb9132873),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3970e939),
	.w1(32'h3a3e64f4),
	.w2(32'h3a778358),
	.w3(32'h384bc400),
	.w4(32'h3a52291a),
	.w5(32'h3a8755d5),
	.w6(32'h3a60eb52),
	.w7(32'h3a443fff),
	.w8(32'h3a605b4d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a138d96),
	.w1(32'hba99cfca),
	.w2(32'hba66d3cc),
	.w3(32'h3a473adf),
	.w4(32'hba650a75),
	.w5(32'hba89dc8e),
	.w6(32'hba885d69),
	.w7(32'hba6cfa65),
	.w8(32'hb8392a6a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d339a3),
	.w1(32'hba856fc0),
	.w2(32'hba494b89),
	.w3(32'hb96fd464),
	.w4(32'hba670ece),
	.w5(32'hba13834e),
	.w6(32'hba956fcf),
	.w7(32'hbab0b87e),
	.w8(32'hba384d61),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba590a54),
	.w1(32'hba5df8e1),
	.w2(32'h393f5933),
	.w3(32'hba3700ad),
	.w4(32'hba144eb5),
	.w5(32'hb94e3187),
	.w6(32'hbab38504),
	.w7(32'hb9a89745),
	.w8(32'hb9c79db7),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e497d8),
	.w1(32'hb93433a2),
	.w2(32'h3af48079),
	.w3(32'h3902c33d),
	.w4(32'hb767cf4b),
	.w5(32'h39f12652),
	.w6(32'hba87fc4b),
	.w7(32'hbae3d34f),
	.w8(32'hba4d119c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8ac1b),
	.w1(32'h3a2db779),
	.w2(32'h3a777e2d),
	.w3(32'h394cbbbc),
	.w4(32'hba0a1171),
	.w5(32'hb8f29246),
	.w6(32'h37e5a88c),
	.w7(32'h3aa5c466),
	.w8(32'h396b9858),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb893a340),
	.w1(32'h39ab39b3),
	.w2(32'h39c9c66c),
	.w3(32'hb9721472),
	.w4(32'h38eb6922),
	.w5(32'h3a02e353),
	.w6(32'h3a2ad678),
	.w7(32'h3a0e393d),
	.w8(32'h3a029a9e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d3bfd),
	.w1(32'h3a9fa11f),
	.w2(32'h3a6277ce),
	.w3(32'h39ff6a2c),
	.w4(32'h3a9fa4cd),
	.w5(32'h3a1b402f),
	.w6(32'h3a86f210),
	.w7(32'h3a629e72),
	.w8(32'h39c50bb2),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384aeb31),
	.w1(32'hb9d75fe8),
	.w2(32'hb8158d89),
	.w3(32'h395b8016),
	.w4(32'hb9348ddb),
	.w5(32'hb90fa736),
	.w6(32'hba41e159),
	.w7(32'hb97e8991),
	.w8(32'hb969288b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c10a47),
	.w1(32'hb9f7f936),
	.w2(32'h3ab29349),
	.w3(32'hb91f9191),
	.w4(32'hbb09176b),
	.w5(32'hbafee731),
	.w6(32'hba06d145),
	.w7(32'hba638ce0),
	.w8(32'hbb050a62),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97df6b),
	.w1(32'h3aa55997),
	.w2(32'h3aa7c6a5),
	.w3(32'hbabe5054),
	.w4(32'h3a88c0c0),
	.w5(32'h3a25176d),
	.w6(32'h3addec5e),
	.w7(32'h3adca6c2),
	.w8(32'h3acf77d3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5566e1),
	.w1(32'hba86f67d),
	.w2(32'hbaa4b399),
	.w3(32'h3a09475a),
	.w4(32'hba1e9e22),
	.w5(32'hb9eac4da),
	.w6(32'hba980725),
	.w7(32'hbad85cb7),
	.w8(32'hba7b3d2e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6433bcf),
	.w1(32'hba5fc30c),
	.w2(32'hba67b5a2),
	.w3(32'hb9fffae2),
	.w4(32'hba47888c),
	.w5(32'hb9ed233c),
	.w6(32'hba1d37d4),
	.w7(32'hba154e77),
	.w8(32'hb9022590),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c0057),
	.w1(32'hb994ab62),
	.w2(32'hbabc7678),
	.w3(32'hba01fe4f),
	.w4(32'hb8e3e6a1),
	.w5(32'hba3c238e),
	.w6(32'h39f684ed),
	.w7(32'hb817b51c),
	.w8(32'hb9ff37ff),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba890c44),
	.w1(32'hb982f2d4),
	.w2(32'h371bf15e),
	.w3(32'hb9c30dd5),
	.w4(32'hb975378f),
	.w5(32'hb9b897a2),
	.w6(32'h39de546a),
	.w7(32'h3a255771),
	.w8(32'h396a35be),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0a10e),
	.w1(32'hb9c56b0a),
	.w2(32'hbaa848e0),
	.w3(32'hb5ffd963),
	.w4(32'h3941943f),
	.w5(32'h38596674),
	.w6(32'hba98bd6b),
	.w7(32'hba934f27),
	.w8(32'hba455981),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12af2e),
	.w1(32'h3a045162),
	.w2(32'h3a246d5b),
	.w3(32'hb9babe23),
	.w4(32'h387f3b6e),
	.w5(32'hb8b74ae0),
	.w6(32'hb89e6d4f),
	.w7(32'h38a2bcbd),
	.w8(32'h39ad226c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a001f0d),
	.w1(32'h3a9c2455),
	.w2(32'h3aaaca38),
	.w3(32'hb9361f40),
	.w4(32'h3a77f3e8),
	.w5(32'h3ab08cb9),
	.w6(32'h3a60d5fc),
	.w7(32'h3a61ff9c),
	.w8(32'h3a08b6ac),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393dd6b7),
	.w1(32'h39544ab6),
	.w2(32'h3960f269),
	.w3(32'h39c77c40),
	.w4(32'hb939053a),
	.w5(32'hb951574e),
	.w6(32'hb8c2a5cc),
	.w7(32'h3975d980),
	.w8(32'h39a33879),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d0710),
	.w1(32'h3a87ee56),
	.w2(32'h3a65a942),
	.w3(32'h37f4fed7),
	.w4(32'h3a94cb8c),
	.w5(32'h3a7334e3),
	.w6(32'h3aa30542),
	.w7(32'h3a93f4ca),
	.w8(32'h3a2769df),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39136fb2),
	.w1(32'h3a1b3360),
	.w2(32'hba935af2),
	.w3(32'h3a37a3a1),
	.w4(32'h3a4fee1e),
	.w5(32'h3a8ce3f7),
	.w6(32'h380ce3da),
	.w7(32'hba3eec1c),
	.w8(32'hbab1271f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d0988),
	.w1(32'hba83a604),
	.w2(32'hba30166d),
	.w3(32'hb91b003a),
	.w4(32'hba440495),
	.w5(32'hba35d72f),
	.w6(32'hba652468),
	.w7(32'hba32d429),
	.w8(32'hb80ae48f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ebdfb),
	.w1(32'hba453975),
	.w2(32'hb9381eb4),
	.w3(32'hb924d854),
	.w4(32'hba3a77ff),
	.w5(32'hba04ca0f),
	.w6(32'hba8032c7),
	.w7(32'hba1a422f),
	.w8(32'hb91e4597),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f0895a),
	.w1(32'hba2885be),
	.w2(32'hb9dd0058),
	.w3(32'hb9c15426),
	.w4(32'hb9c48015),
	.w5(32'hb9d885c4),
	.w6(32'hbab2b503),
	.w7(32'hb9ccacbc),
	.w8(32'hb94cf7a9),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94c13dc),
	.w1(32'h39b948fe),
	.w2(32'hb99d73e5),
	.w3(32'hb5fe737b),
	.w4(32'h3a8f3804),
	.w5(32'h3a150a2d),
	.w6(32'h3a2b31a2),
	.w7(32'h39587ee0),
	.w8(32'h3943a5f0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb803a9ef),
	.w1(32'hb8e5c4fe),
	.w2(32'hb96fc101),
	.w3(32'h3a65fb64),
	.w4(32'hba445554),
	.w5(32'hba98f297),
	.w6(32'hb973a1a4),
	.w7(32'hb822b22b),
	.w8(32'hb9fe03ad),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95040b),
	.w1(32'h3a5cc056),
	.w2(32'h3a707739),
	.w3(32'hba9febc9),
	.w4(32'h3a3eaf27),
	.w5(32'h3911c67b),
	.w6(32'h3a923975),
	.w7(32'h3a8485b3),
	.w8(32'h3a3dbc13),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d636b),
	.w1(32'hbab0e727),
	.w2(32'hba8b0d2b),
	.w3(32'h395627bd),
	.w4(32'hba7a4499),
	.w5(32'hba718560),
	.w6(32'hbb2b9c58),
	.w7(32'hbada7d9c),
	.w8(32'hbae46464),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1ec96),
	.w1(32'h39b7c935),
	.w2(32'h3a09086a),
	.w3(32'hba1df184),
	.w4(32'h3806a889),
	.w5(32'h3866402d),
	.w6(32'h39c65854),
	.w7(32'h39f11ed8),
	.w8(32'h3a18f99b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa012e),
	.w1(32'h39fd330f),
	.w2(32'h39397e9e),
	.w3(32'h39677ebb),
	.w4(32'h39e543d7),
	.w5(32'h39711efb),
	.w6(32'h3a406114),
	.w7(32'h3a0cca76),
	.w8(32'h39dc897c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a939d),
	.w1(32'h3a22f98a),
	.w2(32'h3a2da199),
	.w3(32'h39cc673d),
	.w4(32'h39ec1b8d),
	.w5(32'h39a729e4),
	.w6(32'h3a68fb6d),
	.w7(32'h3a7cd3e5),
	.w8(32'h39e13191),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c66395),
	.w1(32'h3a140cc8),
	.w2(32'h39a402c7),
	.w3(32'h39a94f32),
	.w4(32'h3a761322),
	.w5(32'h3a55e8eb),
	.w6(32'h3a940b01),
	.w7(32'h3a499e47),
	.w8(32'h39aa8301),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b9066),
	.w1(32'h39f248b5),
	.w2(32'h3a3ed5f2),
	.w3(32'h3a53e903),
	.w4(32'hba04eb55),
	.w5(32'hba23e6ba),
	.w6(32'hb8f459ef),
	.w7(32'h387a1267),
	.w8(32'h39ab09a1),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398795cf),
	.w1(32'hba5b4c66),
	.w2(32'h3a9f1581),
	.w3(32'hba046b28),
	.w4(32'hba769d4f),
	.w5(32'hb9d902ec),
	.w6(32'hba490b84),
	.w7(32'hbb056353),
	.w8(32'hbb23b958),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a9f52),
	.w1(32'h3a777050),
	.w2(32'h3a26bbad),
	.w3(32'h3a0f8fe6),
	.w4(32'h3a94d216),
	.w5(32'h3a4702f8),
	.w6(32'h3a9dcf70),
	.w7(32'h3a6c8de1),
	.w8(32'h3a19451b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb798dd39),
	.w1(32'h3a2c1d5d),
	.w2(32'h391ef4cd),
	.w3(32'h3a2fcc03),
	.w4(32'h39538d42),
	.w5(32'hb85af957),
	.w6(32'h39aa92d5),
	.w7(32'h39320cf8),
	.w8(32'h3920ba23),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392cb1d0),
	.w1(32'hba7c49e1),
	.w2(32'hb9700d17),
	.w3(32'hb971063e),
	.w4(32'hba8763ad),
	.w5(32'hba032c97),
	.w6(32'hba602fc0),
	.w7(32'hba5ec8f0),
	.w8(32'hb9a21aaa),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ffc7d1),
	.w1(32'h3aba7ae0),
	.w2(32'h3aa538be),
	.w3(32'hb999a737),
	.w4(32'h3acbcca6),
	.w5(32'h3acf17f3),
	.w6(32'h3aed8053),
	.w7(32'h3adf8424),
	.w8(32'h3a92ee7a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81d234),
	.w1(32'h38244f24),
	.w2(32'hba30bb2e),
	.w3(32'h3ab7c49a),
	.w4(32'hb8e48f2b),
	.w5(32'hba308e42),
	.w6(32'h386d82b3),
	.w7(32'h390631f4),
	.w8(32'hb9545b25),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3302b),
	.w1(32'h39e386e0),
	.w2(32'h3a5b0358),
	.w3(32'hba816eca),
	.w4(32'h39a12b4b),
	.w5(32'h39e45f01),
	.w6(32'h363ce7dd),
	.w7(32'h3a0aab3c),
	.w8(32'h3a3b39cd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a823423),
	.w1(32'h3a227969),
	.w2(32'h3911886f),
	.w3(32'h3a0edc87),
	.w4(32'h39215d14),
	.w5(32'hb9748d63),
	.w6(32'h39c1f8d6),
	.w7(32'h3a014d65),
	.w8(32'h391848f1),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6d977),
	.w1(32'h393bfbdc),
	.w2(32'h3975c2d8),
	.w3(32'hb933dd10),
	.w4(32'h398f7d7e),
	.w5(32'h384e668e),
	.w6(32'hb9818a38),
	.w7(32'h38b550f8),
	.w8(32'h383e1a3e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11c801),
	.w1(32'h397af14a),
	.w2(32'h3a1595a5),
	.w3(32'h39706237),
	.w4(32'hba5aa6bb),
	.w5(32'h36efb925),
	.w6(32'h399eeec9),
	.w7(32'h3a93723e),
	.w8(32'h38931168),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397bf9b4),
	.w1(32'h39f2253b),
	.w2(32'h39a21dc4),
	.w3(32'hb9789fe7),
	.w4(32'h39ef6559),
	.w5(32'h39886e9d),
	.w6(32'h3a0b193a),
	.w7(32'h39caa504),
	.w8(32'h39d395d5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f47618),
	.w1(32'hb9c28620),
	.w2(32'h3a1fa498),
	.w3(32'h38f5985d),
	.w4(32'hb841fb77),
	.w5(32'h3a3e360e),
	.w6(32'hba264121),
	.w7(32'hb9f9d98b),
	.w8(32'hb9ea38bc),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38194b7a),
	.w1(32'h3a26d34b),
	.w2(32'h3a1dbe92),
	.w3(32'h39295c43),
	.w4(32'h3a894d8b),
	.w5(32'h3a860314),
	.w6(32'h3a93efbe),
	.w7(32'h3a94bb60),
	.w8(32'h3a1b6326),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ee52a),
	.w1(32'hb90d8851),
	.w2(32'hb981cdfd),
	.w3(32'h3a6327d5),
	.w4(32'hb90d7146),
	.w5(32'hb8a3ee9f),
	.w6(32'hb955f576),
	.w7(32'hb93c5a6d),
	.w8(32'h397ecd27),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb58764da),
	.w1(32'h3a868a60),
	.w2(32'h3a473ecc),
	.w3(32'hb9172811),
	.w4(32'h3a9389e7),
	.w5(32'h3a8818e4),
	.w6(32'h3ae3b5ba),
	.w7(32'h3ac12f96),
	.w8(32'h3a72019a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a369dc8),
	.w1(32'h3a61757d),
	.w2(32'h3a5fed68),
	.w3(32'h3acef38a),
	.w4(32'h3ac649a6),
	.w5(32'h3abeb558),
	.w6(32'h3aab169a),
	.w7(32'h3a93d2fb),
	.w8(32'h3a2d42fe),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a4ae0),
	.w1(32'hb7b9d038),
	.w2(32'h39ba08e5),
	.w3(32'h3a42364d),
	.w4(32'h38bbefeb),
	.w5(32'h39fdb6c3),
	.w6(32'h3a24edc5),
	.w7(32'h3a407df2),
	.w8(32'h3a107f68),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10ff32),
	.w1(32'h3a3c8255),
	.w2(32'h3a12a4d6),
	.w3(32'h3a3babbe),
	.w4(32'h3a2d4703),
	.w5(32'h39b9108b),
	.w6(32'h3a5bc39a),
	.w7(32'h3a83bc9e),
	.w8(32'h3a7f465c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b0f0f),
	.w1(32'hba5d3eb7),
	.w2(32'hbaf236da),
	.w3(32'h39e9534f),
	.w4(32'hba3615af),
	.w5(32'hbadb7487),
	.w6(32'h364d59b7),
	.w7(32'hb96cb517),
	.w8(32'hba076354),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4ecbf),
	.w1(32'h39a1e9c5),
	.w2(32'h3976602b),
	.w3(32'hbaa55b0f),
	.w4(32'h37543bf9),
	.w5(32'hb99bff73),
	.w6(32'hb9aca51c),
	.w7(32'hb883fc4f),
	.w8(32'h39f5a217),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae5a96),
	.w1(32'hba3a9eae),
	.w2(32'h39c74315),
	.w3(32'hb8f08a2c),
	.w4(32'h3a7e915e),
	.w5(32'h3aa7352e),
	.w6(32'hba3eb3f6),
	.w7(32'hba0f9f82),
	.w8(32'hb999cc9d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67920c),
	.w1(32'h3a49997f),
	.w2(32'h390db658),
	.w3(32'h3aa51abf),
	.w4(32'hb966e3fa),
	.w5(32'hb97eb7a7),
	.w6(32'h39ebb5ee),
	.w7(32'hb96cf33a),
	.w8(32'hba288d93),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c25ff),
	.w1(32'hb8e04117),
	.w2(32'hba328d8b),
	.w3(32'hba33e651),
	.w4(32'hb9e54d48),
	.w5(32'hb9ae7b0d),
	.w6(32'h39acf885),
	.w7(32'hb9916a93),
	.w8(32'hba4b2375),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba358ec5),
	.w1(32'h39f6eba0),
	.w2(32'h3a6923b0),
	.w3(32'hb99201cb),
	.w4(32'h397f7d3b),
	.w5(32'h3a0f5c71),
	.w6(32'hb9a42d46),
	.w7(32'h3937ac6f),
	.w8(32'h3a1b63ab),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae821a),
	.w1(32'h39d60a14),
	.w2(32'h3a4081ee),
	.w3(32'h3a07cdf3),
	.w4(32'hb85a9513),
	.w5(32'h38377360),
	.w6(32'h3a21c2c2),
	.w7(32'h3a4aee4c),
	.w8(32'h3a86d142),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a26c1e),
	.w1(32'hb9514ac3),
	.w2(32'hbac492b7),
	.w3(32'h3857a773),
	.w4(32'h39d0f1b2),
	.w5(32'hba1b17b6),
	.w6(32'hba75d115),
	.w7(32'hbafc2962),
	.w8(32'hba9564bd),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f05704),
	.w1(32'h39863bfd),
	.w2(32'h3ad2c96d),
	.w3(32'hba67d9aa),
	.w4(32'h3950fb10),
	.w5(32'h3a92c627),
	.w6(32'hb93e6bab),
	.w7(32'hb7da348f),
	.w8(32'hba33ded1),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88646ab),
	.w1(32'h3a8a7cc5),
	.w2(32'h3aa146fc),
	.w3(32'h3ae0165d),
	.w4(32'h3ae26977),
	.w5(32'h3ab8da08),
	.w6(32'h3b06cbfe),
	.w7(32'h3ac1b022),
	.w8(32'h3a977312),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7da4c8c),
	.w1(32'h3a213db6),
	.w2(32'h3997c51c),
	.w3(32'h3a86a28b),
	.w4(32'h3a267819),
	.w5(32'h39e083f5),
	.w6(32'h3a6d0c5a),
	.w7(32'h3a0967fb),
	.w8(32'h3a1d6939),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39517852),
	.w1(32'h3a311848),
	.w2(32'h39efeac7),
	.w3(32'h39d388a0),
	.w4(32'h3a5882a6),
	.w5(32'h3a0c4301),
	.w6(32'h3a6b0c97),
	.w7(32'h3a440d6b),
	.w8(32'h3a004d43),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3792a578),
	.w1(32'h39b70132),
	.w2(32'h3a13237e),
	.w3(32'h3a1b055d),
	.w4(32'h392e2c39),
	.w5(32'h3a3993c3),
	.w6(32'h3a2161dc),
	.w7(32'h3a2cf73b),
	.w8(32'h38bc3fba),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39535556),
	.w1(32'h39a3d535),
	.w2(32'h39efbbd0),
	.w3(32'h399cbce3),
	.w4(32'hb8361f64),
	.w5(32'hb8bbb53e),
	.w6(32'hb7829cad),
	.w7(32'h393d2c5b),
	.w8(32'h3a06ea3f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09105c),
	.w1(32'h3a3314e4),
	.w2(32'h39ded9cc),
	.w3(32'h38812fce),
	.w4(32'h3ab1119a),
	.w5(32'h3aae5741),
	.w6(32'h3abdf230),
	.w7(32'h3aafcc42),
	.w8(32'h3a0ffb6c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec707f),
	.w1(32'h3a5b4311),
	.w2(32'h3a143da9),
	.w3(32'h3a917dca),
	.w4(32'h3a861caf),
	.w5(32'h3a2f4073),
	.w6(32'h3a66bff1),
	.w7(32'h3a4bafa2),
	.w8(32'h39fae8bd),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385117ae),
	.w1(32'hba45fb1b),
	.w2(32'hba014ff2),
	.w3(32'h3a1aa91a),
	.w4(32'hb9d649c9),
	.w5(32'hba23bf8e),
	.w6(32'hba85047a),
	.w7(32'hbaaa28eb),
	.w8(32'hb9b560f7),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91dd778),
	.w1(32'h3a2cde60),
	.w2(32'h3a511d86),
	.w3(32'hb9a2071c),
	.w4(32'h39c506de),
	.w5(32'h39493082),
	.w6(32'h3a667664),
	.w7(32'h3a5114f0),
	.w8(32'h39b21f80),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39803b08),
	.w1(32'hba6420a0),
	.w2(32'hbabbced6),
	.w3(32'h39ac4eca),
	.w4(32'hb9cf0877),
	.w5(32'hb90188d1),
	.w6(32'hb9eb486b),
	.w7(32'hbae0a7ef),
	.w8(32'hbaa28177),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43e01c),
	.w1(32'h3a10092b),
	.w2(32'h3a743ae7),
	.w3(32'hb8139da7),
	.w4(32'hb73df106),
	.w5(32'hb8a10c92),
	.w6(32'h3a39fbcb),
	.w7(32'h3a49f39e),
	.w8(32'h3a5f8f92),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb847eb07),
	.w1(32'hb862f556),
	.w2(32'h39980bb2),
	.w3(32'hb9346d71),
	.w4(32'hb9a9e1ef),
	.w5(32'hb875350f),
	.w6(32'hb8f1fe39),
	.w7(32'hb9120637),
	.w8(32'h39b49fbc),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39049df0),
	.w1(32'h39cad406),
	.w2(32'h38893201),
	.w3(32'h38cb4246),
	.w4(32'h3a0a1ea3),
	.w5(32'h38c605a1),
	.w6(32'h39c374b5),
	.w7(32'h38e9ecde),
	.w8(32'hb8e29116),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2bcfc),
	.w1(32'h3a93a699),
	.w2(32'h3a3eda50),
	.w3(32'hb935a91e),
	.w4(32'h3ab17fa4),
	.w5(32'h3a5dabc3),
	.w6(32'h3aab135c),
	.w7(32'h3a92e4f3),
	.w8(32'h3a3396cc),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb602c21f),
	.w1(32'h3a746cc9),
	.w2(32'h3a584670),
	.w3(32'h3a49cc68),
	.w4(32'h3a709858),
	.w5(32'h3a4b2929),
	.w6(32'h3a8c5dc1),
	.w7(32'h3a91cc01),
	.w8(32'h3a526663),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a025e61),
	.w1(32'h3a6c156d),
	.w2(32'h3a4be702),
	.w3(32'h3a5d58dc),
	.w4(32'h3a52082f),
	.w5(32'h3a29b64a),
	.w6(32'h3a96d493),
	.w7(32'h3a9860cf),
	.w8(32'h3a60c58a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f62c0),
	.w1(32'h3935d405),
	.w2(32'h3a4d82ee),
	.w3(32'h3a51f07b),
	.w4(32'h3a512d45),
	.w5(32'h39b80f76),
	.w6(32'hb9b6e288),
	.w7(32'hb971c7ad),
	.w8(32'hb9eba2b4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f620e8),
	.w1(32'hb9845545),
	.w2(32'h39f390f0),
	.w3(32'h3a641e4b),
	.w4(32'hb9e2ec4b),
	.w5(32'hb90fceff),
	.w6(32'hba5a587a),
	.w7(32'h39f54f73),
	.w8(32'h38c6863c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a41729),
	.w1(32'h3987a941),
	.w2(32'hba45c021),
	.w3(32'hb8f782a3),
	.w4(32'h36f31198),
	.w5(32'hb96fbd93),
	.w6(32'h3a62e372),
	.w7(32'h39b82b99),
	.w8(32'h393f7d54),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9949853),
	.w1(32'h39ede0b5),
	.w2(32'h3a03da73),
	.w3(32'hb913d076),
	.w4(32'h39133e74),
	.w5(32'h39c048dd),
	.w6(32'h3a4540bc),
	.w7(32'h3a832e89),
	.w8(32'h398009b0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d5e21d),
	.w1(32'h3a92f95c),
	.w2(32'h3a74533a),
	.w3(32'hb7af626b),
	.w4(32'h3a912844),
	.w5(32'h3a48b57f),
	.w6(32'h3a92e98f),
	.w7(32'h3a93ba08),
	.w8(32'h3a27165a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995646b),
	.w1(32'hb9f7b5c2),
	.w2(32'h3abaca87),
	.w3(32'h3a239ce0),
	.w4(32'h3ac58788),
	.w5(32'h3b0ef54f),
	.w6(32'hba3f339c),
	.w7(32'hba79aadf),
	.w8(32'hbabbc7a6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f4e7a),
	.w1(32'h3a96ba85),
	.w2(32'h3abec7ce),
	.w3(32'h3b1649ad),
	.w4(32'h3a9ee545),
	.w5(32'h3a6f07a3),
	.w6(32'h3ae7f4e8),
	.w7(32'h3ae8f636),
	.w8(32'h3b0299dc),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad65732),
	.w1(32'h3a40edef),
	.w2(32'h3a699abf),
	.w3(32'h3a4f6811),
	.w4(32'h3a827c9c),
	.w5(32'h3ac64775),
	.w6(32'h3ab4fc37),
	.w7(32'h3aef317d),
	.w8(32'h3a43a345),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39763599),
	.w1(32'hba4d8241),
	.w2(32'h3a2eacb9),
	.w3(32'h3a9ee0f0),
	.w4(32'h3c2d50ea),
	.w5(32'h3c2d7890),
	.w6(32'hbbbd63d9),
	.w7(32'hbc015d30),
	.w8(32'hbb00b231),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95f813),
	.w1(32'h3a17e212),
	.w2(32'hbacfd30c),
	.w3(32'hbb0de671),
	.w4(32'hbaa0eb00),
	.w5(32'hbb888ed4),
	.w6(32'h3b6e4ba9),
	.w7(32'h3961d8ac),
	.w8(32'h3b85f995),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule