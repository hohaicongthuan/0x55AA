module layer_10_featuremap_275(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40773a),
	.w1(32'h39a2b799),
	.w2(32'h39c1412c),
	.w3(32'h39a8cf9d),
	.w4(32'h39c6cb48),
	.w5(32'hb83a38c3),
	.w6(32'h3947a230),
	.w7(32'h393949f9),
	.w8(32'hb9e33c55),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa50a89),
	.w1(32'hbb03a80b),
	.w2(32'hbb1e7d4a),
	.w3(32'hba5b53f9),
	.w4(32'hbab2fb2f),
	.w5(32'hb9acff7f),
	.w6(32'hb9291c28),
	.w7(32'hba919862),
	.w8(32'hbaa38935),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39898c29),
	.w1(32'h38306260),
	.w2(32'hb79f6715),
	.w3(32'h3ac6a222),
	.w4(32'h3a87c4c1),
	.w5(32'h381a1812),
	.w6(32'h39dc76a8),
	.w7(32'hb79e26d3),
	.w8(32'h391793fc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35e9f5),
	.w1(32'h39b6bc62),
	.w2(32'h39bed95c),
	.w3(32'h3a048ccd),
	.w4(32'h399c2cf3),
	.w5(32'hba97856a),
	.w6(32'h39507024),
	.w7(32'hb94ec603),
	.w8(32'hbaaea8d6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb1446),
	.w1(32'hbaaea125),
	.w2(32'hbad2ee77),
	.w3(32'hbab1e892),
	.w4(32'hbad91e62),
	.w5(32'hb9fd67c2),
	.w6(32'hbaf92a6d),
	.w7(32'hbb0f71fa),
	.w8(32'hb9eb2127),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac6b00),
	.w1(32'hb9e03489),
	.w2(32'hba213d76),
	.w3(32'hba09ce7e),
	.w4(32'hba36648f),
	.w5(32'hb952dc78),
	.w6(32'hb9e52c68),
	.w7(32'hba0ee3ab),
	.w8(32'hb9924b7f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a507673),
	.w1(32'h3b457873),
	.w2(32'h3b41a460),
	.w3(32'h3a9d7c22),
	.w4(32'h3b882a4f),
	.w5(32'h3bdaff81),
	.w6(32'hba04bbcc),
	.w7(32'h3b4207f1),
	.w8(32'h3be080b4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a799f),
	.w1(32'h3b680259),
	.w2(32'h3b19a277),
	.w3(32'h3a5642fe),
	.w4(32'hbb2cb83c),
	.w5(32'hbbafc401),
	.w6(32'hba06a064),
	.w7(32'hbaa4c28e),
	.w8(32'hbbdb9825),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af3aa3),
	.w1(32'h39caf83a),
	.w2(32'h39807509),
	.w3(32'h39c9fb31),
	.w4(32'h38348bcd),
	.w5(32'hb9ce64f8),
	.w6(32'h3a329c26),
	.w7(32'h39ea4347),
	.w8(32'hb9982f9d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0eec78),
	.w1(32'hba960e9e),
	.w2(32'hba380416),
	.w3(32'hba960c42),
	.w4(32'hba882b14),
	.w5(32'hb99671bc),
	.w6(32'hba7157b0),
	.w7(32'hb8f364eb),
	.w8(32'hb8fa912e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba753195),
	.w1(32'hba4d910d),
	.w2(32'hba5cfa25),
	.w3(32'hba8a1a57),
	.w4(32'hba83ca07),
	.w5(32'hba3cd9d6),
	.w6(32'hba7204eb),
	.w7(32'hba75ece0),
	.w8(32'hb904f850),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fec57),
	.w1(32'h3aed14c6),
	.w2(32'h3b09c2bd),
	.w3(32'h3a33678e),
	.w4(32'h3b030dbf),
	.w5(32'h3b8cf608),
	.w6(32'hbadf8f7d),
	.w7(32'h3a107a5f),
	.w8(32'h3bb550d0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e90d9d),
	.w1(32'h39c5f664),
	.w2(32'h3ab4c4c6),
	.w3(32'hb92693dc),
	.w4(32'h3a354834),
	.w5(32'h3b13e2a9),
	.w6(32'hba0daede),
	.w7(32'h3a54c2b9),
	.w8(32'h3b26e392),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38407c12),
	.w1(32'h3a7e65de),
	.w2(32'h3aee1680),
	.w3(32'hba88a65b),
	.w4(32'h397e5a4e),
	.w5(32'hba87fb79),
	.w6(32'hba4ed331),
	.w7(32'h39a35d76),
	.w8(32'hba9610d0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba876488),
	.w1(32'hbaeaa8f7),
	.w2(32'hbb3e7b4f),
	.w3(32'hbaec8a9e),
	.w4(32'hbb08affb),
	.w5(32'hbb03b668),
	.w6(32'hba6e0f2a),
	.w7(32'hbad87aa1),
	.w8(32'hbaa142f8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9479bc),
	.w1(32'hbb9350a1),
	.w2(32'hbbc0d2e3),
	.w3(32'hbb8867c6),
	.w4(32'hbbd6f55e),
	.w5(32'hbbabebe3),
	.w6(32'hbb26ba7b),
	.w7(32'hbbbd5c01),
	.w8(32'hbbbaf738),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fbf136),
	.w1(32'h39482d92),
	.w2(32'h39187dec),
	.w3(32'h394a0fe4),
	.w4(32'h3702f80b),
	.w5(32'hb9491f8f),
	.w6(32'h3a282461),
	.w7(32'h39cecbf1),
	.w8(32'hb9b2d44c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9ad0e),
	.w1(32'hbada3cdc),
	.w2(32'hb9d84ab4),
	.w3(32'hb9345023),
	.w4(32'hbb7029bb),
	.w5(32'hb9dd0f88),
	.w6(32'hbaaf4558),
	.w7(32'h39a3fbe7),
	.w8(32'hba235bbc),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a1098),
	.w1(32'hba0dba84),
	.w2(32'h39c7db0e),
	.w3(32'hba419eda),
	.w4(32'hba99480a),
	.w5(32'h3b08d142),
	.w6(32'hbabbceb3),
	.w7(32'hba1dd9f4),
	.w8(32'h3b329034),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeda1e3),
	.w1(32'h3aaac228),
	.w2(32'h39a9d358),
	.w3(32'h39e22b0d),
	.w4(32'hb950b47d),
	.w5(32'h3a5b4355),
	.w6(32'h3a9df89a),
	.w7(32'h3a132705),
	.w8(32'h3aaef31c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbf25c),
	.w1(32'h3a845ec4),
	.w2(32'h3995deb1),
	.w3(32'h39c3180d),
	.w4(32'hb9c9b980),
	.w5(32'h3a5c76ce),
	.w6(32'h3a46f1ef),
	.w7(32'hb8d9f45a),
	.w8(32'h3a49bce4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95ec6d),
	.w1(32'h39c4c982),
	.w2(32'h39a6e3d1),
	.w3(32'h3a7bf305),
	.w4(32'h3a06558e),
	.w5(32'h3808a799),
	.w6(32'h3aa2f1c4),
	.w7(32'h3a51a040),
	.w8(32'h393936e6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf9ad7),
	.w1(32'hbb6bd379),
	.w2(32'hbaf5b850),
	.w3(32'hb8ae31e9),
	.w4(32'hba27e9a8),
	.w5(32'hba95756b),
	.w6(32'hba3fb972),
	.w7(32'h3b2b30d7),
	.w8(32'h3b03b045),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bdf74),
	.w1(32'hba99c943),
	.w2(32'hbaedc219),
	.w3(32'hbaa1df30),
	.w4(32'hbaf0d347),
	.w5(32'h3a65d821),
	.w6(32'hba1f3019),
	.w7(32'hba910ada),
	.w8(32'h3a201f6c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a7979),
	.w1(32'hb9482314),
	.w2(32'hba30eb5d),
	.w3(32'h3ab05a14),
	.w4(32'hba8ef57d),
	.w5(32'hbb8eba35),
	.w6(32'h3b4a6a7c),
	.w7(32'h3a80bb6e),
	.w8(32'hbb795d11),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef7fee),
	.w1(32'hb7aa7df9),
	.w2(32'hb8f0468b),
	.w3(32'hb71cf019),
	.w4(32'h37cd327a),
	.w5(32'h39bd8c04),
	.w6(32'h39e0a200),
	.w7(32'h398feb1c),
	.w8(32'h3a73b811),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2582f9),
	.w1(32'h3a4be50a),
	.w2(32'h3a88ba75),
	.w3(32'h3a383db7),
	.w4(32'h3a8cac8e),
	.w5(32'h390a6c1e),
	.w6(32'h3aacb725),
	.w7(32'h3aad6f92),
	.w8(32'h39099ec7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcee4b2),
	.w1(32'h3b88a9cb),
	.w2(32'h3b8463ed),
	.w3(32'h3b0dadd0),
	.w4(32'h3a84c85f),
	.w5(32'h3bd9b576),
	.w6(32'h39dfcac1),
	.w7(32'h3b057cd7),
	.w8(32'h3ba93c9c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f8277),
	.w1(32'h3b22f8b6),
	.w2(32'h3b084809),
	.w3(32'h3afeffde),
	.w4(32'h3af79098),
	.w5(32'hba8f6b0a),
	.w6(32'h3b22710d),
	.w7(32'h3b1dbf12),
	.w8(32'hba917e36),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd987a),
	.w1(32'h39a4c480),
	.w2(32'h3ab155c3),
	.w3(32'h3a7a8c25),
	.w4(32'h3a78af15),
	.w5(32'h3a24f2b9),
	.w6(32'h39f56573),
	.w7(32'h38d13ef1),
	.w8(32'hb920c8f1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88189bf),
	.w1(32'hb8863177),
	.w2(32'h39641ece),
	.w3(32'hbb06ebc2),
	.w4(32'hbaa9b39d),
	.w5(32'h3a56b155),
	.w6(32'hba69e24a),
	.w7(32'hba054d28),
	.w8(32'hb9f8cb85),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba474e9c),
	.w1(32'hb990db37),
	.w2(32'hb8e2a3be),
	.w3(32'h3a9a018a),
	.w4(32'h3aaade7d),
	.w5(32'hba715e2a),
	.w6(32'hb691bd8d),
	.w7(32'h399ad17d),
	.w8(32'hb9a70302),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3f493),
	.w1(32'hb9cd9288),
	.w2(32'h388f8d42),
	.w3(32'hba9f79bf),
	.w4(32'hbace790f),
	.w5(32'hb9dbf1b1),
	.w6(32'hba451e9d),
	.w7(32'hb9174a7b),
	.w8(32'hb9c36723),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab5ada),
	.w1(32'hb9fdb836),
	.w2(32'hba4351a5),
	.w3(32'hba3f3497),
	.w4(32'hba07fb66),
	.w5(32'hbb0a4437),
	.w6(32'hb9d2df2e),
	.w7(32'hb909b981),
	.w8(32'hbae49098),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d6e23),
	.w1(32'hb9478415),
	.w2(32'hb9becb08),
	.w3(32'hba1cc138),
	.w4(32'hb99b2804),
	.w5(32'h39c95845),
	.w6(32'hba16f9af),
	.w7(32'hb9b3ccea),
	.w8(32'h39daccdd),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b74d07),
	.w1(32'h3a3135a9),
	.w2(32'hb9a2521e),
	.w3(32'h3a646082),
	.w4(32'h3a07ed6b),
	.w5(32'hba30cd45),
	.w6(32'h39d8d7b8),
	.w7(32'hb8221760),
	.w8(32'hba2dfb2a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd7e73),
	.w1(32'hbbbac59a),
	.w2(32'hbbf7e7eb),
	.w3(32'hbb3b4e7f),
	.w4(32'hbc4d5975),
	.w5(32'hbc3a8d57),
	.w6(32'hbbf80741),
	.w7(32'hbc126505),
	.w8(32'hbbf69b2f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76353c),
	.w1(32'hba7b8db9),
	.w2(32'hbb382317),
	.w3(32'h3b14a3a1),
	.w4(32'hb9af9a6b),
	.w5(32'hbb8339da),
	.w6(32'h3bc78704),
	.w7(32'h3b20d99e),
	.w8(32'hbb268788),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1505ec),
	.w1(32'h3b9fb32f),
	.w2(32'h3bd26d07),
	.w3(32'h3c01e88c),
	.w4(32'h3c0128af),
	.w5(32'h3bf45aee),
	.w6(32'h3beb5218),
	.w7(32'h3bdae1bb),
	.w8(32'h3bafa707),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390fb38d),
	.w1(32'hbacb0780),
	.w2(32'hbb00841e),
	.w3(32'hba96bbee),
	.w4(32'hbae783b6),
	.w5(32'hba846b97),
	.w6(32'hb9eb84e6),
	.w7(32'hbaa6e4aa),
	.w8(32'hb94093a8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a7896),
	.w1(32'h3ab4c611),
	.w2(32'h3adfacc8),
	.w3(32'h3a96d712),
	.w4(32'h3acda09c),
	.w5(32'h399eeee7),
	.w6(32'h3adb9930),
	.w7(32'h3b03e8b0),
	.w8(32'h39789aa8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb876490f),
	.w1(32'h38f78784),
	.w2(32'h38c5e089),
	.w3(32'h3a02e4e0),
	.w4(32'h39e75e23),
	.w5(32'hba1b5a16),
	.w6(32'h39e68cf6),
	.w7(32'h39c0e2e4),
	.w8(32'hb8a21a48),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f2d3c8),
	.w1(32'hb9a4dd5f),
	.w2(32'hb9a9cdb3),
	.w3(32'hb9ccdbea),
	.w4(32'hba07d56c),
	.w5(32'hbb10b013),
	.w6(32'hb73d6a99),
	.w7(32'hb9da9ade),
	.w8(32'hbb01ca63),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3e9df),
	.w1(32'h3adc45dc),
	.w2(32'hb823051e),
	.w3(32'hba3628d8),
	.w4(32'h3a61b808),
	.w5(32'h3b125a86),
	.w6(32'hbad84199),
	.w7(32'h3a99352c),
	.w8(32'h3b4b833a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7d56e),
	.w1(32'hba0094ae),
	.w2(32'h38320d6f),
	.w3(32'hba4d1e60),
	.w4(32'hba7c0306),
	.w5(32'hba402899),
	.w6(32'h3a78830e),
	.w7(32'h38a0ed9c),
	.w8(32'hb8ddafba),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d17a8),
	.w1(32'hba44d985),
	.w2(32'h38542c61),
	.w3(32'hba6c8e5f),
	.w4(32'hba2db298),
	.w5(32'hbaad041c),
	.w6(32'hb97249b4),
	.w7(32'h37aac381),
	.w8(32'hba2e3e03),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a2f13),
	.w1(32'hba40a7b0),
	.w2(32'hba98aaa4),
	.w3(32'hba277039),
	.w4(32'hba8f0c47),
	.w5(32'hb9af1569),
	.w6(32'h3a88268a),
	.w7(32'h3a75346a),
	.w8(32'h3a62c774),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddb971),
	.w1(32'h39e632ab),
	.w2(32'h3b810b16),
	.w3(32'h3b06e5b4),
	.w4(32'h3ac4a4f6),
	.w5(32'h3b574690),
	.w6(32'hba54b03c),
	.w7(32'h3b2a8b27),
	.w8(32'h3b7a05b8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b87d8),
	.w1(32'h3a118404),
	.w2(32'h39262184),
	.w3(32'h3a14e206),
	.w4(32'h39c58fdd),
	.w5(32'h3a1fe82d),
	.w6(32'h39f3307f),
	.w7(32'h39435f20),
	.w8(32'h3a07f453),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49da58),
	.w1(32'h39f6fe8b),
	.w2(32'h3a3ec520),
	.w3(32'h3a089b79),
	.w4(32'h3a1c281c),
	.w5(32'h3a9b01ed),
	.w6(32'h39e332f3),
	.w7(32'h3a032bb3),
	.w8(32'h3a56415e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6069e0),
	.w1(32'h3a034a99),
	.w2(32'hb9e7d826),
	.w3(32'h3a42115b),
	.w4(32'hb9c6d5de),
	.w5(32'hba131609),
	.w6(32'h39875438),
	.w7(32'hb94e9a7c),
	.w8(32'hb9889547),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6c71a),
	.w1(32'hb9a87fe0),
	.w2(32'hba8583c0),
	.w3(32'hba347b5b),
	.w4(32'hb9d82e31),
	.w5(32'h3b14901a),
	.w6(32'h387480f1),
	.w7(32'h3a0cc9cf),
	.w8(32'h3b282fb9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39961cde),
	.w1(32'h3a81b75d),
	.w2(32'h3a89698d),
	.w3(32'h3ae79842),
	.w4(32'h3ad02884),
	.w5(32'hba8771b3),
	.w6(32'h3afb2b1e),
	.w7(32'h3af3cfb0),
	.w8(32'hbaa287bd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d0879),
	.w1(32'hbab04606),
	.w2(32'h39831532),
	.w3(32'h3a3a0bc9),
	.w4(32'hbab71eb4),
	.w5(32'h3b3b49f3),
	.w6(32'hbb524e16),
	.w7(32'hba3823e4),
	.w8(32'h3b846467),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27d179),
	.w1(32'h3b380b8a),
	.w2(32'h3afd1741),
	.w3(32'h3aa6e870),
	.w4(32'h3a7a5c0c),
	.w5(32'h3982c45d),
	.w6(32'h3b26dbf9),
	.w7(32'h3af47d12),
	.w8(32'hba1270d8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8a4c7),
	.w1(32'hba1c2b99),
	.w2(32'hb99fd4da),
	.w3(32'h3a38c110),
	.w4(32'h3a6a06f7),
	.w5(32'hb781266d),
	.w6(32'h398f5a8d),
	.w7(32'h39d28245),
	.w8(32'h39197946),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392ae8d6),
	.w1(32'h3a50a9a2),
	.w2(32'h3aa83183),
	.w3(32'h3a819a5b),
	.w4(32'h3ac8119e),
	.w5(32'hb9342a23),
	.w6(32'h3a8e404d),
	.w7(32'h3ae2d5ef),
	.w8(32'h39dc050b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a754843),
	.w1(32'h39849346),
	.w2(32'h36e8fbfc),
	.w3(32'hb9b4e6cb),
	.w4(32'hba163d3f),
	.w5(32'h3a365b8c),
	.w6(32'h3a2a2222),
	.w7(32'hb971d3c1),
	.w8(32'h3a36cc88),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ccf76),
	.w1(32'h39cb435c),
	.w2(32'h3a16e63c),
	.w3(32'h39c7c696),
	.w4(32'h39b539c1),
	.w5(32'h3920860a),
	.w6(32'h39de96b2),
	.w7(32'h39aba160),
	.w8(32'hb98f949d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba180e15),
	.w1(32'hb919d10e),
	.w2(32'h3a07ac5f),
	.w3(32'h3a34f088),
	.w4(32'h3abb4997),
	.w5(32'hb7bcf9b3),
	.w6(32'hb9636d90),
	.w7(32'h3aa186eb),
	.w8(32'hb88f15ba),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa886ec),
	.w1(32'hbab07156),
	.w2(32'hb9bfa116),
	.w3(32'hba77459c),
	.w4(32'hba35d48b),
	.w5(32'h3a167ee9),
	.w6(32'hbaf00728),
	.w7(32'hba3f2eb0),
	.w8(32'h3a51e7e9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a2704),
	.w1(32'hb9324b17),
	.w2(32'hbaa790d3),
	.w3(32'hbab3205e),
	.w4(32'hbac7f76c),
	.w5(32'hbac94c5f),
	.w6(32'hb938ee89),
	.w7(32'hb96935c4),
	.w8(32'hba785f1a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f52ef),
	.w1(32'hb7eb1466),
	.w2(32'hba355f4b),
	.w3(32'hba4c450e),
	.w4(32'hba19bdf7),
	.w5(32'hba1edc15),
	.w6(32'hba016cfb),
	.w7(32'hba71c158),
	.w8(32'hb9a29cc6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f8180),
	.w1(32'hb9413459),
	.w2(32'hb7c78df9),
	.w3(32'hb97a80c9),
	.w4(32'h389a37c8),
	.w5(32'hba21e3b6),
	.w6(32'h395103a5),
	.w7(32'h39473589),
	.w8(32'hb82ade61),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b49412),
	.w1(32'h38963d92),
	.w2(32'h3a0781f3),
	.w3(32'hba0af010),
	.w4(32'h39f90697),
	.w5(32'h3ae85be0),
	.w6(32'hb8a9f549),
	.w7(32'h3a0f6356),
	.w8(32'h3b36dade),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2890fe),
	.w1(32'h3b53c378),
	.w2(32'h3b250add),
	.w3(32'h3b0d6742),
	.w4(32'h3b092179),
	.w5(32'h37dd6141),
	.w6(32'h3b6e19ca),
	.w7(32'h3b4bdabe),
	.w8(32'hb8e42886),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe927f5),
	.w1(32'hbb9cbee3),
	.w2(32'hbbdaae27),
	.w3(32'hbaf1e4d7),
	.w4(32'hbba7ef36),
	.w5(32'hbb0a699c),
	.w6(32'hbb9b35f9),
	.w7(32'hbb582ce5),
	.w8(32'hbb234151),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe43ddf),
	.w1(32'hbb75baa8),
	.w2(32'h3a24ab86),
	.w3(32'hbb976358),
	.w4(32'hbbb03c2b),
	.w5(32'hbb5ff03b),
	.w6(32'hbb62ec68),
	.w7(32'hbb39acdd),
	.w8(32'hbb99e59c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395186d7),
	.w1(32'h39e01dc0),
	.w2(32'h39276a76),
	.w3(32'hba871365),
	.w4(32'hb98ab7d2),
	.w5(32'hbb48d172),
	.w6(32'h39195eaa),
	.w7(32'h3b2ed961),
	.w8(32'hbaa5cb34),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964695f),
	.w1(32'hbaf5a3c5),
	.w2(32'hba49b093),
	.w3(32'hbadc25c4),
	.w4(32'hbb19a878),
	.w5(32'hbaff06ef),
	.w6(32'h3b2b90a8),
	.w7(32'h39d22ad6),
	.w8(32'h37e695d3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd3d0f),
	.w1(32'h3a0874ab),
	.w2(32'h39be1c4a),
	.w3(32'h38f4f298),
	.w4(32'h38df7878),
	.w5(32'h39b4332d),
	.w6(32'h3a3faf90),
	.w7(32'h39d93e18),
	.w8(32'h3a00120a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e78aa5),
	.w1(32'hb93adb6c),
	.w2(32'hba058c7f),
	.w3(32'h390447f2),
	.w4(32'hb921a435),
	.w5(32'h394943fe),
	.w6(32'h389b7c09),
	.w7(32'hb9ec24d0),
	.w8(32'h379db73e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26a654),
	.w1(32'hba83e209),
	.w2(32'hba696f89),
	.w3(32'h3a0c74e7),
	.w4(32'h3a1b5eb6),
	.w5(32'hba26220d),
	.w6(32'h392d0420),
	.w7(32'h387e7702),
	.w8(32'hb9f131c4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba760794),
	.w1(32'hba74eba1),
	.w2(32'hba6c8682),
	.w3(32'hbaa29a4d),
	.w4(32'hba8649ba),
	.w5(32'h38ca6b16),
	.w6(32'hbac50971),
	.w7(32'hbaad8c35),
	.w8(32'hb81a8491),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fc49a1),
	.w1(32'hb9e6b1ff),
	.w2(32'hb9dabf13),
	.w3(32'hb9fc3905),
	.w4(32'hb9f4079c),
	.w5(32'hb7b9dc75),
	.w6(32'hb984bb2e),
	.w7(32'hb983a218),
	.w8(32'hb99734b9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40ab98),
	.w1(32'hbae10fc0),
	.w2(32'hba8107ce),
	.w3(32'h38bb79af),
	.w4(32'hba7e08c1),
	.w5(32'hb7c2c4e9),
	.w6(32'hbac194c5),
	.w7(32'h38db94dd),
	.w8(32'h3ab43c6f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55a0b6),
	.w1(32'hba24d972),
	.w2(32'h3a86513e),
	.w3(32'h3a84db94),
	.w4(32'hb9ddb3b8),
	.w5(32'hbafd6e58),
	.w6(32'hba956c4b),
	.w7(32'hb9db2ab8),
	.w8(32'hbae6178a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba510ff9),
	.w1(32'hbaa7e621),
	.w2(32'hbace1b8e),
	.w3(32'hbb059577),
	.w4(32'hbb0f5aac),
	.w5(32'hbb31be80),
	.w6(32'hb7212d9e),
	.w7(32'hba3eb3e0),
	.w8(32'hba9e2c10),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0debea),
	.w1(32'hba0474b5),
	.w2(32'hba87b5f6),
	.w3(32'hba2fb2ec),
	.w4(32'hba8f364f),
	.w5(32'hbb043cfa),
	.w6(32'hba4d8bd2),
	.w7(32'hb9751a63),
	.w8(32'hbb05553a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c484f),
	.w1(32'hbb07f767),
	.w2(32'hbabd1975),
	.w3(32'hba4f3402),
	.w4(32'hbb25bfec),
	.w5(32'hb9822ca0),
	.w6(32'hbaab6752),
	.w7(32'hba4a4f5a),
	.w8(32'h39992ed1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8745ad),
	.w1(32'h3aab269a),
	.w2(32'h3ad350e5),
	.w3(32'h39f8d633),
	.w4(32'h3a96cdb7),
	.w5(32'h391d93a2),
	.w6(32'h3a963371),
	.w7(32'h3adbd664),
	.w8(32'h3a12a539),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa65b6a),
	.w1(32'hb9dbb5f8),
	.w2(32'h39f0d90c),
	.w3(32'h36a59974),
	.w4(32'h39e9dacc),
	.w5(32'h3afa47bc),
	.w6(32'hba8dd736),
	.w7(32'h38c433bb),
	.w8(32'h3a881b21),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fcc08),
	.w1(32'hb996cac5),
	.w2(32'h3a9256fc),
	.w3(32'h39067e34),
	.w4(32'h39821dcd),
	.w5(32'h38c5bfe9),
	.w6(32'h381b1183),
	.w7(32'h39ce6fd3),
	.w8(32'h39838d34),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d1ea07),
	.w1(32'hba246bb9),
	.w2(32'hba089446),
	.w3(32'hba30ac8d),
	.w4(32'hb9dfb229),
	.w5(32'h3b12a126),
	.w6(32'hba03b82b),
	.w7(32'hba0f127f),
	.w8(32'h3a7da7bf),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b58d5),
	.w1(32'hba2e73d7),
	.w2(32'hba2a6833),
	.w3(32'h3adb87d4),
	.w4(32'h39d6664d),
	.w5(32'hb8e7e9ae),
	.w6(32'h3a4cb4a8),
	.w7(32'hba1ed2dd),
	.w8(32'hb9fc7e7d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a523953),
	.w1(32'h3a5d0635),
	.w2(32'h3a2a8c91),
	.w3(32'h3a8e8957),
	.w4(32'h3aae56d9),
	.w5(32'h38e6726a),
	.w6(32'h3a8e3975),
	.w7(32'h3ac4314c),
	.w8(32'h392a351f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabac739),
	.w1(32'hbaefe530),
	.w2(32'hbad4c588),
	.w3(32'hbacce9ce),
	.w4(32'hbaee7d2d),
	.w5(32'hbb3a640a),
	.w6(32'h3915e5dd),
	.w7(32'hbad514f0),
	.w8(32'hbadaa7af),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a335523),
	.w1(32'h39a35b20),
	.w2(32'h392f5349),
	.w3(32'h391328cd),
	.w4(32'hb95c337a),
	.w5(32'hb9c875d8),
	.w6(32'h3921d60c),
	.w7(32'hb915d483),
	.w8(32'hb8fd9536),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6cce8e),
	.w1(32'hba5de2ae),
	.w2(32'hb9c773e1),
	.w3(32'hba990c6e),
	.w4(32'hbb1294ab),
	.w5(32'hbabbf753),
	.w6(32'h39b63309),
	.w7(32'hba9d22fd),
	.w8(32'hbaeace23),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd396e),
	.w1(32'hba675b9a),
	.w2(32'h39487cff),
	.w3(32'h3984d622),
	.w4(32'h39509468),
	.w5(32'h39c3d5f0),
	.w6(32'hba9741b7),
	.w7(32'h3ae608a9),
	.w8(32'h3adfcabe),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba43755),
	.w1(32'h3b605a86),
	.w2(32'h3b29b29a),
	.w3(32'h3b5e85cf),
	.w4(32'h3b422a1b),
	.w5(32'h3b629f17),
	.w6(32'h3b2c7dd3),
	.w7(32'h3b4033ee),
	.w8(32'h3b83bb0a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1dc96),
	.w1(32'hbbadc1e4),
	.w2(32'hbb1ecb78),
	.w3(32'hbb94b193),
	.w4(32'hbbc8097c),
	.w5(32'hbb6a47d3),
	.w6(32'hbb93f16a),
	.w7(32'hbb90ebe2),
	.w8(32'hbb8093db),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39ba35),
	.w1(32'h3add620c),
	.w2(32'h3a42684f),
	.w3(32'h3b49f91f),
	.w4(32'h3b6f32a2),
	.w5(32'h3a18e0d4),
	.w6(32'h3b76cd09),
	.w7(32'h3b6b2020),
	.w8(32'h3ae8d241),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eae52),
	.w1(32'hbb36f97a),
	.w2(32'hbb9abd25),
	.w3(32'hbbc554e9),
	.w4(32'hbbe66988),
	.w5(32'hbbd23b76),
	.w6(32'hbba37537),
	.w7(32'hbbb3d3c4),
	.w8(32'hbbdd7611),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa991ca),
	.w1(32'hbb13fe81),
	.w2(32'hbb285043),
	.w3(32'hbb229d33),
	.w4(32'hbb5921cf),
	.w5(32'hbb091566),
	.w6(32'h39789944),
	.w7(32'hbaccd1a9),
	.w8(32'hbb44e12a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29beea),
	.w1(32'h389211ab),
	.w2(32'hb9ec1a59),
	.w3(32'h3b203618),
	.w4(32'h3a925ade),
	.w5(32'h3a186ba7),
	.w6(32'h3abfbe0b),
	.w7(32'hb97738a5),
	.w8(32'hb9145a1d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae7e1e),
	.w1(32'h3a664933),
	.w2(32'h3a676881),
	.w3(32'h3a86decb),
	.w4(32'h3a88696f),
	.w5(32'hbaf10bed),
	.w6(32'h3a4e2e64),
	.w7(32'h3a6cc525),
	.w8(32'hbaac2976),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21822f),
	.w1(32'hba929eac),
	.w2(32'h388e9ad4),
	.w3(32'hba8cec1e),
	.w4(32'hbaa1acf0),
	.w5(32'hb903543d),
	.w6(32'hbaa78502),
	.w7(32'h39dac4b0),
	.w8(32'h3a81c805),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc0ab4),
	.w1(32'hb9837035),
	.w2(32'h3af11b65),
	.w3(32'hbad2ab18),
	.w4(32'hba48156c),
	.w5(32'hbb57c413),
	.w6(32'hbab2d49a),
	.w7(32'h3b07c20b),
	.w8(32'hba88e467),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbbaa1),
	.w1(32'hbc30b124),
	.w2(32'hbc2ac5fa),
	.w3(32'hbc02edbf),
	.w4(32'hbc628676),
	.w5(32'hbc24f23a),
	.w6(32'hbc299039),
	.w7(32'hbc4198bb),
	.w8(32'hbc1a8715),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94ec4f),
	.w1(32'h3adc4ffe),
	.w2(32'hbb354330),
	.w3(32'h3b4495d9),
	.w4(32'hb98cc8f5),
	.w5(32'hbbaffe23),
	.w6(32'h3b8e4b7d),
	.w7(32'hb94dc1d0),
	.w8(32'hbb840061),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39640506),
	.w1(32'hba0a6fee),
	.w2(32'hba48ebb9),
	.w3(32'hba99a02d),
	.w4(32'hbb3110ca),
	.w5(32'hbb0e3005),
	.w6(32'hb909ef6f),
	.w7(32'hba9ff047),
	.w8(32'hbb36e085),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb72d71),
	.w1(32'hbaaf1ff9),
	.w2(32'hba846dde),
	.w3(32'hbb3c178c),
	.w4(32'hbb006117),
	.w5(32'hbb701c37),
	.w6(32'hbbbec5d6),
	.w7(32'hbb0e3526),
	.w8(32'hbb29e859),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f2376),
	.w1(32'hba662ed0),
	.w2(32'hbb009f87),
	.w3(32'hba161398),
	.w4(32'hbae71270),
	.w5(32'h3acf1ecf),
	.w6(32'hba8930c6),
	.w7(32'hbafb0bb9),
	.w8(32'h3aba3338),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdaba61),
	.w1(32'hbbbd3ff0),
	.w2(32'hbb5d4ed0),
	.w3(32'hbab5696a),
	.w4(32'hbba0d8bf),
	.w5(32'hbb660cc6),
	.w6(32'hbb8f8c2c),
	.w7(32'hbbcca433),
	.w8(32'hbb3f65c9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9027c),
	.w1(32'h3b0ca7a5),
	.w2(32'h3b5c2e4d),
	.w3(32'h3b08539b),
	.w4(32'h3b8f0dd0),
	.w5(32'h3b2eb6c2),
	.w6(32'h3a630e13),
	.w7(32'h3b47ddd5),
	.w8(32'h3b6ea3c4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6cfcb),
	.w1(32'hbaa37437),
	.w2(32'hbb333bdb),
	.w3(32'hbaffb8e9),
	.w4(32'hbae2c766),
	.w5(32'hba5f7792),
	.w6(32'hbad1eebe),
	.w7(32'hbad8f0a1),
	.w8(32'hbac5e184),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5963a),
	.w1(32'hba328aef),
	.w2(32'hbaba6f66),
	.w3(32'hbae33aaa),
	.w4(32'hbaed5ce6),
	.w5(32'hbaf8b679),
	.w6(32'hba43d92a),
	.w7(32'hbb0cba1b),
	.w8(32'hbaf86b26),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44209a),
	.w1(32'hba6e686e),
	.w2(32'h3adcb7ea),
	.w3(32'hbac84b60),
	.w4(32'h3a2f3997),
	.w5(32'hb9f2cfd4),
	.w6(32'hbaeb2a76),
	.w7(32'h3a8c8124),
	.w8(32'hb9f7ecb6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbf2d2),
	.w1(32'hb99d4a08),
	.w2(32'hb931b194),
	.w3(32'hb94c8199),
	.w4(32'hb98c207f),
	.w5(32'hba1338fc),
	.w6(32'h39b447bc),
	.w7(32'hb9f3d4c4),
	.w8(32'hb98212f9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9332b5),
	.w1(32'h3b808f0c),
	.w2(32'h3b75a3da),
	.w3(32'h3b7c1dba),
	.w4(32'h3bb1aea6),
	.w5(32'h3b88bb02),
	.w6(32'h3b894d04),
	.w7(32'h3b9d50ae),
	.w8(32'h3ba8c334),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f87a2),
	.w1(32'h39f9caa6),
	.w2(32'hb9514dbf),
	.w3(32'hb7ad2a4b),
	.w4(32'h39a19de2),
	.w5(32'hba98d046),
	.w6(32'h3a3fa470),
	.w7(32'h3a7496b6),
	.w8(32'hba2dd3b1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0abf8a),
	.w1(32'hba39589e),
	.w2(32'hb9e862ac),
	.w3(32'hbb274ba8),
	.w4(32'hbb93cb65),
	.w5(32'hbb9be9f7),
	.w6(32'h399501cd),
	.w7(32'hbb2ca395),
	.w8(32'hbb303de0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ca5e7),
	.w1(32'hbac16f0a),
	.w2(32'hbb1093a1),
	.w3(32'hbb179d63),
	.w4(32'hbb438b9b),
	.w5(32'hbbd8c3ca),
	.w6(32'hbb1043b7),
	.w7(32'hbb16ad91),
	.w8(32'hbbe87ea2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e5f67),
	.w1(32'hba4ae824),
	.w2(32'hba81ebfd),
	.w3(32'hba457994),
	.w4(32'hba7293de),
	.w5(32'hba9e2f81),
	.w6(32'h3a56299c),
	.w7(32'hb8dadfa2),
	.w8(32'hb9d6cba7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb829025b),
	.w1(32'hb98a6871),
	.w2(32'hb99fd450),
	.w3(32'hba297078),
	.w4(32'hb96dc66e),
	.w5(32'h3aa7dbca),
	.w6(32'hba18480f),
	.w7(32'h3762433c),
	.w8(32'h3aa3ddcd),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96e368),
	.w1(32'h3a338063),
	.w2(32'h3a2a5c41),
	.w3(32'h3a0b406c),
	.w4(32'h39973d5f),
	.w5(32'hba904c9a),
	.w6(32'h3a68336d),
	.w7(32'h3a475691),
	.w8(32'hba8956f2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdbcac),
	.w1(32'hba8f8f69),
	.w2(32'hba448660),
	.w3(32'hba428251),
	.w4(32'hbb12d48d),
	.w5(32'hbaa1b486),
	.w6(32'hb99bd0b1),
	.w7(32'hba5a5ae4),
	.w8(32'hbabc35c6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5cb3d),
	.w1(32'hbaf5ccb8),
	.w2(32'hba766c86),
	.w3(32'hbacea4e9),
	.w4(32'hba56ac9a),
	.w5(32'h3a989168),
	.w6(32'hbab1d302),
	.w7(32'hbaa09b01),
	.w8(32'h3a3a2093),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e7f6f),
	.w1(32'hb9fac372),
	.w2(32'h39da6916),
	.w3(32'hb92a7dce),
	.w4(32'h39500b1c),
	.w5(32'hbab7fa19),
	.w6(32'hba5de3d6),
	.w7(32'h39a49f85),
	.w8(32'hba238f89),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a321a49),
	.w1(32'h3a9dd66b),
	.w2(32'h3ae0709e),
	.w3(32'h396bfc83),
	.w4(32'h3a698cad),
	.w5(32'h39083335),
	.w6(32'hb9a23415),
	.w7(32'h3a9fdd58),
	.w8(32'hb8275279),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba110679),
	.w1(32'hb788a4c6),
	.w2(32'hb82167e2),
	.w3(32'h3a5c36b5),
	.w4(32'h3a1378ca),
	.w5(32'h3ac74ff8),
	.w6(32'h38d6e994),
	.w7(32'h39b37104),
	.w8(32'h3abab3ea),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f454ab),
	.w1(32'hbab837a2),
	.w2(32'hbb10e22b),
	.w3(32'hb9a97ac9),
	.w4(32'hba7cc0b9),
	.w5(32'hbb0937e5),
	.w6(32'h3a91a911),
	.w7(32'h37dfaf09),
	.w8(32'hbac9455e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea2cc9),
	.w1(32'h39289d4f),
	.w2(32'hb97d237e),
	.w3(32'h38127c56),
	.w4(32'h391d7462),
	.w5(32'h39cb3ca0),
	.w6(32'h37d2805f),
	.w7(32'hb98a9788),
	.w8(32'h38b65cc4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c6426),
	.w1(32'h3a4972c3),
	.w2(32'h3a07b986),
	.w3(32'h3894da07),
	.w4(32'h3995102b),
	.w5(32'hb7daa2a5),
	.w6(32'hb9509eee),
	.w7(32'h39b12841),
	.w8(32'hb97bbf89),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95af45),
	.w1(32'hb957328a),
	.w2(32'h3a37b814),
	.w3(32'h3a0af264),
	.w4(32'h3a728d30),
	.w5(32'h39272401),
	.w6(32'hb81477ce),
	.w7(32'h3a8904c8),
	.w8(32'h38aabb64),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d19df),
	.w1(32'hb868c0a0),
	.w2(32'hb9008ba3),
	.w3(32'hb8fea24e),
	.w4(32'hba0591c8),
	.w5(32'hb94ea6c3),
	.w6(32'h3a48bb7f),
	.w7(32'hb9870592),
	.w8(32'h391e1f92),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f8e75),
	.w1(32'h38ef9ad5),
	.w2(32'h3bf57023),
	.w3(32'hbb911fba),
	.w4(32'hbba186e2),
	.w5(32'hb923fb80),
	.w6(32'hbb80d65c),
	.w7(32'hbb226175),
	.w8(32'hbb9fda5c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb371713),
	.w1(32'hba0e099d),
	.w2(32'h3a5d069c),
	.w3(32'hb991eae0),
	.w4(32'hba34ce0f),
	.w5(32'h3a95252c),
	.w6(32'hbb2f933a),
	.w7(32'hba1f91a4),
	.w8(32'h3a64a25f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac336b),
	.w1(32'h391f3340),
	.w2(32'hb7dc2d65),
	.w3(32'h3936ef91),
	.w4(32'hba130605),
	.w5(32'hbacc19d3),
	.w6(32'h3a25d1e8),
	.w7(32'h3988fb4e),
	.w8(32'hba8092a5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89cb65),
	.w1(32'hb805cbe6),
	.w2(32'hba85dc45),
	.w3(32'hbaad9290),
	.w4(32'hbb08a1ba),
	.w5(32'h37a6ebb6),
	.w6(32'hba188eae),
	.w7(32'hba789305),
	.w8(32'hb9aafcad),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f9437),
	.w1(32'h3a001d0a),
	.w2(32'h390e3990),
	.w3(32'h3a02c670),
	.w4(32'hb8f3a6a0),
	.w5(32'hba999eb1),
	.w6(32'h3acaa20c),
	.w7(32'h3a08d5e8),
	.w8(32'hbb292fb4),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aa1ff),
	.w1(32'hbb8b7977),
	.w2(32'hbb731f31),
	.w3(32'hbb45287f),
	.w4(32'hbb52e1ec),
	.w5(32'hbb231d4f),
	.w6(32'hbb907806),
	.w7(32'hbb90264b),
	.w8(32'hbb449e49),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53fe4e),
	.w1(32'hbb10243b),
	.w2(32'hbb238402),
	.w3(32'hbb8768d2),
	.w4(32'hbb897f7c),
	.w5(32'hbb35d2be),
	.w6(32'hbb2b347d),
	.w7(32'hbb74aae9),
	.w8(32'hbb3b0954),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb500a2e),
	.w1(32'hba990bd0),
	.w2(32'h38aac06e),
	.w3(32'h39d8544d),
	.w4(32'hbaf8911d),
	.w5(32'h3b21c8ae),
	.w6(32'hba7d7a12),
	.w7(32'hb9cfdc6c),
	.w8(32'h3b2df4b3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58bb28),
	.w1(32'h39f9b7f2),
	.w2(32'h39fa786e),
	.w3(32'h3a52300c),
	.w4(32'h397d0036),
	.w5(32'hbb0f7432),
	.w6(32'h3b0fe873),
	.w7(32'h3a3f4fd5),
	.w8(32'hbb13d984),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cb89f),
	.w1(32'hbb01b968),
	.w2(32'hbae6104b),
	.w3(32'hbb4f16e0),
	.w4(32'hbb419806),
	.w5(32'hbb239b25),
	.w6(32'hbb20ccdd),
	.w7(32'hbb116501),
	.w8(32'hbb0e8274),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7d13e),
	.w1(32'hba93f687),
	.w2(32'hba36c8ea),
	.w3(32'hb7523680),
	.w4(32'hbaba529c),
	.w5(32'hb903803e),
	.w6(32'hbb58d973),
	.w7(32'hba830432),
	.w8(32'h3a643b5f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb106956),
	.w1(32'hbb060a56),
	.w2(32'hbad75259),
	.w3(32'hbb0bb8a2),
	.w4(32'hbb849317),
	.w5(32'hbb45ba3b),
	.w6(32'h393f0fe1),
	.w7(32'hbb32f2b2),
	.w8(32'hbb596548),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6407e1),
	.w1(32'hbae4fd30),
	.w2(32'hbad1b19b),
	.w3(32'hba9db596),
	.w4(32'hbb069296),
	.w5(32'hb9880c0f),
	.w6(32'hbaea6222),
	.w7(32'hba696db4),
	.w8(32'h39e72d83),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30f0c1),
	.w1(32'hb9a77b80),
	.w2(32'h3916ad4b),
	.w3(32'h3aa9031f),
	.w4(32'h3a8d8954),
	.w5(32'hba89f79a),
	.w6(32'h3a218b2b),
	.w7(32'h39ebe62f),
	.w8(32'hba83c350),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d110d),
	.w1(32'h3aeae457),
	.w2(32'h3a05a1c8),
	.w3(32'h3b5a43f5),
	.w4(32'h3b1c0be1),
	.w5(32'h3a8d41da),
	.w6(32'h3b863b94),
	.w7(32'h3b5aca37),
	.w8(32'hb95f8037),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd5709),
	.w1(32'hba5c595f),
	.w2(32'hba04e96a),
	.w3(32'hb946df3e),
	.w4(32'hb9abeebc),
	.w5(32'h39f51e36),
	.w6(32'h3a4a4fce),
	.w7(32'hb859971e),
	.w8(32'hb797b5eb),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfdf02),
	.w1(32'h3a36a331),
	.w2(32'h3a864abe),
	.w3(32'h3a186af8),
	.w4(32'h39b7a6de),
	.w5(32'h38d932cb),
	.w6(32'h3a2d646c),
	.w7(32'h3978aa33),
	.w8(32'hba5b3e26),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37575f80),
	.w1(32'hba5127dc),
	.w2(32'hba52c691),
	.w3(32'hba3b8277),
	.w4(32'hba70cf3e),
	.w5(32'hb9f21192),
	.w6(32'hba80ce45),
	.w7(32'hbac70400),
	.w8(32'hb9ce2dbd),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0420f4),
	.w1(32'hba9ea962),
	.w2(32'hbb17db0c),
	.w3(32'hba497ce2),
	.w4(32'hba8ee703),
	.w5(32'hbb36ebf3),
	.w6(32'hba9e73b8),
	.w7(32'hbaaf4d2c),
	.w8(32'hbafef2fc),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4625ed),
	.w1(32'hbb49065b),
	.w2(32'hbb4469c8),
	.w3(32'hbb51049f),
	.w4(32'hbb5509f6),
	.w5(32'hba1a53ed),
	.w6(32'hba7130e8),
	.w7(32'hbb29c5f8),
	.w8(32'hb98b23fc),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50b128),
	.w1(32'hb71fede3),
	.w2(32'h3a431c9f),
	.w3(32'h38efd7e8),
	.w4(32'h3a08ad23),
	.w5(32'h39cd20e4),
	.w6(32'hb9479ba4),
	.w7(32'h3a848860),
	.w8(32'h39c802b9),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b5f72e),
	.w1(32'h3a7a6935),
	.w2(32'h3a652a56),
	.w3(32'h399116e8),
	.w4(32'h383e5b29),
	.w5(32'h3aebf72e),
	.w6(32'h3a514440),
	.w7(32'h3a0e8ad7),
	.w8(32'h3ad750c8),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34b16a64),
	.w1(32'h39890a0f),
	.w2(32'h3a3e6a6e),
	.w3(32'h3a679251),
	.w4(32'h3a8529e2),
	.w5(32'hb89bc650),
	.w6(32'h38c1dfab),
	.w7(32'h3aa8d683),
	.w8(32'hb8add9bb),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d41a58),
	.w1(32'h38ced227),
	.w2(32'h3a066208),
	.w3(32'hba219e0d),
	.w4(32'h3a2446ef),
	.w5(32'hb9a428d1),
	.w6(32'hb9837160),
	.w7(32'h3a838a46),
	.w8(32'hba30d5c8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb787b2c),
	.w1(32'hbac2f72e),
	.w2(32'hba2fd681),
	.w3(32'hbad4a226),
	.w4(32'hbb5237d9),
	.w5(32'hbb048234),
	.w6(32'hbae9b9eb),
	.w7(32'hbb40ec33),
	.w8(32'hba9bb96c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9f4df),
	.w1(32'h3aa4da0f),
	.w2(32'h3b2c06b9),
	.w3(32'h3aa05e47),
	.w4(32'h3acef849),
	.w5(32'h3b89a72e),
	.w6(32'h3a8d390c),
	.w7(32'h3b1f22d9),
	.w8(32'h3b63417f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b49f2),
	.w1(32'hba5c1e14),
	.w2(32'hba6bc620),
	.w3(32'hba061276),
	.w4(32'hba7bb491),
	.w5(32'hbaff0de1),
	.w6(32'hb95c0670),
	.w7(32'hba9d5ba6),
	.w8(32'hbb009b68),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77b3dd3),
	.w1(32'hba677e8b),
	.w2(32'hb9ca5e3c),
	.w3(32'hba5522d2),
	.w4(32'hb9d5383e),
	.w5(32'hbac221a7),
	.w6(32'hba24c029),
	.w7(32'hb9f0561e),
	.w8(32'hbadf1dbd),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e3772),
	.w1(32'hbab4feac),
	.w2(32'hba478da3),
	.w3(32'hba9395af),
	.w4(32'hba415b46),
	.w5(32'hbaad23c0),
	.w6(32'hba227ac1),
	.w7(32'hba094bef),
	.w8(32'hba7eee62),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e7026),
	.w1(32'hba04eba9),
	.w2(32'hb9b67451),
	.w3(32'h38c3b018),
	.w4(32'hb962dbae),
	.w5(32'hbabeca28),
	.w6(32'h3a8bb36c),
	.w7(32'h3a246931),
	.w8(32'hba8461c2),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a524176),
	.w1(32'hb876f26a),
	.w2(32'hbac74452),
	.w3(32'h3a5795a2),
	.w4(32'hba031581),
	.w5(32'hbb07671c),
	.w6(32'h3aa5005c),
	.w7(32'hb9d1c9fe),
	.w8(32'hb9c75405),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab10b46),
	.w1(32'hba816b54),
	.w2(32'hb9e3de45),
	.w3(32'hbaa317d0),
	.w4(32'hb9160fc7),
	.w5(32'h3a4fd77d),
	.w6(32'hba83e630),
	.w7(32'hb9a6b1ab),
	.w8(32'h39fd6e87),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5ddbd),
	.w1(32'h3a28b66c),
	.w2(32'h3a05b812),
	.w3(32'h3a792606),
	.w4(32'hb8adebca),
	.w5(32'hb8d85934),
	.w6(32'h3919ea03),
	.w7(32'h3a0a22a5),
	.w8(32'h3a275e3f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa62484),
	.w1(32'h38847381),
	.w2(32'h3a014f7e),
	.w3(32'h3817ca20),
	.w4(32'hba86a319),
	.w5(32'hba41c09f),
	.w6(32'hba9b7486),
	.w7(32'hba9ce574),
	.w8(32'h3824ab56),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3ee40),
	.w1(32'h3a724fd6),
	.w2(32'h38feddec),
	.w3(32'h395193b3),
	.w4(32'h3a715548),
	.w5(32'h3a93de88),
	.w6(32'hb981344e),
	.w7(32'hb8a55c67),
	.w8(32'h3acd5274),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa83c73),
	.w1(32'h3954dd70),
	.w2(32'h3a6664be),
	.w3(32'h3a0bf89b),
	.w4(32'hba45ee5a),
	.w5(32'hbb24c7a2),
	.w6(32'h3a61b15d),
	.w7(32'h3a179030),
	.w8(32'hbade3399),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cdf02),
	.w1(32'hba810360),
	.w2(32'hb9ebe178),
	.w3(32'hbaefc347),
	.w4(32'hba8d61d6),
	.w5(32'h39e75bfd),
	.w6(32'hba8e8ce9),
	.w7(32'hba8c57f9),
	.w8(32'h36c16098),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d20f85),
	.w1(32'h3a071863),
	.w2(32'h3b27a626),
	.w3(32'h3a7d102f),
	.w4(32'h39639598),
	.w5(32'h3ad24071),
	.w6(32'hb988dbb3),
	.w7(32'hb9186382),
	.w8(32'h3a837a40),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c5b64a),
	.w1(32'hb8cbb21d),
	.w2(32'h39c3096b),
	.w3(32'hba422793),
	.w4(32'hb91ac53a),
	.w5(32'h391943a3),
	.w6(32'h39a8dbb4),
	.w7(32'h39b5615c),
	.w8(32'h3a0eddfa),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eb56d),
	.w1(32'h396b6d01),
	.w2(32'h38ccc59d),
	.w3(32'h3886b341),
	.w4(32'h39d91960),
	.w5(32'h39f3a04e),
	.w6(32'hb91c3e8b),
	.w7(32'h375522c8),
	.w8(32'hb9ba9190),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2118b8),
	.w1(32'hb9cb2262),
	.w2(32'hbac79cc0),
	.w3(32'hb91b52b0),
	.w4(32'hba5f9c2e),
	.w5(32'hbaf0dba9),
	.w6(32'h3a27fe82),
	.w7(32'hba0116ba),
	.w8(32'hbaafdf47),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb304d5e),
	.w1(32'hb921bd86),
	.w2(32'h3b04e05e),
	.w3(32'hba85b396),
	.w4(32'hba0a7793),
	.w5(32'h3aee7163),
	.w6(32'hbaa6c7dd),
	.w7(32'h3aa30cca),
	.w8(32'h39cef826),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a41fe8),
	.w1(32'hb90b22d2),
	.w2(32'h3766fd67),
	.w3(32'h392e4dea),
	.w4(32'hb9aeda0c),
	.w5(32'hb8db74a6),
	.w6(32'h3a2bf82d),
	.w7(32'hba33dee9),
	.w8(32'hb872de03),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392158d8),
	.w1(32'hba20eb0b),
	.w2(32'h39391665),
	.w3(32'hba876f77),
	.w4(32'hb90ce43b),
	.w5(32'hb9de4761),
	.w6(32'hb91c3e04),
	.w7(32'h3a080b95),
	.w8(32'hb7907156),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b497e5),
	.w1(32'h39d5d4cd),
	.w2(32'h39bbe2dc),
	.w3(32'hba6bc152),
	.w4(32'h39497739),
	.w5(32'h39b11f65),
	.w6(32'h3a91edd6),
	.w7(32'h398d6964),
	.w8(32'hb905c625),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ec195),
	.w1(32'h39a93e12),
	.w2(32'hbab8b84c),
	.w3(32'hba618eb5),
	.w4(32'hba30504f),
	.w5(32'hb889f196),
	.w6(32'h39cc7e5c),
	.w7(32'h3a4eacd3),
	.w8(32'h3ae61f85),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba895a96),
	.w1(32'h39f9c272),
	.w2(32'hba21fe13),
	.w3(32'hbb08c686),
	.w4(32'hbb0ffad8),
	.w5(32'hbb5b1696),
	.w6(32'hba8f0d50),
	.w7(32'hbaf5b6b2),
	.w8(32'hbb31cf65),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafca894),
	.w1(32'hba7ae8ea),
	.w2(32'hba88026d),
	.w3(32'hba90016a),
	.w4(32'hbaea6c7d),
	.w5(32'h3b6224f9),
	.w6(32'hbaba8fb5),
	.w7(32'hba9bb659),
	.w8(32'h3b3e7fbc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d8113),
	.w1(32'h3ac8bbab),
	.w2(32'h3b03cbb8),
	.w3(32'h3affd86f),
	.w4(32'h3b0ff4d4),
	.w5(32'h3b08c490),
	.w6(32'h3ab0971d),
	.w7(32'h3ad26387),
	.w8(32'h3b0bbc1a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b5a9a),
	.w1(32'h3ae3e670),
	.w2(32'h3acd173f),
	.w3(32'h3a4e45ce),
	.w4(32'h3ab89d0e),
	.w5(32'h39ad3cb1),
	.w6(32'h3a3da7dc),
	.w7(32'h3ab0fdcf),
	.w8(32'hb982d63f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9f6d5),
	.w1(32'h3aacda10),
	.w2(32'h3acf8b19),
	.w3(32'h3aaf613c),
	.w4(32'h3ac8c918),
	.w5(32'hbac1c543),
	.w6(32'h3a98b9c2),
	.w7(32'h3a9dfbb3),
	.w8(32'hbae7c92d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba827b1b),
	.w1(32'hbadcac65),
	.w2(32'hb9acc47c),
	.w3(32'hbad0e9c4),
	.w4(32'h395801af),
	.w5(32'hba1daf56),
	.w6(32'hbad253c1),
	.w7(32'hb98d69d9),
	.w8(32'h39e38c12),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8bdc9),
	.w1(32'hbaf2d3f4),
	.w2(32'hbb1b5857),
	.w3(32'hbabdfa00),
	.w4(32'hbb1178c2),
	.w5(32'hb7f17afb),
	.w6(32'hb8c871ca),
	.w7(32'hbaa250b7),
	.w8(32'hb903b176),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40bb39),
	.w1(32'hbaa42fd3),
	.w2(32'hbb0f04e8),
	.w3(32'hbabee23e),
	.w4(32'hbb0adc60),
	.w5(32'hbb508e0d),
	.w6(32'hbab26877),
	.w7(32'hbae6f57c),
	.w8(32'hbb62814d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba554bd2),
	.w1(32'h39bc2a3f),
	.w2(32'h391ad5b9),
	.w3(32'h398253ec),
	.w4(32'h39793991),
	.w5(32'hb83925d9),
	.w6(32'h3979209c),
	.w7(32'h3962db44),
	.w8(32'h39a866d9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9946af2),
	.w1(32'hb9362613),
	.w2(32'hba3a26b7),
	.w3(32'h392f1fe2),
	.w4(32'hba13b7fc),
	.w5(32'hba0257ff),
	.w6(32'h399ae680),
	.w7(32'hb9677a66),
	.w8(32'h3a3ea032),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b7a82a),
	.w1(32'h3a3f140f),
	.w2(32'h3a5ecbb8),
	.w3(32'hbac675cf),
	.w4(32'hbae57fec),
	.w5(32'h39acdf2e),
	.w6(32'h395a5ab1),
	.w7(32'h387bd241),
	.w8(32'h3a4dc744),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f506b),
	.w1(32'h3ab72e53),
	.w2(32'hba9f49bf),
	.w3(32'hb9c7d024),
	.w4(32'hba6a0043),
	.w5(32'hbb6a9e63),
	.w6(32'hbb167891),
	.w7(32'hb9d86837),
	.w8(32'hbb6138bc),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb396192),
	.w1(32'hba664238),
	.w2(32'hbad9a2a1),
	.w3(32'h3a2a9937),
	.w4(32'hbb5acacc),
	.w5(32'h3aee2c71),
	.w6(32'h39419ef8),
	.w7(32'hbaea4040),
	.w8(32'h3b2332cc),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cbc56),
	.w1(32'h3a537502),
	.w2(32'h3a9996d4),
	.w3(32'h3a716571),
	.w4(32'h3a872599),
	.w5(32'h3afd90d0),
	.w6(32'h3a8b9565),
	.w7(32'h3a59f1dc),
	.w8(32'h3ab3e2e0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61f5ea),
	.w1(32'h3a84124d),
	.w2(32'h3b980417),
	.w3(32'h3a80e11e),
	.w4(32'h3ab8e09c),
	.w5(32'h3b342536),
	.w6(32'h3aa27762),
	.w7(32'h3b572ee3),
	.w8(32'h3b823976),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a120a0c),
	.w1(32'hba43141d),
	.w2(32'hba8e1db5),
	.w3(32'hbb139890),
	.w4(32'hba74006b),
	.w5(32'h39e79b69),
	.w6(32'h3a3b1933),
	.w7(32'h3ad69a93),
	.w8(32'h3a0ea219),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd3152),
	.w1(32'h3a92b5db),
	.w2(32'h3ae80994),
	.w3(32'h3ab7568f),
	.w4(32'h3a9afd82),
	.w5(32'h3a5c304d),
	.w6(32'h3ac65842),
	.w7(32'h3abdd1f6),
	.w8(32'h3aa0c92d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb966dfb3),
	.w1(32'hba089ead),
	.w2(32'hb9e71132),
	.w3(32'hbad71449),
	.w4(32'hbace93d3),
	.w5(32'hb99eacc1),
	.w6(32'hbadb36f0),
	.w7(32'hba799594),
	.w8(32'hb9779642),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a51d2e),
	.w1(32'h39dd1fda),
	.w2(32'h3a2677d3),
	.w3(32'hb95b42f0),
	.w4(32'h39483f56),
	.w5(32'hb99ddf81),
	.w6(32'hb9452300),
	.w7(32'h39be39af),
	.w8(32'h3a03fcf2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39adf4cc),
	.w1(32'h3985a0d2),
	.w2(32'hba31cfb7),
	.w3(32'hb9e8208c),
	.w4(32'hbab26c30),
	.w5(32'h396b0025),
	.w6(32'hba25f1af),
	.w7(32'hba8b8051),
	.w8(32'h3a0b6f34),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e11e39),
	.w1(32'h3a9deaec),
	.w2(32'h3b1a66b8),
	.w3(32'h3a069eac),
	.w4(32'h3a3efe5f),
	.w5(32'h3ac37dfa),
	.w6(32'hba8d8cf1),
	.w7(32'h3a65aa23),
	.w8(32'h3abbb2bd),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b86aa),
	.w1(32'hba9ec0b8),
	.w2(32'hb986c918),
	.w3(32'hbae09a62),
	.w4(32'hba2b4a05),
	.w5(32'hb96bebfe),
	.w6(32'hba114e65),
	.w7(32'hb7e454b3),
	.w8(32'h395ebb64),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386dae95),
	.w1(32'hbb0483da),
	.w2(32'hbabfc026),
	.w3(32'hba998402),
	.w4(32'hba8c1eec),
	.w5(32'hbb56513f),
	.w6(32'h39bf18d9),
	.w7(32'hba6caa09),
	.w8(32'hbb46a11c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3950a5ee),
	.w1(32'hba072d28),
	.w2(32'hba132d2a),
	.w3(32'hba32a403),
	.w4(32'hba7b4e5c),
	.w5(32'hbadcf137),
	.w6(32'h38318528),
	.w7(32'hba16d4c1),
	.w8(32'hba6c829a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dec86),
	.w1(32'hbae2750f),
	.w2(32'hba3689fb),
	.w3(32'hbb373a52),
	.w4(32'hba979322),
	.w5(32'h3a8a1a10),
	.w6(32'hba3362ab),
	.w7(32'hb8df47c8),
	.w8(32'h3b12632a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c35623),
	.w1(32'hba32b815),
	.w2(32'hb99cd624),
	.w3(32'hb842dfc5),
	.w4(32'h39270b85),
	.w5(32'h398dd08f),
	.w6(32'hb95f7fdb),
	.w7(32'hb8b28ba8),
	.w8(32'hb8feb40d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26d68c),
	.w1(32'h3a8052c0),
	.w2(32'h393ade28),
	.w3(32'h3a0c98b0),
	.w4(32'h38c14ba7),
	.w5(32'h38ec46a7),
	.w6(32'h3a0ec360),
	.w7(32'hb92fe8e7),
	.w8(32'h390f50ab),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96921de),
	.w1(32'hb9de8b64),
	.w2(32'hba9de9af),
	.w3(32'hba09bf4c),
	.w4(32'hbaa7d594),
	.w5(32'hba7f29b6),
	.w6(32'hbaa33032),
	.w7(32'hbab4da0d),
	.w8(32'hba9ddbc3),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4441ad),
	.w1(32'h3a3218d0),
	.w2(32'h3a83c9e7),
	.w3(32'h3a76b457),
	.w4(32'h38b239e1),
	.w5(32'hb9ff0eab),
	.w6(32'h3aa5a525),
	.w7(32'h3a8c2a46),
	.w8(32'hba1709cb),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae57790),
	.w1(32'h39bf9c2f),
	.w2(32'h3a9945a9),
	.w3(32'hba0dddef),
	.w4(32'h398ef077),
	.w5(32'h3a64ed5d),
	.w6(32'hb981117c),
	.w7(32'h3a27adfe),
	.w8(32'h3a2f1615),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd8711),
	.w1(32'hbb0f798f),
	.w2(32'hbae2c315),
	.w3(32'hbad1db44),
	.w4(32'hbaf8dd27),
	.w5(32'hbb2c5b62),
	.w6(32'hb988c7f7),
	.w7(32'hba876dcc),
	.w8(32'hba6945ef),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba926135),
	.w1(32'hb9aa814d),
	.w2(32'hb8dad796),
	.w3(32'hba8211b5),
	.w4(32'hb9c311a6),
	.w5(32'hbb772ffd),
	.w6(32'h391c967b),
	.w7(32'h3a02ea8d),
	.w8(32'hbb211cdd),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb150132),
	.w1(32'hbb03fe27),
	.w2(32'hbb20613f),
	.w3(32'hbb1465ad),
	.w4(32'hbb229104),
	.w5(32'h371d49f6),
	.w6(32'hbabc4db4),
	.w7(32'hbb153e4f),
	.w8(32'h391e96ba),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f4a0f),
	.w1(32'hbacb642c),
	.w2(32'hbaca598a),
	.w3(32'hbae0969f),
	.w4(32'hbab6585a),
	.w5(32'hbb3e4c50),
	.w6(32'hb7561bd0),
	.w7(32'hb9932110),
	.w8(32'hbb0ca7f5),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb058acb),
	.w1(32'hbada43ab),
	.w2(32'hbaadbcbb),
	.w3(32'hbb003e0c),
	.w4(32'hbb0046c5),
	.w5(32'h3b0aee3b),
	.w6(32'hbabbca07),
	.w7(32'hbadcfc7b),
	.w8(32'h3b170699),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dae54),
	.w1(32'h3b5e1f99),
	.w2(32'h3b8e4014),
	.w3(32'h3b560bf5),
	.w4(32'h3b8e9015),
	.w5(32'h3a2e76ac),
	.w6(32'h3b8b4f1c),
	.w7(32'h3bb389ea),
	.w8(32'h3ac3536d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7385a8),
	.w1(32'h39b121c2),
	.w2(32'h3a5a568a),
	.w3(32'h3a16787c),
	.w4(32'h3aadd122),
	.w5(32'hba3ae3fa),
	.w6(32'h398c6829),
	.w7(32'h3a56e1fe),
	.w8(32'hb9d99363),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00f593),
	.w1(32'hba4121d7),
	.w2(32'hb99b2e87),
	.w3(32'hba667fe8),
	.w4(32'hba12b82e),
	.w5(32'hbaa77280),
	.w6(32'hba8794ea),
	.w7(32'hb9de9750),
	.w8(32'hba554108),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5ea60),
	.w1(32'hbb083c3a),
	.w2(32'h3a68a8bb),
	.w3(32'hbb563d76),
	.w4(32'hbb46d204),
	.w5(32'h3a19340e),
	.w6(32'hbae2858e),
	.w7(32'hbadc1d03),
	.w8(32'hbace755f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf15a2),
	.w1(32'hbb062b3b),
	.w2(32'h39ce23bf),
	.w3(32'hbab9963e),
	.w4(32'hb817bf1a),
	.w5(32'h391cfa95),
	.w6(32'hbaaaf7d2),
	.w7(32'h3ad0134f),
	.w8(32'hb82d0a7e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadece55),
	.w1(32'hba293dbe),
	.w2(32'hba2e65c3),
	.w3(32'hbad14dbe),
	.w4(32'hbb07b844),
	.w5(32'hbb1b4965),
	.w6(32'h3a0af55b),
	.w7(32'hb9a5c6e0),
	.w8(32'hbb12d1c8),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9aaf9),
	.w1(32'hbb375989),
	.w2(32'hbb024418),
	.w3(32'hbafb4526),
	.w4(32'hbb9d6c42),
	.w5(32'hbb19b203),
	.w6(32'hbb1b02ec),
	.w7(32'hba6d3ed3),
	.w8(32'hbab618f0),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32fded),
	.w1(32'hb8f33d07),
	.w2(32'h392b294f),
	.w3(32'h399c248a),
	.w4(32'h3a4ed859),
	.w5(32'hba397e08),
	.w6(32'hba3e8916),
	.w7(32'h399f5885),
	.w8(32'hba293c3e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa01f63),
	.w1(32'hbaac3bd1),
	.w2(32'hba88a9b0),
	.w3(32'hbaec0d90),
	.w4(32'hbadad64e),
	.w5(32'hba9141f7),
	.w6(32'hbabd9bfb),
	.w7(32'hbae3d24c),
	.w8(32'hbae59894),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b17637),
	.w1(32'h3b6a5c4b),
	.w2(32'h3b596d5e),
	.w3(32'h3b07d3b8),
	.w4(32'h3b0263bf),
	.w5(32'h3bd739c7),
	.w6(32'hbafd09d1),
	.w7(32'hba766551),
	.w8(32'h3b97652f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968b079),
	.w1(32'h3a31b555),
	.w2(32'h3b51e528),
	.w3(32'h39a4af17),
	.w4(32'hb9917995),
	.w5(32'h391a3821),
	.w6(32'h39806395),
	.w7(32'h3ac58ef7),
	.w8(32'h3a9e4b51),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e2629),
	.w1(32'hbb2da00a),
	.w2(32'hbb13441d),
	.w3(32'hbb212866),
	.w4(32'hbafe605b),
	.w5(32'hba6880b3),
	.w6(32'hbb8d368b),
	.w7(32'hbb41c82e),
	.w8(32'hb9f66527),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d8a56),
	.w1(32'h399f8d90),
	.w2(32'hba1102b1),
	.w3(32'h3ac1d8f8),
	.w4(32'h3a5b34fc),
	.w5(32'hba91a0ae),
	.w6(32'h3b3bfa84),
	.w7(32'h3a8c3252),
	.w8(32'hba18f525),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f8d83),
	.w1(32'hba1e3e54),
	.w2(32'hbaa1ba5a),
	.w3(32'hb98175e3),
	.w4(32'hba50939b),
	.w5(32'hbae5624c),
	.w6(32'h3a944bfc),
	.w7(32'hba02db51),
	.w8(32'hba975931),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a2546),
	.w1(32'h3a8f715b),
	.w2(32'h3a81efd6),
	.w3(32'h3942fa91),
	.w4(32'h3995e134),
	.w5(32'hbaad99cd),
	.w6(32'h3aab9db1),
	.w7(32'h3a75b819),
	.w8(32'hbaca3824),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac971e0),
	.w1(32'hbb095e6e),
	.w2(32'hbac2f387),
	.w3(32'hbad718d8),
	.w4(32'hba8d7374),
	.w5(32'h39bef355),
	.w6(32'hbae31aef),
	.w7(32'hba8fcabd),
	.w8(32'h38778257),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9414afd),
	.w1(32'hba2f52e0),
	.w2(32'hb9ff34f5),
	.w3(32'h36a92722),
	.w4(32'hba233c74),
	.w5(32'hb8984f45),
	.w6(32'hba974a65),
	.w7(32'hba53a146),
	.w8(32'h398eecdb),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9404b),
	.w1(32'h3aa312a9),
	.w2(32'h3a8bdc84),
	.w3(32'h3a95234a),
	.w4(32'h3a5a4ea8),
	.w5(32'hb91de12c),
	.w6(32'h3aad10a2),
	.w7(32'h3a826ba6),
	.w8(32'h3905aac8),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa626b),
	.w1(32'h3b05b39d),
	.w2(32'h3b418d42),
	.w3(32'h3a5a2a4f),
	.w4(32'h3b5923a5),
	.w5(32'h3b6d8552),
	.w6(32'hba8404b3),
	.w7(32'h3ab26d88),
	.w8(32'h3af19fbc),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ad481),
	.w1(32'hbb8158a1),
	.w2(32'hbb3d1567),
	.w3(32'hbae4c118),
	.w4(32'hbb674866),
	.w5(32'hbb325f65),
	.w6(32'hbb8237b7),
	.w7(32'hbb07af77),
	.w8(32'hbb3b0e29),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ffc0c),
	.w1(32'hba9ee214),
	.w2(32'hbb13d16e),
	.w3(32'hbb0e3bc1),
	.w4(32'hbad83a80),
	.w5(32'hbaea7587),
	.w6(32'hba3e179b),
	.w7(32'hb9d1cb02),
	.w8(32'hba04efbc),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986a410),
	.w1(32'hba551f4f),
	.w2(32'h3a012702),
	.w3(32'hba8d9e89),
	.w4(32'hb822a2a0),
	.w5(32'h37ae105e),
	.w6(32'h3ab2388c),
	.w7(32'hb89b54f3),
	.w8(32'hba568fe4),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb031284),
	.w1(32'h3a006072),
	.w2(32'h3b1e68ac),
	.w3(32'hbb22f411),
	.w4(32'hbb62430b),
	.w5(32'hbb7095e4),
	.w6(32'hbb9e1f33),
	.w7(32'h3a6848ca),
	.w8(32'hbb0ebdef),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941b21),
	.w1(32'hbbc1891e),
	.w2(32'hbbbfb5ee),
	.w3(32'hbace6726),
	.w4(32'hbb5da98b),
	.w5(32'h3aae71dd),
	.w6(32'hbb7eb1d0),
	.w7(32'hbb2988f9),
	.w8(32'h39ad9203),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b107622),
	.w1(32'hb9da2383),
	.w2(32'h3af610ca),
	.w3(32'h3a7a5647),
	.w4(32'hbad7988b),
	.w5(32'hba801b97),
	.w6(32'hbb654ec7),
	.w7(32'hba2b7424),
	.w8(32'hbb2b28da),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf880cc),
	.w1(32'hba937b92),
	.w2(32'hba897667),
	.w3(32'hb983d1f4),
	.w4(32'hbae0921a),
	.w5(32'hba81913b),
	.w6(32'h397356fa),
	.w7(32'hbb297200),
	.w8(32'h3920b0ec),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf91734),
	.w1(32'hbb979914),
	.w2(32'hbb2a196c),
	.w3(32'hb94849aa),
	.w4(32'hbac99bec),
	.w5(32'h3ab7544c),
	.w6(32'hba189b31),
	.w7(32'hbba815d0),
	.w8(32'h39d24bf8),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bceffc),
	.w1(32'h3970291b),
	.w2(32'h3abb124b),
	.w3(32'hba945918),
	.w4(32'hba1b891d),
	.w5(32'hba52c49e),
	.w6(32'hba21d1e7),
	.w7(32'h39f01c34),
	.w8(32'hb9aad93a),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7dbc8),
	.w1(32'h3a92b4c9),
	.w2(32'h3b029ef0),
	.w3(32'hb87f7eac),
	.w4(32'h3b3197b4),
	.w5(32'hbb02c222),
	.w6(32'h39424878),
	.w7(32'h3b6320fc),
	.w8(32'hbb03fe3f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff69a1),
	.w1(32'hba272442),
	.w2(32'hbb21eca1),
	.w3(32'hbae0e502),
	.w4(32'hbb5c2940),
	.w5(32'h39c04be3),
	.w6(32'hbb08c89c),
	.w7(32'hbb817499),
	.w8(32'hb8482430),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa4261),
	.w1(32'hb81a4a83),
	.w2(32'h39b178cc),
	.w3(32'h3a8ddf6e),
	.w4(32'h3ab3cc01),
	.w5(32'h3a157cd7),
	.w6(32'hbb28121c),
	.w7(32'hba86c71c),
	.w8(32'h39f58037),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79a167),
	.w1(32'hbb08cc41),
	.w2(32'hbb14d977),
	.w3(32'hbb81caf3),
	.w4(32'hba853fdc),
	.w5(32'h3a5b3b01),
	.w6(32'hba0d0465),
	.w7(32'hb9d21255),
	.w8(32'h3b00b888),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1de6b7),
	.w1(32'h3b082f4c),
	.w2(32'h3b25e08c),
	.w3(32'h3b368d26),
	.w4(32'h3a1fa63e),
	.w5(32'hb9bd5217),
	.w6(32'h3b166b4f),
	.w7(32'h39015c37),
	.w8(32'hb9df8f25),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9ad6c),
	.w1(32'h3b038e93),
	.w2(32'h3b5a16a2),
	.w3(32'hb78c1c0a),
	.w4(32'h3adad4f6),
	.w5(32'h3b7fa08b),
	.w6(32'hba02c204),
	.w7(32'h3b1c779d),
	.w8(32'h3bbbf4d5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec449b),
	.w1(32'hbb436987),
	.w2(32'hbb0eef7c),
	.w3(32'hbaabb420),
	.w4(32'hbaa2a6bc),
	.w5(32'h3a9bd4ca),
	.w6(32'hbaca9db8),
	.w7(32'hbac481ef),
	.w8(32'h3aa3836c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa67de6),
	.w1(32'hba337ca9),
	.w2(32'hb9f291f5),
	.w3(32'hbb20f048),
	.w4(32'hba616f30),
	.w5(32'hbb8a22ba),
	.w6(32'h3b52f115),
	.w7(32'h39ace06d),
	.w8(32'hbb6225b2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01e26b),
	.w1(32'hba47b773),
	.w2(32'hba3f819c),
	.w3(32'hbb4e6f73),
	.w4(32'hb971f97a),
	.w5(32'h3a94b339),
	.w6(32'hbb41cf07),
	.w7(32'hb8e178a6),
	.w8(32'hba347bfc),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba684070),
	.w1(32'h39d36a15),
	.w2(32'h3a88e4b6),
	.w3(32'h3b3d8e6f),
	.w4(32'h39aebb49),
	.w5(32'h3a5d49f3),
	.w6(32'h3aadbb20),
	.w7(32'hb9545dd1),
	.w8(32'hb9de7bf3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42b4a6),
	.w1(32'hbaab2d97),
	.w2(32'hbb449755),
	.w3(32'hbb3b7bdc),
	.w4(32'hbb483491),
	.w5(32'hbbe4e684),
	.w6(32'hbbae2483),
	.w7(32'hbb474608),
	.w8(32'hbbd1a9e2),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac9bff),
	.w1(32'hbb89f529),
	.w2(32'hbb84ad13),
	.w3(32'hbb47bb21),
	.w4(32'hbb2c917c),
	.w5(32'h3b1b9c3a),
	.w6(32'hbb461034),
	.w7(32'hbb18c7aa),
	.w8(32'hb995f0e3),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e77cc),
	.w1(32'hbac107de),
	.w2(32'hbb0dc284),
	.w3(32'hba815be8),
	.w4(32'hbab21c7e),
	.w5(32'h3b3769a5),
	.w6(32'h3a5682b8),
	.w7(32'hbaa8d89d),
	.w8(32'h3b45df27),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbb56f),
	.w1(32'h3b926a34),
	.w2(32'h3b366c70),
	.w3(32'h3a5a7a69),
	.w4(32'h394a8c65),
	.w5(32'h39fc7082),
	.w6(32'h3b3b7152),
	.w7(32'h3b1405f9),
	.w8(32'hba8ec44e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae13e85),
	.w1(32'h393a1ab9),
	.w2(32'h3b034031),
	.w3(32'h3af4fbbf),
	.w4(32'h3b63efdc),
	.w5(32'hbabbecc7),
	.w6(32'h3c2ae100),
	.w7(32'h3c012fff),
	.w8(32'h3ab3bc7d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9eddc5),
	.w1(32'h3b30eb12),
	.w2(32'hbaa2424d),
	.w3(32'hba8f41b5),
	.w4(32'hba98647d),
	.w5(32'h3b8c8c32),
	.w6(32'h3840451a),
	.w7(32'hbb218847),
	.w8(32'h3b221b92),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dc5f7),
	.w1(32'h3bb3737a),
	.w2(32'h3bb2effd),
	.w3(32'h3aac0bcd),
	.w4(32'h3b245c7a),
	.w5(32'hbaa2b70c),
	.w6(32'h3c0c3663),
	.w7(32'h3bcd11f7),
	.w8(32'hb94acf57),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57b4cf),
	.w1(32'h39eebd32),
	.w2(32'hbb42344f),
	.w3(32'hbb6ebbfa),
	.w4(32'hbb6429b8),
	.w5(32'hbbd893b2),
	.w6(32'hbb8d95ab),
	.w7(32'hbb65f7cc),
	.w8(32'hbbdb386e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05258b),
	.w1(32'h3a997ec9),
	.w2(32'h3ae24e8c),
	.w3(32'hb9a88e3a),
	.w4(32'h3a6b237c),
	.w5(32'h3a84337d),
	.w6(32'h3b181f3c),
	.w7(32'h3b43b63f),
	.w8(32'h3a2422d7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe5336),
	.w1(32'hbb143131),
	.w2(32'hbb03b552),
	.w3(32'hbb08cdf2),
	.w4(32'hbb219d44),
	.w5(32'hbb184c8f),
	.w6(32'h39eba449),
	.w7(32'hbac62e43),
	.w8(32'hba315799),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule