module layer_10_featuremap_127(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba0416),
	.w1(32'h3ac7e24b),
	.w2(32'h3aac6668),
	.w3(32'hbabddc95),
	.w4(32'h3a93e3e5),
	.w5(32'h3b012991),
	.w6(32'h3b106dd9),
	.w7(32'h3b468470),
	.w8(32'h3b0e9d12),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aded823),
	.w1(32'hb7ce3715),
	.w2(32'h3aae6322),
	.w3(32'h3aa7a629),
	.w4(32'h39c2852d),
	.w5(32'h390cc84f),
	.w6(32'hb8e18071),
	.w7(32'h3a0d7b03),
	.w8(32'h3ac4c5f7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2beae),
	.w1(32'h3a1c22c3),
	.w2(32'h39dff776),
	.w3(32'h3a7ba530),
	.w4(32'hb8ee6dd4),
	.w5(32'hbb26b302),
	.w6(32'h3acf274d),
	.w7(32'hba2b7148),
	.w8(32'h39998d41),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85eb94),
	.w1(32'hbaa907d6),
	.w2(32'hbb2eb825),
	.w3(32'hbaaf9a22),
	.w4(32'hba92dda2),
	.w5(32'hbb8f48e7),
	.w6(32'h3b429b9f),
	.w7(32'h3a9ba389),
	.w8(32'h3bc9de08),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e1d5a),
	.w1(32'hba2932cf),
	.w2(32'h3aeb2221),
	.w3(32'hbab9c2c3),
	.w4(32'hba9bdb12),
	.w5(32'h3aeb8cd6),
	.w6(32'h387ffccd),
	.w7(32'h3b7186c7),
	.w8(32'h3a81a877),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b093f7f),
	.w1(32'h3966212b),
	.w2(32'hbaadb77c),
	.w3(32'hba48ed53),
	.w4(32'hbb563e5f),
	.w5(32'hbb6e491d),
	.w6(32'hbab0f0c6),
	.w7(32'hbb4bf49e),
	.w8(32'hbb6883c1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaede385),
	.w1(32'hb94460b3),
	.w2(32'hba13130d),
	.w3(32'hbb1fdbe1),
	.w4(32'h3a8b16e2),
	.w5(32'h3958c7d1),
	.w6(32'hb8b9ddab),
	.w7(32'hba8b55c1),
	.w8(32'h3b3bc590),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afda306),
	.w1(32'hba49da6d),
	.w2(32'h39cdd8bf),
	.w3(32'h3b173a8e),
	.w4(32'hbb54eb46),
	.w5(32'hba06e3e5),
	.w6(32'hbad7dcad),
	.w7(32'hb9f428bf),
	.w8(32'hba80814e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba387253),
	.w1(32'h3a1de852),
	.w2(32'h3a81d694),
	.w3(32'hba69b0ab),
	.w4(32'hba87c258),
	.w5(32'hb736f455),
	.w6(32'h3a91fe81),
	.w7(32'h3acb0843),
	.w8(32'hbaaa0100),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e871e),
	.w1(32'hbbdfea02),
	.w2(32'hb9ba3438),
	.w3(32'hbab466ad),
	.w4(32'hbbe68183),
	.w5(32'hbb219a3e),
	.w6(32'hbc1f34ed),
	.w7(32'hbb95984b),
	.w8(32'hbaf0b77a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce1f5c),
	.w1(32'h3b91f9b7),
	.w2(32'hba76943c),
	.w3(32'hba993045),
	.w4(32'h3a9a04fc),
	.w5(32'hbb76c13e),
	.w6(32'h3b79ebc4),
	.w7(32'hbb08e200),
	.w8(32'hbb0d558e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06cef3),
	.w1(32'hbad34184),
	.w2(32'hbaca7702),
	.w3(32'hbb285a2e),
	.w4(32'hbb7bd4a0),
	.w5(32'hbb610dbf),
	.w6(32'hbadcad5d),
	.w7(32'hbaaa3cfe),
	.w8(32'h398929e3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3906e196),
	.w1(32'hba5fe571),
	.w2(32'hbaeba6f9),
	.w3(32'hbb98bfa3),
	.w4(32'hbb0fb182),
	.w5(32'hbae1d21e),
	.w6(32'hb916b57f),
	.w7(32'hb9b4ef3f),
	.w8(32'h3ae970ef),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a5fca),
	.w1(32'hbb3cf25f),
	.w2(32'h3a5d9ae6),
	.w3(32'h39c94e10),
	.w4(32'hbb4ae7a4),
	.w5(32'h3a8216b8),
	.w6(32'hbba05cd2),
	.w7(32'hbaee99b9),
	.w8(32'h3a0bf0e8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b693b),
	.w1(32'h3bb6d33f),
	.w2(32'hbad6942b),
	.w3(32'h3b932e44),
	.w4(32'h3aeefa7a),
	.w5(32'hbb15ff8c),
	.w6(32'h3ae7ae5a),
	.w7(32'h3abffcb5),
	.w8(32'h38bddc3e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaadc2d),
	.w1(32'h3af200b7),
	.w2(32'h3b4779d5),
	.w3(32'hbbbbcd39),
	.w4(32'hb89b847a),
	.w5(32'h3abe1578),
	.w6(32'h3b1fddca),
	.w7(32'h3b7ea5af),
	.w8(32'h3af60ab6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad27a7b),
	.w1(32'h3b717c37),
	.w2(32'h3b288c6c),
	.w3(32'h3ab70978),
	.w4(32'h3b88b8c7),
	.w5(32'h3aa03928),
	.w6(32'h39a342a4),
	.w7(32'hb9f3500f),
	.w8(32'hbbc7a1cc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5de43),
	.w1(32'hbaf52c4a),
	.w2(32'h3ad7f61c),
	.w3(32'h3a9de50d),
	.w4(32'hba884ef7),
	.w5(32'h3ac9ebb3),
	.w6(32'hbb279fd8),
	.w7(32'h39b18a26),
	.w8(32'h3add4368),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52f107),
	.w1(32'hb9a68d6f),
	.w2(32'h3abd8ee4),
	.w3(32'h38f18b45),
	.w4(32'hba86cadc),
	.w5(32'h3a07c739),
	.w6(32'hb8ac9a28),
	.w7(32'h39cc3126),
	.w8(32'h3a2d8f2b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba552068),
	.w1(32'hb8b5c98b),
	.w2(32'h3a688252),
	.w3(32'hbb0c1d17),
	.w4(32'hbaf10bc2),
	.w5(32'hb880b539),
	.w6(32'hb913e696),
	.w7(32'h3afe405b),
	.w8(32'hbacf95db),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97fa5b),
	.w1(32'h3b23c28c),
	.w2(32'hbaa7c921),
	.w3(32'hbaad7b32),
	.w4(32'hba4607a3),
	.w5(32'hbb653df4),
	.w6(32'hb93b5531),
	.w7(32'hbb6e4037),
	.w8(32'h3a455beb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ad594),
	.w1(32'hbbbf6cfc),
	.w2(32'hbbcbdccc),
	.w3(32'h3975c658),
	.w4(32'h3ab6c90b),
	.w5(32'hbb6a2c68),
	.w6(32'h3b047c98),
	.w7(32'hbb1d139e),
	.w8(32'h3b513ebf),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0899c),
	.w1(32'h3c107160),
	.w2(32'h3cb96af5),
	.w3(32'hbb8f4f34),
	.w4(32'hbb2b3801),
	.w5(32'h3c35d839),
	.w6(32'h3bb92565),
	.w7(32'h3c818d0b),
	.w8(32'hbb0da7d8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec4abc),
	.w1(32'hb9afcbcd),
	.w2(32'h39f0f097),
	.w3(32'hbbd8c1a1),
	.w4(32'hbb4ba273),
	.w5(32'hba897d3d),
	.w6(32'hba81a309),
	.w7(32'hb9f7e56c),
	.w8(32'hba6ae6e7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12fd5a),
	.w1(32'h3b9276a1),
	.w2(32'h3bb05838),
	.w3(32'hb94a67e5),
	.w4(32'hba9a681f),
	.w5(32'hbab70d19),
	.w6(32'h3b597e74),
	.w7(32'h3b87afba),
	.w8(32'h3ab033f3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca0b1f),
	.w1(32'h3be430b8),
	.w2(32'h3b5cdd85),
	.w3(32'hb96fb70e),
	.w4(32'h3ba7e10b),
	.w5(32'h3bcf330f),
	.w6(32'h3b2d2a5a),
	.w7(32'h39d7ab4f),
	.w8(32'hba0b70e4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0ef69),
	.w1(32'hba308411),
	.w2(32'h3a9c2088),
	.w3(32'h3b2b9058),
	.w4(32'hbb1c57ee),
	.w5(32'hb753ad8a),
	.w6(32'hba24d5ae),
	.w7(32'h3af9d96d),
	.w8(32'hb7c74aee),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c8982),
	.w1(32'h38471c0f),
	.w2(32'hb9f49949),
	.w3(32'hb9cdbf97),
	.w4(32'hbb1bca92),
	.w5(32'hbb7ba69a),
	.w6(32'h3a61dea8),
	.w7(32'hbb01e886),
	.w8(32'hbb159683),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb0412),
	.w1(32'h3c8dcf62),
	.w2(32'h3d178c88),
	.w3(32'hbb7e6f07),
	.w4(32'h3a3d034a),
	.w5(32'h3c9042b6),
	.w6(32'h3b90bf3e),
	.w7(32'h3cb92875),
	.w8(32'hba80f1da),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06bb3b),
	.w1(32'h3b5aeb35),
	.w2(32'hbb97ecce),
	.w3(32'hbafcfc8f),
	.w4(32'h3c457353),
	.w5(32'hba1dee9c),
	.w6(32'h378b8ccc),
	.w7(32'hbc30ea94),
	.w8(32'h3b578f85),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84f97e),
	.w1(32'h39ccea92),
	.w2(32'hb88b9f1b),
	.w3(32'h3c7be8c3),
	.w4(32'hbaddfe74),
	.w5(32'hbab62a4c),
	.w6(32'hba181b13),
	.w7(32'hbb00706f),
	.w8(32'hb86810c1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55be0a),
	.w1(32'h3b0dd74d),
	.w2(32'h3a79f671),
	.w3(32'hb9b8e1af),
	.w4(32'h38dd119e),
	.w5(32'h39e634ae),
	.w6(32'h3aaaa8cb),
	.w7(32'h39c648e2),
	.w8(32'h3ab6f527),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b255034),
	.w1(32'hb9e4a402),
	.w2(32'hbab27059),
	.w3(32'h3a9d196a),
	.w4(32'hb9c42c0b),
	.w5(32'hba091965),
	.w6(32'h3aa05fa4),
	.w7(32'h3b07a5b4),
	.w8(32'h3a37319f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf8b65),
	.w1(32'hba4742f4),
	.w2(32'hba41ab99),
	.w3(32'h3a6cecc6),
	.w4(32'hbb195dab),
	.w5(32'h3b139bdc),
	.w6(32'h399377f2),
	.w7(32'h3b05f870),
	.w8(32'h3ae77b78),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac91ead),
	.w1(32'hbaf552e4),
	.w2(32'h3a4bdf15),
	.w3(32'hbbb0df22),
	.w4(32'hbba54732),
	.w5(32'hbb762aec),
	.w6(32'hbb843276),
	.w7(32'hbb345fdc),
	.w8(32'hbb0683de),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac21f00),
	.w1(32'h39c5ed24),
	.w2(32'h396b9092),
	.w3(32'hbb9b830d),
	.w4(32'hbb2749fd),
	.w5(32'h386cc4ad),
	.w6(32'h39ec9199),
	.w7(32'hb9b61b81),
	.w8(32'hbac0ae64),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9686680),
	.w1(32'hbaf279bb),
	.w2(32'hb9df1d12),
	.w3(32'hbaba04fd),
	.w4(32'hbb52cdec),
	.w5(32'hbb1dd977),
	.w6(32'hbb4535c0),
	.w7(32'hba638253),
	.w8(32'hbace6138),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5c170),
	.w1(32'h39847677),
	.w2(32'h3aff0808),
	.w3(32'hbb5b286b),
	.w4(32'h3aa23ad7),
	.w5(32'h3abb9275),
	.w6(32'h392450af),
	.w7(32'h39be9b72),
	.w8(32'h3afffa54),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ae254),
	.w1(32'h3a79fe7f),
	.w2(32'h3a217f1b),
	.w3(32'h3b959298),
	.w4(32'hbb07c84d),
	.w5(32'hbaf5530f),
	.w6(32'h3a54866f),
	.w7(32'h398e73c7),
	.w8(32'hbac0ae92),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39671aa2),
	.w1(32'hb9a947ae),
	.w2(32'hbaae4ce7),
	.w3(32'hb9d17e91),
	.w4(32'hb8ab172c),
	.w5(32'hbaba634a),
	.w6(32'hb91b4efd),
	.w7(32'hbab06810),
	.w8(32'hb9ce3f60),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a375d6),
	.w1(32'h3bfa09b5),
	.w2(32'hbb245988),
	.w3(32'h397c3a1e),
	.w4(32'h3c6faf74),
	.w5(32'hbb209b77),
	.w6(32'h3b826398),
	.w7(32'hbc23ea5b),
	.w8(32'h3bdf60a3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b804a6c),
	.w1(32'h3b42277e),
	.w2(32'hba781751),
	.w3(32'h3c858cd3),
	.w4(32'hb98685a2),
	.w5(32'hbb4e795d),
	.w6(32'h3ac04db2),
	.w7(32'hbaccd966),
	.w8(32'h3a23e1bb),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae18874),
	.w1(32'h3b0c4aa9),
	.w2(32'hb9bdd55a),
	.w3(32'hba4e8840),
	.w4(32'h3a00fb6e),
	.w5(32'hb9b58efd),
	.w6(32'h3b02d8c3),
	.w7(32'h3ac5a81a),
	.w8(32'h3aad40f1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adea5a8),
	.w1(32'hbc5e21ba),
	.w2(32'hbb5eeb00),
	.w3(32'h3a7225de),
	.w4(32'hbc1ea035),
	.w5(32'hbb5b3e36),
	.w6(32'hbc9be941),
	.w7(32'hbc14ecbd),
	.w8(32'hbb868476),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf824e),
	.w1(32'hbb6e9121),
	.w2(32'h3a0f50d7),
	.w3(32'h3ae8eeb4),
	.w4(32'hbb28be1a),
	.w5(32'hba32b771),
	.w6(32'hbb3e2599),
	.w7(32'h39721260),
	.w8(32'h3a9586d4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf8dcc),
	.w1(32'hb990dfa0),
	.w2(32'h3a8177cb),
	.w3(32'h3afbb4c0),
	.w4(32'hbafd4e1b),
	.w5(32'hbab743b0),
	.w6(32'hb9f64c17),
	.w7(32'hba10adc8),
	.w8(32'h3a0b9f1a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac85582),
	.w1(32'h3a2c2e45),
	.w2(32'h3aea4ab1),
	.w3(32'hbae7cd25),
	.w4(32'h3af381a7),
	.w5(32'h39994ea3),
	.w6(32'h3a8c9a69),
	.w7(32'h3abb2e91),
	.w8(32'h3b8cefe3),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f81bd),
	.w1(32'h3c2e8f98),
	.w2(32'h3cb6a4eb),
	.w3(32'hbb37860e),
	.w4(32'hbb19dc2d),
	.w5(32'h3c543dc4),
	.w6(32'h3b06383c),
	.w7(32'h3c498c87),
	.w8(32'h3a16c2c3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8d377),
	.w1(32'h3aa5eb94),
	.w2(32'h39dfb6d9),
	.w3(32'hbac71791),
	.w4(32'hba20bdf6),
	.w5(32'hb8026f69),
	.w6(32'h3a71c5a3),
	.w7(32'h3a777fb5),
	.w8(32'h39765b10),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace05ac),
	.w1(32'hb94c0654),
	.w2(32'h3aa9e2be),
	.w3(32'h3a25cbd6),
	.w4(32'hbae25b10),
	.w5(32'h39bed01e),
	.w6(32'hba92a9bb),
	.w7(32'h39c554d7),
	.w8(32'hb9ce99c9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a475879),
	.w1(32'h3ab6e249),
	.w2(32'h3bc26895),
	.w3(32'h3a9682aa),
	.w4(32'h3aabc9c5),
	.w5(32'h3bbe75da),
	.w6(32'hb9b4fa44),
	.w7(32'h3b50d16c),
	.w8(32'h3ac5d677),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11f67d),
	.w1(32'h3a496b8b),
	.w2(32'h3ad53a3a),
	.w3(32'h3b351970),
	.w4(32'hbb7f734e),
	.w5(32'hbbb25f7a),
	.w6(32'h3abada93),
	.w7(32'h3b20b57a),
	.w8(32'hb9ef3189),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08082e),
	.w1(32'h3a5c8e63),
	.w2(32'hb8d9ec8a),
	.w3(32'hbb008c1a),
	.w4(32'hbac39383),
	.w5(32'hbb2a7edd),
	.w6(32'h38849ba9),
	.w7(32'h39bedc0d),
	.w8(32'h39fc3064),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d3461),
	.w1(32'hbabbd4be),
	.w2(32'hb9312852),
	.w3(32'h3a8c8297),
	.w4(32'hbb416799),
	.w5(32'h38d7a3d5),
	.w6(32'hba5030cc),
	.w7(32'h3b4d7a98),
	.w8(32'h3b938cdd),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f17d6),
	.w1(32'h39963477),
	.w2(32'h3b456dcc),
	.w3(32'hba62d3c9),
	.w4(32'h39b9e14a),
	.w5(32'h3a83dbf7),
	.w6(32'h3b2d3c7e),
	.w7(32'h3b74649e),
	.w8(32'h3b45cd2f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05526c),
	.w1(32'h3aae5ad6),
	.w2(32'h3c97fb13),
	.w3(32'h39465165),
	.w4(32'h3b8e765c),
	.w5(32'h3c961a18),
	.w6(32'hbc01362c),
	.w7(32'h3bd618af),
	.w8(32'h3a5d8bf0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82e4b5),
	.w1(32'h3a973126),
	.w2(32'h3a39faaa),
	.w3(32'h3c4421b7),
	.w4(32'h3bc84e1d),
	.w5(32'h3ad12e3d),
	.w6(32'h3b5d0f41),
	.w7(32'h3a7bc60c),
	.w8(32'h3bbe4c89),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af01769),
	.w1(32'h390aa3dc),
	.w2(32'hba180c5b),
	.w3(32'h3b97b1e9),
	.w4(32'h3a3b7012),
	.w5(32'h3ac2d226),
	.w6(32'hba77895c),
	.w7(32'hbae417cf),
	.w8(32'hbb2b234c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b3cfe),
	.w1(32'hb8e6ed38),
	.w2(32'h3ab042db),
	.w3(32'hbb5fdf3d),
	.w4(32'h38ba89fc),
	.w5(32'h39a71602),
	.w6(32'h3a6b7f2d),
	.w7(32'h3a66649e),
	.w8(32'h3a11570b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b714af),
	.w1(32'h398789c3),
	.w2(32'h38d5283b),
	.w3(32'h3a64bf3e),
	.w4(32'hbb13833a),
	.w5(32'hbaac5f76),
	.w6(32'h37ab4d6a),
	.w7(32'h392777f1),
	.w8(32'hba9d2108),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b27cd),
	.w1(32'hb9fb3da9),
	.w2(32'h3ad0faac),
	.w3(32'hbaadf648),
	.w4(32'hba6af32a),
	.w5(32'h39b1f9aa),
	.w6(32'hb9bc9f97),
	.w7(32'h39c800e9),
	.w8(32'hb8c7766c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c9db5),
	.w1(32'hba0a3b2d),
	.w2(32'hb8eb0efe),
	.w3(32'hb9cc8695),
	.w4(32'hbb08da67),
	.w5(32'hbb118db7),
	.w6(32'hba0f2638),
	.w7(32'hba3d6ca3),
	.w8(32'hba196f2d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369109f1),
	.w1(32'h3a4d0536),
	.w2(32'hbac72520),
	.w3(32'hb921ac21),
	.w4(32'h39fbfc59),
	.w5(32'hbacb99d2),
	.w6(32'h3ad9be9b),
	.w7(32'h3a712a49),
	.w8(32'hbba2ccff),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab4f48),
	.w1(32'hbc09ec03),
	.w2(32'hbb22edf1),
	.w3(32'hbb118d63),
	.w4(32'hbbd3a8d7),
	.w5(32'hbb41604f),
	.w6(32'hbc3e1078),
	.w7(32'hbbbdb2c2),
	.w8(32'hbb4f0138),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac990c5),
	.w1(32'hba2c2d46),
	.w2(32'h3b2423ff),
	.w3(32'h398c5df8),
	.w4(32'hbab8f42a),
	.w5(32'h388deeca),
	.w6(32'h3985081d),
	.w7(32'h3ae1b7e8),
	.w8(32'hbab7907b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb2f4e),
	.w1(32'hbaf7020a),
	.w2(32'hbab97355),
	.w3(32'hbabdd49a),
	.w4(32'hbb03624f),
	.w5(32'h3aa0af59),
	.w6(32'hbad85313),
	.w7(32'hbaeb8099),
	.w8(32'hba4e36b0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb037f74),
	.w1(32'h3b9abd62),
	.w2(32'hba96f28e),
	.w3(32'hbb1bd092),
	.w4(32'h3c874439),
	.w5(32'h3bea7e0a),
	.w6(32'h3b1fc841),
	.w7(32'hbb96ea3d),
	.w8(32'h3bf4448a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d609e),
	.w1(32'h3bbd6e03),
	.w2(32'h3b5225bc),
	.w3(32'h3c81e8b3),
	.w4(32'h3b823538),
	.w5(32'hba669a9f),
	.w6(32'h3b368820),
	.w7(32'hbb48f0ff),
	.w8(32'h3b4668f6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaed905),
	.w1(32'h3b36c9c1),
	.w2(32'h3b27ed62),
	.w3(32'h3b3bec79),
	.w4(32'h38df378f),
	.w5(32'h3a98131c),
	.w6(32'h3b2e48ff),
	.w7(32'h3b42a911),
	.w8(32'h3b24c903),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e0bef),
	.w1(32'hbb16dad9),
	.w2(32'h3b5799de),
	.w3(32'h3aaf55e2),
	.w4(32'hbb9b4854),
	.w5(32'h3a8904fd),
	.w6(32'hbb87f494),
	.w7(32'h35d3ec7b),
	.w8(32'hba902a78),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5502ea),
	.w1(32'hb9df3e1f),
	.w2(32'h3a2e2f2c),
	.w3(32'hba6d34e2),
	.w4(32'hba012e8e),
	.w5(32'h38328bd3),
	.w6(32'hba8878a0),
	.w7(32'hba61ca1d),
	.w8(32'hb9d3036b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38138a5d),
	.w1(32'h3a8af714),
	.w2(32'h39c4a665),
	.w3(32'h3929c83b),
	.w4(32'hbab250b4),
	.w5(32'hba8996df),
	.w6(32'h3a54e0dc),
	.w7(32'h39aba643),
	.w8(32'hb9008243),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9142948),
	.w1(32'h3a1f3e6c),
	.w2(32'h3a0dd4c6),
	.w3(32'hb7c2f28d),
	.w4(32'hbaed94dd),
	.w5(32'hba6ed474),
	.w6(32'h39b9cb20),
	.w7(32'h3a166859),
	.w8(32'hba5c49ec),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d83492),
	.w1(32'h3b29ea34),
	.w2(32'h3af5ca28),
	.w3(32'hba385f50),
	.w4(32'hba364ab1),
	.w5(32'h39670dba),
	.w6(32'h3a8a4527),
	.w7(32'h394a9d3c),
	.w8(32'h3a00c2c1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dc70a),
	.w1(32'h3a46d126),
	.w2(32'h3b6f46d5),
	.w3(32'h3a80b0ba),
	.w4(32'hbac4cc2a),
	.w5(32'hb91203e4),
	.w6(32'h3a2c43d1),
	.w7(32'h3b0638d0),
	.w8(32'hba5a7d8a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba180905),
	.w1(32'hbb1cf146),
	.w2(32'hbb8bb9de),
	.w3(32'hbad352df),
	.w4(32'hbb1b186f),
	.w5(32'h39e78326),
	.w6(32'hbb8fbc34),
	.w7(32'hbb95b34a),
	.w8(32'hbb35e915),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc0cb9),
	.w1(32'hbbb25d05),
	.w2(32'h3a8b3d95),
	.w3(32'hba9e7708),
	.w4(32'hbbf2749c),
	.w5(32'hba5aef92),
	.w6(32'hbbe34bb4),
	.w7(32'hbae5751a),
	.w8(32'hbb49a4eb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac79408),
	.w1(32'hb9f1ad80),
	.w2(32'h3b1834fb),
	.w3(32'hba667bc2),
	.w4(32'hbaa8a756),
	.w5(32'h3b157e31),
	.w6(32'hb8a905e3),
	.w7(32'h3a61d284),
	.w8(32'hbb321c28),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4112a3),
	.w1(32'h3a7f784a),
	.w2(32'h3af37d78),
	.w3(32'hbb19edf5),
	.w4(32'h397326ed),
	.w5(32'h3b0ad253),
	.w6(32'h3b287d5f),
	.w7(32'h3b6f6f78),
	.w8(32'hb9f2cb2e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f3548),
	.w1(32'h39c23bf3),
	.w2(32'hba50ebf6),
	.w3(32'hb81057e9),
	.w4(32'hbafbde66),
	.w5(32'hbafc3960),
	.w6(32'hba74fab9),
	.w7(32'hbae6af07),
	.w8(32'h39ff90eb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11c04b),
	.w1(32'h3baef7cc),
	.w2(32'h3c407f2a),
	.w3(32'hb9cab517),
	.w4(32'h3b28063d),
	.w5(32'h3bcf0fe7),
	.w6(32'hba694d09),
	.w7(32'h3afc7a66),
	.w8(32'h3b448f05),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ab3be),
	.w1(32'h3af5a4c3),
	.w2(32'hba16a445),
	.w3(32'h3ba2b2f6),
	.w4(32'h3b011cbb),
	.w5(32'hbaa14160),
	.w6(32'h3b243cdd),
	.w7(32'h39a70d6e),
	.w8(32'h3b0c44d9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a606a71),
	.w1(32'h3b9b744c),
	.w2(32'h3bda9964),
	.w3(32'h3b00fb8e),
	.w4(32'h39df2d26),
	.w5(32'h3b14c320),
	.w6(32'h39e6f70a),
	.w7(32'h3ad9c588),
	.w8(32'h38ed03b9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ad337),
	.w1(32'hba8eef98),
	.w2(32'hb8e4c9c9),
	.w3(32'h3b697ad3),
	.w4(32'hba160b82),
	.w5(32'hb989e026),
	.w6(32'hb7c02288),
	.w7(32'h398152d1),
	.w8(32'h392f5c86),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cdfa5d),
	.w1(32'h3baca6c4),
	.w2(32'h3c02fb4d),
	.w3(32'h38f67a47),
	.w4(32'h3953b9fa),
	.w5(32'h3bcfb7ef),
	.w6(32'hbb0afbaf),
	.w7(32'hba348980),
	.w8(32'hbb8083a5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2dc12),
	.w1(32'h3abb7857),
	.w2(32'h3a4a60c2),
	.w3(32'h389683f8),
	.w4(32'h3be23f82),
	.w5(32'h3b922631),
	.w6(32'h3ab0c16d),
	.w7(32'h3960e527),
	.w8(32'h3b83ca77),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c603d),
	.w1(32'h3a80cf2b),
	.w2(32'h3b1c75b8),
	.w3(32'h3bfe5b0c),
	.w4(32'h39e5ccb6),
	.w5(32'h3af76a0d),
	.w6(32'hb977cda8),
	.w7(32'h3ad2265f),
	.w8(32'h389da2cd),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ccce4),
	.w1(32'h3a975465),
	.w2(32'h3a1b4255),
	.w3(32'hba13c1c7),
	.w4(32'hba22fb2c),
	.w5(32'hb9fbf87a),
	.w6(32'hb9e78faa),
	.w7(32'hba8b9456),
	.w8(32'h397e21cf),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5b964),
	.w1(32'h3b09614e),
	.w2(32'h3b800107),
	.w3(32'h3a1995dc),
	.w4(32'h3af03395),
	.w5(32'h3ac6a01f),
	.w6(32'h3b6a5701),
	.w7(32'h3b8c5118),
	.w8(32'h3bae740c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c1ae2),
	.w1(32'h3b238a88),
	.w2(32'h3b13f777),
	.w3(32'h3b12a2f7),
	.w4(32'h399279c8),
	.w5(32'h3aa13ef0),
	.w6(32'h3aa8b4b0),
	.w7(32'h382d9a64),
	.w8(32'h3b0ed4cf),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24cfd7),
	.w1(32'h3b40a282),
	.w2(32'h3887b7cf),
	.w3(32'h3a9ca196),
	.w4(32'hb987913a),
	.w5(32'hbaf3ba9d),
	.w6(32'h3a2dba48),
	.w7(32'hbb12dab9),
	.w8(32'hba2b8cf3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99046a),
	.w1(32'hbba89963),
	.w2(32'hba713655),
	.w3(32'hba35ccc9),
	.w4(32'hba2cf39e),
	.w5(32'h3b07a655),
	.w6(32'hbbba15ef),
	.w7(32'hbb11d83f),
	.w8(32'h3b242bc2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3faa0f),
	.w1(32'hb9877d83),
	.w2(32'h3987fea2),
	.w3(32'h3bb61922),
	.w4(32'hbae0d8f8),
	.w5(32'hbafd5c38),
	.w6(32'hbaf624a7),
	.w7(32'hba428009),
	.w8(32'hba49a415),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a10dc),
	.w1(32'h3bc9ed3c),
	.w2(32'h3cc546e3),
	.w3(32'hba31fd8c),
	.w4(32'h3ad69dcc),
	.w5(32'h3c657f59),
	.w6(32'hb98428a8),
	.w7(32'h3c7f6f90),
	.w8(32'hba2c739b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab756e0),
	.w1(32'h3b2a8b9a),
	.w2(32'h3b696e8a),
	.w3(32'h3a5fdf8a),
	.w4(32'hb98ff91f),
	.w5(32'hba88408a),
	.w6(32'h3b33e544),
	.w7(32'h3b135b0b),
	.w8(32'h3b068700),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b227cdc),
	.w1(32'h3b2c1384),
	.w2(32'hb9bec286),
	.w3(32'hba828597),
	.w4(32'hb98bc231),
	.w5(32'hba905796),
	.w6(32'h3a6264ce),
	.w7(32'hbb1b2dd4),
	.w8(32'h3a84524b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b2377),
	.w1(32'h3c21a738),
	.w2(32'h3c533161),
	.w3(32'hbb0323ec),
	.w4(32'h3b074cde),
	.w5(32'h3c0a5215),
	.w6(32'h3c2aa3dd),
	.w7(32'h3c277d25),
	.w8(32'h3a9b6714),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9391d5),
	.w1(32'h3b06f126),
	.w2(32'hbb83c776),
	.w3(32'hbb871e32),
	.w4(32'h39efef92),
	.w5(32'hbc433bb5),
	.w6(32'h3a4662ca),
	.w7(32'hbc021152),
	.w8(32'hbb00a0d4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5538eb),
	.w1(32'h3aae57a7),
	.w2(32'hb9d4d4e9),
	.w3(32'hbb9460da),
	.w4(32'h38575a40),
	.w5(32'hbafce7f1),
	.w6(32'h3abc7e10),
	.w7(32'hba108d7e),
	.w8(32'h3b07a6aa),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba588602),
	.w1(32'h3ab6e33f),
	.w2(32'hb9b14744),
	.w3(32'h39bda885),
	.w4(32'hbab75e3e),
	.w5(32'hbb29ddec),
	.w6(32'hbb2f4138),
	.w7(32'hbac88436),
	.w8(32'hbab0a49f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac32f0e),
	.w1(32'hba11f994),
	.w2(32'hbb9ef8c3),
	.w3(32'hbb030280),
	.w4(32'h3aae4753),
	.w5(32'hbb868b57),
	.w6(32'hba642565),
	.w7(32'hbb9baa4d),
	.w8(32'hbb17056a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7527d6),
	.w1(32'h3a85fc3d),
	.w2(32'hbb5db2e2),
	.w3(32'hbb837900),
	.w4(32'hbb14565c),
	.w5(32'hbb1f95ab),
	.w6(32'h3ac82c6a),
	.w7(32'hb9c2c841),
	.w8(32'hbaa25afc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a9c85a),
	.w1(32'hbbe026ec),
	.w2(32'h3a997537),
	.w3(32'hb98172dc),
	.w4(32'hbc1a9b09),
	.w5(32'hba9b709f),
	.w6(32'hbc20037c),
	.w7(32'hbb28fcef),
	.w8(32'hbb9b9e61),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30bfff),
	.w1(32'h3a1f72b9),
	.w2(32'h3b016822),
	.w3(32'hb8e181e9),
	.w4(32'hbab1d930),
	.w5(32'h3994336b),
	.w6(32'h3a4c35c9),
	.w7(32'h3aa34a71),
	.w8(32'h396d8007),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13f54f),
	.w1(32'hbb92d511),
	.w2(32'h39e9a65f),
	.w3(32'hba809bfe),
	.w4(32'hbbad4744),
	.w5(32'hba5f17d9),
	.w6(32'hbbb2df86),
	.w7(32'hbaa7e8bb),
	.w8(32'hbad4b7fe),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9afcb),
	.w1(32'hba9bdc76),
	.w2(32'hb9f58e60),
	.w3(32'hba3b3b7c),
	.w4(32'hbb68e220),
	.w5(32'hba6b3472),
	.w6(32'hba8ac550),
	.w7(32'h392f818d),
	.w8(32'hbb2d3fb0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4edaa),
	.w1(32'h3ae87dc7),
	.w2(32'h3a85fce4),
	.w3(32'hbb1368ed),
	.w4(32'hbb0537d1),
	.w5(32'hbb81fc04),
	.w6(32'h3b22740d),
	.w7(32'h3a59f8df),
	.w8(32'h39de0c5b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cea30),
	.w1(32'h3b633124),
	.w2(32'h3ab8d593),
	.w3(32'hbb471579),
	.w4(32'hba612267),
	.w5(32'hbb2065d9),
	.w6(32'hb9b0a83c),
	.w7(32'hbb56b053),
	.w8(32'hba18dfc7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08f11f),
	.w1(32'hbb64e8cd),
	.w2(32'h3a2ba8ff),
	.w3(32'hba9258bf),
	.w4(32'hbbaedbe8),
	.w5(32'hba5a83c6),
	.w6(32'hbbab7516),
	.w7(32'hbb023714),
	.w8(32'hbb27b529),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba863316),
	.w1(32'hb9ef634d),
	.w2(32'h3ab4077f),
	.w3(32'hb98251d4),
	.w4(32'hbac1abc6),
	.w5(32'h3a1c08c6),
	.w6(32'hb928c024),
	.w7(32'h3a698e25),
	.w8(32'hba909012),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ecf6b),
	.w1(32'h3adb2309),
	.w2(32'h3b78da2d),
	.w3(32'h3a671236),
	.w4(32'hbb0fa3df),
	.w5(32'h3a8e5cb4),
	.w6(32'h3aa716df),
	.w7(32'h3b5b558a),
	.w8(32'h397e6e97),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0099ad),
	.w1(32'hbb5e5061),
	.w2(32'hb989e902),
	.w3(32'h38c6383b),
	.w4(32'hbba3f25a),
	.w5(32'hbb1e133b),
	.w6(32'hbbb0a219),
	.w7(32'hbab5d9ab),
	.w8(32'hbb6feba0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbdacb),
	.w1(32'h3b171fcc),
	.w2(32'h3b594520),
	.w3(32'hba12c20c),
	.w4(32'hba8120b9),
	.w5(32'h3a9b83ca),
	.w6(32'h3b1dda03),
	.w7(32'h3b7eb0f7),
	.w8(32'h3aa76943),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b023b66),
	.w1(32'h3b090211),
	.w2(32'h3b20f662),
	.w3(32'h3ab02178),
	.w4(32'h3a0c02d8),
	.w5(32'h392eec22),
	.w6(32'h3ac2dc00),
	.w7(32'h3a90b703),
	.w8(32'hb9cb7333),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addbf82),
	.w1(32'h3b174d96),
	.w2(32'h3b3598c3),
	.w3(32'hba11eb09),
	.w4(32'h3903d26e),
	.w5(32'h3b534262),
	.w6(32'h3b1c78cd),
	.w7(32'h3ba56007),
	.w8(32'h3aa66665),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79cfc1),
	.w1(32'hbba25178),
	.w2(32'h3a7db3c3),
	.w3(32'h3acee86d),
	.w4(32'hbbecc2e7),
	.w5(32'hba989e0f),
	.w6(32'hbbf2dcb0),
	.w7(32'hbb0e2415),
	.w8(32'hbb846566),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08f313),
	.w1(32'hba59a15a),
	.w2(32'hb9738143),
	.w3(32'hb975ba14),
	.w4(32'hbb4dd0b6),
	.w5(32'hbb18ddfb),
	.w6(32'hbb14233c),
	.w7(32'hbaf2c7a0),
	.w8(32'hbb4930a9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf9f6d),
	.w1(32'hba92652b),
	.w2(32'hb88b3b58),
	.w3(32'hbab0b47f),
	.w4(32'hbb944197),
	.w5(32'hbb41e1a2),
	.w6(32'hbb3a1212),
	.w7(32'hbacd3e54),
	.w8(32'hbb7cca1a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb118aa9),
	.w1(32'hba953bfa),
	.w2(32'hbad96faf),
	.w3(32'hbb0cf1b6),
	.w4(32'hbb88b894),
	.w5(32'hbbd31b46),
	.w6(32'h3789a5e9),
	.w7(32'hbb02876c),
	.w8(32'hbb37036a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f24a26),
	.w1(32'h39bfa01a),
	.w2(32'h3c2db46a),
	.w3(32'hbb53a58c),
	.w4(32'hbb280c81),
	.w5(32'h3c1e7110),
	.w6(32'hba92aca8),
	.w7(32'h3bed690e),
	.w8(32'hbb40308d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71ed16),
	.w1(32'h3ac73f0a),
	.w2(32'h3b3bfd66),
	.w3(32'hbbcd27b7),
	.w4(32'hbb56b6fe),
	.w5(32'h3a003a17),
	.w6(32'h39982ad7),
	.w7(32'h3ae07def),
	.w8(32'hba5e203b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a824cf),
	.w1(32'h3a99301f),
	.w2(32'h39cde4db),
	.w3(32'hbb189aa5),
	.w4(32'hbb35a2e4),
	.w5(32'hbb2c3af9),
	.w6(32'h3a64e63c),
	.w7(32'h3aa63eac),
	.w8(32'hba40e18c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb974d7ca),
	.w1(32'h3793e335),
	.w2(32'h3a52c9c5),
	.w3(32'hbb3690e4),
	.w4(32'hbb4ae3b5),
	.w5(32'hbaaee986),
	.w6(32'hb97ddc86),
	.w7(32'hba6dec02),
	.w8(32'hba957d88),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9521ed0),
	.w1(32'h3962fa6b),
	.w2(32'hba57de80),
	.w3(32'hb99f038f),
	.w4(32'hbaea9d86),
	.w5(32'hbb2f6a67),
	.w6(32'hbad23729),
	.w7(32'hbb49a90f),
	.w8(32'hbb5486ad),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a35d3),
	.w1(32'h3b0a5769),
	.w2(32'hbaba1940),
	.w3(32'hbb0dc722),
	.w4(32'hbad51d16),
	.w5(32'hbb87d196),
	.w6(32'hba0c47c3),
	.w7(32'hbb00ca7d),
	.w8(32'hbb01f9a9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c50cf),
	.w1(32'h3b0d6ccf),
	.w2(32'h3a60c9cf),
	.w3(32'hba67fe20),
	.w4(32'hbb49c2cc),
	.w5(32'hbadb47db),
	.w6(32'hbae28587),
	.w7(32'hbad6c2ea),
	.w8(32'hbab12b09),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe04db),
	.w1(32'h3acd5f7f),
	.w2(32'h3b587a1e),
	.w3(32'hba5fdb57),
	.w4(32'h3a986843),
	.w5(32'h3af1164e),
	.w6(32'hb98581fa),
	.w7(32'hba3d5f27),
	.w8(32'h3a2b579b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add596e),
	.w1(32'h3a90c76f),
	.w2(32'h3a9396d1),
	.w3(32'h3a5b9bef),
	.w4(32'h3a6b7a12),
	.w5(32'h3a99ccd1),
	.w6(32'h3abea635),
	.w7(32'h3a86dd33),
	.w8(32'h3b0a1376),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a526ed1),
	.w1(32'hb9a75ee2),
	.w2(32'hbb1ee7b9),
	.w3(32'h3a33bcfb),
	.w4(32'h3b0e51eb),
	.w5(32'h37ab7446),
	.w6(32'hbafa0310),
	.w7(32'hba42ee95),
	.w8(32'h3a94274e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d7809),
	.w1(32'hbac0ba0c),
	.w2(32'hbb50220a),
	.w3(32'h3ac7c97a),
	.w4(32'hba19f09d),
	.w5(32'hbb3f3c7a),
	.w6(32'hba3b13d8),
	.w7(32'hbafa9dc0),
	.w8(32'hb95f615e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba863a63),
	.w1(32'h3ac6bbf6),
	.w2(32'h3b801266),
	.w3(32'hb9468bcf),
	.w4(32'hba6c81bd),
	.w5(32'hba1a00b3),
	.w6(32'h3b02cd71),
	.w7(32'hb9e66ffe),
	.w8(32'hbb455e36),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b756cd),
	.w1(32'h3a454deb),
	.w2(32'h3ba771e2),
	.w3(32'hbb04e65d),
	.w4(32'h3b4d5470),
	.w5(32'hb811fe54),
	.w6(32'h3b9ce655),
	.w7(32'h3bd40c67),
	.w8(32'h3b38f895),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55fdbb),
	.w1(32'hbb3a7568),
	.w2(32'h3b320aec),
	.w3(32'hbb533ef0),
	.w4(32'hbb525481),
	.w5(32'h3b2a0b58),
	.w6(32'hbb61ed7a),
	.w7(32'hbabc32bb),
	.w8(32'hbb216cff),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac88b5e),
	.w1(32'h3b6af2d6),
	.w2(32'h3b4d8ecd),
	.w3(32'h3a515960),
	.w4(32'h38dc5c9d),
	.w5(32'h3a9ce31b),
	.w6(32'h3b6266ee),
	.w7(32'h3ba5f254),
	.w8(32'h3b41f2ea),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a823ea9),
	.w1(32'h3aa5c786),
	.w2(32'h3a93ac95),
	.w3(32'h3a6e9ca6),
	.w4(32'h3b00f42b),
	.w5(32'h3b101b5d),
	.w6(32'h3a1e7d97),
	.w7(32'h3a03c71d),
	.w8(32'h3b4c79e0),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c68cf),
	.w1(32'h3aeeb3f1),
	.w2(32'hb6d98b58),
	.w3(32'h3aac4df9),
	.w4(32'h3a841410),
	.w5(32'hb9c3b8ea),
	.w6(32'h3afb3d2d),
	.w7(32'hb975b147),
	.w8(32'h39fb98bf),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcc465),
	.w1(32'h3a856a79),
	.w2(32'h3b687ccc),
	.w3(32'hb68477fe),
	.w4(32'hb9979e59),
	.w5(32'h3b902aad),
	.w6(32'h3ad3cdab),
	.w7(32'h3b3703da),
	.w8(32'h3b56bae1),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5b6b4),
	.w1(32'h38c7de28),
	.w2(32'h3abea58b),
	.w3(32'h3ad57901),
	.w4(32'hbb22e1c2),
	.w5(32'hbac68063),
	.w6(32'h3b78cd8a),
	.w7(32'h3b90d3c9),
	.w8(32'h3a1eec01),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb141a23),
	.w1(32'hb9f27253),
	.w2(32'hbbb1c49e),
	.w3(32'hba2b9161),
	.w4(32'hbb782c11),
	.w5(32'hbc013729),
	.w6(32'h3ad49b0c),
	.w7(32'hbb9cf3c7),
	.w8(32'hbbb71f79),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4629f),
	.w1(32'h3bbe69c8),
	.w2(32'hbab6d017),
	.w3(32'hbbf94cbb),
	.w4(32'h3b4f0a79),
	.w5(32'hbacb8706),
	.w6(32'h3bf040b5),
	.w7(32'hba557522),
	.w8(32'h3a6fe249),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba561992),
	.w1(32'hbac1d288),
	.w2(32'hbb0ff51b),
	.w3(32'hbb2892c1),
	.w4(32'hbadf9f46),
	.w5(32'hbb117687),
	.w6(32'hbb0add75),
	.w7(32'hbb34c9ba),
	.w8(32'hbb31cdf7),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6889c2),
	.w1(32'h3b89f8a0),
	.w2(32'hba8a32c8),
	.w3(32'hbb04e51c),
	.w4(32'h3ab5a065),
	.w5(32'hbb3d88ab),
	.w6(32'h3b876a3e),
	.w7(32'hb80d249e),
	.w8(32'hba5ed38e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba917cb6),
	.w1(32'h3951d5c5),
	.w2(32'hbb153c2b),
	.w3(32'hba570746),
	.w4(32'h3ad7ea12),
	.w5(32'h3a25a970),
	.w6(32'h3823c478),
	.w7(32'hba7de6a7),
	.w8(32'h3a909cbe),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e32a5),
	.w1(32'h3a3d869c),
	.w2(32'hb98098ac),
	.w3(32'h3941acca),
	.w4(32'h3a3b3382),
	.w5(32'h39a4a4f0),
	.w6(32'h3af4dc98),
	.w7(32'h39acf861),
	.w8(32'h3a8cbe3a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98328ce),
	.w1(32'h3b772378),
	.w2(32'h3c9efd56),
	.w3(32'hba2fe7c8),
	.w4(32'hbc3308d5),
	.w5(32'h3c8e77e4),
	.w6(32'hbc932a72),
	.w7(32'h3bc3f1d5),
	.w8(32'hbc78deed),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a019e),
	.w1(32'hbaf59991),
	.w2(32'h3a20863c),
	.w3(32'h3bf85479),
	.w4(32'h39ab661e),
	.w5(32'hb98294dd),
	.w6(32'hb9a77a00),
	.w7(32'h39620f5c),
	.w8(32'h3b26b131),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2a6ad),
	.w1(32'hbabf615c),
	.w2(32'h39203468),
	.w3(32'h3b20f447),
	.w4(32'hbacf612c),
	.w5(32'hbaa2d626),
	.w6(32'hba903974),
	.w7(32'hba95a310),
	.w8(32'hba20723b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e50128),
	.w1(32'hba29d3eb),
	.w2(32'h39e25c8d),
	.w3(32'hbb28d81e),
	.w4(32'hbb1193dc),
	.w5(32'h3a5cd37e),
	.w6(32'h3a288fc3),
	.w7(32'h3a7bddc5),
	.w8(32'h3afb2833),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb17d2),
	.w1(32'h3a9a0a61),
	.w2(32'h3afc471c),
	.w3(32'hba9b93c8),
	.w4(32'h3aaa40aa),
	.w5(32'h3a829cf1),
	.w6(32'hbb17fed6),
	.w7(32'hbab42236),
	.w8(32'h3aac3f0e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81eb20),
	.w1(32'hb9faff54),
	.w2(32'hbb792f2d),
	.w3(32'hb8b6b0ae),
	.w4(32'hbb884e41),
	.w5(32'hbbf8b9c4),
	.w6(32'hba8edfa4),
	.w7(32'hbb106155),
	.w8(32'h3a2145e5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e69c9),
	.w1(32'h3bb8b57d),
	.w2(32'h3c849289),
	.w3(32'hbbccbd44),
	.w4(32'hbc0dc4bc),
	.w5(32'hbb18e3f9),
	.w6(32'hbb521720),
	.w7(32'h3b274421),
	.w8(32'hbb4bb320),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b0cdd),
	.w1(32'h3a7d74e9),
	.w2(32'hb9deb6ea),
	.w3(32'hbc4a1a2f),
	.w4(32'h3a924d5b),
	.w5(32'h38a7c93a),
	.w6(32'h3abcaed9),
	.w7(32'hb9f8d841),
	.w8(32'h3ab97313),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4491b1),
	.w1(32'h3af1ab6f),
	.w2(32'h3ae9c088),
	.w3(32'h3a1d7278),
	.w4(32'h3a5d64b9),
	.w5(32'h3b3e071f),
	.w6(32'hb9c6df2f),
	.w7(32'hb957dda1),
	.w8(32'hbb28702b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7f87a),
	.w1(32'h3bf200cf),
	.w2(32'hbae6b9eb),
	.w3(32'h3af80ed9),
	.w4(32'hbc6de406),
	.w5(32'h3b2e4115),
	.w6(32'hbb80d4ca),
	.w7(32'hbc17e582),
	.w8(32'hbcaceb86),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58b810),
	.w1(32'hba7f6678),
	.w2(32'hbb0bc965),
	.w3(32'hbb204439),
	.w4(32'hbb0c96cf),
	.w5(32'hbaab47c5),
	.w6(32'hb96cb97f),
	.w7(32'hba4bc001),
	.w8(32'hba01d2ff),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb233e2d),
	.w1(32'hbb129b9f),
	.w2(32'h3a675d98),
	.w3(32'hbb3053b3),
	.w4(32'hba5dfa7a),
	.w5(32'hbaeb5e79),
	.w6(32'h3b2c25f7),
	.w7(32'h3aa40e3e),
	.w8(32'h3a862701),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86bdca),
	.w1(32'hbabb8364),
	.w2(32'h3b88f74c),
	.w3(32'hb959cdff),
	.w4(32'hbb9adddc),
	.w5(32'hba3fda20),
	.w6(32'hbc258efa),
	.w7(32'h3aabce1e),
	.w8(32'hba81806d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb25eb9),
	.w1(32'hbbb9051b),
	.w2(32'h3c876810),
	.w3(32'hbae31714),
	.w4(32'h3c1c749e),
	.w5(32'h3cdd94cf),
	.w6(32'hbcca5af5),
	.w7(32'h3b4f4f33),
	.w8(32'h3bbdf2fb),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c955534),
	.w1(32'hba98acd8),
	.w2(32'hbb0cfb0f),
	.w3(32'h3d029ed8),
	.w4(32'h3960e058),
	.w5(32'hba5d68a3),
	.w6(32'hbb0483b7),
	.w7(32'hbb3397dd),
	.w8(32'hb9f00ad5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9043ae9),
	.w1(32'h3a84844b),
	.w2(32'h3939735c),
	.w3(32'hba25d04f),
	.w4(32'hba29b537),
	.w5(32'hba51250a),
	.w6(32'hbad0dc34),
	.w7(32'hbacab8f3),
	.w8(32'hbab306f9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb810be5f),
	.w1(32'hbc0b8bb5),
	.w2(32'hbaa2e6b4),
	.w3(32'hbaf4d197),
	.w4(32'hbc448639),
	.w5(32'hbb9ff102),
	.w6(32'hbb31b014),
	.w7(32'h3b3fa040),
	.w8(32'hbb0dc3db),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52698c),
	.w1(32'hbb230707),
	.w2(32'hbbdc5ba0),
	.w3(32'hbb218618),
	.w4(32'h3b6b820a),
	.w5(32'hbb70334d),
	.w6(32'hb992685c),
	.w7(32'h3b0e497d),
	.w8(32'hb9ae9be0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e8f6f),
	.w1(32'h3b1e3ba6),
	.w2(32'h3b2129a2),
	.w3(32'hbc51a9cc),
	.w4(32'h3a992bbd),
	.w5(32'h3a993c22),
	.w6(32'h3aeb03c8),
	.w7(32'h3b1cfbd8),
	.w8(32'h3a386104),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d4d26),
	.w1(32'hb807c3bd),
	.w2(32'hbb410ac6),
	.w3(32'h3afbeb7b),
	.w4(32'hba2da3e3),
	.w5(32'hbaa13473),
	.w6(32'h3a36093e),
	.w7(32'hbaef8228),
	.w8(32'hb9bcda3e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae01a35),
	.w1(32'hbb08533d),
	.w2(32'h3812a063),
	.w3(32'hbaa234d7),
	.w4(32'hbab329f2),
	.w5(32'h3ae30ef5),
	.w6(32'hbb0fbbdb),
	.w7(32'hba339340),
	.w8(32'h3a70470d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370fa0ba),
	.w1(32'hb8fe0ecc),
	.w2(32'h39e3399d),
	.w3(32'h3ab9c172),
	.w4(32'h3aeaf956),
	.w5(32'h3a831835),
	.w6(32'hb921eb95),
	.w7(32'h39850a8d),
	.w8(32'h3a7f06b8),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eedcd0),
	.w1(32'h3ab24881),
	.w2(32'h394dec6f),
	.w3(32'h3ade6be1),
	.w4(32'h3ae74afa),
	.w5(32'h3a192ce0),
	.w6(32'h3b04c9cc),
	.w7(32'h3a3a1ec9),
	.w8(32'h3b262646),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4be3a),
	.w1(32'h3a236f82),
	.w2(32'hb9d7203c),
	.w3(32'h3ad1a0f0),
	.w4(32'h3adc3789),
	.w5(32'h39de6999),
	.w6(32'h3aab6672),
	.w7(32'hb7a5b1f0),
	.w8(32'h39b08033),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac306ae),
	.w1(32'hbc843b02),
	.w2(32'h3bd10e91),
	.w3(32'hba36e1de),
	.w4(32'h3c44e594),
	.w5(32'h3cb4d0f7),
	.w6(32'hbcea2cd8),
	.w7(32'h3b61a96b),
	.w8(32'h3c042901),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26c562),
	.w1(32'h3aec8b12),
	.w2(32'h3ae27c3c),
	.w3(32'h3ce5ad6a),
	.w4(32'h3a99de79),
	.w5(32'h3ab41679),
	.w6(32'h3b0832eb),
	.w7(32'h3a1b96cc),
	.w8(32'h3a9564b2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28d8f2),
	.w1(32'hbb2e942f),
	.w2(32'hba377731),
	.w3(32'h39bc775a),
	.w4(32'hbb8f89bd),
	.w5(32'hbacfbfa6),
	.w6(32'hbb64aaae),
	.w7(32'hbaa7f0be),
	.w8(32'hbb30dd92),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab59f8c),
	.w1(32'h3a999bc7),
	.w2(32'h3a06bdff),
	.w3(32'hbb4798db),
	.w4(32'hbb75c3b2),
	.w5(32'hbbb25376),
	.w6(32'h3b740792),
	.w7(32'h3b99e2fa),
	.w8(32'h3a70edf6),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8acb2),
	.w1(32'h3ab75ef4),
	.w2(32'h3b11db66),
	.w3(32'hb9694b86),
	.w4(32'h3b88e93d),
	.w5(32'h3b297f53),
	.w6(32'h3b78b14c),
	.w7(32'h3bb6dde1),
	.w8(32'h3a0f5d40),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb520b28),
	.w1(32'hbaf24e6d),
	.w2(32'hbaa0e502),
	.w3(32'hbacbe765),
	.w4(32'h3a5f6a0c),
	.w5(32'hbaeaadf6),
	.w6(32'h3a6b8374),
	.w7(32'hba4a5c7b),
	.w8(32'h3a052e49),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae760f7),
	.w1(32'hb9030e49),
	.w2(32'hbb2927d2),
	.w3(32'hba8947d2),
	.w4(32'hb91de6bc),
	.w5(32'hb8909538),
	.w6(32'hbac0d100),
	.w7(32'hbb30eeec),
	.w8(32'h3adf78eb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d26cc),
	.w1(32'h3bd886c0),
	.w2(32'h3cb20673),
	.w3(32'hbab61785),
	.w4(32'hbafb6883),
	.w5(32'h3c804d99),
	.w6(32'hbbfe8bb8),
	.w7(32'h3c68cd89),
	.w8(32'h3ad0949a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bcafa),
	.w1(32'hbb2b1993),
	.w2(32'hbacf2e2c),
	.w3(32'hba658bc2),
	.w4(32'hbb8fefa3),
	.w5(32'hbad7a568),
	.w6(32'hbb4b1186),
	.w7(32'hbac67c3b),
	.w8(32'hbb1ef3a5),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf38b75),
	.w1(32'h39961368),
	.w2(32'hbb229f35),
	.w3(32'hbb552126),
	.w4(32'h3a63186e),
	.w5(32'hbb0cd101),
	.w6(32'h3a125e57),
	.w7(32'hbb280cb4),
	.w8(32'hb9dd8780),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59a8a8),
	.w1(32'h3b56e6f3),
	.w2(32'h3924b518),
	.w3(32'hba016b25),
	.w4(32'h3a68844b),
	.w5(32'hbb15b038),
	.w6(32'h3b9bf4b4),
	.w7(32'hb9803ac9),
	.w8(32'hb9f5be11),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7c5c6),
	.w1(32'h3b25cecd),
	.w2(32'hbaa265a5),
	.w3(32'hbaf01f6f),
	.w4(32'h38aac61e),
	.w5(32'hbbb68cad),
	.w6(32'h3b63f941),
	.w7(32'hba871e35),
	.w8(32'h3b299351),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38e2a5),
	.w1(32'h3ae37a9a),
	.w2(32'h397c1db0),
	.w3(32'hbaaa927f),
	.w4(32'hbab76868),
	.w5(32'hbaa4afe1),
	.w6(32'hba658e7e),
	.w7(32'h3aaa15ee),
	.w8(32'hb9c3b4b3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc3997),
	.w1(32'hb9771a6f),
	.w2(32'h3b8c4abe),
	.w3(32'hbb221801),
	.w4(32'hba9eb042),
	.w5(32'h3bba98b2),
	.w6(32'h3b1e4a57),
	.w7(32'h3b244dd5),
	.w8(32'h39e7ffcd),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f4c785),
	.w1(32'h3aa615ae),
	.w2(32'h3c03e0cd),
	.w3(32'hb92cff52),
	.w4(32'hbbe06982),
	.w5(32'h3b6f926d),
	.w6(32'hbb7e0d0b),
	.w7(32'h3add0bd8),
	.w8(32'hbc4a8110),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8567b2),
	.w1(32'hbd0ea154),
	.w2(32'hbcd48e3f),
	.w3(32'hbbc5712d),
	.w4(32'h3af936f7),
	.w5(32'h3a0ac7d2),
	.w6(32'hbd08413e),
	.w7(32'hbcaa3170),
	.w8(32'h3c7f2bd0),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b553a07),
	.w1(32'hbbc25f63),
	.w2(32'hba3ba313),
	.w3(32'h3ce87bca),
	.w4(32'hbb5ba53b),
	.w5(32'hbb67407c),
	.w6(32'hbbe82288),
	.w7(32'hb9f8d59c),
	.w8(32'hbad35ccd),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0db770),
	.w1(32'h3b039c64),
	.w2(32'h3af46e41),
	.w3(32'hbb9c2656),
	.w4(32'h39ed9fec),
	.w5(32'hb95842b0),
	.w6(32'h3b7a1c68),
	.w7(32'h3abf8417),
	.w8(32'h3b818fd0),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb5332),
	.w1(32'h3ac38b3e),
	.w2(32'hbab7283a),
	.w3(32'h3a540ebe),
	.w4(32'h3b086cdd),
	.w5(32'hbb055150),
	.w6(32'h3b2dcb93),
	.w7(32'h3aadb3e8),
	.w8(32'h3b329243),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac49d58),
	.w1(32'h3abcd5aa),
	.w2(32'h3ac7e5eb),
	.w3(32'hbb2eb0ce),
	.w4(32'h3a9fb688),
	.w5(32'h3b3d53ed),
	.w6(32'h3abebed7),
	.w7(32'h3ad44cf4),
	.w8(32'h3b914c04),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16171e),
	.w1(32'hbb02f9fa),
	.w2(32'hbb1bbeba),
	.w3(32'h3ad4e7ac),
	.w4(32'hb98c5e37),
	.w5(32'hba3185d7),
	.w6(32'h3a491d0b),
	.w7(32'hbb0712af),
	.w8(32'hbae46755),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389c60ab),
	.w1(32'hbab35085),
	.w2(32'hba38e36a),
	.w3(32'hb947c05f),
	.w4(32'h3991bddc),
	.w5(32'h3a0b183c),
	.w6(32'h3a347b31),
	.w7(32'hb9247161),
	.w8(32'h3a2782cb),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a092b94),
	.w1(32'h3adb781e),
	.w2(32'h3ac7e190),
	.w3(32'h3a91c816),
	.w4(32'h38f8e390),
	.w5(32'hbafcba72),
	.w6(32'h3a874cca),
	.w7(32'h3ac336be),
	.w8(32'h3a02a105),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55fd62),
	.w1(32'h3a598df6),
	.w2(32'h39897e80),
	.w3(32'hba24628a),
	.w4(32'hbb1dc38e),
	.w5(32'hbb62df64),
	.w6(32'h3b36b8b3),
	.w7(32'h3b5378cf),
	.w8(32'h39dde01a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb636cbd),
	.w1(32'hba9715f6),
	.w2(32'h3a29c7ab),
	.w3(32'h37ecf0bc),
	.w4(32'hbab20133),
	.w5(32'hbad592ca),
	.w6(32'h3884cbb9),
	.w7(32'h3acfc8ab),
	.w8(32'h3a0f4e4f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a578796),
	.w1(32'h3b049291),
	.w2(32'h3aee19bf),
	.w3(32'hb9b7d79b),
	.w4(32'h3a2ceef0),
	.w5(32'hba83fab5),
	.w6(32'h3b97c4a1),
	.w7(32'h3af493c9),
	.w8(32'h3b205d11),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46385e),
	.w1(32'hbc1c4851),
	.w2(32'hba22c6f0),
	.w3(32'hb8d42d0f),
	.w4(32'h3c32dca2),
	.w5(32'h3c45b022),
	.w6(32'hbc661efe),
	.w7(32'h395c6a1d),
	.w8(32'h3c84c421),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4737ea),
	.w1(32'h3c04b6ad),
	.w2(32'h3d06b471),
	.w3(32'h3d0a673e),
	.w4(32'h3b548bae),
	.w5(32'h3c9704aa),
	.w6(32'hbc4efc85),
	.w7(32'h3c54275d),
	.w8(32'h3a7a9d5b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb66261),
	.w1(32'h3ad1ba36),
	.w2(32'hb93c73a9),
	.w3(32'hbae85e28),
	.w4(32'h3a036066),
	.w5(32'hba0bf1d2),
	.w6(32'h3ac4636a),
	.w7(32'hb9bd9e4f),
	.w8(32'hb897c693),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba093047),
	.w1(32'hbb1ad684),
	.w2(32'hbb7dcaf2),
	.w3(32'hba9dfe94),
	.w4(32'hbb255ac7),
	.w5(32'hbbc466f8),
	.w6(32'h3b36a53e),
	.w7(32'hbb421ea8),
	.w8(32'h3b261470),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba819890),
	.w1(32'hbaae1ad2),
	.w2(32'hba7bcb23),
	.w3(32'hb9d9f589),
	.w4(32'h3a3d16af),
	.w5(32'hba966287),
	.w6(32'hbb07f08f),
	.w7(32'hba81bc79),
	.w8(32'h3ae74420),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75e232),
	.w1(32'h3aab4e63),
	.w2(32'h3a43056b),
	.w3(32'h3b1c280b),
	.w4(32'h3ae1c788),
	.w5(32'h3a7caf08),
	.w6(32'h3acd0d77),
	.w7(32'h39af91ed),
	.w8(32'h3ad5c016),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a2478),
	.w1(32'h3a769ec1),
	.w2(32'h39a1fa8a),
	.w3(32'h3a37ffb3),
	.w4(32'h3aa87a87),
	.w5(32'h3a3d2e12),
	.w6(32'h3b0099de),
	.w7(32'h3a42ff1d),
	.w8(32'h3b06aaff),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac4094),
	.w1(32'h3a94e914),
	.w2(32'hba5d2900),
	.w3(32'h3abcd5dc),
	.w4(32'hba9eb5cf),
	.w5(32'hbb05f033),
	.w6(32'hbb144654),
	.w7(32'hbb1274c8),
	.w8(32'hbaabc8cf),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0adfe),
	.w1(32'h3a893263),
	.w2(32'hba9dbd1b),
	.w3(32'hbb0ec874),
	.w4(32'h3add702a),
	.w5(32'hbab3dc04),
	.w6(32'h3a9704b3),
	.w7(32'hba7956a3),
	.w8(32'h39f2f6b8),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1cb02),
	.w1(32'h39d5b01b),
	.w2(32'hbc039545),
	.w3(32'hba56ec98),
	.w4(32'hbb39f4c6),
	.w5(32'hba1983b9),
	.w6(32'h3b42b885),
	.w7(32'hbba67f5a),
	.w8(32'hbbcb7cb2),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb986e08),
	.w1(32'h3a4a0824),
	.w2(32'h3968561e),
	.w3(32'h3b953fd8),
	.w4(32'hbae99940),
	.w5(32'hbb249914),
	.w6(32'h3afcf3f6),
	.w7(32'h3ab5bb40),
	.w8(32'h3a5ddf4a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d21ad0),
	.w1(32'hb8220136),
	.w2(32'h3afc8d53),
	.w3(32'h3922bebb),
	.w4(32'hb93bddcd),
	.w5(32'h3ac07366),
	.w6(32'hba61c677),
	.w7(32'hba21f94e),
	.w8(32'hb88650a7),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cef5c),
	.w1(32'h3bbb4e36),
	.w2(32'h3c5e177e),
	.w3(32'h39ba2dde),
	.w4(32'hbc8e6257),
	.w5(32'h3bddd22d),
	.w6(32'hbb8c4c62),
	.w7(32'h3b006baa),
	.w8(32'hbcc4dd87),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b289b92),
	.w1(32'hba0cc9ac),
	.w2(32'hbaff208f),
	.w3(32'hbbdb5a01),
	.w4(32'h3a717fbb),
	.w5(32'hbac5d77e),
	.w6(32'hbb1fb492),
	.w7(32'hbb81684a),
	.w8(32'h39d7fb8f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f1ae3),
	.w1(32'hbcb13258),
	.w2(32'hbc1f3ad8),
	.w3(32'hbad62385),
	.w4(32'h3afbcd65),
	.w5(32'h3b9e1177),
	.w6(32'hbc843459),
	.w7(32'h3b665414),
	.w8(32'h3c8f829f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953d0cf),
	.w1(32'hb9e53dec),
	.w2(32'h399b4755),
	.w3(32'h3bb9fd0b),
	.w4(32'h3997cc5d),
	.w5(32'h3a931caa),
	.w6(32'hba97c4bc),
	.w7(32'hb97d65a8),
	.w8(32'hba872a75),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c1c57),
	.w1(32'hbb5671be),
	.w2(32'hb96f1da1),
	.w3(32'hb931ee0c),
	.w4(32'hbab71676),
	.w5(32'h3b787a2e),
	.w6(32'hbbdd3a1d),
	.w7(32'hbac5ab9e),
	.w8(32'hbb412327),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adeda42),
	.w1(32'hb9f7230c),
	.w2(32'hba30af04),
	.w3(32'h3b8c4f36),
	.w4(32'h3ad9d4af),
	.w5(32'h3a830ec1),
	.w6(32'hba094c03),
	.w7(32'hb9b51a10),
	.w8(32'hb99a7b90),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2a18a),
	.w1(32'hbc0d231c),
	.w2(32'hbb8e49f3),
	.w3(32'h3a8715bf),
	.w4(32'h3adefce7),
	.w5(32'h3a5d8f97),
	.w6(32'hbc408cfc),
	.w7(32'hbb22828d),
	.w8(32'h3bdb5ff1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72df9f),
	.w1(32'hbba55947),
	.w2(32'hbae4f698),
	.w3(32'hba090ab4),
	.w4(32'hbacbf290),
	.w5(32'h3905c66b),
	.w6(32'hbbd0f742),
	.w7(32'hbae144da),
	.w8(32'h3b86026e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babaef3),
	.w1(32'h3ba00fff),
	.w2(32'h3ae01d71),
	.w3(32'h3c214cb3),
	.w4(32'h3ab697d7),
	.w5(32'h3b1aa7e9),
	.w6(32'h3b140276),
	.w7(32'h3b1b372f),
	.w8(32'h3af39d8c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb933c775),
	.w1(32'hbaac4bf4),
	.w2(32'hbb26d8fa),
	.w3(32'hba1494c3),
	.w4(32'h3a11efe2),
	.w5(32'hba611f5d),
	.w6(32'hbb197ad4),
	.w7(32'hbb41c341),
	.w8(32'hba121e03),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c6aaf),
	.w1(32'h398e284f),
	.w2(32'h3b74e9fa),
	.w3(32'hba0b541d),
	.w4(32'hbb9f3402),
	.w5(32'h39bd682a),
	.w6(32'hbb8f50a5),
	.w7(32'h39a90f0e),
	.w8(32'hbc0be9f0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2327ce),
	.w1(32'hba7bd3eb),
	.w2(32'hba68519d),
	.w3(32'hbba2aa12),
	.w4(32'h3aac4897),
	.w5(32'hb96d7b52),
	.w6(32'hbb52dec0),
	.w7(32'hbb7abdd3),
	.w8(32'h379430f8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82890b2),
	.w1(32'h39976b51),
	.w2(32'h3ab38b26),
	.w3(32'hba9f8d93),
	.w4(32'hbab4b5e0),
	.w5(32'h3a56b67d),
	.w6(32'hbb5938ad),
	.w7(32'hbadba0a0),
	.w8(32'hbaab6590),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba819433),
	.w1(32'hbb076e7b),
	.w2(32'h3ad06387),
	.w3(32'hbb15348b),
	.w4(32'hb9c8eccb),
	.w5(32'h3ab887ad),
	.w6(32'hba8e5602),
	.w7(32'h3b257f0d),
	.w8(32'h3a0cb203),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9b348),
	.w1(32'hbb756450),
	.w2(32'hbb2eda0d),
	.w3(32'h3acae568),
	.w4(32'hbb580d77),
	.w5(32'hbb27d3d9),
	.w6(32'hbb9e915a),
	.w7(32'hbaaf01de),
	.w8(32'hbb27da98),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba332989),
	.w1(32'hbca75bca),
	.w2(32'hbc4aadc3),
	.w3(32'hb90838ef),
	.w4(32'hba277ed0),
	.w5(32'hba748449),
	.w6(32'hbc94a53f),
	.w7(32'hba951b89),
	.w8(32'h3c31ff3c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d6019),
	.w1(32'h3b108a40),
	.w2(32'h3b5bfe6a),
	.w3(32'h3a03717c),
	.w4(32'hba092a78),
	.w5(32'hba37e734),
	.w6(32'hb99c716a),
	.w7(32'hbb771bcb),
	.w8(32'hbb625a52),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82003b),
	.w1(32'h3b0e384a),
	.w2(32'h391a77a1),
	.w3(32'hbae70d10),
	.w4(32'h3a1e9801),
	.w5(32'h3ad29ca9),
	.w6(32'h3aa38a42),
	.w7(32'hb9cc292b),
	.w8(32'hba8d68d3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c106f),
	.w1(32'h3c17f2a4),
	.w2(32'h3c36be6d),
	.w3(32'hb92cb0be),
	.w4(32'hbbb06542),
	.w5(32'hbca7fbee),
	.w6(32'hbafbd2b2),
	.w7(32'hbc49d59e),
	.w8(32'hbbbf45c2),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb7fcf5),
	.w1(32'hba9fd656),
	.w2(32'h3b257fc5),
	.w3(32'hbc3ed715),
	.w4(32'hbb01cd72),
	.w5(32'hbbbe1428),
	.w6(32'h3b0b2396),
	.w7(32'h3bb06ace),
	.w8(32'h3abedc89),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb016366),
	.w1(32'hbac5425b),
	.w2(32'hba55fdb6),
	.w3(32'hbb835e84),
	.w4(32'hba84bdc7),
	.w5(32'h38601398),
	.w6(32'hbb068a82),
	.w7(32'hb928113f),
	.w8(32'h388ed22c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fbdad1),
	.w1(32'hba9cf0a0),
	.w2(32'hbac971e3),
	.w3(32'hba60f57c),
	.w4(32'hbab89b5f),
	.w5(32'h39a2a4ca),
	.w6(32'hbb8f07a9),
	.w7(32'hba5f4fad),
	.w8(32'h3aae2348),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00c17f),
	.w1(32'hba0fa1c0),
	.w2(32'h3b36e8e2),
	.w3(32'h3b2cedf7),
	.w4(32'hbb3b6c87),
	.w5(32'hbb6ec0fd),
	.w6(32'h3a215eb9),
	.w7(32'h3ac78773),
	.w8(32'hb9eca03a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7da976),
	.w1(32'hb9b9f002),
	.w2(32'hbb6576aa),
	.w3(32'hbbb4a105),
	.w4(32'hba3648ef),
	.w5(32'hbad9b1c9),
	.w6(32'hba944f43),
	.w7(32'hbbcf2db5),
	.w8(32'hbb48d81f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0a905),
	.w1(32'h3989d90d),
	.w2(32'h39466919),
	.w3(32'h3992ab98),
	.w4(32'hbb2f9b23),
	.w5(32'hbb451ad6),
	.w6(32'h3b1eecce),
	.w7(32'h3b191521),
	.w8(32'h3b067cae),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d5ed3),
	.w1(32'h3a235a77),
	.w2(32'h3ad9c0b5),
	.w3(32'h38921e7e),
	.w4(32'h3a2690b4),
	.w5(32'h3ab12240),
	.w6(32'h3a9c365a),
	.w7(32'h3aa88328),
	.w8(32'h3b332702),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac005e9),
	.w1(32'h3a047d40),
	.w2(32'h3793857a),
	.w3(32'hb81a54d6),
	.w4(32'hbaa2170c),
	.w5(32'hbaf1ff94),
	.w6(32'h3ab6043b),
	.w7(32'h3a8d28a3),
	.w8(32'h3a1fa6af),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d344b),
	.w1(32'hbae20757),
	.w2(32'h39f69e72),
	.w3(32'hb8dad2f1),
	.w4(32'hbb2bacb9),
	.w5(32'h3ac4c003),
	.w6(32'h3a36c108),
	.w7(32'h3aee37df),
	.w8(32'h3a9c1342),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d7180),
	.w1(32'h3a5fb818),
	.w2(32'h3ac09652),
	.w3(32'hbaa382b0),
	.w4(32'hb9bf7408),
	.w5(32'hba78c784),
	.w6(32'h3a26933a),
	.w7(32'h399056b4),
	.w8(32'hbb0c85df),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9d1bf),
	.w1(32'hba89ab6d),
	.w2(32'h398467e5),
	.w3(32'hbb31a72a),
	.w4(32'hb8b712a8),
	.w5(32'h3a6a7e75),
	.w6(32'hbb453ae9),
	.w7(32'hbb005dcc),
	.w8(32'hba44dd21),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05e15e),
	.w1(32'h3a38e9b0),
	.w2(32'h39987a76),
	.w3(32'hb9e7c928),
	.w4(32'hba874cb8),
	.w5(32'hbadacc1e),
	.w6(32'h3ac36ccc),
	.w7(32'h3a9bbd9e),
	.w8(32'h3a641b64),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9030504),
	.w1(32'h3b17b8c2),
	.w2(32'h39cd935b),
	.w3(32'h399291ab),
	.w4(32'h3b61f214),
	.w5(32'h3a8d937c),
	.w6(32'h3bf01798),
	.w7(32'h3b51c024),
	.w8(32'h3a19b4d0),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e183b),
	.w1(32'h3b502dba),
	.w2(32'h39a8422a),
	.w3(32'hba8fa9e9),
	.w4(32'h3b22a82f),
	.w5(32'hb8d60ed1),
	.w6(32'h3b884102),
	.w7(32'h3aa444a1),
	.w8(32'h3b1c09e5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a625817),
	.w1(32'h3a8dc6da),
	.w2(32'hba8e5a07),
	.w3(32'h398615a6),
	.w4(32'h39a69a59),
	.w5(32'h3aa82494),
	.w6(32'h3a594285),
	.w7(32'h395f83ad),
	.w8(32'h3aa6a614),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d503e),
	.w1(32'h3b274285),
	.w2(32'h38ed58b5),
	.w3(32'hba4ff03a),
	.w4(32'h3ad96846),
	.w5(32'hb98c12b2),
	.w6(32'h3b4953d0),
	.w7(32'h3a2e4b41),
	.w8(32'h3b0d426e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4a537),
	.w1(32'h3b1c862c),
	.w2(32'h3a167dc4),
	.w3(32'hba349376),
	.w4(32'hb8c5e84e),
	.w5(32'hbb3e9b05),
	.w6(32'h3a44ccb2),
	.w7(32'hba629fb3),
	.w8(32'h3aaac149),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27950a),
	.w1(32'hbac7f6b3),
	.w2(32'h3a8ac2c9),
	.w3(32'hbae36d56),
	.w4(32'hbb80e877),
	.w5(32'hbab51790),
	.w6(32'hbb4fe41a),
	.w7(32'hba1039a4),
	.w8(32'hbb8302e4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba161de2),
	.w1(32'h3a64a301),
	.w2(32'h398fe5e0),
	.w3(32'hbb77e935),
	.w4(32'hbaec81c4),
	.w5(32'hbb2a321b),
	.w6(32'h3b07e46e),
	.w7(32'h3ad8fd02),
	.w8(32'h3a8b7684),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b86909),
	.w1(32'hb908becc),
	.w2(32'h3a30caea),
	.w3(32'h39835c8e),
	.w4(32'h39eb7bad),
	.w5(32'h39d937b5),
	.w6(32'h38d9f0aa),
	.w7(32'h3ab11065),
	.w8(32'h3a9ff028),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a664f55),
	.w1(32'h3a1e0d34),
	.w2(32'h3a165379),
	.w3(32'h3abfdd2c),
	.w4(32'hb9896bf1),
	.w5(32'hb904315d),
	.w6(32'h3a606d52),
	.w7(32'h3af7496f),
	.w8(32'h3ab0858b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9b500),
	.w1(32'h3ac1b4c5),
	.w2(32'hbaea87fe),
	.w3(32'h3ac43065),
	.w4(32'h3af7ff99),
	.w5(32'hba99b8a7),
	.w6(32'h3b9baade),
	.w7(32'h3ad5fb02),
	.w8(32'hbb3882bb),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb853795),
	.w1(32'hba63548a),
	.w2(32'h3b5b4434),
	.w3(32'hbb22dac9),
	.w4(32'hb93b7330),
	.w5(32'hbb084e27),
	.w6(32'hbac46ab5),
	.w7(32'h3933db74),
	.w8(32'hb9bd9249),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac89f1d),
	.w1(32'h3b24f57a),
	.w2(32'h3b33ece4),
	.w3(32'hbb14e03f),
	.w4(32'h3adad677),
	.w5(32'h3aae7dc4),
	.w6(32'hb94727ac),
	.w7(32'h39a58944),
	.w8(32'hba6744e5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88efab),
	.w1(32'h3addf6a1),
	.w2(32'h3a89404c),
	.w3(32'hbaf48bbe),
	.w4(32'h399ee802),
	.w5(32'hba4776f2),
	.w6(32'h3a646a2e),
	.w7(32'h39ae742b),
	.w8(32'h3a96739d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad41f0),
	.w1(32'h3aab6859),
	.w2(32'hb9cdcca8),
	.w3(32'hbaa43fd2),
	.w4(32'h3ac377cd),
	.w5(32'hb8e1df5d),
	.w6(32'h3ac29719),
	.w7(32'hb9b54a78),
	.w8(32'h3aa54706),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13d55c),
	.w1(32'h3b9c8096),
	.w2(32'h3b52c905),
	.w3(32'h3a1f9658),
	.w4(32'h3b9a72fc),
	.w5(32'h3aa2ab64),
	.w6(32'h3b54f614),
	.w7(32'h3aa1c903),
	.w8(32'h3b19290f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36ec3f),
	.w1(32'hbb11dd5a),
	.w2(32'hbb1f965a),
	.w3(32'hb9e0ac2f),
	.w4(32'hbb649630),
	.w5(32'hbb40019c),
	.w6(32'hbb4b83c8),
	.w7(32'h3a313452),
	.w8(32'h3a730b82),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb338c15),
	.w1(32'hba302522),
	.w2(32'hbb203e84),
	.w3(32'hbb1f8593),
	.w4(32'h3a327e68),
	.w5(32'hba7026cd),
	.w6(32'hbb00930f),
	.w7(32'hbb0f4155),
	.w8(32'hba025ccb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c2a37),
	.w1(32'hb9ea8b69),
	.w2(32'hb92f50b0),
	.w3(32'hbae27f51),
	.w4(32'hba254cbe),
	.w5(32'hba0d5c88),
	.w6(32'hb98e9b33),
	.w7(32'h3983ca46),
	.w8(32'h39cbd36d),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a422a),
	.w1(32'hb9ad67ad),
	.w2(32'h38b41c82),
	.w3(32'h372ac4ac),
	.w4(32'hb90be3a8),
	.w5(32'hba17f14e),
	.w6(32'hb9807bbb),
	.w7(32'hb75a2e1a),
	.w8(32'h366aadfa),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule