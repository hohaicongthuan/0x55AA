module layer_10_featuremap_404(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b610e37),
	.w1(32'h3c3c3111),
	.w2(32'h3c450f07),
	.w3(32'h3b480d7b),
	.w4(32'h3c8fb401),
	.w5(32'h3c694448),
	.w6(32'hbbfb1e24),
	.w7(32'h3bb5f1bf),
	.w8(32'h398cab7d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e0607),
	.w1(32'h39d44bac),
	.w2(32'hba083097),
	.w3(32'hbc764f70),
	.w4(32'hbb371c5a),
	.w5(32'hbb9a8390),
	.w6(32'hbc0495d4),
	.w7(32'hbb380504),
	.w8(32'hbba8547d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c8b3e),
	.w1(32'hb9cfa4f9),
	.w2(32'hbab2e182),
	.w3(32'hbb34f7e6),
	.w4(32'h39cd445c),
	.w5(32'hbb9ab699),
	.w6(32'hb9e514ed),
	.w7(32'h3a779002),
	.w8(32'h39793758),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9b0ff),
	.w1(32'hbabdc262),
	.w2(32'hbbcea9ab),
	.w3(32'hbb204736),
	.w4(32'h3aeb8418),
	.w5(32'hb99d89dd),
	.w6(32'h3ae1be3c),
	.w7(32'hb9d51df4),
	.w8(32'hbc384502),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61d85b),
	.w1(32'h3be52cd8),
	.w2(32'h3b852283),
	.w3(32'hbbc478b2),
	.w4(32'h3bf7cd27),
	.w5(32'h3ba58223),
	.w6(32'hb99a80cb),
	.w7(32'h3bb6449f),
	.w8(32'h3ab7282e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad39c86),
	.w1(32'hbb758b75),
	.w2(32'hbbc29679),
	.w3(32'h3b56e487),
	.w4(32'h3a99560e),
	.w5(32'hbc580f46),
	.w6(32'hbade6cf5),
	.w7(32'h3b6ff41d),
	.w8(32'h3c468108),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bd9fd),
	.w1(32'hbbd8f7f0),
	.w2(32'hbb7d5c66),
	.w3(32'hba36dbc7),
	.w4(32'hbb947f86),
	.w5(32'h3ba6ccc7),
	.w6(32'h3b81f674),
	.w7(32'h3b11c318),
	.w8(32'h3c14f4cb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac67aa2),
	.w1(32'hbc00b9ef),
	.w2(32'h3b7ee9c7),
	.w3(32'hbbba654a),
	.w4(32'hbb9f2535),
	.w5(32'h3b49115b),
	.w6(32'hbb03e69c),
	.w7(32'hbb89d23a),
	.w8(32'h3bebdd19),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0891fe),
	.w1(32'hbae7daed),
	.w2(32'h3b24faf0),
	.w3(32'hbb570e75),
	.w4(32'hbb3fbdaa),
	.w5(32'hbb80a194),
	.w6(32'hbb41c3d2),
	.w7(32'hbb0e4a6f),
	.w8(32'hbbabb67a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7eaa4e),
	.w1(32'h3b98c9b7),
	.w2(32'h39c77a6a),
	.w3(32'hbb286115),
	.w4(32'h3b0c1ea3),
	.w5(32'hba71e0e8),
	.w6(32'hbb245e79),
	.w7(32'h39c5d1a1),
	.w8(32'h3b31bbca),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb004d40),
	.w1(32'h3a8ade12),
	.w2(32'hbb62ed33),
	.w3(32'h3b8e38ed),
	.w4(32'hbbb60c9b),
	.w5(32'hbbd98650),
	.w6(32'h3b0dae32),
	.w7(32'hbb0dc2e4),
	.w8(32'hbbcd112b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0991b8),
	.w1(32'h3b06cb35),
	.w2(32'hbc0e7ee5),
	.w3(32'hbb206445),
	.w4(32'h39b7729c),
	.w5(32'hbc32cc1a),
	.w6(32'hbb36e2d4),
	.w7(32'h3a41b3a5),
	.w8(32'h3b99a26c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9786d1),
	.w1(32'hbb98fde6),
	.w2(32'hbbebb73f),
	.w3(32'h3c431f6c),
	.w4(32'hbbaaf7b0),
	.w5(32'hbb8ef042),
	.w6(32'h3bcc13bf),
	.w7(32'hbae06948),
	.w8(32'h3b62220a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bf2ce),
	.w1(32'hbab66147),
	.w2(32'h3b6b4a8a),
	.w3(32'h3c694982),
	.w4(32'hbacfcb90),
	.w5(32'hbbe09eb8),
	.w6(32'h3b95cdc8),
	.w7(32'hbbe09b1f),
	.w8(32'hbc1f375a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add78d6),
	.w1(32'hba99731c),
	.w2(32'hbb7f14e8),
	.w3(32'h3b47b150),
	.w4(32'hbb21f543),
	.w5(32'hbbcf0c71),
	.w6(32'hbb16f829),
	.w7(32'h3a3edc41),
	.w8(32'hba3d527f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50a9a4),
	.w1(32'hbb8dda1f),
	.w2(32'hbbc71b09),
	.w3(32'hb8ae53cd),
	.w4(32'hbbc6d58e),
	.w5(32'hba192a7e),
	.w6(32'hbb0ef4f9),
	.w7(32'hba4d0be4),
	.w8(32'h3aea7210),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb335444),
	.w1(32'hbb0d9b61),
	.w2(32'hbae3661c),
	.w3(32'h3baae516),
	.w4(32'hbaf68731),
	.w5(32'hbb9a4dd8),
	.w6(32'h3b1e633f),
	.w7(32'hba90c86c),
	.w8(32'hbbd77432),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb512380),
	.w1(32'h3c2fb5a2),
	.w2(32'h3c474536),
	.w3(32'hba576fbf),
	.w4(32'h3c5b9d67),
	.w5(32'h3b26551d),
	.w6(32'h39b7faae),
	.w7(32'h3bb435b2),
	.w8(32'hbb7bd96a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29a7f8),
	.w1(32'h3a95f9c6),
	.w2(32'hbc150f7c),
	.w3(32'hbcc21641),
	.w4(32'hbb1b1aa0),
	.w5(32'hbc18a101),
	.w6(32'hbc66996d),
	.w7(32'h3a7e248c),
	.w8(32'h3b30eb0e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5d783),
	.w1(32'h3adffeb2),
	.w2(32'hba6853e5),
	.w3(32'h3b32f24a),
	.w4(32'hba6490b2),
	.w5(32'hbbabf1e0),
	.w6(32'hbb88ac4d),
	.w7(32'h3ac72fbe),
	.w8(32'hbc3eced8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d647b),
	.w1(32'hbbe31b69),
	.w2(32'hbc2af710),
	.w3(32'hbb90a895),
	.w4(32'hbc09bb9a),
	.w5(32'hbc86dbca),
	.w6(32'hbb78e0d5),
	.w7(32'hbc3011b6),
	.w8(32'h3adf31bb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fd14d),
	.w1(32'hbbdba13b),
	.w2(32'hbb15f973),
	.w3(32'h3c700e18),
	.w4(32'hbbd35afc),
	.w5(32'h3b08100a),
	.w6(32'h3c11ef62),
	.w7(32'hbbe19674),
	.w8(32'h3b09b306),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2e203),
	.w1(32'hba459677),
	.w2(32'hbb6cfd70),
	.w3(32'hbc20a1ee),
	.w4(32'hbbb2cb9f),
	.w5(32'hbc12d6e5),
	.w6(32'hbc4fb8c2),
	.w7(32'hbbeee0be),
	.w8(32'h3a5eb5b8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f9605),
	.w1(32'h3aba0b97),
	.w2(32'hbb6bf207),
	.w3(32'hbb5104dd),
	.w4(32'h3c4f9690),
	.w5(32'h3b764393),
	.w6(32'h3b775384),
	.w7(32'hba229f1c),
	.w8(32'hbc22d1df),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb632f7b),
	.w1(32'hbc0ea594),
	.w2(32'hbba5fa7b),
	.w3(32'h3b65ae01),
	.w4(32'hbc4c5eaf),
	.w5(32'hbaaf3631),
	.w6(32'hbb99d81c),
	.w7(32'hbc02d0c5),
	.w8(32'hbbd5bece),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89aee1),
	.w1(32'hbbafba61),
	.w2(32'h3bb37672),
	.w3(32'hb9886c8b),
	.w4(32'h3b33e508),
	.w5(32'h3ba40a9f),
	.w6(32'hbb9b0ba1),
	.w7(32'hb9441405),
	.w8(32'h3ae66759),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe007a7),
	.w1(32'hba891f36),
	.w2(32'hbbb208f0),
	.w3(32'hbb5e98fe),
	.w4(32'hbbac079f),
	.w5(32'hbbe90938),
	.w6(32'hbb5cbc75),
	.w7(32'hbc3400aa),
	.w8(32'hbbf071dd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ee7d3),
	.w1(32'h3a606c94),
	.w2(32'h3b52bde4),
	.w3(32'hba4abddd),
	.w4(32'hbb3ebb5b),
	.w5(32'h3bbe4ba1),
	.w6(32'hbc288151),
	.w7(32'hba66893a),
	.w8(32'hbbac2e38),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f59cb4),
	.w1(32'hbbdb766c),
	.w2(32'h3b151e28),
	.w3(32'hbb329783),
	.w4(32'hbb4019db),
	.w5(32'hbb87034f),
	.w6(32'h391aaf6a),
	.w7(32'hbb4f4d61),
	.w8(32'h3b17a39a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c1b0a),
	.w1(32'hbc2c7d27),
	.w2(32'hbb91dca4),
	.w3(32'hbb9ffcb8),
	.w4(32'hbc8623e9),
	.w5(32'hbbbba4cc),
	.w6(32'hbb345623),
	.w7(32'hb9b15625),
	.w8(32'h3c8ce45a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c195ae2),
	.w1(32'h3acb3f6e),
	.w2(32'h3c069070),
	.w3(32'h3c6427a3),
	.w4(32'h3b73182b),
	.w5(32'hbc042f0d),
	.w6(32'h3c8bf9e1),
	.w7(32'h3b4b2797),
	.w8(32'h3b38c910),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee4667),
	.w1(32'h3a330525),
	.w2(32'hbb1ecfa3),
	.w3(32'hbc14e665),
	.w4(32'hbbc877b9),
	.w5(32'hbbaf014f),
	.w6(32'h3b0b25da),
	.w7(32'hbbf4233e),
	.w8(32'hbb0819f7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9d353),
	.w1(32'hbb462791),
	.w2(32'hbb8118ff),
	.w3(32'hbbf81c2a),
	.w4(32'hbb6b4d3f),
	.w5(32'h3b307729),
	.w6(32'hbb232e2a),
	.w7(32'hbb28a9f3),
	.w8(32'h3a2eecf5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba658b98),
	.w1(32'h3af77bc0),
	.w2(32'h3bd3bfbf),
	.w3(32'h3b2831a9),
	.w4(32'h3b3c27c5),
	.w5(32'h3c49f5b0),
	.w6(32'hba47927a),
	.w7(32'hba10944f),
	.w8(32'hbab98fe5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17d558),
	.w1(32'hbb080a13),
	.w2(32'h3bc3d422),
	.w3(32'hbbca0020),
	.w4(32'hbb7df6e2),
	.w5(32'hbad1c805),
	.w6(32'hba5d173b),
	.w7(32'hb9f181a4),
	.w8(32'h3ba3a199),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e44b48),
	.w1(32'h39971534),
	.w2(32'hba39bfa8),
	.w3(32'hbb66c649),
	.w4(32'h3bca390f),
	.w5(32'hbb6d8f42),
	.w6(32'hb7ad6b2c),
	.w7(32'hbb666fef),
	.w8(32'hbc48ff1d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb410b6c),
	.w1(32'h3a5f1b07),
	.w2(32'hbb4f298e),
	.w3(32'hbb878505),
	.w4(32'hbb46463a),
	.w5(32'hbba9ea50),
	.w6(32'hbbcc0481),
	.w7(32'h3c01e7e8),
	.w8(32'hbb99e709),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8de7d91),
	.w1(32'hbab211bf),
	.w2(32'hbb4e34fe),
	.w3(32'hbb897ac7),
	.w4(32'h3b8bf00b),
	.w5(32'hbbf82e50),
	.w6(32'hbc2dce7f),
	.w7(32'hba8224c3),
	.w8(32'hbada76e4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98acad),
	.w1(32'hbabc6000),
	.w2(32'h3b1c4dea),
	.w3(32'h39e0ded6),
	.w4(32'h3b6fc160),
	.w5(32'h3c4c7679),
	.w6(32'h3b5157b0),
	.w7(32'hbaea5163),
	.w8(32'hbc2fcd61),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba982540),
	.w1(32'h3b3472db),
	.w2(32'h3a9ace71),
	.w3(32'hbbb46951),
	.w4(32'h3bededd9),
	.w5(32'h3bf99922),
	.w6(32'hbbb8a599),
	.w7(32'h3b1e0db6),
	.w8(32'hbbc1fdd7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba908959),
	.w1(32'hbbc3838b),
	.w2(32'hbb0d4a26),
	.w3(32'hbb47db8c),
	.w4(32'h3bc47c1a),
	.w5(32'hbb92ee42),
	.w6(32'hbae8ab7f),
	.w7(32'hbb1c9170),
	.w8(32'hbc1c5686),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf3897),
	.w1(32'hbb9133dc),
	.w2(32'hbc6f86ef),
	.w3(32'hbae89e52),
	.w4(32'hbbbd1819),
	.w5(32'hbbe31adb),
	.w6(32'hbb48909d),
	.w7(32'hbb0a4cab),
	.w8(32'hbb89cee2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a0c50),
	.w1(32'h3bc6affb),
	.w2(32'hbaba2c33),
	.w3(32'h39aab009),
	.w4(32'h3b261a66),
	.w5(32'h3b671040),
	.w6(32'hbc01c8cc),
	.w7(32'h3af58af1),
	.w8(32'hbbb90c2d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddea7b),
	.w1(32'hbc4c45ee),
	.w2(32'hbb0a65d9),
	.w3(32'hbb1a2dfc),
	.w4(32'hbb697d8b),
	.w5(32'h3c44e628),
	.w6(32'hbbda1b7f),
	.w7(32'hbc07e386),
	.w8(32'hbc485e0d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba579b9),
	.w1(32'h3b1f7c75),
	.w2(32'h3a9c9175),
	.w3(32'hbc82d2d2),
	.w4(32'h3b221cd6),
	.w5(32'hba7b0270),
	.w6(32'hbc67a385),
	.w7(32'h3b74eac0),
	.w8(32'h3b062c8e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce04bd),
	.w1(32'hbaa706ba),
	.w2(32'hbb9102cf),
	.w3(32'hbbce2338),
	.w4(32'hbc0ad18a),
	.w5(32'hba078298),
	.w6(32'hbb659128),
	.w7(32'hbb80a92f),
	.w8(32'hbae7d426),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab2a8e),
	.w1(32'h3b11dcb9),
	.w2(32'hbb5ebaa1),
	.w3(32'h3c2a00e0),
	.w4(32'hbb6ec48d),
	.w5(32'hbb9b9e90),
	.w6(32'h3bbe09e9),
	.w7(32'hbb61a8b8),
	.w8(32'h3ade152b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b033f8b),
	.w1(32'h3a3b1361),
	.w2(32'h3bad9e8f),
	.w3(32'h3b96c6f7),
	.w4(32'h3a94ab60),
	.w5(32'h3c435ad2),
	.w6(32'h3b8f4f87),
	.w7(32'h3a243c1d),
	.w8(32'h3bf68f6b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a914a27),
	.w1(32'hbbea0a12),
	.w2(32'hbb5eaf55),
	.w3(32'hbb2c7667),
	.w4(32'hbbcca4b4),
	.w5(32'hbb7140c7),
	.w6(32'hbb92cce7),
	.w7(32'hbc196120),
	.w8(32'hbb8fe9e3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb515d45),
	.w1(32'hbbea9eb8),
	.w2(32'hbb264ad8),
	.w3(32'h3b61246e),
	.w4(32'hbbdc095f),
	.w5(32'hbb08000e),
	.w6(32'hba40eafd),
	.w7(32'hbc2effbc),
	.w8(32'hbbb231fa),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf4df1),
	.w1(32'h3c04efb2),
	.w2(32'h3b922d71),
	.w3(32'h3b039ecd),
	.w4(32'h3ca4e332),
	.w5(32'hbc5ad796),
	.w6(32'hbb752d01),
	.w7(32'hbb592223),
	.w8(32'hbbe2f535),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7f461),
	.w1(32'h39e2b973),
	.w2(32'hbc19e61d),
	.w3(32'h3c8f0324),
	.w4(32'hbbd7bae3),
	.w5(32'hbc5e0586),
	.w6(32'h3c0b2063),
	.w7(32'hba36b288),
	.w8(32'hbc401167),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb710d48),
	.w1(32'hbba97e58),
	.w2(32'h3b22ca85),
	.w3(32'hba372280),
	.w4(32'hbaf7dbb6),
	.w5(32'hbb1b19a4),
	.w6(32'hbb1f38e6),
	.w7(32'hbb13c39e),
	.w8(32'h3b3f528f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74a800),
	.w1(32'h3955d266),
	.w2(32'h3b56c829),
	.w3(32'hbc1a68ed),
	.w4(32'h3a8001bf),
	.w5(32'hbba864fa),
	.w6(32'hbb94aab5),
	.w7(32'hbacfba2c),
	.w8(32'h39d07105),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79ff18),
	.w1(32'hbaaeabff),
	.w2(32'hbb488654),
	.w3(32'hbad6d704),
	.w4(32'hba7d83d0),
	.w5(32'hbb58d667),
	.w6(32'hbad92a79),
	.w7(32'hbb50d9d4),
	.w8(32'hbb02c507),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9997d7),
	.w1(32'h3b55eb4c),
	.w2(32'hbb0ea264),
	.w3(32'hbb17b4e6),
	.w4(32'h3beb5144),
	.w5(32'hbb7d4d5c),
	.w6(32'hba85ec28),
	.w7(32'hbb51895b),
	.w8(32'hbbd3d1a1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47064e),
	.w1(32'h3c339ca1),
	.w2(32'hbab397b3),
	.w3(32'hbbb60961),
	.w4(32'h3bed512c),
	.w5(32'hbc53006c),
	.w6(32'hbb86da5a),
	.w7(32'h3badacc9),
	.w8(32'h3bfb83ff),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2239eb),
	.w1(32'hbb845532),
	.w2(32'hbb5c08e9),
	.w3(32'h3cc4eaad),
	.w4(32'hbb6b41d2),
	.w5(32'h3b10db96),
	.w6(32'h3c248a89),
	.w7(32'hbb76b977),
	.w8(32'hbbcda76d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4ab27),
	.w1(32'h39387090),
	.w2(32'hbbebdcce),
	.w3(32'hbb737bdb),
	.w4(32'h39739628),
	.w5(32'hbbb294aa),
	.w6(32'hbbb5893c),
	.w7(32'hb98c7f13),
	.w8(32'hbb8f729f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8bd98),
	.w1(32'hbba1f487),
	.w2(32'hbbc72cda),
	.w3(32'h39a75eb3),
	.w4(32'hb897e7b0),
	.w5(32'h3bbf264b),
	.w6(32'h3af7484f),
	.w7(32'h3b908168),
	.w8(32'h3bfa5d0c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5271f),
	.w1(32'h3ad6e5be),
	.w2(32'h3a3e3288),
	.w3(32'hbb9ff41a),
	.w4(32'hbc144ba5),
	.w5(32'hb9658547),
	.w6(32'h385950b5),
	.w7(32'hbc316370),
	.w8(32'h3ba73dce),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f43f5),
	.w1(32'h3b1605e2),
	.w2(32'hbb6880be),
	.w3(32'h3c14446b),
	.w4(32'hbb1fa1bf),
	.w5(32'hbb7ce652),
	.w6(32'hba466af1),
	.w7(32'h39d4efb3),
	.w8(32'hb98a00f7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad8c47),
	.w1(32'h3bc1f2f2),
	.w2(32'h3aa1002a),
	.w3(32'hbb2586f1),
	.w4(32'h3c458d33),
	.w5(32'h3b6dee0b),
	.w6(32'hb9959e7e),
	.w7(32'hbb149ebc),
	.w8(32'hbc704d44),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc173e83),
	.w1(32'h3bf849f9),
	.w2(32'hbc05ea44),
	.w3(32'hbc62bb6c),
	.w4(32'h3b051959),
	.w5(32'hbc44542e),
	.w6(32'hbc185f01),
	.w7(32'h3bc65804),
	.w8(32'h3c31a1d9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b876cd2),
	.w1(32'h3babe4e5),
	.w2(32'h3b94b729),
	.w3(32'h3c8a51e6),
	.w4(32'h3c00dd68),
	.w5(32'h3a820659),
	.w6(32'h3c11455a),
	.w7(32'h3aaf35fc),
	.w8(32'h3a151562),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d3825),
	.w1(32'h3afaaa0d),
	.w2(32'h3b0fdd48),
	.w3(32'h3baddc24),
	.w4(32'h3ad182c2),
	.w5(32'h3c2c38a1),
	.w6(32'h3ba71cbf),
	.w7(32'h3b734707),
	.w8(32'hbc0c9db6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b401249),
	.w1(32'h3c2b2178),
	.w2(32'hbb47aa1f),
	.w3(32'hbac1a0e9),
	.w4(32'h3b8cacac),
	.w5(32'hbc553198),
	.w6(32'hbc04d5eb),
	.w7(32'h3b81ce16),
	.w8(32'hb60a6d7f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ec9f7),
	.w1(32'hbbbdc0fd),
	.w2(32'h3ae7e35a),
	.w3(32'h3bd145f1),
	.w4(32'hbc041d7f),
	.w5(32'h3ba9def6),
	.w6(32'h3af1cb63),
	.w7(32'hbbbb3455),
	.w8(32'h3c20c289),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09344d),
	.w1(32'hbc7a3d6d),
	.w2(32'h3a9f6d63),
	.w3(32'h3bd5fff7),
	.w4(32'hbc38991f),
	.w5(32'h3bd06752),
	.w6(32'h3b9340df),
	.w7(32'hbc274d15),
	.w8(32'hbbac9525),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb376b1d),
	.w1(32'hb8088494),
	.w2(32'hb84a322b),
	.w3(32'hbbaa91f5),
	.w4(32'hb80ac402),
	.w5(32'hb78c6ee0),
	.w6(32'hbb901490),
	.w7(32'hb80a82be),
	.w8(32'hb6f6423a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378a9452),
	.w1(32'h370fdddb),
	.w2(32'h371e2f29),
	.w3(32'h3746c3ed),
	.w4(32'h36aad443),
	.w5(32'hb5acd0e9),
	.w6(32'h369ca93d),
	.w7(32'hb5e53164),
	.w8(32'h363bb5ed),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a63ec1),
	.w1(32'h370063e9),
	.w2(32'hb713c2cc),
	.w3(32'h36ae807f),
	.w4(32'h372b4829),
	.w5(32'hb6860a65),
	.w6(32'h37296c6a),
	.w7(32'hb5f6f53d),
	.w8(32'h3538a0ff),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374bc80f),
	.w1(32'hb65f0f9d),
	.w2(32'h3714e66c),
	.w3(32'hb66082b1),
	.w4(32'hb3ae79d4),
	.w5(32'h373ef1d5),
	.w6(32'hb69320af),
	.w7(32'h36739ad4),
	.w8(32'h36dd3720),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3793ef8a),
	.w1(32'h36df1d75),
	.w2(32'h3784e314),
	.w3(32'h37a2ad93),
	.w4(32'h3703e163),
	.w5(32'h372ed852),
	.w6(32'h37985756),
	.w7(32'h36503fb4),
	.w8(32'h3659261d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb682b3c4),
	.w1(32'h36495eaa),
	.w2(32'hb6a898d2),
	.w3(32'h35ef362b),
	.w4(32'h35fc91f3),
	.w5(32'h36605199),
	.w6(32'h36368d9d),
	.w7(32'h37a71ce1),
	.w8(32'h37a7e4cb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35cb2bd0),
	.w1(32'h37a79de9),
	.w2(32'h36f67d08),
	.w3(32'hb46383ef),
	.w4(32'h3812e9b8),
	.w5(32'h37f71f29),
	.w6(32'h36686f9e),
	.w7(32'h3611b9ad),
	.w8(32'hb78c0149),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7eeaa66),
	.w1(32'h385970dd),
	.w2(32'h3809e25c),
	.w3(32'hb7b1debb),
	.w4(32'h37d0d04e),
	.w5(32'h37e33195),
	.w6(32'hb875e420),
	.w7(32'hb736bb8b),
	.w8(32'h3652fc07),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7914d42),
	.w1(32'hb7be25c9),
	.w2(32'hb61bc0f2),
	.w3(32'h345c5b98),
	.w4(32'hb722c9bc),
	.w5(32'h36bc0f25),
	.w6(32'hb72ca29d),
	.w7(32'hb5169fa6),
	.w8(32'h37c13e90),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372916c0),
	.w1(32'h37e80c74),
	.w2(32'h3841106c),
	.w3(32'h368032db),
	.w4(32'h37ef1819),
	.w5(32'h37cc74ff),
	.w6(32'h37899122),
	.w7(32'h379ee5d4),
	.w8(32'h38184549),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3747a7ed),
	.w1(32'h384607b7),
	.w2(32'h38784588),
	.w3(32'h37a03dde),
	.w4(32'h37a44348),
	.w5(32'h38047d76),
	.w6(32'hb5be6a78),
	.w7(32'h378b25f3),
	.w8(32'h37ce2fdb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c9b28d),
	.w1(32'hb7477766),
	.w2(32'hb6abe682),
	.w3(32'h3758ccd0),
	.w4(32'hb607b3ec),
	.w5(32'hb71d863b),
	.w6(32'h3746391e),
	.w7(32'hb586606a),
	.w8(32'hb6484734),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a7059b),
	.w1(32'h37e9c87b),
	.w2(32'h3823c575),
	.w3(32'hb4b83af3),
	.w4(32'h37d0ac17),
	.w5(32'h369fc0f6),
	.w6(32'hb7493abd),
	.w7(32'hb6722bee),
	.w8(32'hb79b8d1c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368bc04f),
	.w1(32'h35bcf72d),
	.w2(32'h3709f6da),
	.w3(32'h359ccfd2),
	.w4(32'h37086e6f),
	.w5(32'h36802dab),
	.w6(32'h36b0cd24),
	.w7(32'h369d8810),
	.w8(32'hb61b2966),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a1c57b),
	.w1(32'h37976baa),
	.w2(32'h3734fd10),
	.w3(32'hb744757a),
	.w4(32'h36c6b771),
	.w5(32'hb6d41f16),
	.w6(32'hb7a910e5),
	.w7(32'hb6e02e14),
	.w8(32'hb5a8e4f0),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69d9f9c),
	.w1(32'hb66637e8),
	.w2(32'hb640122b),
	.w3(32'hb653562c),
	.w4(32'hb70e37ff),
	.w5(32'h362c2470),
	.w6(32'h37dce8d8),
	.w7(32'hb6c9c369),
	.w8(32'h330e8392),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7012758),
	.w1(32'hb6983d1a),
	.w2(32'h369f1e23),
	.w3(32'hb6a7fb4e),
	.w4(32'hb705867d),
	.w5(32'h366736cc),
	.w6(32'h36607b28),
	.w7(32'hb63bbfb4),
	.w8(32'h37308983),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81919c0),
	.w1(32'hb7d91004),
	.w2(32'hb7e38cff),
	.w3(32'hb759cc66),
	.w4(32'hb6f2aaac),
	.w5(32'hb6f8476c),
	.w6(32'hb609c117),
	.w7(32'h37c238c6),
	.w8(32'h3731f45e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6118165),
	.w1(32'hb68c3602),
	.w2(32'h34f487e9),
	.w3(32'hb5e845ee),
	.w4(32'hb61fa078),
	.w5(32'hb6ce867e),
	.w6(32'hb76aa78e),
	.w7(32'h3711b993),
	.w8(32'hb6c2a74a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c406c7),
	.w1(32'h36c26605),
	.w2(32'h3715ae40),
	.w3(32'h369c799c),
	.w4(32'h37d4c9e8),
	.w5(32'h37da3e2d),
	.w6(32'hb6082402),
	.w7(32'hb6788d98),
	.w8(32'h36f4faac),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3703bbc4),
	.w1(32'h383b1e9a),
	.w2(32'h375fd92b),
	.w3(32'hb511ca29),
	.w4(32'h3851aef6),
	.w5(32'h35ff0a78),
	.w6(32'hb7a713e3),
	.w7(32'hb6965f79),
	.w8(32'hb7cdaae9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7008345),
	.w1(32'hb7b139ed),
	.w2(32'hb852dc6a),
	.w3(32'h368e48a9),
	.w4(32'hb7e17052),
	.w5(32'hb8497d50),
	.w6(32'h36563440),
	.w7(32'hb787cf7d),
	.w8(32'hb845378d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388915c3),
	.w1(32'h391146eb),
	.w2(32'h38ec715b),
	.w3(32'h37c62371),
	.w4(32'h38d81bcc),
	.w5(32'h39018820),
	.w6(32'hb71ce342),
	.w7(32'h38df2621),
	.w8(32'h38ff4f3a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h356c9680),
	.w1(32'h36ab01e6),
	.w2(32'hb6ef140d),
	.w3(32'h377690a0),
	.w4(32'hb7cb07bc),
	.w5(32'hb7860c43),
	.w6(32'h37bf937e),
	.w7(32'hb7a5d978),
	.w8(32'hb7867a2b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380398ce),
	.w1(32'h387252b4),
	.w2(32'h38a5feca),
	.w3(32'h37ba2e90),
	.w4(32'h38807246),
	.w5(32'h38688dca),
	.w6(32'h3701c22d),
	.w7(32'h3807343e),
	.w8(32'h37f76291),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79a7e88),
	.w1(32'h3784a3c5),
	.w2(32'h36db4718),
	.w3(32'h38058dd0),
	.w4(32'h37d8c10d),
	.w5(32'h37c89818),
	.w6(32'h37ff0620),
	.w7(32'h381d6d6a),
	.w8(32'h3820000e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e4d03f),
	.w1(32'hb7e8ada9),
	.w2(32'hb83ceddb),
	.w3(32'h37e8fbdf),
	.w4(32'hb7903953),
	.w5(32'h367f0e11),
	.w6(32'h3763319d),
	.w7(32'hb6cb646b),
	.w8(32'h37b1a9d4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36808415),
	.w1(32'hb647025b),
	.w2(32'h3592cb3d),
	.w3(32'hb6491777),
	.w4(32'h360f3b5e),
	.w5(32'h369bd5e6),
	.w6(32'h37194c8a),
	.w7(32'hb701bd0d),
	.w8(32'hb612229f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aeb90c),
	.w1(32'h383354b2),
	.w2(32'h3881d5bb),
	.w3(32'h37b39c08),
	.w4(32'h38419b8c),
	.w5(32'h381fdb1e),
	.w6(32'h3720c9fa),
	.w7(32'h378b8b12),
	.w8(32'h35b18412),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38882b70),
	.w1(32'h38afdd62),
	.w2(32'h38391f96),
	.w3(32'h383db128),
	.w4(32'h386d3b60),
	.w5(32'h370b2b6d),
	.w6(32'h37030296),
	.w7(32'h387dfc34),
	.w8(32'h37704658),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb869239a),
	.w1(32'hb73c314c),
	.w2(32'h387a4fdb),
	.w3(32'hb8e7e9b0),
	.w4(32'hb82ba64e),
	.w5(32'h3892936c),
	.w6(32'hb8d0e84f),
	.w7(32'hb7216934),
	.w8(32'h37a2a850),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37485976),
	.w1(32'hb83a46c8),
	.w2(32'hb8a89b5b),
	.w3(32'hb738846c),
	.w4(32'hb8394af4),
	.w5(32'hb84fdebb),
	.w6(32'h380b37e5),
	.w7(32'hb76ba1ed),
	.w8(32'hb76b2740),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79e388b),
	.w1(32'hb6e8a745),
	.w2(32'hb6d37dae),
	.w3(32'h37b491ab),
	.w4(32'h36e9af2f),
	.w5(32'h37aa1d85),
	.w6(32'h379e6540),
	.w7(32'hb766ddc5),
	.w8(32'h37a2cc4a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3736b678),
	.w1(32'h388ff20c),
	.w2(32'h3872e6e2),
	.w3(32'hb82e8265),
	.w4(32'h382a7bd0),
	.w5(32'h37c9a550),
	.w6(32'hb84adbbf),
	.w7(32'h389ff6ff),
	.w8(32'hb52cce05),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b3b4ce),
	.w1(32'hb6ad3b7f),
	.w2(32'hb2b08471),
	.w3(32'hb7e6e4f5),
	.w4(32'hb68c52b7),
	.w5(32'h372ff313),
	.w6(32'hb7df95bb),
	.w7(32'h35dab04e),
	.w8(32'h379f4f2f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9006990),
	.w1(32'h372d7cac),
	.w2(32'h38e33604),
	.w3(32'hb81649d8),
	.w4(32'h372239d0),
	.w5(32'h39029670),
	.w6(32'hb8d159d8),
	.w7(32'h363c2a4e),
	.w8(32'h37c3f7d3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb698de0c),
	.w1(32'h34985ec4),
	.w2(32'hb790d8bc),
	.w3(32'hb732d181),
	.w4(32'hb74b42d4),
	.w5(32'hb7eaa8e4),
	.w6(32'h365dd81a),
	.w7(32'h35e8ec17),
	.w8(32'hb80610c7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361d89b2),
	.w1(32'h35634198),
	.w2(32'h3733625c),
	.w3(32'hb6b9f228),
	.w4(32'hb66a391d),
	.w5(32'h36ce6610),
	.w6(32'hb6623813),
	.w7(32'hb74d5bef),
	.w8(32'hb5b26e7c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e9327d),
	.w1(32'hb749a894),
	.w2(32'h3797f234),
	.w3(32'hb6143f31),
	.w4(32'hb7778d25),
	.w5(32'h3765ce80),
	.w6(32'hb7972137),
	.w7(32'hb63c3151),
	.w8(32'h37b45d73),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b7e226),
	.w1(32'h380126d3),
	.w2(32'h3853db86),
	.w3(32'h37d50a23),
	.w4(32'h383e7c28),
	.w5(32'h38320bc5),
	.w6(32'h36eb3c7c),
	.w7(32'h37ddd515),
	.w8(32'h37ec414b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6299f90),
	.w1(32'h36d7fd40),
	.w2(32'h360cd368),
	.w3(32'h36d63388),
	.w4(32'hb70f89af),
	.w5(32'h37948e1c),
	.w6(32'hb6748c96),
	.w7(32'h36499783),
	.w8(32'h379b2830),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37292126),
	.w1(32'hb67154e9),
	.w2(32'hb8617bbf),
	.w3(32'h37c4918d),
	.w4(32'h33e57691),
	.w5(32'hb7f9cb10),
	.w6(32'h3780228b),
	.w7(32'hb638621e),
	.w8(32'hb757aef7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b1da95),
	.w1(32'hb7a47856),
	.w2(32'hb718b984),
	.w3(32'h370aac0b),
	.w4(32'h363c4075),
	.w5(32'h37081187),
	.w6(32'hb5defd29),
	.w7(32'hb7366e84),
	.w8(32'h36ff78cf),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80cc4bb),
	.w1(32'hb8081975),
	.w2(32'hb7d51aab),
	.w3(32'hb84244d0),
	.w4(32'hb7ab0113),
	.w5(32'h37a82f37),
	.w6(32'hb82808b2),
	.w7(32'hb6fd7fce),
	.w8(32'h3728e24a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3710306b),
	.w1(32'h36358b70),
	.w2(32'h38476e81),
	.w3(32'h346eac45),
	.w4(32'h378bf673),
	.w5(32'h38a9462d),
	.w6(32'hb73b16b4),
	.w7(32'hb5fed2c4),
	.w8(32'h383283f7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d79efb),
	.w1(32'hb5c3937f),
	.w2(32'h374b138f),
	.w3(32'hb681229e),
	.w4(32'h3624e3e7),
	.w5(32'h370844a8),
	.w6(32'hb71373b1),
	.w7(32'hb6f38bb5),
	.w8(32'hb63a9106),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c29242),
	.w1(32'h35ce45f4),
	.w2(32'h37013eac),
	.w3(32'h359b3f64),
	.w4(32'h36a4440d),
	.w5(32'hb5c29d77),
	.w6(32'hb6a81e39),
	.w7(32'h37356f6b),
	.w8(32'h3700a7bc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb617eedf),
	.w1(32'h36526232),
	.w2(32'hb68b961a),
	.w3(32'h36528708),
	.w4(32'hb58bca67),
	.w5(32'h374e2603),
	.w6(32'h3709a07d),
	.w7(32'hb732d8e7),
	.w8(32'hb6402f91),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3783e509),
	.w1(32'h37a2efee),
	.w2(32'h378bd44d),
	.w3(32'h371ee397),
	.w4(32'h3662b80c),
	.w5(32'hb58ba153),
	.w6(32'h3659a9ad),
	.w7(32'hb73f11f3),
	.w8(32'hb5c3dfc8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a8cfcd),
	.w1(32'hb59a726a),
	.w2(32'hb70c1b8f),
	.w3(32'h37a054aa),
	.w4(32'hb6961dd5),
	.w5(32'hb71a01f0),
	.w6(32'h368a3bf9),
	.w7(32'h3717c0da),
	.w8(32'hb6899908),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7054026),
	.w1(32'hb79ef2ce),
	.w2(32'hb78857a4),
	.w3(32'h35f6cbc6),
	.w4(32'hb72549be),
	.w5(32'hb5c0e3dd),
	.w6(32'h36cc0764),
	.w7(32'hb653a571),
	.w8(32'hb7a27580),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3700b411),
	.w1(32'h35e30719),
	.w2(32'hb51d23ca),
	.w3(32'h36d387bf),
	.w4(32'hb632e666),
	.w5(32'hb5a46e9e),
	.w6(32'h361aaf59),
	.w7(32'h36d54c39),
	.w8(32'hb3670ded),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb633ebb4),
	.w1(32'h37ca4127),
	.w2(32'h37839d9c),
	.w3(32'h36806b9c),
	.w4(32'h37641892),
	.w5(32'h33bda197),
	.w6(32'h36d67340),
	.w7(32'hb46f9ae5),
	.w8(32'hb5fc2ffa),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fb8b60),
	.w1(32'hb7957420),
	.w2(32'hb82eb232),
	.w3(32'hb779c228),
	.w4(32'hb742b4b8),
	.w5(32'hb75212d1),
	.w6(32'hb6d2e568),
	.w7(32'hb7dd18d9),
	.w8(32'hb6321407),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f3f80c),
	.w1(32'h36dba91c),
	.w2(32'hb6b19135),
	.w3(32'hb6d5b07b),
	.w4(32'h367e8e42),
	.w5(32'h36d85067),
	.w6(32'hb549c912),
	.w7(32'h36ed5871),
	.w8(32'h366745d0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6400c47),
	.w1(32'h3780f830),
	.w2(32'h36227227),
	.w3(32'hb6f243be),
	.w4(32'h376e0cea),
	.w5(32'h36f9b3d9),
	.w6(32'h35653128),
	.w7(32'hb6a5334a),
	.w8(32'h375e7913),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371de82a),
	.w1(32'h361879d1),
	.w2(32'hb67fdb9a),
	.w3(32'hb5a84853),
	.w4(32'hb5b5c806),
	.w5(32'h3303fdc4),
	.w6(32'hb549c355),
	.w7(32'h3552c8c3),
	.w8(32'h36dc682b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f56daa),
	.w1(32'hb6363c12),
	.w2(32'h376268ac),
	.w3(32'hb5dd9007),
	.w4(32'hb6c6704a),
	.w5(32'h36994d42),
	.w6(32'h37314abc),
	.w7(32'h36851b1e),
	.w8(32'h35f291dd),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6db0140),
	.w1(32'h3894065a),
	.w2(32'h380b4052),
	.w3(32'hb8846f1e),
	.w4(32'h38b3fce8),
	.w5(32'h38a0e91d),
	.w6(32'hb6dc0c59),
	.w7(32'h3846fa3a),
	.w8(32'h37de27e9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3808736e),
	.w1(32'h386a06a9),
	.w2(32'h38acc69d),
	.w3(32'h37f6fdb8),
	.w4(32'h383309b0),
	.w5(32'h3803813a),
	.w6(32'h37a2bb48),
	.w7(32'h37c64034),
	.w8(32'h373674c8),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64cbb7a),
	.w1(32'h365d7741),
	.w2(32'h374a0b05),
	.w3(32'hb6787fd2),
	.w4(32'h370d281d),
	.w5(32'hb6693f59),
	.w6(32'hb7026613),
	.w7(32'h3754b343),
	.w8(32'hb6c2c1ed),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36478b32),
	.w1(32'h3735b17b),
	.w2(32'hb72f848d),
	.w3(32'hb71c9abd),
	.w4(32'h374c38b3),
	.w5(32'h37855406),
	.w6(32'hb7ad883b),
	.w7(32'hb80b6bf6),
	.w8(32'hb76a9e0c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ea5cbb),
	.w1(32'hb716e82c),
	.w2(32'hb77beb4a),
	.w3(32'h37cd73a6),
	.w4(32'hb7204ef8),
	.w5(32'hb68ee234),
	.w6(32'h36dca2b1),
	.w7(32'hb7834f91),
	.w8(32'h36abb5a4),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d14bab),
	.w1(32'h379c24b3),
	.w2(32'h37ef8b9f),
	.w3(32'hb64088c3),
	.w4(32'h377e1804),
	.w5(32'h379ac746),
	.w6(32'hb7653ab8),
	.w7(32'h36cc4979),
	.w8(32'h377570e4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d17a6c),
	.w1(32'h36b9d60c),
	.w2(32'h37825ccb),
	.w3(32'hb7a1422f),
	.w4(32'h37aebfbe),
	.w5(32'h378c07bf),
	.w6(32'hb7d8c45c),
	.w7(32'h36997f0f),
	.w8(32'h37dcc65a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d874bc),
	.w1(32'h38745590),
	.w2(32'h38aa41c4),
	.w3(32'hb73079dc),
	.w4(32'h386bd86c),
	.w5(32'h37ac6397),
	.w6(32'h36c4463f),
	.w7(32'h37bda691),
	.w8(32'h3782cc18),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7066518),
	.w1(32'hb76ba943),
	.w2(32'hb38be546),
	.w3(32'h37418131),
	.w4(32'h34c5765f),
	.w5(32'h3787356c),
	.w6(32'h36c90184),
	.w7(32'h36d0a575),
	.w8(32'h37b7118c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370e97ca),
	.w1(32'hb7448d23),
	.w2(32'h37dc3c75),
	.w3(32'h37a1cd11),
	.w4(32'h36d9b651),
	.w5(32'h37d9f9b2),
	.w6(32'h37644d99),
	.w7(32'h3739ebf3),
	.w8(32'h379659e1),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360d36af),
	.w1(32'h387a4dd2),
	.w2(32'h3834233d),
	.w3(32'hb7669bc1),
	.w4(32'h3883cc62),
	.w5(32'h37e9c914),
	.w6(32'hb7814954),
	.w7(32'h37808597),
	.w8(32'hb6dc1667),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b08a1e),
	.w1(32'hb6b01ae7),
	.w2(32'hb7390d1c),
	.w3(32'hb7714585),
	.w4(32'h36d7faf5),
	.w5(32'h37dba19b),
	.w6(32'hb66bbd11),
	.w7(32'hb71522b5),
	.w8(32'h37457b12),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66f53e9),
	.w1(32'h3831dc39),
	.w2(32'h385e9317),
	.w3(32'hb64862fe),
	.w4(32'h37c9ebd9),
	.w5(32'h37ad57e8),
	.w6(32'h351664e5),
	.w7(32'h37d7c553),
	.w8(32'h37ab2944),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4a4a87c),
	.w1(32'hb68c320e),
	.w2(32'h3776eb13),
	.w3(32'h371cacb4),
	.w4(32'h36c960bc),
	.w5(32'h375597d5),
	.w6(32'h376bc065),
	.w7(32'h36f96ea8),
	.w8(32'h37abd219),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e449d3),
	.w1(32'hb718718f),
	.w2(32'hb8453320),
	.w3(32'h372a89c4),
	.w4(32'h372c0d8a),
	.w5(32'hb7b7f2c4),
	.w6(32'h36c63dc0),
	.w7(32'h37cbbd94),
	.w8(32'hb70ff563),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70f7c0d),
	.w1(32'h378860c2),
	.w2(32'hb73dbb79),
	.w3(32'hb69c802d),
	.w4(32'h36c6f97f),
	.w5(32'hb6efa946),
	.w6(32'hb753cff4),
	.w7(32'hb68f59bc),
	.w8(32'hb71c7c4b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d9382d),
	.w1(32'h36e06159),
	.w2(32'h3715a416),
	.w3(32'h36151713),
	.w4(32'hb4c18c2a),
	.w5(32'h343b303c),
	.w6(32'h365f6cf1),
	.w7(32'hb5aa31cc),
	.w8(32'h3659ce41),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36936d52),
	.w1(32'h36a37e42),
	.w2(32'hb6b579fd),
	.w3(32'h3687f2b7),
	.w4(32'hb6b50c48),
	.w5(32'h35a76042),
	.w6(32'h37843e1b),
	.w7(32'h3704bc05),
	.w8(32'h36685dad),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6be2d45),
	.w1(32'h376ed025),
	.w2(32'h36bda626),
	.w3(32'h34fa0476),
	.w4(32'h372ff175),
	.w5(32'h3743fef8),
	.w6(32'h37077075),
	.w7(32'h37653b6a),
	.w8(32'h36c82c7a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ca5259),
	.w1(32'hb7ec25a9),
	.w2(32'hb7f9bf56),
	.w3(32'h3699a1f5),
	.w4(32'hb719e45c),
	.w5(32'h3701efa8),
	.w6(32'hb739fd53),
	.w7(32'hb773e5e4),
	.w8(32'h37882a86),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f363c1),
	.w1(32'h3770c32d),
	.w2(32'h37b0b7a1),
	.w3(32'h3665b86b),
	.w4(32'hb780f05a),
	.w5(32'h37a34881),
	.w6(32'hb76f0e08),
	.w7(32'hb72ec5b0),
	.w8(32'hb58b2fe3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6aabdf7),
	.w1(32'h371cf967),
	.w2(32'h35ab3860),
	.w3(32'h371142fc),
	.w4(32'hb617c479),
	.w5(32'hb66a1eff),
	.w6(32'h375c07e7),
	.w7(32'hb7090099),
	.w8(32'hb6ba6720),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f1b5b4),
	.w1(32'h381bff01),
	.w2(32'h3868e22d),
	.w3(32'h3812ba64),
	.w4(32'h37f9f8e8),
	.w5(32'h381ddc78),
	.w6(32'h364c7db4),
	.w7(32'h36ff955e),
	.w8(32'h360ffbf4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f99bd7),
	.w1(32'h36dd3fbd),
	.w2(32'h37d8b2dd),
	.w3(32'h3790c466),
	.w4(32'h37e44d61),
	.w5(32'h3801d2de),
	.w6(32'h369151eb),
	.w7(32'h3667d274),
	.w8(32'h3746edf7),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38013748),
	.w1(32'h3843be7b),
	.w2(32'h389f080b),
	.w3(32'hb5d54880),
	.w4(32'h37e709ee),
	.w5(32'h38339c67),
	.w6(32'hb7b3971c),
	.w7(32'h38075579),
	.w8(32'h38221a9c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb658be22),
	.w1(32'hb7417bfc),
	.w2(32'hb88ec530),
	.w3(32'h379584aa),
	.w4(32'hb69cf313),
	.w5(32'hb801e465),
	.w6(32'h361718c2),
	.w7(32'hb7e194ac),
	.w8(32'hb7f9e58f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3716fd04),
	.w1(32'hb78a1c40),
	.w2(32'hb73be6a7),
	.w3(32'h361a4344),
	.w4(32'hb67825d9),
	.w5(32'hb646189a),
	.w6(32'hb5decb6a),
	.w7(32'hb71d66e7),
	.w8(32'hb612b279),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3731a173),
	.w1(32'h35a2e989),
	.w2(32'hb7a04dbf),
	.w3(32'hb6f0321e),
	.w4(32'h36939904),
	.w5(32'hb6a70c76),
	.w6(32'hb655a561),
	.w7(32'h374a28bb),
	.w8(32'h35a27e19),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374bdcbd),
	.w1(32'h376d9e0d),
	.w2(32'h36c4e80f),
	.w3(32'h378811d8),
	.w4(32'h3709944a),
	.w5(32'h3763133a),
	.w6(32'h37ab36ae),
	.w7(32'h3702a658),
	.w8(32'h362df935),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36460e97),
	.w1(32'hb78bf7c8),
	.w2(32'hb7e16062),
	.w3(32'hb58447aa),
	.w4(32'hb6023839),
	.w5(32'hb6b9432c),
	.w6(32'h3590bee2),
	.w7(32'h374ad344),
	.w8(32'hb6924c64),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369c051d),
	.w1(32'hb6fdb045),
	.w2(32'hb7d7f13c),
	.w3(32'hb728d3e3),
	.w4(32'hb76e5bb4),
	.w5(32'hb797091d),
	.w6(32'hb708a644),
	.w7(32'hb79d7217),
	.w8(32'hb73153f8),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3626f0be),
	.w1(32'h37ac7596),
	.w2(32'h37704c61),
	.w3(32'h360949a1),
	.w4(32'h375fc84a),
	.w5(32'h364cfca1),
	.w6(32'hb61b7550),
	.w7(32'h375ebe5f),
	.w8(32'hb66ddc9b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d59046),
	.w1(32'hb78c1dd0),
	.w2(32'hb768d4f2),
	.w3(32'hb69fee8e),
	.w4(32'hb6d9d9cc),
	.w5(32'hb719b5a5),
	.w6(32'hb731bca6),
	.w7(32'hb73a9cad),
	.w8(32'hb7aba5a4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37532a2a),
	.w1(32'h37357a6a),
	.w2(32'h38254037),
	.w3(32'h376145df),
	.w4(32'h37fa68c1),
	.w5(32'h372b46ff),
	.w6(32'hb6bae893),
	.w7(32'h37def3b1),
	.w8(32'h366fbb1a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66e28bd),
	.w1(32'hb6c87057),
	.w2(32'hb6f2b8da),
	.w3(32'h3532e54c),
	.w4(32'hb6cff4dc),
	.w5(32'hb721ff13),
	.w6(32'h36ce915a),
	.w7(32'hb63cd15a),
	.w8(32'hb76a7a86),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71757e6),
	.w1(32'h376c66ca),
	.w2(32'h359f4047),
	.w3(32'hb6aa2a8f),
	.w4(32'h37bb5f82),
	.w5(32'hb6f124f2),
	.w6(32'h35cf3b85),
	.w7(32'h37af8c5f),
	.w8(32'hb570bf0b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3630d19d),
	.w1(32'h35f8382c),
	.w2(32'h37488cd5),
	.w3(32'hb7a10b1a),
	.w4(32'hb6788a5c),
	.w5(32'h361e3037),
	.w6(32'hb79c4043),
	.w7(32'h36142853),
	.w8(32'h376ad482),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3699862d),
	.w1(32'h35c0e9e1),
	.w2(32'h36c47812),
	.w3(32'hb799bcd8),
	.w4(32'h36c16877),
	.w5(32'h372c2bca),
	.w6(32'hb7094f42),
	.w7(32'h37380ab7),
	.w8(32'h3759aaf6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4807467),
	.w1(32'hb75ee602),
	.w2(32'hb41069fb),
	.w3(32'h3709e959),
	.w4(32'hb6ab8ff9),
	.w5(32'hb6bdddf0),
	.w6(32'h372b6183),
	.w7(32'h367b3922),
	.w8(32'hb6644677),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3607e449),
	.w1(32'hb6b2ffae),
	.w2(32'h35a0fc5c),
	.w3(32'h36026329),
	.w4(32'hb78dde6d),
	.w5(32'h36cbb9cc),
	.w6(32'h3764bd17),
	.w7(32'hb61018b5),
	.w8(32'h36d8e409),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb677dfe5),
	.w1(32'hb7556932),
	.w2(32'hb70de369),
	.w3(32'h35a8c7c3),
	.w4(32'hb5698e6d),
	.w5(32'hb6d15224),
	.w6(32'h374d10bd),
	.w7(32'h3768735d),
	.w8(32'h370e1fc5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7496772),
	.w1(32'h389ca671),
	.w2(32'h38175bc8),
	.w3(32'hb7934e3b),
	.w4(32'h3891ec63),
	.w5(32'h381d7c54),
	.w6(32'hb7c37654),
	.w7(32'h386e2849),
	.w8(32'hb6075565),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374bf24c),
	.w1(32'hb53a45ea),
	.w2(32'hb7052314),
	.w3(32'hb7a80e41),
	.w4(32'hb7917d2c),
	.w5(32'hb746f69c),
	.w6(32'hb729c0e9),
	.w7(32'h36d0e6c3),
	.w8(32'hb6cd0612),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76ce33c),
	.w1(32'hb7e3d2d3),
	.w2(32'hb725c0ad),
	.w3(32'h371f0ec7),
	.w4(32'hb69cd46e),
	.w5(32'h3638921c),
	.w6(32'hb654d09f),
	.w7(32'hb628b356),
	.w8(32'h378e7d13),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb756adcb),
	.w1(32'h35df5f24),
	.w2(32'hb70ff594),
	.w3(32'hb623cc14),
	.w4(32'h36e42695),
	.w5(32'h36a6876a),
	.w6(32'hb62e6ae8),
	.w7(32'h36dd829a),
	.w8(32'h37ad0132),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381bd02e),
	.w1(32'h38094480),
	.w2(32'h386ae95b),
	.w3(32'h37e5e09d),
	.w4(32'h3812700e),
	.w5(32'h3719d8a0),
	.w6(32'h384650cb),
	.w7(32'h377e2988),
	.w8(32'h36bdea7e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5423c35),
	.w1(32'h38020c6d),
	.w2(32'h382b7e86),
	.w3(32'h36807092),
	.w4(32'h3795fba4),
	.w5(32'h37b8d5bc),
	.w6(32'h372f2783),
	.w7(32'h3711f360),
	.w8(32'h37be43bf),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a6bcc0),
	.w1(32'h385d111f),
	.w2(32'h3896b3e8),
	.w3(32'h37ae987e),
	.w4(32'h3803c933),
	.w5(32'h3814f477),
	.w6(32'h37cf06ce),
	.w7(32'h37a7ab8e),
	.w8(32'h37bea1ad),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e6ec77),
	.w1(32'hb7608826),
	.w2(32'h36895704),
	.w3(32'hb5e95558),
	.w4(32'hb79525a6),
	.w5(32'hb6c46c6b),
	.w6(32'hb64253a6),
	.w7(32'hb6cd4864),
	.w8(32'hb67767af),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a48b80),
	.w1(32'h3713c299),
	.w2(32'h374822eb),
	.w3(32'h3785c5f2),
	.w4(32'h37a216f3),
	.w5(32'h3771bf2d),
	.w6(32'h35219bd4),
	.w7(32'h3744ee13),
	.w8(32'h374d9a08),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3599bfeb),
	.w1(32'h376b98f0),
	.w2(32'hb685e415),
	.w3(32'h367b3ca0),
	.w4(32'h3795ad7e),
	.w5(32'hb6a3b564),
	.w6(32'hb56709e8),
	.w7(32'h378392b7),
	.w8(32'hb74732df),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a1efeb),
	.w1(32'h36c9b144),
	.w2(32'h3794db64),
	.w3(32'h377824b5),
	.w4(32'h36b012c6),
	.w5(32'h37628fb4),
	.w6(32'h36235e7b),
	.w7(32'hb6ced14a),
	.w8(32'hb7818601),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3770d5b2),
	.w1(32'hb703af28),
	.w2(32'hb38519a0),
	.w3(32'h368f07e2),
	.w4(32'hb7d87fcb),
	.w5(32'hb62be68a),
	.w6(32'hb6b19fc2),
	.w7(32'hb73285b9),
	.w8(32'h37342dad),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372bd2c5),
	.w1(32'h37e9342b),
	.w2(32'h3824b707),
	.w3(32'h379cf59c),
	.w4(32'h37f6a19a),
	.w5(32'h37fb9fbe),
	.w6(32'h376c2d39),
	.w7(32'h3816a053),
	.w8(32'h3803b0ba),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35108fdb),
	.w1(32'hb7b61210),
	.w2(32'hb4017574),
	.w3(32'hb364584d),
	.w4(32'hb71eaff5),
	.w5(32'hb6b5f1d6),
	.w6(32'h36bc5cac),
	.w7(32'h34d2e50e),
	.w8(32'h36d515b2),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb56f993c),
	.w1(32'hb705d28f),
	.w2(32'hb618d19d),
	.w3(32'hb64224b2),
	.w4(32'hb671afd2),
	.w5(32'hb6f2d828),
	.w6(32'hb729b3fe),
	.w7(32'h36c15a42),
	.w8(32'hb5688f16),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb744fdae),
	.w1(32'hb714f352),
	.w2(32'hb6884421),
	.w3(32'hb78e50db),
	.w4(32'h37472213),
	.w5(32'h3707b78f),
	.w6(32'hb7437946),
	.w7(32'h376f17a1),
	.w8(32'h37880093),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb736b4b6),
	.w1(32'hb51fb6af),
	.w2(32'h37d55c76),
	.w3(32'hb7dc6843),
	.w4(32'hb6c8c381),
	.w5(32'h36dce230),
	.w6(32'hb7aea41f),
	.w7(32'h37559d2f),
	.w8(32'hb6a88a34),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fb35fe),
	.w1(32'hb7c4dc55),
	.w2(32'h3799fcab),
	.w3(32'h3710cb1d),
	.w4(32'hb714c5a4),
	.w5(32'h37fc1bf5),
	.w6(32'hb80d0516),
	.w7(32'hb7d88ec0),
	.w8(32'h379f34ea),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5351fe7),
	.w1(32'h37184b50),
	.w2(32'h362eda20),
	.w3(32'hb64f64e0),
	.w4(32'h37022742),
	.w5(32'hb67526fd),
	.w6(32'h36a173e8),
	.w7(32'h3717b4f0),
	.w8(32'h36c67c6c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e0d754),
	.w1(32'h38b69f51),
	.w2(32'h39169f8a),
	.w3(32'h387d4b1e),
	.w4(32'h3851b0e4),
	.w5(32'h387b8eb0),
	.w6(32'h38742cc5),
	.w7(32'h3805bf80),
	.w8(32'h37365334),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb738a3f9),
	.w1(32'h37585666),
	.w2(32'hb809a3cb),
	.w3(32'h3813d0b4),
	.w4(32'h381770d5),
	.w5(32'h37a2f9e3),
	.w6(32'h35a05f03),
	.w7(32'h3831eaf4),
	.w8(32'h38251054),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb477237e),
	.w1(32'h374b81f2),
	.w2(32'h3732dc8e),
	.w3(32'h37b6b635),
	.w4(32'h36b5d636),
	.w5(32'h37395137),
	.w6(32'h36bac50e),
	.w7(32'h3780b1ca),
	.w8(32'h36f6f5dd),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b93d67),
	.w1(32'h36710876),
	.w2(32'hb70530f4),
	.w3(32'h3459ee03),
	.w4(32'h375369bc),
	.w5(32'hb66805cc),
	.w6(32'hb7025479),
	.w7(32'h3784a715),
	.w8(32'hb6ef65c4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36167308),
	.w1(32'h361340c4),
	.w2(32'h36aeb422),
	.w3(32'hb655bf50),
	.w4(32'h34a717a3),
	.w5(32'h35ef1c3a),
	.w6(32'hb740c75c),
	.w7(32'h36fc942a),
	.w8(32'h371dbc2f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35243afa),
	.w1(32'h32994cd9),
	.w2(32'hb5f13d25),
	.w3(32'hb4bc9cdf),
	.w4(32'h36c9a05e),
	.w5(32'h345a4187),
	.w6(32'h36f15d89),
	.w7(32'h3676de9c),
	.w8(32'h3617e4ef),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3660e86c),
	.w1(32'h37303d58),
	.w2(32'h3667cff5),
	.w3(32'hb6035bf6),
	.w4(32'hb7086ec0),
	.w5(32'h36557fbe),
	.w6(32'hb6fd2e5c),
	.w7(32'h376022f6),
	.w8(32'h37330d41),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80106b6),
	.w1(32'h36259c8f),
	.w2(32'h37b097d4),
	.w3(32'h3536f983),
	.w4(32'h37bc9db6),
	.w5(32'h379555b4),
	.w6(32'h37d1eeff),
	.w7(32'h37c8691e),
	.w8(32'h37a311a4),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7881162),
	.w1(32'hb7c21b8e),
	.w2(32'hb6ac752a),
	.w3(32'h37753f87),
	.w4(32'h36c630cc),
	.w5(32'h37772e9b),
	.w6(32'hb788a007),
	.w7(32'h363f4b45),
	.w8(32'h37870c1b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ca0a2b),
	.w1(32'hb579482f),
	.w2(32'h368e4780),
	.w3(32'h36889582),
	.w4(32'h371e4ea8),
	.w5(32'h374d8d5c),
	.w6(32'hb6e34f83),
	.w7(32'h37baf6bf),
	.w8(32'h36f2e073),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38020c1d),
	.w1(32'hbb325159),
	.w2(32'hbb15bfce),
	.w3(32'h366ad6a9),
	.w4(32'hbb041dc5),
	.w5(32'hbb6b101a),
	.w6(32'hb6d1dc2f),
	.w7(32'hbb0cf6f2),
	.w8(32'h3b8f0e60),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c4803),
	.w1(32'hb95a5fbc),
	.w2(32'h393e1388),
	.w3(32'hbb53bfcd),
	.w4(32'hbb00512f),
	.w5(32'hbad69934),
	.w6(32'hbae1796a),
	.w7(32'hb9d8b292),
	.w8(32'h3a7e2f6d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcb6b4),
	.w1(32'hbb3dd78b),
	.w2(32'h3a312a9e),
	.w3(32'hbb38b515),
	.w4(32'hbbeca511),
	.w5(32'h3bb7ac13),
	.w6(32'hbb3b3684),
	.w7(32'hbadc17eb),
	.w8(32'hbad52e81),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ff2fb),
	.w1(32'h3afe3190),
	.w2(32'h3a3dd364),
	.w3(32'h3a55864f),
	.w4(32'hbb00df49),
	.w5(32'hbb062959),
	.w6(32'hbab09ee8),
	.w7(32'hbb887ed6),
	.w8(32'hb8082554),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c12a93),
	.w1(32'h3a85fec5),
	.w2(32'h389e58bf),
	.w3(32'h3b32146c),
	.w4(32'h3bb2edba),
	.w5(32'h3ad3c6a9),
	.w6(32'hb9a153da),
	.w7(32'h3b3469af),
	.w8(32'h3aeb47fe),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb893192),
	.w1(32'h3b8d12af),
	.w2(32'hbb51993c),
	.w3(32'hbb85f008),
	.w4(32'h3a76d570),
	.w5(32'h3bc96386),
	.w6(32'hba0878de),
	.w7(32'hbb072e79),
	.w8(32'hba515e18),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53bb0a),
	.w1(32'h3a31441a),
	.w2(32'hbb82dc46),
	.w3(32'h3b956bc4),
	.w4(32'h3ad61701),
	.w5(32'h3b8ac32e),
	.w6(32'h3c0531f3),
	.w7(32'h3b6b1f1c),
	.w8(32'h3b9349f4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab593ce),
	.w1(32'hba0f74f4),
	.w2(32'h3b2a169c),
	.w3(32'h3b2bb187),
	.w4(32'hbb5469c7),
	.w5(32'hbb2fde3e),
	.w6(32'h3bd19807),
	.w7(32'hbab6d3f2),
	.w8(32'h3b1e4e9c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb872136),
	.w1(32'hbb23d216),
	.w2(32'hbc072d7b),
	.w3(32'hb9a4e09d),
	.w4(32'h3c45b789),
	.w5(32'h3cc03638),
	.w6(32'hbaebc475),
	.w7(32'hbc2939c4),
	.w8(32'hb98ac108),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdacfb7),
	.w1(32'hbb473c3a),
	.w2(32'hbb7c7e7a),
	.w3(32'hbb57db3a),
	.w4(32'h3b76f2e6),
	.w5(32'h3c06458d),
	.w6(32'h3b8e58c1),
	.w7(32'h39eaa069),
	.w8(32'h3b649539),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06c4d9),
	.w1(32'hbb13b5a5),
	.w2(32'h39156f5b),
	.w3(32'h3aec0148),
	.w4(32'hbc1068c7),
	.w5(32'hb90994da),
	.w6(32'h3b7b8db7),
	.w7(32'hbc13e3b0),
	.w8(32'hbc0e0cf8),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba070190),
	.w1(32'h3c3baa6f),
	.w2(32'h3b9bbd54),
	.w3(32'hb8eaff5b),
	.w4(32'h3a8c634d),
	.w5(32'h3b99da88),
	.w6(32'hbbce8ca1),
	.w7(32'hbb171409),
	.w8(32'hbb397bd2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b302930),
	.w1(32'h3abc8adc),
	.w2(32'hbaf860cd),
	.w3(32'h3b772c86),
	.w4(32'h39c3661e),
	.w5(32'hba9545f6),
	.w6(32'hba6a5b5e),
	.w7(32'hbb1c09d9),
	.w8(32'hbb018658),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16064f),
	.w1(32'hbb7c89cb),
	.w2(32'hbb33428f),
	.w3(32'hb8c05946),
	.w4(32'hbb36459c),
	.w5(32'hbb393be2),
	.w6(32'hbb191ebd),
	.w7(32'hbb1fad92),
	.w8(32'hbbaeabde),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97eb6bb),
	.w1(32'hbb88ef08),
	.w2(32'hbb188601),
	.w3(32'h3b7ea660),
	.w4(32'hbbc674b1),
	.w5(32'hbbd006f8),
	.w6(32'hbb0339f4),
	.w7(32'hbb4a5836),
	.w8(32'hbaaf784f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c096552),
	.w1(32'h3af181c5),
	.w2(32'h3b4a0996),
	.w3(32'hbb2003c4),
	.w4(32'hba8edbd7),
	.w5(32'h3b95c849),
	.w6(32'h3b52e379),
	.w7(32'hbb755de6),
	.w8(32'h3a8534cb),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c98b4),
	.w1(32'h3aa786d4),
	.w2(32'hbb1f78a7),
	.w3(32'h3b7cae2d),
	.w4(32'h3aec8705),
	.w5(32'h3ba7e84f),
	.w6(32'hbacf13ea),
	.w7(32'hbaa072fe),
	.w8(32'h3ba8efad),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97cdadf),
	.w1(32'hbbd2f10a),
	.w2(32'hbc4c0c0e),
	.w3(32'h3ad1658d),
	.w4(32'h3c3b22e7),
	.w5(32'h3c59ddc3),
	.w6(32'h3c02b2d1),
	.w7(32'hbaa5ac01),
	.w8(32'h3b4a8bed),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb8622),
	.w1(32'hb99f0e67),
	.w2(32'hbb6e5eb2),
	.w3(32'hbb40f02e),
	.w4(32'h3c72968c),
	.w5(32'h3c0c4142),
	.w6(32'h3b70270b),
	.w7(32'h3ae895a8),
	.w8(32'h3bd70bbb),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80ba56),
	.w1(32'hbb5b725d),
	.w2(32'hbaf4380b),
	.w3(32'h3a7ac30c),
	.w4(32'hbb793c4a),
	.w5(32'h3b2e1f7c),
	.w6(32'h3c1de572),
	.w7(32'hbb5d1dd8),
	.w8(32'hbb92ccd5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0f161),
	.w1(32'hbb340476),
	.w2(32'hbb4c4498),
	.w3(32'h3aec4b40),
	.w4(32'h3bdba11e),
	.w5(32'h3c11dd9b),
	.w6(32'hbb809e86),
	.w7(32'h3bdc1c5f),
	.w8(32'h3bb5e1c0),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8db521),
	.w1(32'h3b77f5ee),
	.w2(32'hba45be2c),
	.w3(32'hba01f806),
	.w4(32'h3b7016e9),
	.w5(32'h3a81ac69),
	.w6(32'h393d7e44),
	.w7(32'h39a52357),
	.w8(32'h3b20e957),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b293a),
	.w1(32'h3b304a9f),
	.w2(32'h3b8b07bb),
	.w3(32'hba273016),
	.w4(32'hbb02f0d6),
	.w5(32'hbb8012bc),
	.w6(32'h3ab35fb3),
	.w7(32'h3689e6d8),
	.w8(32'hbafdde52),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c378e7),
	.w1(32'h39cb8f0a),
	.w2(32'h3bb50a90),
	.w3(32'hbbbd17d5),
	.w4(32'hbc22e6b2),
	.w5(32'hbb8a16cb),
	.w6(32'h3b3cc067),
	.w7(32'hb9f7a35c),
	.w8(32'hbba53cb6),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bf77c),
	.w1(32'hb9a11977),
	.w2(32'h3a51b54d),
	.w3(32'h3bb666c2),
	.w4(32'hb80b7cc1),
	.w5(32'hbad42b1b),
	.w6(32'hbc032593),
	.w7(32'h3b545aea),
	.w8(32'h38fa2752),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f71ea),
	.w1(32'hbb1a6d72),
	.w2(32'hbb126d43),
	.w3(32'hbb25c36e),
	.w4(32'hbb7e35bd),
	.w5(32'hbb04f349),
	.w6(32'hbab59da3),
	.w7(32'hbbaecd42),
	.w8(32'hbc2362c6),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb676228),
	.w1(32'hbb0520e9),
	.w2(32'h3af15b2e),
	.w3(32'h3b58808c),
	.w4(32'hbbb33c08),
	.w5(32'hbc821b2b),
	.w6(32'hbb847049),
	.w7(32'h3bd0e437),
	.w8(32'hbaab79ef),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19dd04),
	.w1(32'hbb1706e5),
	.w2(32'h3ac2bd4d),
	.w3(32'hbc0d5812),
	.w4(32'hbb9033c2),
	.w5(32'hbc1bd49f),
	.w6(32'hbb2880b1),
	.w7(32'hbb3ec8f8),
	.w8(32'h3a957615),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae924e3),
	.w1(32'hbab896df),
	.w2(32'hbb21f0f7),
	.w3(32'hbb503794),
	.w4(32'h3befdfaa),
	.w5(32'hbadc41dc),
	.w6(32'h3a441664),
	.w7(32'h3b272a3b),
	.w8(32'h3b823e83),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914ad2c),
	.w1(32'hbb5c9522),
	.w2(32'hbb29986d),
	.w3(32'hbb735d3c),
	.w4(32'h3b81cca0),
	.w5(32'hbb1afae9),
	.w6(32'hbac3f614),
	.w7(32'h3be263d8),
	.w8(32'h3be7a838),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb226c06),
	.w1(32'hbb7c3490),
	.w2(32'h3b2f99c3),
	.w3(32'hbb23d22e),
	.w4(32'hbb0b8d6b),
	.w5(32'hbbb9a0d0),
	.w6(32'hb9c60afc),
	.w7(32'hba6614f0),
	.w8(32'h3b9b4897),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b621173),
	.w1(32'hbb16cbf7),
	.w2(32'hbb26e66c),
	.w3(32'hbbf5c7e5),
	.w4(32'h3b7284e2),
	.w5(32'hb992102f),
	.w6(32'h39c66b2b),
	.w7(32'h3b72a727),
	.w8(32'h3b48a678),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e0dc1),
	.w1(32'hbb598908),
	.w2(32'h39060490),
	.w3(32'hbb77cdc2),
	.w4(32'hbb682c67),
	.w5(32'hbae9acbe),
	.w6(32'hbaf32624),
	.w7(32'h3b0ba372),
	.w8(32'h3abd2bc8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8c54a),
	.w1(32'hb9c378b8),
	.w2(32'hbb0b400e),
	.w3(32'h3b3bfee8),
	.w4(32'h3c28d9f5),
	.w5(32'hbb60c15e),
	.w6(32'hbbbca7cc),
	.w7(32'h3bc8b0d6),
	.w8(32'h3b00972f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed1abe),
	.w1(32'hbb8490e4),
	.w2(32'hbb65c10f),
	.w3(32'hbb2f29c0),
	.w4(32'h3a4507c7),
	.w5(32'h3b7e6f57),
	.w6(32'h3b939ab2),
	.w7(32'h39dc9844),
	.w8(32'h3ba05728),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafff6c6),
	.w1(32'h3b24ca0c),
	.w2(32'h3b9e0933),
	.w3(32'h3b75873b),
	.w4(32'hbc035b06),
	.w5(32'hb9954de7),
	.w6(32'h3a8dfbf4),
	.w7(32'hb91a4269),
	.w8(32'hbb8279c4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30a073),
	.w1(32'h3b20cfff),
	.w2(32'h3ae72f4b),
	.w3(32'h3ba1bd8e),
	.w4(32'hba56569e),
	.w5(32'hbb010694),
	.w6(32'hbb6c8215),
	.w7(32'hbab6a3d4),
	.w8(32'hbbad19b3),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c6fde),
	.w1(32'hbbb26746),
	.w2(32'hbbc9015e),
	.w3(32'hbaf9866e),
	.w4(32'hba981e85),
	.w5(32'hba427078),
	.w6(32'hbb0d9db0),
	.w7(32'hba51b2a2),
	.w8(32'hbaecc458),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93e087),
	.w1(32'h3b3a19bf),
	.w2(32'hbaf02824),
	.w3(32'hbb1a33b9),
	.w4(32'h37bb7c89),
	.w5(32'hb90f3b4a),
	.w6(32'hbb35e56a),
	.w7(32'h3a42a692),
	.w8(32'hba4445f3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eae024),
	.w1(32'hbae9e0ef),
	.w2(32'h3a8ea1b0),
	.w3(32'hbb8d4fab),
	.w4(32'hbb835431),
	.w5(32'hbb85af1b),
	.w6(32'hbb4eaf79),
	.w7(32'hba84679c),
	.w8(32'hbbaef154),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c0c48),
	.w1(32'h3b15764f),
	.w2(32'h3ba1ec99),
	.w3(32'h3aa71210),
	.w4(32'hbc1bd73d),
	.w5(32'h3a5d1dad),
	.w6(32'hbbbab088),
	.w7(32'h3b14b7e6),
	.w8(32'hbaec86d2),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e34ca),
	.w1(32'hbb9ec3bf),
	.w2(32'h393bfd35),
	.w3(32'h3b8a3a15),
	.w4(32'h3a44b5cb),
	.w5(32'hba29cd9d),
	.w6(32'hbbcfdf5c),
	.w7(32'h3acdf3bb),
	.w8(32'h3b139365),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d93cd),
	.w1(32'h3a0d0972),
	.w2(32'h3b95e5ce),
	.w3(32'h3b184387),
	.w4(32'hbb5be5b5),
	.w5(32'hbb4267e4),
	.w6(32'h38c03546),
	.w7(32'hba9c6c84),
	.w8(32'hbb949570),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84bff9),
	.w1(32'h3b39f2d8),
	.w2(32'h3b1e7ba6),
	.w3(32'hbad4bfb1),
	.w4(32'h3a90d6b8),
	.w5(32'hbc214b91),
	.w6(32'hbb619cb1),
	.w7(32'h3a021984),
	.w8(32'hba9f337a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fbe26),
	.w1(32'hba0d778a),
	.w2(32'hb8d5023c),
	.w3(32'hbb95233c),
	.w4(32'h3a9ea40b),
	.w5(32'h3c123dc4),
	.w6(32'hbb83d3c3),
	.w7(32'h3aa3a43f),
	.w8(32'h3b4ba397),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d1d2b),
	.w1(32'hbb325cc5),
	.w2(32'hbb4b458c),
	.w3(32'h3b72fd20),
	.w4(32'h38ec92c7),
	.w5(32'hbb4fd7c9),
	.w6(32'h3b43b769),
	.w7(32'h393b9085),
	.w8(32'hba61996c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2568f),
	.w1(32'h3ab5c451),
	.w2(32'hb9ea6447),
	.w3(32'hbb918515),
	.w4(32'h3b1881f5),
	.w5(32'h3b52576d),
	.w6(32'hbaff43ca),
	.w7(32'h3b2c9b00),
	.w8(32'h3ac0870d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a764b8),
	.w1(32'h3bf57904),
	.w2(32'h3b04565d),
	.w3(32'h382abb30),
	.w4(32'hbb36c869),
	.w5(32'hbba37e9f),
	.w6(32'h3b007fe1),
	.w7(32'h3b608f28),
	.w8(32'hba7ea2e6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82bc3d),
	.w1(32'hbabba8e9),
	.w2(32'h3b7ce5f4),
	.w3(32'h3b0da9f9),
	.w4(32'hbbb5086c),
	.w5(32'hbb43cc25),
	.w6(32'hba22b56a),
	.w7(32'hbb0b966f),
	.w8(32'hbaadaf88),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba36a87),
	.w1(32'hbae56a2c),
	.w2(32'hbb8495d1),
	.w3(32'hb906a505),
	.w4(32'h3bfda5e9),
	.w5(32'h3c22f71e),
	.w6(32'hbb94ff6c),
	.w7(32'h3ae1e4cd),
	.w8(32'h3b64a794),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01f7fd),
	.w1(32'h3a196d43),
	.w2(32'h3b0674d6),
	.w3(32'h3ad120a6),
	.w4(32'h3ad948b8),
	.w5(32'hbad16ea3),
	.w6(32'h3bf74ac4),
	.w7(32'h3bec0428),
	.w8(32'h3a1d713b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f1b1f),
	.w1(32'hb90ff119),
	.w2(32'hba2d98c0),
	.w3(32'hbb0cdfd5),
	.w4(32'hbb61d4f1),
	.w5(32'h3a03493b),
	.w6(32'h3a1e3060),
	.w7(32'hbae80e96),
	.w8(32'h3b31fa53),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38041142),
	.w1(32'h3bec16d9),
	.w2(32'h3bb0725f),
	.w3(32'h3ba2d437),
	.w4(32'hb792e10b),
	.w5(32'hbb1fe48d),
	.w6(32'hba926314),
	.w7(32'h3b5def75),
	.w8(32'h3bb49656),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7cc51),
	.w1(32'h3b83805d),
	.w2(32'h3b40fdb0),
	.w3(32'h390177e2),
	.w4(32'h3ae91159),
	.w5(32'hbb94a59e),
	.w6(32'h3bfa7949),
	.w7(32'hbb9e884a),
	.w8(32'hb9064a8f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa91dd),
	.w1(32'h3bf3cbd3),
	.w2(32'h3bbee1ef),
	.w3(32'h39fab35f),
	.w4(32'hbbb80af8),
	.w5(32'hbbfe6b63),
	.w6(32'h373be22b),
	.w7(32'h3ab1e70c),
	.w8(32'hbaf4503e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee0730),
	.w1(32'h3a1856de),
	.w2(32'h3b60f80b),
	.w3(32'hba8fc892),
	.w4(32'hbc14280b),
	.w5(32'h3ba3b580),
	.w6(32'hbc1e5836),
	.w7(32'h3ae97264),
	.w8(32'hb96fc890),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba626556),
	.w1(32'hbba92dc0),
	.w2(32'hbbcda57b),
	.w3(32'h3bca4bcb),
	.w4(32'hbbd114f2),
	.w5(32'h3ad09c69),
	.w6(32'hbbaeced6),
	.w7(32'hbaed3132),
	.w8(32'h3a1e3dc6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9843b5f),
	.w1(32'hbb9f586b),
	.w2(32'hbb207f79),
	.w3(32'hb8e6c845),
	.w4(32'hbb40fe97),
	.w5(32'hbb71b03c),
	.w6(32'hbb475808),
	.w7(32'hbb949cde),
	.w8(32'hba20c2b0),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ba059),
	.w1(32'hbb87903b),
	.w2(32'hbb05ec02),
	.w3(32'hbb5dc924),
	.w4(32'hbae603fd),
	.w5(32'hba019173),
	.w6(32'h3a8a8302),
	.w7(32'h3ad78b66),
	.w8(32'h3a86dee3),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule