module layer_10_featuremap_279(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f2c93),
	.w1(32'h3a6ab84a),
	.w2(32'h3a5ee77f),
	.w3(32'h3a8d130c),
	.w4(32'h3a7dd212),
	.w5(32'h39ed53fd),
	.w6(32'h3a90e54f),
	.w7(32'h3a2e0f68),
	.w8(32'h3a150faf),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15208b),
	.w1(32'h3a01d0ff),
	.w2(32'h39e26bcf),
	.w3(32'h3a04a2fb),
	.w4(32'h3a269793),
	.w5(32'h387af1a0),
	.w6(32'h39d0c916),
	.w7(32'h3a028b01),
	.w8(32'h379c98c1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39293f7b),
	.w1(32'hb9d7426b),
	.w2(32'h39925078),
	.w3(32'hba13a221),
	.w4(32'h39b19574),
	.w5(32'h3861765b),
	.w6(32'hb9b37d97),
	.w7(32'h39dbca76),
	.w8(32'h39ac5c09),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3948899b),
	.w1(32'h3987af55),
	.w2(32'hb95701f0),
	.w3(32'h392d73b0),
	.w4(32'hb9468651),
	.w5(32'h3986581e),
	.w6(32'h39dddb43),
	.w7(32'hb8ea40ca),
	.w8(32'h39b13f77),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07eeff),
	.w1(32'hb9770935),
	.w2(32'h39d57c92),
	.w3(32'hb9ed098b),
	.w4(32'h37a6706b),
	.w5(32'hba2683a8),
	.w6(32'hb990ea73),
	.w7(32'h39a30f40),
	.w8(32'hba03a783),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cdd93),
	.w1(32'hb9af306a),
	.w2(32'hb9bd17d5),
	.w3(32'hb9a92462),
	.w4(32'hb9af0dcc),
	.w5(32'hb90305f0),
	.w6(32'hb891eca2),
	.w7(32'hb989bbb8),
	.w8(32'hb835d3b7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6a13b),
	.w1(32'hb9542f9c),
	.w2(32'hb931abff),
	.w3(32'hb6a6ec5c),
	.w4(32'hb9958f83),
	.w5(32'h37f9f751),
	.w6(32'h39e46af7),
	.w7(32'h3811e49b),
	.w8(32'hb8bec698),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a474f5),
	.w1(32'hb9a8aff1),
	.w2(32'hb9a2d054),
	.w3(32'hb8d40308),
	.w4(32'h38e4e403),
	.w5(32'h3a058aba),
	.w6(32'h39f6024e),
	.w7(32'hb953df1d),
	.w8(32'h39f2fd43),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397794d1),
	.w1(32'h39d4912a),
	.w2(32'h39d49560),
	.w3(32'h3a446671),
	.w4(32'h3a10f87e),
	.w5(32'hba0fab13),
	.w6(32'h3a18ed4e),
	.w7(32'h3a0013bf),
	.w8(32'hb9f13aaa),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30d9d5),
	.w1(32'hba239c11),
	.w2(32'hba04d03e),
	.w3(32'hb9ed17b7),
	.w4(32'hba121a68),
	.w5(32'h395a39ca),
	.w6(32'hb978eb33),
	.w7(32'hba00f344),
	.w8(32'h39ac75c7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2d2ac),
	.w1(32'h39a4e692),
	.w2(32'h38e880f4),
	.w3(32'h3a0e2a5d),
	.w4(32'h3977cce3),
	.w5(32'hb9397068),
	.w6(32'h3a2cf61d),
	.w7(32'h39487532),
	.w8(32'hb884ee22),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d8da7d),
	.w1(32'hb938246b),
	.w2(32'hb7be3b9c),
	.w3(32'hba06afe2),
	.w4(32'hb94b03f9),
	.w5(32'hb89f0e48),
	.w6(32'hba2979e4),
	.w7(32'hb9bb8a29),
	.w8(32'h3995de56),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9bbb9),
	.w1(32'h391889f0),
	.w2(32'h3a00a4f2),
	.w3(32'hb959ecb2),
	.w4(32'hb95eb3e1),
	.w5(32'h3a4a621a),
	.w6(32'hb9f7c552),
	.w7(32'hb8a3e540),
	.w8(32'h39c41d4a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e3b25),
	.w1(32'h3a2d5a55),
	.w2(32'h3a8fff49),
	.w3(32'h3a36caa4),
	.w4(32'h3a36d67a),
	.w5(32'hb8f66f03),
	.w6(32'h39c9cca6),
	.w7(32'h3a15da46),
	.w8(32'h3924c5cb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39161e4d),
	.w1(32'h384a7b91),
	.w2(32'hb616fcc1),
	.w3(32'hb8952bb5),
	.w4(32'hb9a552e7),
	.w5(32'hb91a57da),
	.w6(32'h3959ec67),
	.w7(32'h39016f1a),
	.w8(32'hb9e4b32d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d73d15),
	.w1(32'hb728282d),
	.w2(32'hb8e62f7e),
	.w3(32'h3967c2f3),
	.w4(32'hb7ab7b6c),
	.w5(32'h39427d0e),
	.w6(32'hb3852e6b),
	.w7(32'hb9af8036),
	.w8(32'h39d5ae88),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e15ddc),
	.w1(32'h3934de1f),
	.w2(32'h39de15e5),
	.w3(32'h39e4fc08),
	.w4(32'h391d41c1),
	.w5(32'hba559a19),
	.w6(32'h3984f286),
	.w7(32'h38cbabb4),
	.w8(32'hba287f14),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fea7f),
	.w1(32'hb9ef0dbf),
	.w2(32'hb951ac82),
	.w3(32'hba15e93f),
	.w4(32'hb9ba288a),
	.w5(32'hb912f187),
	.w6(32'hb9c1500a),
	.w7(32'hb7e069a0),
	.w8(32'h396fe01b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38909b12),
	.w1(32'hba152b84),
	.w2(32'hb9b22058),
	.w3(32'hb999ec81),
	.w4(32'h39f6f244),
	.w5(32'h3841c2f0),
	.w6(32'h392a349c),
	.w7(32'h397141d0),
	.w8(32'hb950ad5a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8873899),
	.w1(32'hb8523306),
	.w2(32'h39fc051e),
	.w3(32'h3926321b),
	.w4(32'h39370a7e),
	.w5(32'h3a58c7f5),
	.w6(32'hb93efa8b),
	.w7(32'h389aeb3f),
	.w8(32'h3a050e2f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a127d95),
	.w1(32'h3a9664c9),
	.w2(32'h39fd3900),
	.w3(32'h3a967f0e),
	.w4(32'h3a454260),
	.w5(32'hb9e6fecb),
	.w6(32'h3a79c0db),
	.w7(32'h39f77ff1),
	.w8(32'hb9c87ddb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfd814),
	.w1(32'hb95583d9),
	.w2(32'hb9747953),
	.w3(32'hb9eff7c7),
	.w4(32'hba0600e2),
	.w5(32'hb8f44802),
	.w6(32'hb99b3b5a),
	.w7(32'hb9c930ea),
	.w8(32'hb8b83f75),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369990f4),
	.w1(32'hb934cd26),
	.w2(32'hb95a6fb7),
	.w3(32'hb9368c8b),
	.w4(32'hb934407a),
	.w5(32'h39c4a1e5),
	.w6(32'hb94269c0),
	.w7(32'h383e2abd),
	.w8(32'h39a1ef1b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca00ce),
	.w1(32'h391d97cd),
	.w2(32'hb91aee82),
	.w3(32'h3a74a5d2),
	.w4(32'h39b7f19c),
	.w5(32'hb5e303f2),
	.w6(32'h3a3e3f2b),
	.w7(32'h34ed2064),
	.w8(32'hba006c05),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86d6a2),
	.w1(32'hba655893),
	.w2(32'hba1b1d39),
	.w3(32'hb92124f1),
	.w4(32'h38fdc5c2),
	.w5(32'hb89a0115),
	.w6(32'h385f80d5),
	.w7(32'h38e65cc1),
	.w8(32'hb969cb39),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f9895),
	.w1(32'hb980e6bb),
	.w2(32'hb92a2f18),
	.w3(32'hb8f45190),
	.w4(32'hb9ae2751),
	.w5(32'hba5a3b46),
	.w6(32'h39ac7f26),
	.w7(32'hb880bccb),
	.w8(32'hba7f5087),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba469f0a),
	.w1(32'hbaaeb4e2),
	.w2(32'hba48b655),
	.w3(32'hbaa64679),
	.w4(32'hba5d701d),
	.w5(32'h38a395f5),
	.w6(32'hbaa59a95),
	.w7(32'hba819734),
	.w8(32'hb7963036),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb950c64b),
	.w1(32'h383d2671),
	.w2(32'h39af3038),
	.w3(32'h38a90d60),
	.w4(32'h3999b387),
	.w5(32'h39de0b97),
	.w6(32'hb881e6d5),
	.w7(32'h39d0c79c),
	.w8(32'h39135124),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c39ebb),
	.w1(32'hb982dcef),
	.w2(32'h395f95a4),
	.w3(32'h3a2167f9),
	.w4(32'h348f2f1f),
	.w5(32'h3874bbef),
	.w6(32'h3a1dd4fe),
	.w7(32'h38bf348d),
	.w8(32'hb85c80d7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92da6f0),
	.w1(32'h373abf87),
	.w2(32'h3a0e3269),
	.w3(32'h3994e4ee),
	.w4(32'h3a031960),
	.w5(32'hb8bacc98),
	.w6(32'hb9073d02),
	.w7(32'h3955f948),
	.w8(32'hba2f5955),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e2f84b),
	.w1(32'hb8e8055b),
	.w2(32'h39ae4929),
	.w3(32'hba637fb9),
	.w4(32'hba1c9605),
	.w5(32'hb7e8c603),
	.w6(32'hb9a14c2a),
	.w7(32'hb9a394fa),
	.w8(32'h38bfa98f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a85b33),
	.w1(32'hb81bb182),
	.w2(32'h39b24c5b),
	.w3(32'hb96cdf7f),
	.w4(32'h38f2e2ab),
	.w5(32'hba64d1ec),
	.w6(32'hb95bf0c3),
	.w7(32'h393b13e7),
	.w8(32'hbabe10d0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba548e05),
	.w1(32'hba77d14b),
	.w2(32'hba661510),
	.w3(32'hba3ee1b3),
	.w4(32'hba01c4c7),
	.w5(32'hba85ed32),
	.w6(32'hba3e03db),
	.w7(32'hbaa3f76d),
	.w8(32'hba54c242),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5691e9),
	.w1(32'hba193ba3),
	.w2(32'hb9a2beb4),
	.w3(32'hb9c678b4),
	.w4(32'hb9160722),
	.w5(32'h39d65c55),
	.w6(32'hba2240b7),
	.w7(32'hb9cf0241),
	.w8(32'h39300676),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ea7b8),
	.w1(32'hb9be383e),
	.w2(32'hb9bdfe6e),
	.w3(32'hb7d068fa),
	.w4(32'hb8ff3ef2),
	.w5(32'h39825441),
	.w6(32'hb9468c09),
	.w7(32'hb9050fe7),
	.w8(32'hb8686547),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7636a),
	.w1(32'hba35fe45),
	.w2(32'hbab98449),
	.w3(32'h3933dde7),
	.w4(32'hb900a807),
	.w5(32'hb9efa152),
	.w6(32'hb9523d4e),
	.w7(32'hba3f9685),
	.w8(32'hba85f357),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba885f9f),
	.w1(32'hba789c7a),
	.w2(32'hba332ead),
	.w3(32'hba9c0d3f),
	.w4(32'hba8b4f01),
	.w5(32'hba2b385a),
	.w6(32'hba9322e8),
	.w7(32'hbab86a16),
	.w8(32'hba49805b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b722d9),
	.w1(32'hb983b574),
	.w2(32'h38f1a4cc),
	.w3(32'hb8ec7608),
	.w4(32'h397e16aa),
	.w5(32'h3a2d74c4),
	.w6(32'hb84fdd78),
	.w7(32'h3816908a),
	.w8(32'h3a24d68e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ba76e),
	.w1(32'h39669b12),
	.w2(32'h39c0f905),
	.w3(32'h398d39b5),
	.w4(32'h3a4fcff0),
	.w5(32'h3a8b5fc4),
	.w6(32'h3811aa86),
	.w7(32'h3a2312c7),
	.w8(32'h3a756521),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d7da1),
	.w1(32'h3a1261ee),
	.w2(32'hb9a30322),
	.w3(32'h3a453bf5),
	.w4(32'hb8507eec),
	.w5(32'h3912a4bf),
	.w6(32'h3a8cd461),
	.w7(32'hb93e083a),
	.w8(32'h38b34ef3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9de47),
	.w1(32'h39cb5785),
	.w2(32'h39a8234f),
	.w3(32'h39eb8aec),
	.w4(32'h3921eb53),
	.w5(32'hb9d7e2f1),
	.w6(32'hb79c7029),
	.w7(32'h38fffeff),
	.w8(32'hb9bf601d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5c11f),
	.w1(32'hb9e18a84),
	.w2(32'hba07ab19),
	.w3(32'hb9bd9c59),
	.w4(32'hba349530),
	.w5(32'h3a1a3bed),
	.w6(32'h3960e33b),
	.w7(32'hb9cba869),
	.w8(32'h3a0a710a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397805c8),
	.w1(32'hb9ce010a),
	.w2(32'h397e8b32),
	.w3(32'h39c4b521),
	.w4(32'h3a8c4e58),
	.w5(32'hb9de546b),
	.w6(32'hb8b1c3bd),
	.w7(32'h3a817282),
	.w8(32'hbaaaaa9e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86bd5b),
	.w1(32'hbb08933d),
	.w2(32'hba16a238),
	.w3(32'hbab1775b),
	.w4(32'hba224e8d),
	.w5(32'hb9cbf10d),
	.w6(32'hbb29997f),
	.w7(32'hbab054e7),
	.w8(32'hba045efe),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03f588),
	.w1(32'hb95e9302),
	.w2(32'hba0ade8d),
	.w3(32'hb95778ba),
	.w4(32'hb9fd6c9a),
	.w5(32'h3a3ee3fc),
	.w6(32'hb8c9e8fc),
	.w7(32'hba09e9ef),
	.w8(32'h39ab0596),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39636d68),
	.w1(32'h399c40eb),
	.w2(32'h394c3fe7),
	.w3(32'h397ef654),
	.w4(32'h39879e6d),
	.w5(32'hb96b39f0),
	.w6(32'h3a1319e1),
	.w7(32'h3987a99c),
	.w8(32'hba14d727),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a221ed),
	.w1(32'hb961dee8),
	.w2(32'hb93508c1),
	.w3(32'hb98bc4b0),
	.w4(32'h38dbf299),
	.w5(32'h3a8bd80e),
	.w6(32'hba003153),
	.w7(32'hb9bd632d),
	.w8(32'h3aa5c29c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a762d95),
	.w1(32'h3aa24740),
	.w2(32'h3a8a20be),
	.w3(32'h3a6a1b35),
	.w4(32'h3a18a602),
	.w5(32'h39d74982),
	.w6(32'h3a96ca1e),
	.w7(32'h3a518b40),
	.w8(32'h3a209f70),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c0302),
	.w1(32'h3a08afe6),
	.w2(32'h3a0d1b7c),
	.w3(32'h39d6f58c),
	.w4(32'h398bcac6),
	.w5(32'hb697b989),
	.w6(32'h39af76da),
	.w7(32'h39b84276),
	.w8(32'h398b0a9f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a2d76d),
	.w1(32'h3995f45a),
	.w2(32'h394001b6),
	.w3(32'h394cb5f1),
	.w4(32'hb711a9c9),
	.w5(32'hb9b9ac40),
	.w6(32'h3a3835b8),
	.w7(32'h390dcf62),
	.w8(32'hb9f326b7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904d474),
	.w1(32'hba6d184c),
	.w2(32'hba1e8bf1),
	.w3(32'hbaab4a65),
	.w4(32'hba3109ea),
	.w5(32'h3923bb53),
	.w6(32'hba958b9f),
	.w7(32'hba4bb595),
	.w8(32'hb9040518),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e07d6a),
	.w1(32'hb9b77e10),
	.w2(32'h3a207b01),
	.w3(32'h394b4525),
	.w4(32'h39c9e3c5),
	.w5(32'h393af36f),
	.w6(32'h398492a8),
	.w7(32'h3a466353),
	.w8(32'h39e2ac5a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a362817),
	.w1(32'h3a184ce0),
	.w2(32'h39987d77),
	.w3(32'h3a1ce9ce),
	.w4(32'h39eee598),
	.w5(32'hb91d91b5),
	.w6(32'h3a47ca80),
	.w7(32'h39e9326c),
	.w8(32'hb955eab3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba741577),
	.w1(32'hba760076),
	.w2(32'hba72bdb0),
	.w3(32'hba683a3f),
	.w4(32'hbac41b64),
	.w5(32'hb9b6232b),
	.w6(32'hba21dd8d),
	.w7(32'hbadabbb2),
	.w8(32'h37474043),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988a19f),
	.w1(32'h3801bf00),
	.w2(32'h3945be2b),
	.w3(32'hb9a830e7),
	.w4(32'hb989fd0c),
	.w5(32'h3a145587),
	.w6(32'hb91ba274),
	.w7(32'hb9561298),
	.w8(32'h3a2cbbb6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386faa03),
	.w1(32'h38996bce),
	.w2(32'h38eb6add),
	.w3(32'h3a1b6e9e),
	.w4(32'h3a1243dc),
	.w5(32'hb9805e78),
	.w6(32'h3a1ade7e),
	.w7(32'h39c64687),
	.w8(32'hb9ecbd9d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db6197),
	.w1(32'hb8995668),
	.w2(32'h395a04c7),
	.w3(32'hb8940baf),
	.w4(32'h38ec94ff),
	.w5(32'hb8bf7dd3),
	.w6(32'hb9ede3f1),
	.w7(32'h3786bbd0),
	.w8(32'hb739e27f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38905c9b),
	.w1(32'h39184e06),
	.w2(32'h39e80033),
	.w3(32'h380ccc9d),
	.w4(32'h39e5136f),
	.w5(32'hb8c0b837),
	.w6(32'hb92ef3ed),
	.w7(32'hb975e181),
	.w8(32'h38c56fbe),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76cc260),
	.w1(32'h38e2742d),
	.w2(32'h38f0cd32),
	.w3(32'h397f9a2a),
	.w4(32'hb8299981),
	.w5(32'hba3bad42),
	.w6(32'h3a65f97f),
	.w7(32'h3990b27b),
	.w8(32'hba906ec3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f60a6),
	.w1(32'hba6ef043),
	.w2(32'hb99c02aa),
	.w3(32'hbad3b4a0),
	.w4(32'hba204a5a),
	.w5(32'h3a282942),
	.w6(32'hbaae7ef5),
	.w7(32'hb99feead),
	.w8(32'h3a2064be),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e9870),
	.w1(32'h395315b0),
	.w2(32'h39e70f8c),
	.w3(32'h39a13c08),
	.w4(32'h39822b09),
	.w5(32'h39f9b35a),
	.w6(32'h39fe3286),
	.w7(32'h3a0d0df0),
	.w8(32'h3a402946),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e78cf1),
	.w1(32'h39928723),
	.w2(32'h3984ffe2),
	.w3(32'h39d708a2),
	.w4(32'h397b0577),
	.w5(32'h39b830de),
	.w6(32'h3aa61116),
	.w7(32'h3a462d8d),
	.w8(32'h39ab80cb),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4e8af),
	.w1(32'hb97b0e01),
	.w2(32'h38bd6ea2),
	.w3(32'hba05bd53),
	.w4(32'hb96da239),
	.w5(32'hba13762d),
	.w6(32'hb86570df),
	.w7(32'h39ef742c),
	.w8(32'hb9fdb088),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2aaf45),
	.w1(32'hba38800b),
	.w2(32'hba07c465),
	.w3(32'hba3d124d),
	.w4(32'hb9e52cef),
	.w5(32'h3845146d),
	.w6(32'hba5c19ff),
	.w7(32'hba01327f),
	.w8(32'h3968e54f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961a00b),
	.w1(32'h39235a5a),
	.w2(32'h3a08429f),
	.w3(32'hb88dfe0b),
	.w4(32'h3a0f0491),
	.w5(32'hb9849897),
	.w6(32'h378938be),
	.w7(32'h39c765c9),
	.w8(32'h399d453e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2654f3),
	.w1(32'h3a096cbe),
	.w2(32'h39e81f51),
	.w3(32'hb94a962c),
	.w4(32'h373075e5),
	.w5(32'h3a4ac82f),
	.w6(32'h3a0cdde4),
	.w7(32'h3a267f30),
	.w8(32'h3a6d072b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a367ca),
	.w1(32'hb8c7dc71),
	.w2(32'hb87eb807),
	.w3(32'h3a206828),
	.w4(32'h3903a196),
	.w5(32'h390a98ae),
	.w6(32'h39ac4183),
	.w7(32'hb988e237),
	.w8(32'h3929788f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a7051),
	.w1(32'h39ddb2d7),
	.w2(32'h3a02e148),
	.w3(32'h37c76b80),
	.w4(32'h39852431),
	.w5(32'hb98d2c1d),
	.w6(32'h35863d37),
	.w7(32'h39ff3442),
	.w8(32'hb9aa2e19),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bbb21),
	.w1(32'hba0b6370),
	.w2(32'h38b1757a),
	.w3(32'hb9e2e4c3),
	.w4(32'hb8d3e954),
	.w5(32'hba290b02),
	.w6(32'hb99dfa58),
	.w7(32'hb96a2370),
	.w8(32'hba61f5fb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ab9ee),
	.w1(32'hba48a35b),
	.w2(32'h3853a2ee),
	.w3(32'hb99c1959),
	.w4(32'h3a380ae1),
	.w5(32'h38c7f610),
	.w6(32'hbaeab3c8),
	.w7(32'hb9fdbd01),
	.w8(32'hb88fc18c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392cb1e5),
	.w1(32'hb9ab4779),
	.w2(32'h395fd1c9),
	.w3(32'hb9392188),
	.w4(32'h39046968),
	.w5(32'h39976374),
	.w6(32'hb9aba77c),
	.w7(32'h39976208),
	.w8(32'h39734181),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca2751),
	.w1(32'h3a88bdaa),
	.w2(32'h398cd5c6),
	.w3(32'h3a4a5656),
	.w4(32'h39eed131),
	.w5(32'h3a01fe95),
	.w6(32'h3a81834c),
	.w7(32'h3a05bfca),
	.w8(32'h3a86b58b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a334f3e),
	.w1(32'h3a12e41c),
	.w2(32'h3a100d0e),
	.w3(32'h3a25d5ef),
	.w4(32'h3a0eb6d2),
	.w5(32'hba92f5f3),
	.w6(32'h3a846315),
	.w7(32'h3a75025f),
	.w8(32'hba96c00f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4c286),
	.w1(32'hba7811a4),
	.w2(32'hb8615bea),
	.w3(32'hba3d7198),
	.w4(32'h38cf4dce),
	.w5(32'h39a06b8b),
	.w6(32'hba62a24f),
	.w7(32'h3993ba3f),
	.w8(32'h39ff2765),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b17a58),
	.w1(32'h3a023bdd),
	.w2(32'h39a8ec25),
	.w3(32'h3a22d92e),
	.w4(32'h39d30c1c),
	.w5(32'h398fdd4c),
	.w6(32'h398c5309),
	.w7(32'hb852e57f),
	.w8(32'h39b61fe3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a9bea),
	.w1(32'h399761b9),
	.w2(32'h39b0daa9),
	.w3(32'h3939d236),
	.w4(32'h39df9837),
	.w5(32'hb944e792),
	.w6(32'h376f91e8),
	.w7(32'h39a87d6f),
	.w8(32'hb9af95ed),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381a4a2d),
	.w1(32'h38533c35),
	.w2(32'h37dffadb),
	.w3(32'hb8ad3a98),
	.w4(32'h39056c14),
	.w5(32'h39baa34e),
	.w6(32'h39a296fa),
	.w7(32'h394e33df),
	.w8(32'h39d275a3),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984121e),
	.w1(32'h398c2470),
	.w2(32'h3844fcc2),
	.w3(32'h39cbbb8b),
	.w4(32'h392713b9),
	.w5(32'h3974de83),
	.w6(32'h39ed166d),
	.w7(32'hb990d870),
	.w8(32'h390f970a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a3b0e),
	.w1(32'hb9688ba5),
	.w2(32'hb8e11fbb),
	.w3(32'h391813bf),
	.w4(32'hb91e831d),
	.w5(32'h3927ff04),
	.w6(32'h399dacfb),
	.w7(32'hb90962f0),
	.w8(32'h39cb5e74),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd07bc),
	.w1(32'hb7a8ac0a),
	.w2(32'hb9100d3b),
	.w3(32'hb7e05bde),
	.w4(32'hb99cecb0),
	.w5(32'hb960557e),
	.w6(32'h38ad142c),
	.w7(32'hb9ba5ec0),
	.w8(32'hba17252d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe6816),
	.w1(32'hba3419bb),
	.w2(32'hb726840f),
	.w3(32'hba38272a),
	.w4(32'hb9e7e6d8),
	.w5(32'hba2faece),
	.w6(32'hba8882c4),
	.w7(32'hba102245),
	.w8(32'hba2de5fc),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8260a0),
	.w1(32'hba17ef17),
	.w2(32'hb95ea3f3),
	.w3(32'hb9c20bfc),
	.w4(32'h38cad077),
	.w5(32'h3964ddbd),
	.w6(32'hb9d1a740),
	.w7(32'h392168fa),
	.w8(32'h39aa6c42),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb6709),
	.w1(32'h38d238c1),
	.w2(32'h39542a31),
	.w3(32'h3a0381ae),
	.w4(32'h3a73e9d2),
	.w5(32'hba40ec4e),
	.w6(32'h39b6fe64),
	.w7(32'h39341d8f),
	.w8(32'hb9e22427),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5c0d3),
	.w1(32'hb9e35f8e),
	.w2(32'hba8e33ce),
	.w3(32'hba49e619),
	.w4(32'hbab3cfbd),
	.w5(32'h39f3394c),
	.w6(32'hba0d0978),
	.w7(32'hbacb628d),
	.w8(32'h39ed7b9b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983379a),
	.w1(32'hb72736dd),
	.w2(32'h384a7c80),
	.w3(32'h3a01d038),
	.w4(32'h3a112138),
	.w5(32'h3a97f35d),
	.w6(32'h39de680b),
	.w7(32'h394d26a3),
	.w8(32'h3a72478f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a564474),
	.w1(32'h3a077956),
	.w2(32'h3a6a81e0),
	.w3(32'h3a7c0393),
	.w4(32'h3a9425d4),
	.w5(32'hb8fe1ad9),
	.w6(32'h3a9c5c8c),
	.w7(32'h3ab94fa9),
	.w8(32'hb9c25b6d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ed0483),
	.w1(32'hba59a4cc),
	.w2(32'hb9e64193),
	.w3(32'hb9aa2a50),
	.w4(32'h38875ffc),
	.w5(32'hb81c544f),
	.w6(32'hba644593),
	.w7(32'hba5ec2b6),
	.w8(32'hb8f64a71),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acf60f),
	.w1(32'h396766eb),
	.w2(32'h3a06d4ef),
	.w3(32'h39343a81),
	.w4(32'h39b70b20),
	.w5(32'hb8fd362a),
	.w6(32'h399508f4),
	.w7(32'h3a16e86f),
	.w8(32'hb81f38ed),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940586c),
	.w1(32'hb85cd639),
	.w2(32'h3868f24c),
	.w3(32'h38e34919),
	.w4(32'hb7b9d924),
	.w5(32'h3a65a607),
	.w6(32'h3a18b057),
	.w7(32'h3719b803),
	.w8(32'h39b776a5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ad5e8d),
	.w1(32'h399f9f81),
	.w2(32'h39b9b1eb),
	.w3(32'h3a88bd39),
	.w4(32'h3987ffff),
	.w5(32'h3a6938fc),
	.w6(32'h3a099e1a),
	.w7(32'h39e4f320),
	.w8(32'h3aa84a55),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77db74),
	.w1(32'h39c24ac2),
	.w2(32'hb9332625),
	.w3(32'h3a1481b9),
	.w4(32'h36d998f2),
	.w5(32'h3937cd98),
	.w6(32'h39a464a5),
	.w7(32'h3690f8b1),
	.w8(32'hb8b8bed9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba265637),
	.w1(32'h36943a67),
	.w2(32'hb8262290),
	.w3(32'h3a4c4650),
	.w4(32'hb805fa90),
	.w5(32'hba5508db),
	.w6(32'hb8acb92c),
	.w7(32'hb9c59d1f),
	.w8(32'hbaab18ae),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91b695),
	.w1(32'hbaedeb81),
	.w2(32'hba69d0f5),
	.w3(32'hba555717),
	.w4(32'hba828b25),
	.w5(32'hb9f44b6e),
	.w6(32'hbaea0210),
	.w7(32'hbaa67b22),
	.w8(32'hb9b9ef8d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d3a67),
	.w1(32'hba2e6809),
	.w2(32'hba1bd641),
	.w3(32'hb9f27eba),
	.w4(32'hba35d165),
	.w5(32'hb93209ca),
	.w6(32'hb906c6d8),
	.w7(32'hb9eff394),
	.w8(32'hb971e4c2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e9fea),
	.w1(32'hb955fb3d),
	.w2(32'hb9511150),
	.w3(32'h3943f6e8),
	.w4(32'h395e0724),
	.w5(32'hb7693de4),
	.w6(32'hb53fd7f8),
	.w7(32'hb85f9a2c),
	.w8(32'h37d8b08e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3713cb68),
	.w1(32'hb981a47e),
	.w2(32'hb93e1bb5),
	.w3(32'h38762801),
	.w4(32'h3a0f49b3),
	.w5(32'h392bf4d3),
	.w6(32'hb9436b39),
	.w7(32'h39fcdd1c),
	.w8(32'h3719bd1a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dd2eb3),
	.w1(32'h39113ad6),
	.w2(32'hba173b6c),
	.w3(32'h3849881d),
	.w4(32'h38b5d68f),
	.w5(32'h396d748a),
	.w6(32'h39c882e9),
	.w7(32'h383bd703),
	.w8(32'hb6d2ce1d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1df8b0),
	.w1(32'h397092fa),
	.w2(32'h399baa5a),
	.w3(32'h38f214aa),
	.w4(32'hb79e3f5e),
	.w5(32'hbb6fa216),
	.w6(32'h39939987),
	.w7(32'hb924c5a5),
	.w8(32'hb6271e4e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd1763),
	.w1(32'h3bd1b7b0),
	.w2(32'h3c13e3e0),
	.w3(32'hbbaae0f3),
	.w4(32'h3aa82743),
	.w5(32'hbbdfbf97),
	.w6(32'hbaf40ea2),
	.w7(32'h3b845119),
	.w8(32'hbba5eb99),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99492a8),
	.w1(32'hbb58b79d),
	.w2(32'h3b8f7ad3),
	.w3(32'h3a78cee8),
	.w4(32'hb8d6bbcf),
	.w5(32'hbc48c0f6),
	.w6(32'h3a243188),
	.w7(32'h3a85f1c3),
	.w8(32'hbc03e598),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dd76a),
	.w1(32'h3c6b6687),
	.w2(32'h3c33e91d),
	.w3(32'hbc78c1d1),
	.w4(32'hbc0313e3),
	.w5(32'hbb3cf272),
	.w6(32'hb9c7635c),
	.w7(32'hbaf7ef77),
	.w8(32'hba8c0ddc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59f89c),
	.w1(32'hb924d21e),
	.w2(32'h3abfd080),
	.w3(32'h39f8480c),
	.w4(32'hbbce4d01),
	.w5(32'hbb753def),
	.w6(32'h3ad4ffb6),
	.w7(32'hbbbc4dd0),
	.w8(32'hba81b7dd),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9711ea),
	.w1(32'hbb8dde99),
	.w2(32'hbafd303d),
	.w3(32'h3b2655cc),
	.w4(32'hbb5bf269),
	.w5(32'hb9f933be),
	.w6(32'h3b24a48c),
	.w7(32'hbb5324b5),
	.w8(32'hbab3258c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfebbdb),
	.w1(32'hbb99e003),
	.w2(32'hbb9121b3),
	.w3(32'hbb056df0),
	.w4(32'hba8b5da1),
	.w5(32'hbc6348ee),
	.w6(32'h3a1acf24),
	.w7(32'h3a1ab3e8),
	.w8(32'hb8ca8ac4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47bd09),
	.w1(32'h3c57c8f5),
	.w2(32'h3c2ff248),
	.w3(32'hbc2284c5),
	.w4(32'hbc3f2300),
	.w5(32'hbb65e052),
	.w6(32'h3a9ce06a),
	.w7(32'hbabb8a80),
	.w8(32'hb88d8900),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e84595),
	.w1(32'hbb46a196),
	.w2(32'hbb271e78),
	.w3(32'h3b675db4),
	.w4(32'h3affcc71),
	.w5(32'hbbd82d91),
	.w6(32'hbad2ee29),
	.w7(32'hbaecf5f9),
	.w8(32'hbc33308b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14a650),
	.w1(32'hbc314478),
	.w2(32'h3b57976f),
	.w3(32'hbc874f08),
	.w4(32'hbc600ca4),
	.w5(32'h3bda33d5),
	.w6(32'hbc9c02c4),
	.w7(32'hbc60725d),
	.w8(32'h39b347d8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c17a6),
	.w1(32'hbc0d2fa3),
	.w2(32'hbc07937a),
	.w3(32'h3c7346c6),
	.w4(32'hba92df98),
	.w5(32'hbaf77292),
	.w6(32'h3bb9a123),
	.w7(32'h3a16f777),
	.w8(32'h3a95e5a8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c44da),
	.w1(32'h3c865df2),
	.w2(32'h3c803fa1),
	.w3(32'h39e62a8f),
	.w4(32'h3b7ab177),
	.w5(32'h3ba590e1),
	.w6(32'h3b5d5dca),
	.w7(32'h3c0e9c3c),
	.w8(32'h3b73d189),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9ec5a),
	.w1(32'hbc3807c3),
	.w2(32'hbc88cacb),
	.w3(32'h3c44c55e),
	.w4(32'h3b36db7d),
	.w5(32'hbb1743b0),
	.w6(32'h3b9a3620),
	.w7(32'h39bff252),
	.w8(32'h3b2977bb),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ab1ae),
	.w1(32'hbb620e67),
	.w2(32'hbaec9600),
	.w3(32'h3aabbef8),
	.w4(32'h3af67268),
	.w5(32'h3b703305),
	.w6(32'h3b27e177),
	.w7(32'hb949e99c),
	.w8(32'hbac93745),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc85f6d),
	.w1(32'hbbb4ebd8),
	.w2(32'h3bf68ed6),
	.w3(32'h3bc22c94),
	.w4(32'h3ab183fa),
	.w5(32'h3baac308),
	.w6(32'hb8f19275),
	.w7(32'hb8bcfef5),
	.w8(32'h3af33e6a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87dba5),
	.w1(32'hbb6acb70),
	.w2(32'hbc27d3f1),
	.w3(32'h3c2fdb88),
	.w4(32'hbb24ab6a),
	.w5(32'hbaa6347c),
	.w6(32'hbb488657),
	.w7(32'hbc4f6116),
	.w8(32'hbab4ba4c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55ebb7),
	.w1(32'h3a8dc8ad),
	.w2(32'h3a65fdd3),
	.w3(32'hba05f964),
	.w4(32'h39b876af),
	.w5(32'h3bb408e8),
	.w6(32'h3bd663d4),
	.w7(32'h3b872f7c),
	.w8(32'hbbbe28de),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e990f),
	.w1(32'hbc073b87),
	.w2(32'h3b83ec75),
	.w3(32'hbc36cf6d),
	.w4(32'hbaf0f8e6),
	.w5(32'h3b2072ca),
	.w6(32'hbac3e3f2),
	.w7(32'hba69bf14),
	.w8(32'h3af52e8f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf7808),
	.w1(32'hbba391cf),
	.w2(32'h3b90863b),
	.w3(32'h3b386901),
	.w4(32'h3ace5108),
	.w5(32'h390dc634),
	.w6(32'h3b3bc5e1),
	.w7(32'hbbb34712),
	.w8(32'h3bac5b14),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ebd75),
	.w1(32'h3c6194ea),
	.w2(32'h3c1e8e6d),
	.w3(32'hbb3de1c6),
	.w4(32'h3ac681d0),
	.w5(32'hbc06b976),
	.w6(32'h3c2f52ad),
	.w7(32'h3c19ecad),
	.w8(32'hbb69fdf4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12774b),
	.w1(32'h3c688c34),
	.w2(32'h3bb01193),
	.w3(32'hbb801226),
	.w4(32'hbbce4129),
	.w5(32'hbc0f93eb),
	.w6(32'hbbf61728),
	.w7(32'hba81bc45),
	.w8(32'hbb6137c8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e7d77),
	.w1(32'h3986ebeb),
	.w2(32'hbabb56ff),
	.w3(32'hbc044bb8),
	.w4(32'hbbe1b1d2),
	.w5(32'hbc26c0a6),
	.w6(32'h3923bc57),
	.w7(32'hbad62b37),
	.w8(32'hbc07ea72),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc23120),
	.w1(32'h3ab4e5a5),
	.w2(32'h3ba8111b),
	.w3(32'hbc6007f6),
	.w4(32'hbbd70048),
	.w5(32'hbaf6306e),
	.w6(32'hbc6bc674),
	.w7(32'hbb85e502),
	.w8(32'h39edb89b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ad1ca),
	.w1(32'hb9fde57c),
	.w2(32'hbb101631),
	.w3(32'h392de071),
	.w4(32'h3b1e7773),
	.w5(32'h3a8146f5),
	.w6(32'h3c0a9708),
	.w7(32'hbb6bc1ca),
	.w8(32'h3b3e6dd5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9679f9),
	.w1(32'hbc13dd37),
	.w2(32'hbc25f740),
	.w3(32'h3c383ae2),
	.w4(32'h3922fdb4),
	.w5(32'h3b9f39cb),
	.w6(32'h3acfddb8),
	.w7(32'hbbf9dab6),
	.w8(32'h3b805c2a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe06a3a),
	.w1(32'hbc2d727e),
	.w2(32'h3846ab77),
	.w3(32'h3c2c9ddb),
	.w4(32'h3b851f2f),
	.w5(32'h3bcde036),
	.w6(32'hbb4dc6d5),
	.w7(32'hbc0bc20b),
	.w8(32'hbb6bc3ff),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87eb6b),
	.w1(32'hbbbc0786),
	.w2(32'hbc394a58),
	.w3(32'h3c8144ed),
	.w4(32'hb9171856),
	.w5(32'h3b6914e0),
	.w6(32'h3a872a51),
	.w7(32'hbb7f4886),
	.w8(32'h3bd00088),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb974c5a),
	.w1(32'hbc42d7db),
	.w2(32'hbb839413),
	.w3(32'h3a020c9e),
	.w4(32'h3c117854),
	.w5(32'hbb50db33),
	.w6(32'h3bc28f1e),
	.w7(32'h3a2342b2),
	.w8(32'hbb1013b2),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b39dc),
	.w1(32'hbb6408b9),
	.w2(32'hba69556b),
	.w3(32'h3b685b83),
	.w4(32'hbb8531c8),
	.w5(32'h3bf50ceb),
	.w6(32'h3b76531e),
	.w7(32'h3bd91735),
	.w8(32'h3bcf2f27),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b7b85),
	.w1(32'h3b5ec8d0),
	.w2(32'hbbf4098e),
	.w3(32'h3c49f0ac),
	.w4(32'h3ae2b477),
	.w5(32'hba154eaa),
	.w6(32'h3bc8cfbc),
	.w7(32'h3a310a9a),
	.w8(32'hbb629b57),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef16d8),
	.w1(32'hbb91a60e),
	.w2(32'h3c298ee4),
	.w3(32'hbba6565b),
	.w4(32'hbbae6801),
	.w5(32'h3c37c1c9),
	.w6(32'hbbb3cef5),
	.w7(32'h3c2a3229),
	.w8(32'h3bde441c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc182f60),
	.w1(32'hbcb263d7),
	.w2(32'hbccb31ae),
	.w3(32'h3cc62d6b),
	.w4(32'h3be4798a),
	.w5(32'h3ba01b91),
	.w6(32'h3816d8a1),
	.w7(32'hbc04eb39),
	.w8(32'hbb84cc18),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93ae5e),
	.w1(32'h3a9aec23),
	.w2(32'h3a9a5ace),
	.w3(32'h3c101731),
	.w4(32'hbbfad47e),
	.w5(32'hbb9f79ba),
	.w6(32'h395b4f5f),
	.w7(32'hbb580fb0),
	.w8(32'hbac6255e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb069eaa),
	.w1(32'hbbcd6840),
	.w2(32'hbb904e32),
	.w3(32'hbc54ddf3),
	.w4(32'hbb020969),
	.w5(32'hbbaab12f),
	.w6(32'h3c069e12),
	.w7(32'hbbab1462),
	.w8(32'hbb21adb4),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60e397),
	.w1(32'h3bcf5abe),
	.w2(32'h3bb84684),
	.w3(32'hbb948012),
	.w4(32'hb84b894e),
	.w5(32'hbac64e7d),
	.w6(32'h3b4736c9),
	.w7(32'h3b22e46e),
	.w8(32'hbbed8ae7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8c23c),
	.w1(32'h3a2b3192),
	.w2(32'hbb98eeaa),
	.w3(32'h3bcb0f00),
	.w4(32'hbba72e35),
	.w5(32'h3a665cd9),
	.w6(32'hbc08bce7),
	.w7(32'hbbe88e5f),
	.w8(32'h3b605f46),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6b7ad),
	.w1(32'h3919289e),
	.w2(32'hbb517553),
	.w3(32'h3b8bd7a3),
	.w4(32'hba387e55),
	.w5(32'hbb3ab8e2),
	.w6(32'h3c0b6f8d),
	.w7(32'h3b85ef67),
	.w8(32'hb751e894),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4989c8),
	.w1(32'h3c00b900),
	.w2(32'h3b61cfb5),
	.w3(32'hbbc24754),
	.w4(32'hbb6c865e),
	.w5(32'hbb5c6021),
	.w6(32'h3b513f47),
	.w7(32'h3be86053),
	.w8(32'h3b393487),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca719a),
	.w1(32'h391ae4b3),
	.w2(32'hbb22e4c1),
	.w3(32'hba0617a0),
	.w4(32'h3b109985),
	.w5(32'h3b8742af),
	.w6(32'h3c411e4d),
	.w7(32'h3b285d82),
	.w8(32'hbb0eb814),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba887f71),
	.w1(32'hba918b19),
	.w2(32'hbb90aeaf),
	.w3(32'h3b9a4148),
	.w4(32'hba19d73d),
	.w5(32'h3abb9ca2),
	.w6(32'h3add7c1a),
	.w7(32'hbb2fcd18),
	.w8(32'h3af27e08),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928b394),
	.w1(32'hbabf9d62),
	.w2(32'hbba540fe),
	.w3(32'h3ae2f1d3),
	.w4(32'hbb85bc81),
	.w5(32'h3a172c84),
	.w6(32'h3b714279),
	.w7(32'h3a4d3c9a),
	.w8(32'h3a188f89),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bdde3),
	.w1(32'h3919189d),
	.w2(32'hbac1f75e),
	.w3(32'h3acb4cd9),
	.w4(32'h3a68f516),
	.w5(32'h3b654bcd),
	.w6(32'h3bdb247d),
	.w7(32'h3b9a1236),
	.w8(32'hbbffc2cf),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc3bec),
	.w1(32'h3ab41b59),
	.w2(32'hbacd0dae),
	.w3(32'hbc26618f),
	.w4(32'h3b3d98bc),
	.w5(32'h3bb49b00),
	.w6(32'h3bb2ae71),
	.w7(32'hbb913740),
	.w8(32'hbb04f3bd),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb863e6f),
	.w1(32'hbc713435),
	.w2(32'hbc5bbea8),
	.w3(32'h3c5f1551),
	.w4(32'hbaaecc66),
	.w5(32'h3a6dca74),
	.w6(32'hbc219284),
	.w7(32'hbc7ce063),
	.w8(32'hba7f2d75),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a969a0f),
	.w1(32'hbbf2efc2),
	.w2(32'hb930a0e6),
	.w3(32'h3c0a961b),
	.w4(32'h3ab2b57b),
	.w5(32'hbb239475),
	.w6(32'hbbd11772),
	.w7(32'h3aeb76d6),
	.w8(32'h3ada7781),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa406c),
	.w1(32'hbae5c93b),
	.w2(32'hbb31945f),
	.w3(32'hbb5c9fb8),
	.w4(32'hbafae273),
	.w5(32'hb9cf0b3d),
	.w6(32'h3b4c679e),
	.w7(32'hbaab3ca4),
	.w8(32'h3a5c08d1),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80d00e),
	.w1(32'hbc003ce5),
	.w2(32'hbc12c65a),
	.w3(32'h3c5830b0),
	.w4(32'hbb20770e),
	.w5(32'h3c737e06),
	.w6(32'hbc48a4b3),
	.w7(32'hbc259f3a),
	.w8(32'h3b399a26),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f21625),
	.w1(32'hba979cdc),
	.w2(32'hbbc4eae1),
	.w3(32'h3cae427a),
	.w4(32'h3b8546e8),
	.w5(32'hbad6bf6b),
	.w6(32'h3c40adc4),
	.w7(32'h3a4753ff),
	.w8(32'hbb131c3a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377457db),
	.w1(32'hbb2b6e15),
	.w2(32'hbb7b047a),
	.w3(32'h3a4988cc),
	.w4(32'h3abf7010),
	.w5(32'hbbe1eda7),
	.w6(32'hbaf74c74),
	.w7(32'hba06d7ce),
	.w8(32'hbb3c1159),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4dc10a),
	.w1(32'h3bb23df5),
	.w2(32'hba4c8eae),
	.w3(32'hbb945d2d),
	.w4(32'hba11888e),
	.w5(32'hba9c30a9),
	.w6(32'h3b31a7e3),
	.w7(32'h3bc42db1),
	.w8(32'h3a880e41),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b920a4c),
	.w1(32'hbada3255),
	.w2(32'hbaca1009),
	.w3(32'h3bf1975c),
	.w4(32'hb98f85de),
	.w5(32'h3b638a17),
	.w6(32'hb9178626),
	.w7(32'h3a1ab32e),
	.w8(32'hba23200e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39653b9b),
	.w1(32'hbbdb48b9),
	.w2(32'hbc8c6eea),
	.w3(32'h3c9cb448),
	.w4(32'h3bc7215d),
	.w5(32'h3ac52a9d),
	.w6(32'hbc25547d),
	.w7(32'hbc27b91c),
	.w8(32'h3bf1d247),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3188cd),
	.w1(32'h3c79591c),
	.w2(32'h3c4696dd),
	.w3(32'h38d229c2),
	.w4(32'h3b133475),
	.w5(32'hbab31aa3),
	.w6(32'h3c542d2e),
	.w7(32'h3c099d14),
	.w8(32'h3b22febf),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e1ba7),
	.w1(32'hbba945f2),
	.w2(32'hbbe06c2f),
	.w3(32'hbb02d3b4),
	.w4(32'hbb78c49e),
	.w5(32'h3c179e81),
	.w6(32'h3b26a877),
	.w7(32'hbbe13ce1),
	.w8(32'h3b3964d5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8908f1),
	.w1(32'hbc9f55c6),
	.w2(32'hbc150594),
	.w3(32'h3c87830e),
	.w4(32'hbb11a8ec),
	.w5(32'h3a5c9116),
	.w6(32'hbc9058da),
	.w7(32'hbba43493),
	.w8(32'hba2ab2b3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dbfb4),
	.w1(32'h3b692a69),
	.w2(32'h3b6b0aec),
	.w3(32'hbbbff567),
	.w4(32'hb95afa2f),
	.w5(32'hbbd03e58),
	.w6(32'h396e9259),
	.w7(32'hbac2c1af),
	.w8(32'hb9e10e99),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd326fb),
	.w1(32'h3ae0e521),
	.w2(32'hbbf0c6ac),
	.w3(32'h3abaa71a),
	.w4(32'hbb5fd146),
	.w5(32'hbc1a0923),
	.w6(32'h3bd18683),
	.w7(32'h3ab1e022),
	.w8(32'hbb4aec5e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d3c10),
	.w1(32'h3c6eb6d9),
	.w2(32'h3c5ce4fa),
	.w3(32'hbc106443),
	.w4(32'h39aef433),
	.w5(32'h3bf40f01),
	.w6(32'h3bd1013e),
	.w7(32'h3be764a2),
	.w8(32'h3b69fd4a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6dfb8),
	.w1(32'hbc336cfc),
	.w2(32'hbc890701),
	.w3(32'h3c75ff04),
	.w4(32'h3afb9753),
	.w5(32'h3a436ff1),
	.w6(32'hba9669c6),
	.w7(32'hbb5b2389),
	.w8(32'h3b67369b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b9f19),
	.w1(32'hbaf33226),
	.w2(32'hbba57d9c),
	.w3(32'h3b2d673b),
	.w4(32'hbbadbcb3),
	.w5(32'h3bdce867),
	.w6(32'hbb010e47),
	.w7(32'h3aa2323f),
	.w8(32'h3af04b5b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c9911),
	.w1(32'hbb86aad3),
	.w2(32'hbb82e127),
	.w3(32'h3c59c344),
	.w4(32'h39d39d36),
	.w5(32'hbb543a87),
	.w6(32'hbb7ac4fc),
	.w7(32'hbbe79db4),
	.w8(32'hbbf2bd24),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d119b),
	.w1(32'h3b4e368b),
	.w2(32'h3a8d42cb),
	.w3(32'hbbcbd213),
	.w4(32'hbb775b47),
	.w5(32'h3b908f87),
	.w6(32'hbc3f6462),
	.w7(32'hbaa1fc38),
	.w8(32'hbb6c3fbe),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde1a68),
	.w1(32'hbbf4851a),
	.w2(32'h3ad0e5fa),
	.w3(32'hbbac786b),
	.w4(32'h39f8c0db),
	.w5(32'hbb22ba8f),
	.w6(32'h38871a17),
	.w7(32'hbc62b430),
	.w8(32'hbc085817),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b0770),
	.w1(32'h3b65dd7b),
	.w2(32'h3c4b8f91),
	.w3(32'hbacab132),
	.w4(32'hbbae762e),
	.w5(32'hbb1d0296),
	.w6(32'hbbad2b03),
	.w7(32'h3bf1f9eb),
	.w8(32'hba87784e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b0940),
	.w1(32'hbb7fdd50),
	.w2(32'hbc0531f7),
	.w3(32'h3bb5bd1f),
	.w4(32'hbb9abb41),
	.w5(32'h3ab04869),
	.w6(32'hbbadf5d6),
	.w7(32'hbbd847e4),
	.w8(32'h3acd50df),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3c7d5),
	.w1(32'hbb3a402c),
	.w2(32'hbb4c790c),
	.w3(32'h3b60678d),
	.w4(32'h3b6e1144),
	.w5(32'hbb62ebc5),
	.w6(32'hbaaa7612),
	.w7(32'hb9f1f4a1),
	.w8(32'h3b90a07e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b682542),
	.w1(32'hbb814e93),
	.w2(32'hbbade89e),
	.w3(32'h3bb86e45),
	.w4(32'h3a8a70fe),
	.w5(32'hbb87cd30),
	.w6(32'h3b50ab0d),
	.w7(32'h3a6b4d2f),
	.w8(32'hba60a2f5),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b8612),
	.w1(32'h3c4b4b3c),
	.w2(32'h3aea7dde),
	.w3(32'hba2bcfba),
	.w4(32'hba5880c3),
	.w5(32'hbb918688),
	.w6(32'hbbe71dcf),
	.w7(32'hbba02a57),
	.w8(32'hbba68fe1),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd94cd),
	.w1(32'h3bac7d79),
	.w2(32'h3bf952ee),
	.w3(32'hbc81a449),
	.w4(32'hbbab9a1b),
	.w5(32'h3bb666b1),
	.w6(32'hbb9c1374),
	.w7(32'h3b948cb1),
	.w8(32'hbba49a48),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d949d5),
	.w1(32'hbaeeca50),
	.w2(32'hbb90f2be),
	.w3(32'h3c3cd7ec),
	.w4(32'h3b3dac86),
	.w5(32'h3ba3d26f),
	.w6(32'hbbaef38f),
	.w7(32'hba18e387),
	.w8(32'h3c09e692),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2eb0b7),
	.w1(32'h3c03323c),
	.w2(32'h3bf9a5e3),
	.w3(32'h3b941726),
	.w4(32'h3a4c10d6),
	.w5(32'h38843828),
	.w6(32'h3ba1b705),
	.w7(32'h3b6c8f20),
	.w8(32'h3a114ecf),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5446ad),
	.w1(32'h3a53d075),
	.w2(32'h3a886b85),
	.w3(32'hb87ddb3a),
	.w4(32'h3aaca2cd),
	.w5(32'hbb32a69e),
	.w6(32'h3bbdfc53),
	.w7(32'hba8ac535),
	.w8(32'hbb916f08),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5725e),
	.w1(32'h3c0db396),
	.w2(32'hbb34d1fa),
	.w3(32'hbaf73cd3),
	.w4(32'hbb68fac2),
	.w5(32'hbb4f51a7),
	.w6(32'h3b0b9db2),
	.w7(32'hbb9da859),
	.w8(32'hbc0fedce),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adebcf2),
	.w1(32'h3b80e1da),
	.w2(32'h3ada203f),
	.w3(32'hbbaae173),
	.w4(32'hbaf18876),
	.w5(32'hbb1925da),
	.w6(32'hbbbbd0f2),
	.w7(32'hba471383),
	.w8(32'hbc0cffb7),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a0251),
	.w1(32'h3bafe774),
	.w2(32'h3b2bc340),
	.w3(32'hbb71b4c5),
	.w4(32'hbb589635),
	.w5(32'hbc3dd14c),
	.w6(32'h3b86804c),
	.w7(32'hb9d402d5),
	.w8(32'hbbc0c67c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4df1a),
	.w1(32'h3bee8334),
	.w2(32'h3b8f8865),
	.w3(32'hbc531f58),
	.w4(32'hbc1d1b8d),
	.w5(32'hba617a37),
	.w6(32'hbb749477),
	.w7(32'hbb59868c),
	.w8(32'h3a784814),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8c7e6),
	.w1(32'hbc500691),
	.w2(32'hbc5c1fa8),
	.w3(32'h3b970228),
	.w4(32'h3aac04ab),
	.w5(32'hbc0c1945),
	.w6(32'h3ab417cd),
	.w7(32'h3b02f1ea),
	.w8(32'hbb80e148),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba267f1d),
	.w1(32'h3a0137fc),
	.w2(32'h38eeed7a),
	.w3(32'hbc08d55e),
	.w4(32'hbbf7aeae),
	.w5(32'h3c4ff172),
	.w6(32'hbb2cb434),
	.w7(32'hbb5727ef),
	.w8(32'h3b92910c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b539cbf),
	.w1(32'h3a91a371),
	.w2(32'hbb82fb89),
	.w3(32'h3c0f44df),
	.w4(32'h3b1d6fbe),
	.w5(32'hbac91e18),
	.w6(32'h3b308bf5),
	.w7(32'hbb407161),
	.w8(32'hbb8e9da6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0a1a1),
	.w1(32'hbc845c95),
	.w2(32'hbc4db81e),
	.w3(32'h3b9a6af7),
	.w4(32'hbb4db9f3),
	.w5(32'hbace0d24),
	.w6(32'hbc5d65ad),
	.w7(32'hbc529ac4),
	.w8(32'h3bca160d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f64c6),
	.w1(32'h3c4695a9),
	.w2(32'h3bec3faa),
	.w3(32'hbb0715f4),
	.w4(32'hba9f87b6),
	.w5(32'h39075617),
	.w6(32'h3c120b61),
	.w7(32'h3b2fd5df),
	.w8(32'hbbd457ba),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadbc18),
	.w1(32'hbb470a66),
	.w2(32'h3b8daeed),
	.w3(32'hbb135792),
	.w4(32'hbacf0b40),
	.w5(32'hbb4b7057),
	.w6(32'hbb0dbb57),
	.w7(32'hb9266760),
	.w8(32'hbb7f08da),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba98636),
	.w1(32'h3aa526bd),
	.w2(32'hbad09662),
	.w3(32'hbbdd63b6),
	.w4(32'hbb0e86bc),
	.w5(32'hb991c90e),
	.w6(32'hba5655e1),
	.w7(32'hbb73a623),
	.w8(32'hbb7f5b4b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef5265),
	.w1(32'hbbd030f4),
	.w2(32'hba827f85),
	.w3(32'h3b755bdb),
	.w4(32'h3b9c7ae0),
	.w5(32'hbb8aac24),
	.w6(32'h3b03fbf6),
	.w7(32'hbb1cc745),
	.w8(32'h3bb8cfee),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4a6f9),
	.w1(32'h3c33f05c),
	.w2(32'hbc0e3f24),
	.w3(32'h3b9d77af),
	.w4(32'h3b927317),
	.w5(32'h3ab3b7ee),
	.w6(32'h3aee46b1),
	.w7(32'hbbcb4b16),
	.w8(32'h3b807ae2),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc73cbb),
	.w1(32'h39239a14),
	.w2(32'hba87559f),
	.w3(32'h3b3b6de8),
	.w4(32'h39ab1f77),
	.w5(32'h3bb97c62),
	.w6(32'hbb11d294),
	.w7(32'hba3df844),
	.w8(32'hba8bb4f2),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee0667),
	.w1(32'hbba81b42),
	.w2(32'hbb601463),
	.w3(32'h3abff4b1),
	.w4(32'h39ded1f6),
	.w5(32'h3ab34222),
	.w6(32'hbb310f98),
	.w7(32'h3b439b43),
	.w8(32'h39cb2698),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b628da4),
	.w1(32'hb9819881),
	.w2(32'h3a3ccbe1),
	.w3(32'hbb31eb51),
	.w4(32'hbb0a8734),
	.w5(32'hbb5314f3),
	.w6(32'h3b0c984f),
	.w7(32'h381738a4),
	.w8(32'h3b2cb0a5),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc5f45),
	.w1(32'hbb4a8adf),
	.w2(32'h3b33bdc8),
	.w3(32'h3bac2888),
	.w4(32'hba982e2e),
	.w5(32'hbbc3c518),
	.w6(32'hbc12efd4),
	.w7(32'hbba813af),
	.w8(32'h3a437c89),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b1e82),
	.w1(32'h3c10b4b2),
	.w2(32'h3ae9478e),
	.w3(32'hbbe00646),
	.w4(32'hbb72ade3),
	.w5(32'h3aeea223),
	.w6(32'h3bde1bac),
	.w7(32'h3b25bfab),
	.w8(32'h39b629ec),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22fb29),
	.w1(32'h3c758894),
	.w2(32'h3c75e381),
	.w3(32'hbc9df06c),
	.w4(32'h3c153600),
	.w5(32'h3a9fc068),
	.w6(32'h3c0472f3),
	.w7(32'h3ccb56de),
	.w8(32'h3b2d3dac),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb962e38),
	.w1(32'hbaaa36f7),
	.w2(32'hbb100982),
	.w3(32'h3bf26ec0),
	.w4(32'h3b9ec077),
	.w5(32'h3bb6450d),
	.w6(32'hbb03d9f8),
	.w7(32'h3ac157be),
	.w8(32'h3bd6edcc),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8ac50),
	.w1(32'hbb92827d),
	.w2(32'hbc26ba16),
	.w3(32'h3c7841bb),
	.w4(32'h3b234527),
	.w5(32'hbaea9c39),
	.w6(32'h3c0af7b7),
	.w7(32'hb9d6a07e),
	.w8(32'h39a2d547),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e3cc5),
	.w1(32'h3b36d594),
	.w2(32'h3ae7fe40),
	.w3(32'h3b323bfb),
	.w4(32'h3b015a47),
	.w5(32'hbb5589e3),
	.w6(32'hb9b33469),
	.w7(32'h3a83865c),
	.w8(32'h391e3fe2),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f17e2),
	.w1(32'hbba1a825),
	.w2(32'hbbc65c00),
	.w3(32'hba023703),
	.w4(32'hb99d02c4),
	.w5(32'h3b01e695),
	.w6(32'hbbb231c0),
	.w7(32'hbb2473ee),
	.w8(32'hbb568966),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace0600),
	.w1(32'hbb7750e6),
	.w2(32'hbb371101),
	.w3(32'h3c38475b),
	.w4(32'h3bb49ff2),
	.w5(32'h391f283d),
	.w6(32'hbb53570e),
	.w7(32'h3aa28312),
	.w8(32'hba322169),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeaae4a),
	.w1(32'h3b363d71),
	.w2(32'h3b8607fc),
	.w3(32'hbb091b5a),
	.w4(32'hb9d00a04),
	.w5(32'hbac2be29),
	.w6(32'h396cb9cd),
	.w7(32'hb9916857),
	.w8(32'h3bd12918),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ade4a),
	.w1(32'hbc1fd19e),
	.w2(32'hbc4b6c6e),
	.w3(32'h3b839e69),
	.w4(32'h3bc334c4),
	.w5(32'h3beb670d),
	.w6(32'h3c4f3c37),
	.w7(32'hbb6bc885),
	.w8(32'hbbaecadf),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb015c7),
	.w1(32'hbc0e7676),
	.w2(32'hbbb90efa),
	.w3(32'h3bd7e08c),
	.w4(32'hb971c1e4),
	.w5(32'h3a2cfe31),
	.w6(32'hbc429c77),
	.w7(32'hbc09387a),
	.w8(32'h393b68a8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8ac24),
	.w1(32'hbc242617),
	.w2(32'h3bc3c555),
	.w3(32'h3c08d3b6),
	.w4(32'hba2bb6a5),
	.w5(32'h39fd0a03),
	.w6(32'hbb6caa47),
	.w7(32'h3bad70dc),
	.w8(32'h3b84cc5e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1389d9),
	.w1(32'h3c13908f),
	.w2(32'h3c149047),
	.w3(32'hbb435e58),
	.w4(32'h3b426883),
	.w5(32'hbc0755fc),
	.w6(32'h3beec029),
	.w7(32'h3b3bdd5c),
	.w8(32'hbbbb6bc4),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d3fa7),
	.w1(32'h3c0f364e),
	.w2(32'h3bd6d276),
	.w3(32'hbbae2d08),
	.w4(32'hb9a4a359),
	.w5(32'h3be595b4),
	.w6(32'hbade80dd),
	.w7(32'h3b38eebf),
	.w8(32'h3b4db23c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae73df7),
	.w1(32'hbc828a6d),
	.w2(32'hbc35e8e1),
	.w3(32'h3c7ae82c),
	.w4(32'hba9318ec),
	.w5(32'h3c2db361),
	.w6(32'hbba2680d),
	.w7(32'hbc06ce6b),
	.w8(32'hbb1e37d8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd79db5),
	.w1(32'hbc5e7202),
	.w2(32'hbc07bef3),
	.w3(32'h3c10d6f3),
	.w4(32'h3bad8554),
	.w5(32'hbb94d7de),
	.w6(32'h3ab811f1),
	.w7(32'h3a6f5893),
	.w8(32'hbb3f855a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05cd26),
	.w1(32'h3bb8f7ca),
	.w2(32'hbc014f51),
	.w3(32'h3beba294),
	.w4(32'hbab349fa),
	.w5(32'h3b8fed6a),
	.w6(32'hbb31a5bd),
	.w7(32'hbc05d69a),
	.w8(32'h3b290169),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd02479),
	.w1(32'hbc3ff4a3),
	.w2(32'hbc288932),
	.w3(32'h3c443d3d),
	.w4(32'h3bfd413c),
	.w5(32'h3c556ec6),
	.w6(32'h3bc567db),
	.w7(32'hbad42441),
	.w8(32'h3b7b989e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b085863),
	.w1(32'hbc35dfa9),
	.w2(32'hbc5372ad),
	.w3(32'h3c416f4d),
	.w4(32'h3c069da7),
	.w5(32'hbb8245fc),
	.w6(32'hbab4e819),
	.w7(32'hbb451f4c),
	.w8(32'hbb15f542),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5842e6),
	.w1(32'hbb00abb8),
	.w2(32'h3b045059),
	.w3(32'hbb2a1bd9),
	.w4(32'hba3893ec),
	.w5(32'h39dd74db),
	.w6(32'h3b771713),
	.w7(32'h3ac2287e),
	.w8(32'hbac80250),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44d2fc),
	.w1(32'h3b0add73),
	.w2(32'h3b06f13e),
	.w3(32'hbb909bbe),
	.w4(32'hbb4bcb57),
	.w5(32'hbba2cbe6),
	.w6(32'hbaa21de0),
	.w7(32'hbbb2abb9),
	.w8(32'h3b50aedf),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7d824),
	.w1(32'hbc51bcac),
	.w2(32'hbbc35770),
	.w3(32'h3bbc7c35),
	.w4(32'h3b78c61d),
	.w5(32'h3bc6ab80),
	.w6(32'h3ae6ad5b),
	.w7(32'hbb8f28f8),
	.w8(32'h3bd914d0),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48f180),
	.w1(32'hbb823fc2),
	.w2(32'hbc08c5cd),
	.w3(32'h3c8496b4),
	.w4(32'hba1b668a),
	.w5(32'hbb031a19),
	.w6(32'h3bddb1a6),
	.w7(32'hbb7cd126),
	.w8(32'h3aec15d2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37ff1f),
	.w1(32'h3b2905f8),
	.w2(32'hba1a5f18),
	.w3(32'hbad7018d),
	.w4(32'hba1dff5a),
	.w5(32'hbb6eb8c4),
	.w6(32'h3b3e1fa8),
	.w7(32'hbb3642b3),
	.w8(32'hb9fa1fa4),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8874e8),
	.w1(32'hbb9adfb9),
	.w2(32'hbb9d4efd),
	.w3(32'h3a9cb75e),
	.w4(32'h3ae1e9d3),
	.w5(32'hbb5f22e3),
	.w6(32'hbb876002),
	.w7(32'hbacd24fb),
	.w8(32'h39c5516d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae237b),
	.w1(32'hbbf80682),
	.w2(32'hba137af3),
	.w3(32'h3b5bb1ee),
	.w4(32'hbb3374b2),
	.w5(32'h3b230832),
	.w6(32'h3b866d87),
	.w7(32'hbbae032f),
	.w8(32'h3b290900),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0763f2),
	.w1(32'h39fe455c),
	.w2(32'h3b14cb68),
	.w3(32'h3b9f8995),
	.w4(32'h3b847ff0),
	.w5(32'hbb72044e),
	.w6(32'h3bd26683),
	.w7(32'h3bdd82c1),
	.w8(32'h3c011d3f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42f8d0),
	.w1(32'hbaa33537),
	.w2(32'hbb09abe2),
	.w3(32'hba89c0a5),
	.w4(32'hbb65c627),
	.w5(32'h3c0c10b5),
	.w6(32'h3c4aa607),
	.w7(32'h3a7a6ccd),
	.w8(32'h3b969669),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb999992),
	.w1(32'hbc0e0341),
	.w2(32'hbc368646),
	.w3(32'h3c8281ae),
	.w4(32'h3c88c155),
	.w5(32'hbb967b5d),
	.w6(32'h3c30edd4),
	.w7(32'h3c0905e7),
	.w8(32'hbab903e3),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2f7e6),
	.w1(32'h3b304528),
	.w2(32'hb9ce286b),
	.w3(32'hbc2b3332),
	.w4(32'hb9811faa),
	.w5(32'h392bacfb),
	.w6(32'hbb651401),
	.w7(32'h35aa001e),
	.w8(32'hbb3782b5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803706),
	.w1(32'hb9ba248b),
	.w2(32'hbb67aa2f),
	.w3(32'h3b6f3f8b),
	.w4(32'hb95a9560),
	.w5(32'hbb12011b),
	.w6(32'hbb567a1a),
	.w7(32'hbb4a4fd8),
	.w8(32'h3a29afc8),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a824ac2),
	.w1(32'h3bc6fbf7),
	.w2(32'h3a1ba69c),
	.w3(32'h3a7fb377),
	.w4(32'hbbd9f7f7),
	.w5(32'h3c0080e0),
	.w6(32'h3bee70ca),
	.w7(32'hb80f78a9),
	.w8(32'hba473414),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5da4a4),
	.w1(32'hbc90528a),
	.w2(32'hbc1fddb3),
	.w3(32'h3c93fc3e),
	.w4(32'hbb712fee),
	.w5(32'hba8e7b9f),
	.w6(32'hbaa7ca35),
	.w7(32'hbbd071e6),
	.w8(32'h3a9000cd),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e84ae8),
	.w1(32'hbc8a5691),
	.w2(32'hbc3dbf15),
	.w3(32'h3c51dc5d),
	.w4(32'h3a12a387),
	.w5(32'h3b2d76a2),
	.w6(32'hbc0951e2),
	.w7(32'hbbdad833),
	.w8(32'hbbdae97a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf795b8),
	.w1(32'h3a0d3051),
	.w2(32'h3b3b4dcf),
	.w3(32'h3b7a1ecd),
	.w4(32'h3b4aee44),
	.w5(32'hbbdb6204),
	.w6(32'hbb44faf6),
	.w7(32'h3b55d98b),
	.w8(32'hbbeda359),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba99d05),
	.w1(32'hbac4d3c9),
	.w2(32'h3c36b19c),
	.w3(32'hbbc14c73),
	.w4(32'hbb3e77cb),
	.w5(32'hbbb1fec7),
	.w6(32'hbc26dac3),
	.w7(32'hbae98323),
	.w8(32'h39db24bf),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8122124),
	.w1(32'hbaa97199),
	.w2(32'h3985cb73),
	.w3(32'hbb5cf121),
	.w4(32'hbb76f3ab),
	.w5(32'h3bc5498b),
	.w6(32'h3aa10480),
	.w7(32'h3a55c071),
	.w8(32'h3be84a94),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954c55a),
	.w1(32'hbbc994a2),
	.w2(32'hbbfb1c6f),
	.w3(32'h3b9f110f),
	.w4(32'hba6a28ee),
	.w5(32'hbbb6d10d),
	.w6(32'hbb1bede8),
	.w7(32'hbb8a9294),
	.w8(32'hbc3af28a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a55b5b),
	.w1(32'hbb48e940),
	.w2(32'h3b0a794a),
	.w3(32'hbc76e48d),
	.w4(32'h3b8fa1e3),
	.w5(32'h3bc384fa),
	.w6(32'hbae0bc2e),
	.w7(32'hbc174a39),
	.w8(32'h3a9bf19d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed3a7f),
	.w1(32'hbc35e110),
	.w2(32'hbc199146),
	.w3(32'hbb8a4023),
	.w4(32'h3b06f2a8),
	.w5(32'h3c06f3df),
	.w6(32'hbb58ca43),
	.w7(32'h3a54e112),
	.w8(32'hbb5409ed),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb1d4e),
	.w1(32'hbb2500fd),
	.w2(32'h3b84ee7e),
	.w3(32'h3b13815f),
	.w4(32'hbbf488e2),
	.w5(32'hba7b778a),
	.w6(32'hbb91687a),
	.w7(32'h3bc56898),
	.w8(32'hba54f797),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bb79a),
	.w1(32'hba6c7d99),
	.w2(32'hb8ad79e0),
	.w3(32'hba885147),
	.w4(32'hb9a94f48),
	.w5(32'h38c3e053),
	.w6(32'hba964d34),
	.w7(32'hb9a40986),
	.w8(32'h39ffaf25),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b13691),
	.w1(32'hb9a42b61),
	.w2(32'hba078b50),
	.w3(32'h39b74d9e),
	.w4(32'hba367af4),
	.w5(32'h39d8457b),
	.w6(32'h3a13e710),
	.w7(32'hba07f10f),
	.w8(32'hb90715d3),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba078723),
	.w1(32'h37823053),
	.w2(32'h3a1433bb),
	.w3(32'hb834efd4),
	.w4(32'h39f9e40b),
	.w5(32'h3b6b88ec),
	.w6(32'hba2d2a0c),
	.w7(32'h3a003d3b),
	.w8(32'h3b85dc3d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b163429),
	.w1(32'h3ad59fe6),
	.w2(32'hba6c6064),
	.w3(32'h3aa9cc36),
	.w4(32'hbadd8494),
	.w5(32'h3ac3f162),
	.w6(32'h3aec9d3f),
	.w7(32'hba86cb76),
	.w8(32'h3b192996),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b6e01),
	.w1(32'h3b58b7b9),
	.w2(32'h397c8402),
	.w3(32'h3b3a7544),
	.w4(32'h39719907),
	.w5(32'hba6d5f07),
	.w6(32'h3b2b669f),
	.w7(32'h3a8229d2),
	.w8(32'hba49dbda),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87daeb),
	.w1(32'h3888ffd0),
	.w2(32'hb90288d6),
	.w3(32'hb9dca68b),
	.w4(32'hba1a4ec6),
	.w5(32'hba31c934),
	.w6(32'hb951f71a),
	.w7(32'hb9c51499),
	.w8(32'hba3631f1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961810a),
	.w1(32'hb9b36cf6),
	.w2(32'hba471bcd),
	.w3(32'h3913d830),
	.w4(32'h3a330952),
	.w5(32'h3992670f),
	.w6(32'h38be251b),
	.w7(32'h38cb70f8),
	.w8(32'h38accd80),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b52f53),
	.w1(32'h39859640),
	.w2(32'hb817578a),
	.w3(32'h3a8a847f),
	.w4(32'hb75899f6),
	.w5(32'hbaaceb91),
	.w6(32'h3a1a640a),
	.w7(32'hb902f138),
	.w8(32'hba985f14),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89197b),
	.w1(32'h3a457771),
	.w2(32'h3a264e09),
	.w3(32'h39ddc49c),
	.w4(32'h3aa27d81),
	.w5(32'h3a565602),
	.w6(32'h3a95ce11),
	.w7(32'h3acf2d6f),
	.w8(32'h3a76c6c1),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58d7d0),
	.w1(32'h39c999eb),
	.w2(32'h36f84a13),
	.w3(32'h3a17867f),
	.w4(32'hb85c41e1),
	.w5(32'hb9855384),
	.w6(32'h3a4b5427),
	.w7(32'h39064da2),
	.w8(32'hb9b51062),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba037975),
	.w1(32'hb9722ded),
	.w2(32'h3a5b8a61),
	.w3(32'hb9b017d3),
	.w4(32'h39c0f954),
	.w5(32'hb98f9c38),
	.w6(32'hb9dc8f47),
	.w7(32'h39ba6588),
	.w8(32'hb9d76afb),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9304361),
	.w1(32'hb940ee6b),
	.w2(32'h39a2bff0),
	.w3(32'h3942d3a0),
	.w4(32'h3a34edbb),
	.w5(32'h3a4d2e9a),
	.w6(32'hb94e16d2),
	.w7(32'h3892da6c),
	.w8(32'h3a0cffe3),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e48058),
	.w1(32'h39aed393),
	.w2(32'hb9014e5e),
	.w3(32'h3a1d235a),
	.w4(32'h3991161a),
	.w5(32'hbb08308e),
	.w6(32'h39f3e7af),
	.w7(32'h39d34ce9),
	.w8(32'hbb134f5f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab25fac),
	.w1(32'hbb493e88),
	.w2(32'hbb09d3b1),
	.w3(32'hbb675b6d),
	.w4(32'hbb0839eb),
	.w5(32'h38f0cf8b),
	.w6(32'hbac2ed91),
	.w7(32'hbb39b83c),
	.w8(32'hb8b6608a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7996110),
	.w1(32'hb8a1fd36),
	.w2(32'h3854a7a8),
	.w3(32'h3a154b41),
	.w4(32'h3a17be6b),
	.w5(32'hba134729),
	.w6(32'hb94b2ed3),
	.w7(32'hb9ae4d4f),
	.w8(32'hba3bfbac),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25567a),
	.w1(32'h3a9d6b4a),
	.w2(32'h3b4f65e4),
	.w3(32'hb9fe22d2),
	.w4(32'hb8fbc5c7),
	.w5(32'hba0e0cfa),
	.w6(32'hba149e05),
	.w7(32'h3a94ba16),
	.w8(32'hb86198b0),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ec694),
	.w1(32'hba10ee86),
	.w2(32'hba031a39),
	.w3(32'hba5110b7),
	.w4(32'h38c1b07e),
	.w5(32'hbac9ca70),
	.w6(32'hba34abd1),
	.w7(32'hba24bf27),
	.w8(32'hbaa42f2c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aaa22a),
	.w1(32'hbaaf7fe1),
	.w2(32'hbae53e2e),
	.w3(32'hbaa5985b),
	.w4(32'hba0448ef),
	.w5(32'h3a2146cb),
	.w6(32'hb950ea60),
	.w7(32'hbaa84c46),
	.w8(32'h39c3114f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5013e),
	.w1(32'hb9c2fdfe),
	.w2(32'hb9d6ce63),
	.w3(32'hb933b8b9),
	.w4(32'hb9c36d33),
	.w5(32'hba1aca7b),
	.w6(32'hb9fad0b6),
	.w7(32'hba2f832a),
	.w8(32'hb9f70ee9),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd707a),
	.w1(32'hb9a7ce9b),
	.w2(32'hba141eb7),
	.w3(32'hba9cb910),
	.w4(32'hba90def5),
	.w5(32'hbb068a90),
	.w6(32'hb8903581),
	.w7(32'hb98e19c4),
	.w8(32'hbacc5ffd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e900a),
	.w1(32'hb99eb1ec),
	.w2(32'hb88b7251),
	.w3(32'hba375f0d),
	.w4(32'hb7d07699),
	.w5(32'hba01383f),
	.w6(32'hb8e72702),
	.w7(32'hb8ad8aa9),
	.w8(32'hb9bb5fd5),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c0f12),
	.w1(32'hba0d3600),
	.w2(32'hba19c749),
	.w3(32'hb9a0c4f9),
	.w4(32'hb9e73dc2),
	.w5(32'hbaa4856d),
	.w6(32'hba318dcc),
	.w7(32'hb9b3673b),
	.w8(32'hbb0d80d9),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad241de),
	.w1(32'hbad02a8e),
	.w2(32'hbb793c96),
	.w3(32'hbb044226),
	.w4(32'hba11690d),
	.w5(32'h3a6a003d),
	.w6(32'h3a1d5b2c),
	.w7(32'hbb02a1e4),
	.w8(32'h3a7c83df),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e2651),
	.w1(32'hb67510e9),
	.w2(32'hb83b3f82),
	.w3(32'hb7a27279),
	.w4(32'hb8009256),
	.w5(32'h3981dedc),
	.w6(32'h39279dd5),
	.w7(32'h3977f793),
	.w8(32'hb770392d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f85706),
	.w1(32'h39b5f0fe),
	.w2(32'hb9222cf3),
	.w3(32'h3a0d034f),
	.w4(32'h39a9d527),
	.w5(32'h39aa1a6d),
	.w6(32'h39aab9e1),
	.w7(32'hb985f245),
	.w8(32'h39612f35),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905956d),
	.w1(32'hba41c6a4),
	.w2(32'hb9cc38b6),
	.w3(32'h3995e63d),
	.w4(32'hb778c771),
	.w5(32'h39aee860),
	.w6(32'hb9a36aa4),
	.w7(32'h37d04d3e),
	.w8(32'h3890e8ab),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de4a10),
	.w1(32'h3a1d4ce4),
	.w2(32'h3a00f8c8),
	.w3(32'h3a67aa59),
	.w4(32'h3a968bd3),
	.w5(32'h3aecf81c),
	.w6(32'h39e28f9c),
	.w7(32'h3a0859b2),
	.w8(32'hba1d157c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5db5f1),
	.w1(32'hbb2d796b),
	.w2(32'hba7afe79),
	.w3(32'hba239cb1),
	.w4(32'hbb08555d),
	.w5(32'h3938f4ff),
	.w6(32'hba49b2c0),
	.w7(32'hbb2f0a1d),
	.w8(32'h3987328c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91aabb9),
	.w1(32'hb9534968),
	.w2(32'hb8e61c9a),
	.w3(32'h39ada1bc),
	.w4(32'h39e10e27),
	.w5(32'h3950ccfa),
	.w6(32'h396d268c),
	.w7(32'h3892364b),
	.w8(32'hb74a37ea),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e36cf),
	.w1(32'hb9b63e15),
	.w2(32'h3a179b36),
	.w3(32'hba189e3d),
	.w4(32'hb8b5174d),
	.w5(32'hb9b5f8d1),
	.w6(32'h39a396b9),
	.w7(32'h37811141),
	.w8(32'hb9edd908),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule