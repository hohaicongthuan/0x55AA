module layer_10_featuremap_317(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1e8ef),
	.w1(32'h35e8a0ae),
	.w2(32'h3a226095),
	.w3(32'hba80edea),
	.w4(32'hb9cfbdea),
	.w5(32'h3ab418d3),
	.w6(32'hb9f00769),
	.w7(32'h39720ada),
	.w8(32'hba5ae769),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d2b56),
	.w1(32'h3b18eec2),
	.w2(32'h3b6a3667),
	.w3(32'h3b39ae4a),
	.w4(32'h3b22cf17),
	.w5(32'h3af14e0e),
	.w6(32'h3afbf4ec),
	.w7(32'h3a8d172d),
	.w8(32'h3abfb974),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4e0d8),
	.w1(32'hb9bd435d),
	.w2(32'h383f14a5),
	.w3(32'h371cfb47),
	.w4(32'h3a07e0e5),
	.w5(32'h3937f5e2),
	.w6(32'hb9928db0),
	.w7(32'h39e615d8),
	.w8(32'h39fcb5b8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7585b25),
	.w1(32'hb926ca34),
	.w2(32'h39f9355b),
	.w3(32'hb9ac6a97),
	.w4(32'hb95e2016),
	.w5(32'hbab3b331),
	.w6(32'h39bacb7a),
	.w7(32'h39acc5d4),
	.w8(32'hbb332a39),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef4eee),
	.w1(32'hbadcfbef),
	.w2(32'hbb0dbbbb),
	.w3(32'hba939147),
	.w4(32'hb9d62a0f),
	.w5(32'hbab6e06b),
	.w6(32'hbb1bc606),
	.w7(32'hbb01a91e),
	.w8(32'hba987885),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e1a09),
	.w1(32'hba96b8a4),
	.w2(32'hba8224e2),
	.w3(32'hbac5673d),
	.w4(32'hba7d5ed0),
	.w5(32'hba459239),
	.w6(32'hba9a8df8),
	.w7(32'hba8442ab),
	.w8(32'hba1bdffd),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3920fc4d),
	.w1(32'hb9a99595),
	.w2(32'hb9070b7e),
	.w3(32'hba19ac4f),
	.w4(32'h39fb22ac),
	.w5(32'hba760cd6),
	.w6(32'hba9c8788),
	.w7(32'hba65a35b),
	.w8(32'hbacd6aa0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bf6d7),
	.w1(32'hbbc3fa18),
	.w2(32'hbb8bc426),
	.w3(32'hbbc12485),
	.w4(32'hbb9a3b64),
	.w5(32'hba2a05fc),
	.w6(32'hbbb6a2de),
	.w7(32'hbb4b6315),
	.w8(32'hba1f5635),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e85d6),
	.w1(32'hb8b5ce44),
	.w2(32'h39969bd4),
	.w3(32'hb9e52350),
	.w4(32'h3a0390f6),
	.w5(32'hbaf41748),
	.w6(32'hb974928f),
	.w7(32'h397b1e68),
	.w8(32'hbaf9f8f2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c78b9),
	.w1(32'hb9dca566),
	.w2(32'h3a5122f7),
	.w3(32'hbb55ba12),
	.w4(32'hba50cf32),
	.w5(32'hbab053af),
	.w6(32'hbb1d964a),
	.w7(32'hba9f7d1c),
	.w8(32'hbb0dde86),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab364f9),
	.w1(32'hbad86696),
	.w2(32'hbabc5250),
	.w3(32'hbad4cffb),
	.w4(32'hba7fa1cd),
	.w5(32'hb8363b47),
	.w6(32'hbaa5583a),
	.w7(32'hba75f907),
	.w8(32'h39c6f5a2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d16bb),
	.w1(32'hba87a027),
	.w2(32'hbaf12fe8),
	.w3(32'h39cccf59),
	.w4(32'h3aacb75d),
	.w5(32'h39d95ec0),
	.w6(32'hb9e3e6a7),
	.w7(32'h39657044),
	.w8(32'hb9dc5844),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e7497),
	.w1(32'h3a893e6a),
	.w2(32'h3a0394e8),
	.w3(32'hb95c344e),
	.w4(32'hb79fffb4),
	.w5(32'hbb2254a8),
	.w6(32'h3a0a0d12),
	.w7(32'hbac1f087),
	.w8(32'hbb23029f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95bc081),
	.w1(32'h3a74bdf9),
	.w2(32'hb92cf8af),
	.w3(32'hba63e306),
	.w4(32'hb9bfa9e9),
	.w5(32'hba5a51b0),
	.w6(32'hb92c1e12),
	.w7(32'hba3db54f),
	.w8(32'hba5b5ad9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a900ffa),
	.w1(32'h3afe1828),
	.w2(32'h3b10ca87),
	.w3(32'h3a261e3e),
	.w4(32'h3b121a81),
	.w5(32'h3a99265d),
	.w6(32'h3ab68e7e),
	.w7(32'h3afd083e),
	.w8(32'h3a13b661),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fa7f3),
	.w1(32'h3a0a927a),
	.w2(32'h3a6e9f36),
	.w3(32'hba54c2cf),
	.w4(32'hb7563d3a),
	.w5(32'hb71bd512),
	.w6(32'hba792e9f),
	.w7(32'hba635fb3),
	.w8(32'hba0239bd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900658e),
	.w1(32'h3a7e2e7f),
	.w2(32'h3a41cc2a),
	.w3(32'h39ba3df4),
	.w4(32'h3a0a9a9f),
	.w5(32'h39220e37),
	.w6(32'h3a6a35bc),
	.w7(32'h3948145a),
	.w8(32'h3857c214),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b8e5a),
	.w1(32'hbbdcd495),
	.w2(32'hbc012274),
	.w3(32'hbb9678d2),
	.w4(32'hbbec2503),
	.w5(32'hbbf07100),
	.w6(32'hbbb9d6a0),
	.w7(32'hbbf2028c),
	.w8(32'hbbb1edb6),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe9f63),
	.w1(32'hbb81a403),
	.w2(32'hbb403ce1),
	.w3(32'hbb8342f8),
	.w4(32'hbba54e89),
	.w5(32'hbb95ac76),
	.w6(32'hbb8d9824),
	.w7(32'hbb972575),
	.w8(32'hbb522c8f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b36186),
	.w1(32'h39842cc3),
	.w2(32'hba054d4c),
	.w3(32'hb9f93182),
	.w4(32'h3a03959e),
	.w5(32'hb9332d9a),
	.w6(32'h3a76e3cf),
	.w7(32'hb7ff195f),
	.w8(32'hb9aae33a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfb5f4),
	.w1(32'h39f6f547),
	.w2(32'h393cfda4),
	.w3(32'h39ce1e69),
	.w4(32'hb8c7527b),
	.w5(32'h3a8dea81),
	.w6(32'h3a9ad85d),
	.w7(32'hb92e707d),
	.w8(32'h3aa3c2d6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac031d0),
	.w1(32'h3a7b3a75),
	.w2(32'h3a68907e),
	.w3(32'h3aab9bea),
	.w4(32'h3ac75b09),
	.w5(32'h39bd91f2),
	.w6(32'h39f577d4),
	.w7(32'h3aa73c55),
	.w8(32'h3a07b757),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb265a97),
	.w1(32'hbbdc6fd5),
	.w2(32'hbbccbfb7),
	.w3(32'hbb90aac9),
	.w4(32'hbbbf365e),
	.w5(32'hbbcb851e),
	.w6(32'hbbf6b9d4),
	.w7(32'hbbfb2c9b),
	.w8(32'hbb8a2ccf),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90597eb),
	.w1(32'h3accb80d),
	.w2(32'h3b3d86d0),
	.w3(32'hb9a89d07),
	.w4(32'h3ad8c083),
	.w5(32'h3b11663e),
	.w6(32'hb86b7683),
	.w7(32'h3abaef38),
	.w8(32'hb8cf8c03),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987e236),
	.w1(32'h3a980b88),
	.w2(32'h3ab9f187),
	.w3(32'h3aa91674),
	.w4(32'h3b3f0fce),
	.w5(32'h3ae41682),
	.w6(32'h3a1ececf),
	.w7(32'h3aa57a8a),
	.w8(32'h3a8c9efc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6aa5a5),
	.w1(32'h3aad7720),
	.w2(32'h39f51a27),
	.w3(32'hb9c1ce70),
	.w4(32'h39dcebcf),
	.w5(32'h3a446856),
	.w6(32'h39d75b02),
	.w7(32'h3a1a1521),
	.w8(32'h3aa40438),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a138b25),
	.w1(32'h39c38503),
	.w2(32'h399f5f7c),
	.w3(32'h39b4c213),
	.w4(32'h3a84b07a),
	.w5(32'h3907947b),
	.w6(32'h3a310bf3),
	.w7(32'h3a7d9998),
	.w8(32'hb958bdc1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79827d),
	.w1(32'h3a901b85),
	.w2(32'h3a41b1cf),
	.w3(32'h3a373e4e),
	.w4(32'h3a04c143),
	.w5(32'h39c8956b),
	.w6(32'h3b0db991),
	.w7(32'h39700fed),
	.w8(32'hba8113f1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bf051),
	.w1(32'hba86e359),
	.w2(32'hbac6deca),
	.w3(32'hba300d4b),
	.w4(32'h39646b2d),
	.w5(32'h3a60fb83),
	.w6(32'h37ea995b),
	.w7(32'hba79113a),
	.w8(32'h3a34e656),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb884cd96),
	.w1(32'h3b2488e9),
	.w2(32'h3b401dc7),
	.w3(32'hb984de21),
	.w4(32'h3ac755e6),
	.w5(32'h3a6be19c),
	.w6(32'h3af07b1f),
	.w7(32'h3ac3d4c6),
	.w8(32'h39858a9f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11c80f),
	.w1(32'hba40ff7f),
	.w2(32'hbab13102),
	.w3(32'hba3d6a77),
	.w4(32'hb6d3e259),
	.w5(32'h3a64998a),
	.w6(32'hba901f97),
	.w7(32'h3a1f2e03),
	.w8(32'h3afe12f7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09a9ca),
	.w1(32'h3aa4ee3c),
	.w2(32'hb994851d),
	.w3(32'h3a5443a3),
	.w4(32'h3a563371),
	.w5(32'h39e3c5f7),
	.w6(32'h3a143495),
	.w7(32'h3a081cec),
	.w8(32'h3b183def),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade1bdc),
	.w1(32'h3aa890c0),
	.w2(32'h3aa00933),
	.w3(32'hba1bfb0a),
	.w4(32'h39cdc074),
	.w5(32'h390b4c15),
	.w6(32'hb90df91a),
	.w7(32'h3ac72157),
	.w8(32'hba6e7cf0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbf383),
	.w1(32'h3a0bf784),
	.w2(32'h3a03a1d9),
	.w3(32'hb7f818ca),
	.w4(32'h39883af3),
	.w5(32'h39a24a02),
	.w6(32'h39c9ada1),
	.w7(32'hba4c33bf),
	.w8(32'hba9a5188),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd5f9b),
	.w1(32'hba745d9c),
	.w2(32'hba3e2614),
	.w3(32'hb9c3710d),
	.w4(32'hb994ffc1),
	.w5(32'hba4c600e),
	.w6(32'h3a4a9296),
	.w7(32'hba1bff81),
	.w8(32'hbb087f18),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a05cf),
	.w1(32'hba9fe5a7),
	.w2(32'hba0f385f),
	.w3(32'hba3b3b2b),
	.w4(32'hb9fcdde5),
	.w5(32'hb9a51cf0),
	.w6(32'hbae6f5a9),
	.w7(32'hba98b33f),
	.w8(32'hba67c6a1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba363997),
	.w1(32'hba063862),
	.w2(32'hba7ea874),
	.w3(32'hbaa5851a),
	.w4(32'hba6f6e06),
	.w5(32'hba040478),
	.w6(32'hbb4aa52a),
	.w7(32'hb9fe1e21),
	.w8(32'hbaf1843f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8eda42),
	.w1(32'h3aac8c00),
	.w2(32'h3b07ab0a),
	.w3(32'h3b68bb56),
	.w4(32'h3bd7111e),
	.w5(32'h3bdc9ecc),
	.w6(32'h3b9660ac),
	.w7(32'h3bad9a7a),
	.w8(32'h3b5cde95),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e36da),
	.w1(32'h3bbe979a),
	.w2(32'h3b69c40d),
	.w3(32'h3bcb6a61),
	.w4(32'h3be140de),
	.w5(32'h3b3ac6c1),
	.w6(32'h3bc77daa),
	.w7(32'h3b8fac71),
	.w8(32'h3a2012b0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab00703),
	.w1(32'h39d71e9c),
	.w2(32'h3a5a5b28),
	.w3(32'h3a5471b4),
	.w4(32'h3a45a63a),
	.w5(32'h3a6223c8),
	.w6(32'h396e89ad),
	.w7(32'h3a7f3871),
	.w8(32'h392b8bc8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac411a7),
	.w1(32'hb990a9d2),
	.w2(32'h38feb17e),
	.w3(32'hba9cef22),
	.w4(32'hbaad7a17),
	.w5(32'hba185dcf),
	.w6(32'h381e98f2),
	.w7(32'hba8299fb),
	.w8(32'hb8a1a3d8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23a82a),
	.w1(32'h39f08502),
	.w2(32'h38e95f02),
	.w3(32'hb9d2f44d),
	.w4(32'hb9c7346b),
	.w5(32'h3a055902),
	.w6(32'h38dbf86b),
	.w7(32'hb96717b5),
	.w8(32'h3a9c3026),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a633eb3),
	.w1(32'h38bb6961),
	.w2(32'h383aa585),
	.w3(32'hb8bf14d2),
	.w4(32'h3a3d30b4),
	.w5(32'hbb22b71a),
	.w6(32'h3a7eda61),
	.w7(32'hb895bb72),
	.w8(32'hbb8a0fb2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f704b),
	.w1(32'hbb4eaf2c),
	.w2(32'hbb3908a0),
	.w3(32'hbb876f90),
	.w4(32'hbb30831a),
	.w5(32'hbad4ad87),
	.w6(32'hbb356b1e),
	.w7(32'hbb4b068b),
	.w8(32'hba684c25),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da0961),
	.w1(32'h3ae4aab3),
	.w2(32'h3acec9dc),
	.w3(32'hbad91ea7),
	.w4(32'h39efc02f),
	.w5(32'h3a146306),
	.w6(32'h39b754b5),
	.w7(32'h3a53972a),
	.w8(32'hb9b28059),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3874fb4c),
	.w1(32'h3b1d9573),
	.w2(32'h3b864699),
	.w3(32'h3a149752),
	.w4(32'h3a92316b),
	.w5(32'h3abaaf65),
	.w6(32'hb9383644),
	.w7(32'h3a9dee80),
	.w8(32'h3a152eed),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39419823),
	.w1(32'h3a575620),
	.w2(32'h3a6b6323),
	.w3(32'h3a2b29b4),
	.w4(32'h39d31bb7),
	.w5(32'h3af9c446),
	.w6(32'hba968b6e),
	.w7(32'hb94a0f8c),
	.w8(32'h3ad45de0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ba5d1),
	.w1(32'hbbc7d0fa),
	.w2(32'hbbf7c4e9),
	.w3(32'hbb625ae0),
	.w4(32'hbbbb4cc2),
	.w5(32'hbbe3454f),
	.w6(32'hbbca9e2e),
	.w7(32'hbbcbd547),
	.w8(32'hbbc54df0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395defaa),
	.w1(32'h3a6fd958),
	.w2(32'h3a588c9d),
	.w3(32'h3ad3c755),
	.w4(32'h3ac5630a),
	.w5(32'h3ab5c38e),
	.w6(32'h3ae4cd7e),
	.w7(32'h3abe7468),
	.w8(32'h3acd65c9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade9fc9),
	.w1(32'h396f5e8d),
	.w2(32'h3aad61a0),
	.w3(32'h392c77fa),
	.w4(32'h3a9a38b8),
	.w5(32'hbacfc730),
	.w6(32'hba7ac9be),
	.w7(32'h39dae766),
	.w8(32'hba86c7c0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d5929),
	.w1(32'hb8e54ae4),
	.w2(32'hba4b3f90),
	.w3(32'h391a86d7),
	.w4(32'hba23ad40),
	.w5(32'hba567974),
	.w6(32'h394c7397),
	.w7(32'hba0116dc),
	.w8(32'hb9960c9e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb483a74),
	.w1(32'hbb3f2d68),
	.w2(32'hba999a19),
	.w3(32'hbb1d0a56),
	.w4(32'hbaeabea0),
	.w5(32'hb9f5d328),
	.w6(32'hbaec1826),
	.w7(32'hba87badb),
	.w8(32'hba6b8ae6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c191a),
	.w1(32'hba8d8a0a),
	.w2(32'hba4db2d1),
	.w3(32'hba6227a3),
	.w4(32'hbb0ad197),
	.w5(32'hba81364b),
	.w6(32'hba9f2c1f),
	.w7(32'hba8424d1),
	.w8(32'hbad549eb),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8e7ef),
	.w1(32'hbb5264fd),
	.w2(32'hbad07823),
	.w3(32'hbb4177ca),
	.w4(32'hba62421a),
	.w5(32'hbb2b316c),
	.w6(32'hbad35032),
	.w7(32'hbaebac97),
	.w8(32'hbb283d8c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac12496),
	.w1(32'hbb01fee0),
	.w2(32'hbb243a12),
	.w3(32'hb9c3bfc9),
	.w4(32'hb9c53615),
	.w5(32'hba92455b),
	.w6(32'hba1a63a4),
	.w7(32'hba512739),
	.w8(32'hbaf26a1e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16c4ec),
	.w1(32'hba8c6fd6),
	.w2(32'hba54d1d3),
	.w3(32'hbabcb05f),
	.w4(32'hba6198a4),
	.w5(32'h3a6cd6b2),
	.w6(32'h3a0bb7ea),
	.w7(32'hbab5bf29),
	.w8(32'h3a06f7cb),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d7cee),
	.w1(32'h3a94adea),
	.w2(32'h3a5efcf3),
	.w3(32'h398b2af3),
	.w4(32'h3a11f942),
	.w5(32'hb974a996),
	.w6(32'h3ab66bb3),
	.w7(32'h396ef905),
	.w8(32'hb9cb4d4a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba056c3d),
	.w1(32'hbaa12954),
	.w2(32'h399f5711),
	.w3(32'hba926ce8),
	.w4(32'hb749a6e5),
	.w5(32'h3a5d1a7c),
	.w6(32'hba4f316b),
	.w7(32'h3859cab7),
	.w8(32'h3acd1f76),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b111af0),
	.w1(32'h3a4ddd74),
	.w2(32'h3aa8057f),
	.w3(32'h39663cf3),
	.w4(32'h3aef6979),
	.w5(32'h3aa5b7cf),
	.w6(32'hba077426),
	.w7(32'h3a721a5f),
	.w8(32'h3aa44578),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1f67a),
	.w1(32'h3a959b79),
	.w2(32'h3ae7887d),
	.w3(32'h3b025f00),
	.w4(32'h3aa88f0a),
	.w5(32'h3841833c),
	.w6(32'hb898e1c3),
	.w7(32'h3aa8d1ad),
	.w8(32'hb9d094d0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba535ca0),
	.w1(32'hbaea1aee),
	.w2(32'hbb0d126c),
	.w3(32'hbaf5d00e),
	.w4(32'hbae9e3f3),
	.w5(32'hbb1ee75b),
	.w6(32'hbb195503),
	.w7(32'hbb142c7a),
	.w8(32'hbb11b74e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14cba3),
	.w1(32'hbad7b64d),
	.w2(32'hbadebb2a),
	.w3(32'hbb6ac1b0),
	.w4(32'hbb1200b6),
	.w5(32'hbb543bac),
	.w6(32'hbb2054c1),
	.w7(32'hbb10647f),
	.w8(32'hbb2bef90),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb4a28),
	.w1(32'hbaf30cc9),
	.w2(32'hbb14e3ae),
	.w3(32'hba83a3dc),
	.w4(32'hba770748),
	.w5(32'hb9f64d22),
	.w6(32'hbab3073f),
	.w7(32'hbad14dd0),
	.w8(32'hbadcd77a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae392d7),
	.w1(32'hba0f7dd8),
	.w2(32'hb9b5171b),
	.w3(32'hbab5f15d),
	.w4(32'hba6006f5),
	.w5(32'hb9db9816),
	.w6(32'h3954b87a),
	.w7(32'hba922a87),
	.w8(32'hba9bf783),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe261f),
	.w1(32'hba952660),
	.w2(32'hba8b36a6),
	.w3(32'hba2ba94f),
	.w4(32'hb9f41ef2),
	.w5(32'h3802edd6),
	.w6(32'h390ff6f0),
	.w7(32'hba5658f4),
	.w8(32'hba5e86f7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71cfd5),
	.w1(32'hbab6c731),
	.w2(32'hbab9cdab),
	.w3(32'h3968ad09),
	.w4(32'h37fcb9f3),
	.w5(32'hba4dc874),
	.w6(32'hbaaf469f),
	.w7(32'hb91cfd33),
	.w8(32'hba598d15),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f89f58),
	.w1(32'hba79e61d),
	.w2(32'hba4c4694),
	.w3(32'h39e46218),
	.w4(32'h37a70239),
	.w5(32'hbab11c54),
	.w6(32'hba0c710f),
	.w7(32'hba507cdd),
	.w8(32'hbb0afb2b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb031d9e),
	.w1(32'h39559f83),
	.w2(32'h3aa67f7b),
	.w3(32'h39e24ef8),
	.w4(32'h3a8de31f),
	.w5(32'hba371a33),
	.w6(32'hb945dc5d),
	.w7(32'h3a7341dc),
	.w8(32'hbb08564b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24ad0a),
	.w1(32'hbb5647b0),
	.w2(32'hbb8357f8),
	.w3(32'hbaea1eb1),
	.w4(32'hbb0a01e3),
	.w5(32'hbb877493),
	.w6(32'hbb3e3bf8),
	.w7(32'hbb6b565a),
	.w8(32'hbb5d3a70),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9295b99),
	.w1(32'h3a598a20),
	.w2(32'h3aab05d9),
	.w3(32'h3b0d5e6b),
	.w4(32'h3b8571dc),
	.w5(32'h3b2e3a90),
	.w6(32'h3ac352bb),
	.w7(32'h3a4ed08e),
	.w8(32'h3b1a53e5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a927268),
	.w1(32'h3a001bcd),
	.w2(32'h39e3db50),
	.w3(32'h39a3ae21),
	.w4(32'h3877a3fa),
	.w5(32'hb9e83f9c),
	.w6(32'h3a066c09),
	.w7(32'h3a1d5d7d),
	.w8(32'hba67f861),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba675c41),
	.w1(32'h396e452a),
	.w2(32'hba0eee2a),
	.w3(32'hb98458fb),
	.w4(32'hb9ad76f7),
	.w5(32'h39323454),
	.w6(32'hba270aca),
	.w7(32'hb965fceb),
	.w8(32'hb9c68524),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39924fa4),
	.w1(32'h3a208da0),
	.w2(32'h3a839770),
	.w3(32'h3a876d74),
	.w4(32'h3a69e9bb),
	.w5(32'h3a07c190),
	.w6(32'h390833fa),
	.w7(32'h3a22fcbc),
	.w8(32'hba08f9b0),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae522f),
	.w1(32'hbac9c3bd),
	.w2(32'hbb17780c),
	.w3(32'hba948cff),
	.w4(32'hbb25a47c),
	.w5(32'hbb02f064),
	.w6(32'hbac10288),
	.w7(32'hbb41d287),
	.w8(32'hbb0021a0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ae133),
	.w1(32'hba2c5d94),
	.w2(32'h3a4417ce),
	.w3(32'h39b43837),
	.w4(32'h3a52d159),
	.w5(32'h3a0631d8),
	.w6(32'h3955c16e),
	.w7(32'h3a743e54),
	.w8(32'hb810ec2e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3c577),
	.w1(32'hbb171c6a),
	.w2(32'hbb1a024f),
	.w3(32'hb9b00a90),
	.w4(32'hbb469acd),
	.w5(32'hbab5e047),
	.w6(32'hba571315),
	.w7(32'hbb6fb759),
	.w8(32'hba1f80ff),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd90b2),
	.w1(32'hbb84a1bc),
	.w2(32'hbb93c72d),
	.w3(32'hbb40288a),
	.w4(32'hbbe24e68),
	.w5(32'hbb875d9d),
	.w6(32'hbb9d09b8),
	.w7(32'hbbb0d664),
	.w8(32'hbb786547),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb033352),
	.w1(32'hba88313d),
	.w2(32'h3a047c3d),
	.w3(32'hbae8dbd6),
	.w4(32'hba29ab17),
	.w5(32'hba097e54),
	.w6(32'hb9a55940),
	.w7(32'hba246bbd),
	.w8(32'hba07dbc2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d250c),
	.w1(32'hb9b2085a),
	.w2(32'hb8eaa206),
	.w3(32'h38bb18c0),
	.w4(32'hb95b03a6),
	.w5(32'hb996759a),
	.w6(32'hba8276f7),
	.w7(32'hb8dcdf11),
	.w8(32'hbaa78744),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa9b4f),
	.w1(32'h3980c6a2),
	.w2(32'h3a7b9308),
	.w3(32'h3a13b370),
	.w4(32'h3a0e7d5b),
	.w5(32'h3ac0cfc9),
	.w6(32'h390c025f),
	.w7(32'h38949e78),
	.w8(32'h3a8fce4a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9763c8),
	.w1(32'h3ac38721),
	.w2(32'h3acdcfb8),
	.w3(32'h3983b639),
	.w4(32'h3b05d0fc),
	.w5(32'h3a420422),
	.w6(32'h3a5c58e6),
	.w7(32'h3aeb3b4b),
	.w8(32'h38e1f982),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55c4eb),
	.w1(32'hbb10b33c),
	.w2(32'hbb3c7aee),
	.w3(32'hbacc1603),
	.w4(32'hbb3af061),
	.w5(32'hbb0255ca),
	.w6(32'hbb04f0a6),
	.w7(32'hbb65af29),
	.w8(32'hbb147481),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a6156),
	.w1(32'hba2ef33d),
	.w2(32'hba67a9bb),
	.w3(32'h38d114f5),
	.w4(32'hb9e16a29),
	.w5(32'h3a4af2a7),
	.w6(32'hba2d81b9),
	.w7(32'hba3f3bfb),
	.w8(32'h3a57e9d9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981582f),
	.w1(32'h38badc42),
	.w2(32'hb977b43f),
	.w3(32'h3a54fc27),
	.w4(32'h3a737d6d),
	.w5(32'h3a43cfd0),
	.w6(32'h3a3fa670),
	.w7(32'h3a7a145c),
	.w8(32'h396698be),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96edecf),
	.w1(32'hba41e4cf),
	.w2(32'hb9ff7800),
	.w3(32'h39b755c5),
	.w4(32'hb9bac9d0),
	.w5(32'h392cdbd8),
	.w6(32'hba3541fe),
	.w7(32'hba1a2d73),
	.w8(32'hb9cf7de9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992e2d8),
	.w1(32'h3a4b9fd7),
	.w2(32'hba8827c8),
	.w3(32'h39f44421),
	.w4(32'hba6a6f24),
	.w5(32'hba2853c9),
	.w6(32'hb93a2df4),
	.w7(32'hba486436),
	.w8(32'hb98bbbd0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54802e),
	.w1(32'h3a9212dc),
	.w2(32'h3b3a1d92),
	.w3(32'h3ad92426),
	.w4(32'h3b9a4f5f),
	.w5(32'h3b392cbe),
	.w6(32'h3ae1d9a6),
	.w7(32'h3b4abfc0),
	.w8(32'h3a8a0974),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d4305),
	.w1(32'hba180311),
	.w2(32'hba19b165),
	.w3(32'hb9cbcf7d),
	.w4(32'hb93f437a),
	.w5(32'hb9720b83),
	.w6(32'hba17d198),
	.w7(32'hb93941a0),
	.w8(32'h3698ae32),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac79c39),
	.w1(32'h3a987db3),
	.w2(32'h3a6b3b99),
	.w3(32'h3a3c9076),
	.w4(32'h3aa61ff4),
	.w5(32'h3847ee29),
	.w6(32'h3a38c8aa),
	.w7(32'h39c40f85),
	.w8(32'hb9a18ba3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb896172),
	.w1(32'hbbb39155),
	.w2(32'hbb8ce134),
	.w3(32'hbbfd86d9),
	.w4(32'hbbbe8da9),
	.w5(32'hbb58db83),
	.w6(32'hbc025fd1),
	.w7(32'hbbf0a71b),
	.w8(32'hbb1ec765),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3886af),
	.w1(32'h3aaaf8f5),
	.w2(32'h3a0f0d1d),
	.w3(32'h3aad063d),
	.w4(32'h3ab4af7c),
	.w5(32'h398db000),
	.w6(32'h3a7d9599),
	.w7(32'h3a201108),
	.w8(32'hb9945305),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41a281),
	.w1(32'h3a922f97),
	.w2(32'hb9de24a5),
	.w3(32'h395e9a40),
	.w4(32'h39d79812),
	.w5(32'h3ac4d40b),
	.w6(32'hb97fd3f6),
	.w7(32'hb82c5e77),
	.w8(32'hb809b352),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a368c67),
	.w1(32'h3b053738),
	.w2(32'h398d2b51),
	.w3(32'hb8019ec0),
	.w4(32'h3b0d79c2),
	.w5(32'h3aa068f6),
	.w6(32'h3b49d4fd),
	.w7(32'h3a33c3bf),
	.w8(32'h3a4c6b5e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39961bd6),
	.w1(32'h3a668d7e),
	.w2(32'h3a1cfc6a),
	.w3(32'h3aae090f),
	.w4(32'h3a1c366a),
	.w5(32'hb99b849e),
	.w6(32'h3a87d6a9),
	.w7(32'hb929c302),
	.w8(32'hbb090c20),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab28a2d),
	.w1(32'h3ab9a728),
	.w2(32'h3ac80e13),
	.w3(32'h3b0833af),
	.w4(32'h3b0a2cff),
	.w5(32'h3b20eb38),
	.w6(32'h3aeb8353),
	.w7(32'h3abb2cc9),
	.w8(32'h3b6ffe7b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa48588),
	.w1(32'h3aebb478),
	.w2(32'h3ac17109),
	.w3(32'h3b04ce4c),
	.w4(32'h3b8f8ccb),
	.w5(32'h3b3166ab),
	.w6(32'h3b50c001),
	.w7(32'h3b2c0aef),
	.w8(32'h3af2a786),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3870a1db),
	.w1(32'h3a177a90),
	.w2(32'h3ad5aa01),
	.w3(32'h396eaf4d),
	.w4(32'hba2a488b),
	.w5(32'h3a7a167e),
	.w6(32'hba1aacc2),
	.w7(32'hb93fcc62),
	.w8(32'h3ade13a9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08c3d7),
	.w1(32'h3acaccb1),
	.w2(32'hb9f2110c),
	.w3(32'hba5413a8),
	.w4(32'hba2d8ffb),
	.w5(32'hba830e00),
	.w6(32'h3a719e44),
	.w7(32'hb979123f),
	.w8(32'hba89f21f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a760d47),
	.w1(32'h3a909fb3),
	.w2(32'h3a784b54),
	.w3(32'h3b35f561),
	.w4(32'h3b382a6d),
	.w5(32'h3b1aef30),
	.w6(32'h3a77439a),
	.w7(32'h39768764),
	.w8(32'hb9c8aee9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31d9ef),
	.w1(32'hbb8492a0),
	.w2(32'hbb7ab200),
	.w3(32'hbb7fdc40),
	.w4(32'hbba6b64f),
	.w5(32'hbb79b7fd),
	.w6(32'hbbb23d11),
	.w7(32'hbb9a4d20),
	.w8(32'hbaff3d66),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e2f81),
	.w1(32'h3be1a5b2),
	.w2(32'h3ba4c87b),
	.w3(32'h3bd24806),
	.w4(32'h3c1e4306),
	.w5(32'h3bf98e2f),
	.w6(32'h3ba9cb46),
	.w7(32'h3be685ce),
	.w8(32'h3b37d0ee),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b426a8),
	.w1(32'h3b1cb653),
	.w2(32'h3b60be73),
	.w3(32'h39af1d2f),
	.w4(32'h3af4e28b),
	.w5(32'h3a8f852b),
	.w6(32'h3a639370),
	.w7(32'h3a8f5091),
	.w8(32'h3a2f3bf1),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ee9f1),
	.w1(32'h3a84518d),
	.w2(32'hba3339e5),
	.w3(32'h3ace3e98),
	.w4(32'h3abd624c),
	.w5(32'h3970c7ac),
	.w6(32'hb95c6319),
	.w7(32'hb9ad7058),
	.w8(32'hbb08f680),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6277b9),
	.w1(32'h3a133668),
	.w2(32'hb9fbb8f8),
	.w3(32'h39c4ec7c),
	.w4(32'h3a7e40e7),
	.w5(32'h39d0cf1d),
	.w6(32'h39555a6c),
	.w7(32'h39fbe287),
	.w8(32'h39ff75e3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ccb21),
	.w1(32'hbbeb9bed),
	.w2(32'hbbf33a5d),
	.w3(32'hbb58fb9d),
	.w4(32'hbbdb41e1),
	.w5(32'hbb6b2a67),
	.w6(32'hbb9c45b8),
	.w7(32'hbbd44c1f),
	.w8(32'hbb7ec4dd),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a83bee),
	.w1(32'h373c0739),
	.w2(32'h38a70250),
	.w3(32'h3a32df4d),
	.w4(32'h39b4f93f),
	.w5(32'hba365fbc),
	.w6(32'h39d76917),
	.w7(32'h3a0f243b),
	.w8(32'hb9b9e1c2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cbb810),
	.w1(32'h38290835),
	.w2(32'hb89fa151),
	.w3(32'h390af677),
	.w4(32'h38cc4ae7),
	.w5(32'hb85f2533),
	.w6(32'h389374e4),
	.w7(32'h37bd81d5),
	.w8(32'hb839c74f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f5015c),
	.w1(32'h39f3a606),
	.w2(32'h39c6bf20),
	.w3(32'h398cef7b),
	.w4(32'h39d84c3a),
	.w5(32'hb8acce8f),
	.w6(32'hb9b7ee79),
	.w7(32'hb955efc6),
	.w8(32'h399e6409),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b672b),
	.w1(32'h3a8c839f),
	.w2(32'h3a65af6b),
	.w3(32'hb8db38d3),
	.w4(32'hb80fbaee),
	.w5(32'hba0791e9),
	.w6(32'h39b17b2a),
	.w7(32'hb9245a5e),
	.w8(32'hba002cd1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44f9b1),
	.w1(32'h3aad93bb),
	.w2(32'h3afe93d2),
	.w3(32'h3aac9cd7),
	.w4(32'h3aeef5b1),
	.w5(32'h3a63e71c),
	.w6(32'h3adb3e63),
	.w7(32'h3b02a438),
	.w8(32'h3a82bbf0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7de52b8),
	.w1(32'h3a284455),
	.w2(32'h389d6229),
	.w3(32'h3a3af4ab),
	.w4(32'h3a81603c),
	.w5(32'hb9c1eda9),
	.w6(32'h3a9ac4fe),
	.w7(32'hb9540fe0),
	.w8(32'hb91ffdba),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999dd05),
	.w1(32'h3a3b994e),
	.w2(32'h3aa97137),
	.w3(32'h37feed54),
	.w4(32'h3a59e7a4),
	.w5(32'h3a45907c),
	.w6(32'h39aeee40),
	.w7(32'h3959c6a0),
	.w8(32'hb931847b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6218a9),
	.w1(32'hb9536d78),
	.w2(32'h398421c6),
	.w3(32'hba3b4fa3),
	.w4(32'hba304a43),
	.w5(32'h3a17eda9),
	.w6(32'hba3b43a9),
	.w7(32'h39ae8942),
	.w8(32'h39b9eb0a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98836b8),
	.w1(32'h39b4971c),
	.w2(32'h39c695ac),
	.w3(32'hba785c3c),
	.w4(32'h380d4252),
	.w5(32'hba08aedd),
	.w6(32'hba9f14e5),
	.w7(32'hba4a3342),
	.w8(32'hba95a38e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e531e7),
	.w1(32'h39998522),
	.w2(32'h3a871ec0),
	.w3(32'hb98ac408),
	.w4(32'h3a1d3ca6),
	.w5(32'h3a16df82),
	.w6(32'h39891c91),
	.w7(32'h3a35a0f8),
	.w8(32'h38c4caeb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89a0f03),
	.w1(32'hb79da136),
	.w2(32'h3753938a),
	.w3(32'hb8f478ac),
	.w4(32'hb83daad9),
	.w5(32'h37807d56),
	.w6(32'hb8eff907),
	.w7(32'hb8496f99),
	.w8(32'h37740de8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3797809c),
	.w1(32'h38a99378),
	.w2(32'h3806b190),
	.w3(32'h38403593),
	.w4(32'h3830ca74),
	.w5(32'h388265fd),
	.w6(32'h38364228),
	.w7(32'h3763a9b3),
	.w8(32'hb85679b3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cfdf1a),
	.w1(32'h351132a0),
	.w2(32'h383d368d),
	.w3(32'h38ec45ae),
	.w4(32'h38c5b731),
	.w5(32'h38540ef4),
	.w6(32'h38caed70),
	.w7(32'h38b6c569),
	.w8(32'h38c5dc09),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aafe0a),
	.w1(32'h39de3d26),
	.w2(32'h3a0df50a),
	.w3(32'h3956d5e5),
	.w4(32'h398a8ce7),
	.w5(32'h39e1a576),
	.w6(32'h38263feb),
	.w7(32'h3883996a),
	.w8(32'h38d57540),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907213c),
	.w1(32'h3aaf35d8),
	.w2(32'h3b177984),
	.w3(32'h38d0c59f),
	.w4(32'h3a992f17),
	.w5(32'h3a9a239e),
	.w6(32'h3a032a24),
	.w7(32'h3a38633d),
	.w8(32'h3a2dc80e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c2676),
	.w1(32'h38de71b1),
	.w2(32'hb9253302),
	.w3(32'h39923e77),
	.w4(32'h39efc96d),
	.w5(32'h392c3ff5),
	.w6(32'h39cbb005),
	.w7(32'h39ef20e4),
	.w8(32'hb6ffadd7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfdcfd),
	.w1(32'hba8e6f54),
	.w2(32'hba8f73ed),
	.w3(32'hba20da7c),
	.w4(32'hba8fef00),
	.w5(32'hba740b0c),
	.w6(32'hba9d54f6),
	.w7(32'hbaa333d4),
	.w8(32'hba9d5e53),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99e80b),
	.w1(32'h3b3058b7),
	.w2(32'h3b1bf703),
	.w3(32'h3afbe3e4),
	.w4(32'h3b1e4857),
	.w5(32'h3b01e0f4),
	.w6(32'h3b1e24a4),
	.w7(32'h3ad203ad),
	.w8(32'h3a901bed),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c526f6),
	.w1(32'h38c111a1),
	.w2(32'h368495bf),
	.w3(32'h38af8474),
	.w4(32'hb64aef56),
	.w5(32'hb92ebbd2),
	.w6(32'h38b280e2),
	.w7(32'hb8be52b4),
	.w8(32'hb8da1ee4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390561d9),
	.w1(32'h392c38a5),
	.w2(32'h388f8371),
	.w3(32'h3912507a),
	.w4(32'h38cc9782),
	.w5(32'hb78b8c5a),
	.w6(32'h38612f7c),
	.w7(32'h38b72381),
	.w8(32'hb88bc9de),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f46f7f),
	.w1(32'hb4f10a83),
	.w2(32'h36afca28),
	.w3(32'h37c74773),
	.w4(32'h37dfa841),
	.w5(32'h368289c3),
	.w6(32'hb6407425),
	.w7(32'h35b89518),
	.w8(32'hb69532be),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a33ca),
	.w1(32'h3a68ada7),
	.w2(32'h39d1ce47),
	.w3(32'h3a4a63e9),
	.w4(32'h3a282b01),
	.w5(32'h3809c6cc),
	.w6(32'h3a43811f),
	.w7(32'h3a0b7abc),
	.w8(32'h39aa606c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1ee06),
	.w1(32'hba0786cd),
	.w2(32'h3a8c3e34),
	.w3(32'hbad878b6),
	.w4(32'hbaba73db),
	.w5(32'h39087996),
	.w6(32'hbaf3ebac),
	.w7(32'hba3ea13a),
	.w8(32'hb8a6db74),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa04233),
	.w1(32'h3a4a62b2),
	.w2(32'h3816afb5),
	.w3(32'h39d4e5f4),
	.w4(32'h39833049),
	.w5(32'hba0b02ef),
	.w6(32'h38dcc43a),
	.w7(32'h37faf04f),
	.w8(32'hb9cd2cfb),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380d8d1b),
	.w1(32'hba389074),
	.w2(32'hba5d545f),
	.w3(32'hb94cf32e),
	.w4(32'hba2a3133),
	.w5(32'hba334b9f),
	.w6(32'hba209ee8),
	.w7(32'hba529ae6),
	.w8(32'hba27579c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba236221),
	.w1(32'hba0f8eb5),
	.w2(32'hb9bcea76),
	.w3(32'hb9e9efbb),
	.w4(32'hba3b63d3),
	.w5(32'h39951e5d),
	.w6(32'hba7ae26a),
	.w7(32'hb98e346a),
	.w8(32'hb8b23b1b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea163b),
	.w1(32'h3a36ffac),
	.w2(32'h3a1d943d),
	.w3(32'h3a309efe),
	.w4(32'h3a5d623c),
	.w5(32'h3a117ed1),
	.w6(32'h3a157121),
	.w7(32'h39f4540f),
	.w8(32'h38bbe7a6),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3856837e),
	.w1(32'h39a6531e),
	.w2(32'h39828536),
	.w3(32'hb934709a),
	.w4(32'h3914aeb7),
	.w5(32'h38aea061),
	.w6(32'hb95d4c50),
	.w7(32'hb8b7cd6b),
	.w8(32'h38446b98),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa580b5),
	.w1(32'h3b35b01b),
	.w2(32'h3b7892f9),
	.w3(32'h3aa4975e),
	.w4(32'h3b377db0),
	.w5(32'h3b3d1def),
	.w6(32'h3acd4b8d),
	.w7(32'h3b19bebe),
	.w8(32'h3b03f6c0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4abf4b),
	.w1(32'hbb3d85dd),
	.w2(32'hbb38eb7b),
	.w3(32'hbb259baf),
	.w4(32'hbb42bc02),
	.w5(32'hbb1facc3),
	.w6(32'hbb73cb85),
	.w7(32'hbb6c505e),
	.w8(32'hbb06cf6f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce7281),
	.w1(32'h3ade4d11),
	.w2(32'h3aa634fd),
	.w3(32'h3b04920b),
	.w4(32'h3b092e81),
	.w5(32'h3a7caab4),
	.w6(32'h3b1eefd2),
	.w7(32'h3aae2618),
	.w8(32'h3a6e2057),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afe8ae),
	.w1(32'h39c64759),
	.w2(32'hb9f8b51a),
	.w3(32'h3a4fc2a8),
	.w4(32'h3afc4120),
	.w5(32'h39f58731),
	.w6(32'h39bff418),
	.w7(32'h3a2420cb),
	.w8(32'hba4c6c61),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63db1c),
	.w1(32'hbaa971d3),
	.w2(32'hba8ab10c),
	.w3(32'hba588691),
	.w4(32'hba4217ff),
	.w5(32'h3852a3a2),
	.w6(32'hba866c2b),
	.w7(32'hba73a714),
	.w8(32'h3918c345),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c53197),
	.w1(32'h3a8f1c0b),
	.w2(32'h3aa9eebd),
	.w3(32'h3a2a268a),
	.w4(32'h3a74dad7),
	.w5(32'h3a502092),
	.w6(32'h39effed3),
	.w7(32'h3a1744ff),
	.w8(32'h3a8124b4),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb893f5ec),
	.w1(32'h39d2c315),
	.w2(32'h3a1bb3e9),
	.w3(32'hb9a8451e),
	.w4(32'hb718b638),
	.w5(32'hb9025569),
	.w6(32'hb8fd407e),
	.w7(32'h3875bfe8),
	.w8(32'hb98bbff9),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371d978f),
	.w1(32'h3991a6c9),
	.w2(32'h39acd76f),
	.w3(32'hb8e019a3),
	.w4(32'h3934fe8b),
	.w5(32'h38da7d42),
	.w6(32'hb80e08c6),
	.w7(32'h392f84e9),
	.w8(32'h3849e9e1),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cefe8),
	.w1(32'h3b3a7ab4),
	.w2(32'h3b2dfde8),
	.w3(32'h3b7bb032),
	.w4(32'h3b6fd99b),
	.w5(32'h3b15b672),
	.w6(32'h3b917dbd),
	.w7(32'h3b1b5aa4),
	.w8(32'h3a16169c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfcc66),
	.w1(32'h3a99396a),
	.w2(32'h39cc8f8e),
	.w3(32'h3aa0667b),
	.w4(32'h3aa0839d),
	.w5(32'h39f037ab),
	.w6(32'h3a843464),
	.w7(32'h3a694f21),
	.w8(32'h3a238c56),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c8fc15),
	.w1(32'hb65c55d9),
	.w2(32'h36d26d0d),
	.w3(32'h35a87287),
	.w4(32'hb703d3a4),
	.w5(32'hb64b6ec8),
	.w6(32'h37619d53),
	.w7(32'h37928e56),
	.w8(32'h378a48ee),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7719bbe),
	.w1(32'hb7d2bc28),
	.w2(32'hb6adc057),
	.w3(32'h374eca79),
	.w4(32'h3728b25d),
	.w5(32'h371d29a2),
	.w6(32'h377a0922),
	.w7(32'h371a271e),
	.w8(32'h3745b2af),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a8bb7a),
	.w1(32'hb8879fda),
	.w2(32'h39895582),
	.w3(32'h391da7aa),
	.w4(32'hb7c3b700),
	.w5(32'h38e3daec),
	.w6(32'h3988a339),
	.w7(32'h3992c5ed),
	.w8(32'h38456143),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85f5bf),
	.w1(32'h3b1de6da),
	.w2(32'h3a96326b),
	.w3(32'h3b2a6553),
	.w4(32'h3b1291d8),
	.w5(32'h3a8ef816),
	.w6(32'h3b21ea22),
	.w7(32'h3aa01490),
	.w8(32'h3a5a35ca),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb165338),
	.w1(32'hba609cb1),
	.w2(32'h3992573d),
	.w3(32'hbadde7c2),
	.w4(32'hbacd6c55),
	.w5(32'hba572363),
	.w6(32'hb9f4007c),
	.w7(32'hbae26e41),
	.w8(32'hba61fcb2),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6879fa4),
	.w1(32'h351fcab6),
	.w2(32'h371ee368),
	.w3(32'hb79648a3),
	.w4(32'hb6c55e27),
	.w5(32'hb7091268),
	.w6(32'hb74cf0a4),
	.w7(32'hb748a0e8),
	.w8(32'hb5d9da23),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3884e323),
	.w1(32'h3a07085e),
	.w2(32'h3aa6bdf1),
	.w3(32'hb890bb1b),
	.w4(32'h396a438d),
	.w5(32'h39c19351),
	.w6(32'hb8da6ceb),
	.w7(32'hb801c00b),
	.w8(32'hb9a41d2e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a142b),
	.w1(32'h3a5020dc),
	.w2(32'h3abe612c),
	.w3(32'h3a27644d),
	.w4(32'h39daf780),
	.w5(32'h3911ca84),
	.w6(32'h3a3b52c1),
	.w7(32'h396e1a29),
	.w8(32'hb9326778),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ec4e9),
	.w1(32'hbaf9fdf0),
	.w2(32'hbb323665),
	.w3(32'hbb136d8f),
	.w4(32'hbb20861c),
	.w5(32'hbb3f3dc8),
	.w6(32'hbb5755e6),
	.w7(32'hbb778f35),
	.w8(32'hbb73c913),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e8a59),
	.w1(32'h3a28c1df),
	.w2(32'h3a0d7b2c),
	.w3(32'h3a1c876e),
	.w4(32'h3b076812),
	.w5(32'h3a8d6fe1),
	.w6(32'h3aa22119),
	.w7(32'h3a898f8a),
	.w8(32'h39ec206c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af38f07),
	.w1(32'h3b16c022),
	.w2(32'h3b0c7039),
	.w3(32'h3b00202d),
	.w4(32'h3b2c72aa),
	.w5(32'h3af69894),
	.w6(32'h3b1c2d4a),
	.w7(32'h3af3c9be),
	.w8(32'h3ab69143),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a518baf),
	.w1(32'h38f83db1),
	.w2(32'hb9156812),
	.w3(32'h3aa88730),
	.w4(32'h3a8d96a1),
	.w5(32'h39b60011),
	.w6(32'h3a81367f),
	.w7(32'h3a530cce),
	.w8(32'h39d33ff7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3ebb8),
	.w1(32'hba4ee33b),
	.w2(32'hb85298ab),
	.w3(32'hba968328),
	.w4(32'hb94e57e5),
	.w5(32'hb9811bf9),
	.w6(32'hba6614c7),
	.w7(32'h39343382),
	.w8(32'hb9be1b7b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69aa34),
	.w1(32'h3b77674c),
	.w2(32'h3b4d56eb),
	.w3(32'h3bb19278),
	.w4(32'h3b9cc270),
	.w5(32'h3b6694c5),
	.w6(32'h3b9fa284),
	.w7(32'h3b41a817),
	.w8(32'h3b02b56a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aa666f),
	.w1(32'h3a375a8b),
	.w2(32'h3a51620d),
	.w3(32'h3a0ebc40),
	.w4(32'h3a8568a4),
	.w5(32'h3a86450b),
	.w6(32'h39d5f083),
	.w7(32'h3a40e26e),
	.w8(32'h3a4ab9e9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953eff5),
	.w1(32'hba6d0f08),
	.w2(32'hba19a93f),
	.w3(32'hba2747a4),
	.w4(32'hba5371c4),
	.w5(32'hb9fe3494),
	.w6(32'hba7a01c9),
	.w7(32'hba92b607),
	.w8(32'hb9c96251),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3880db9f),
	.w1(32'h3911310b),
	.w2(32'h3902a595),
	.w3(32'h39377f1d),
	.w4(32'h39345ab8),
	.w5(32'h38ab482b),
	.w6(32'h395d4dd2),
	.w7(32'h394866a9),
	.w8(32'h38f395f0),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997d7d4),
	.w1(32'h38458877),
	.w2(32'h393737a4),
	.w3(32'h38cd2f28),
	.w4(32'h398cc3ff),
	.w5(32'h393d993d),
	.w6(32'hb9f85460),
	.w7(32'hb8afda2c),
	.w8(32'h39b1e4c5),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6316843),
	.w1(32'hb89ad71a),
	.w2(32'hb839e938),
	.w3(32'h391d37a3),
	.w4(32'h392ecfbf),
	.w5(32'h390f4e1a),
	.w6(32'h3863584c),
	.w7(32'h38f01187),
	.w8(32'h377b3618),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f78d74),
	.w1(32'h39c1896e),
	.w2(32'h3a48e99f),
	.w3(32'hba18d93c),
	.w4(32'h3a07c4dc),
	.w5(32'h39b2f412),
	.w6(32'hb886c8a9),
	.w7(32'h3a5c0d94),
	.w8(32'h39dbafe0),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b5d03b),
	.w1(32'h37ee29de),
	.w2(32'hb97eafb0),
	.w3(32'h397f2ed9),
	.w4(32'h39629cc1),
	.w5(32'hb854a4d0),
	.w6(32'h387cada3),
	.w7(32'h3912d713),
	.w8(32'hb908788a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374a8c94),
	.w1(32'h38dcb254),
	.w2(32'h39b144ed),
	.w3(32'h3a3d67ce),
	.w4(32'h3a9df163),
	.w5(32'h3a91679f),
	.w6(32'hb84c3934),
	.w7(32'h3a0fa357),
	.w8(32'h39a8b296),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38db5954),
	.w1(32'h3912083a),
	.w2(32'h38fa6f9a),
	.w3(32'h38adaac3),
	.w4(32'h391e0a88),
	.w5(32'h3952bd96),
	.w6(32'h381baccf),
	.w7(32'h3901b0a0),
	.w8(32'h395d56b1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39579838),
	.w1(32'hb988daf4),
	.w2(32'hb9c55954),
	.w3(32'h39460d96),
	.w4(32'hb8ed50e9),
	.w5(32'hb96f447f),
	.w6(32'h38a192ae),
	.w7(32'hb97be2ea),
	.w8(32'hb9c4691e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91a3a4),
	.w1(32'h3b0bd28f),
	.w2(32'h3aa93fc9),
	.w3(32'h3ad4a733),
	.w4(32'h3b34b7d0),
	.w5(32'h3aa2d8c5),
	.w6(32'h3b16ade0),
	.w7(32'h3b2591d4),
	.w8(32'h3a98e269),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f794b0),
	.w1(32'h38c994a9),
	.w2(32'hb953da23),
	.w3(32'hbaa4b505),
	.w4(32'hba9e3188),
	.w5(32'hba041f96),
	.w6(32'hbb812fe4),
	.w7(32'hbb0f33d0),
	.w8(32'hbae8cb5c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d2c6b5),
	.w1(32'h3977c8be),
	.w2(32'hb86b00c5),
	.w3(32'h39572db0),
	.w4(32'h39a801a1),
	.w5(32'h3902de68),
	.w6(32'h397e6b94),
	.w7(32'h392c91e9),
	.w8(32'h39747807),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d0a4c),
	.w1(32'h3a51ebc5),
	.w2(32'h3a437a39),
	.w3(32'hb9347e6c),
	.w4(32'h3a693627),
	.w5(32'hb8d32a29),
	.w6(32'h3a646b46),
	.w7(32'h3926b7b2),
	.w8(32'hba1a0067),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a320d2),
	.w1(32'h39a78b58),
	.w2(32'h391eed68),
	.w3(32'h3a12c9b5),
	.w4(32'h3a075b31),
	.w5(32'h39661099),
	.w6(32'h3a12052c),
	.w7(32'h398795b3),
	.w8(32'h38f90912),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3973d2f2),
	.w1(32'h3a66c02f),
	.w2(32'hb8e47efa),
	.w3(32'h3a5f6ee2),
	.w4(32'h3a4c52cb),
	.w5(32'hb9a6ea77),
	.w6(32'h3a99d609),
	.w7(32'hb85b59a3),
	.w8(32'hb9daa326),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a0d55),
	.w1(32'hba20924c),
	.w2(32'hba75cde1),
	.w3(32'hb97c41b3),
	.w4(32'hb7722ca3),
	.w5(32'hb992eb6a),
	.w6(32'hba83a1df),
	.w7(32'hba4260c7),
	.w8(32'hba39506c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96f403),
	.w1(32'hba015211),
	.w2(32'hb993ced7),
	.w3(32'hbb1da5ba),
	.w4(32'hbaa6c81e),
	.w5(32'hba9e68ae),
	.w6(32'hbb350b48),
	.w7(32'hbb0152a4),
	.w8(32'hbaf3d486),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea79cc),
	.w1(32'h39efae2a),
	.w2(32'h39d08945),
	.w3(32'h3a19cb51),
	.w4(32'h3a3b90ea),
	.w5(32'h3a11f4ed),
	.w6(32'h39e19491),
	.w7(32'h3a560008),
	.w8(32'h3a39e4bc),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2dda3),
	.w1(32'h3ad71574),
	.w2(32'h3a8aacbd),
	.w3(32'h3abedd30),
	.w4(32'h3ae5c15c),
	.w5(32'h3a4476d6),
	.w6(32'h3ab46905),
	.w7(32'h3aaa26f4),
	.w8(32'h39960bc9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375eb154),
	.w1(32'h37919aaa),
	.w2(32'h37ddec64),
	.w3(32'h37b25d4e),
	.w4(32'hb64b419b),
	.w5(32'h3813da9d),
	.w6(32'h385b616f),
	.w7(32'h37a2a610),
	.w8(32'h3814b729),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af1f03),
	.w1(32'hb82da389),
	.w2(32'hb8fe72da),
	.w3(32'hb9e9738b),
	.w4(32'h3797045f),
	.w5(32'h3767a2b1),
	.w6(32'hb9e7a73e),
	.w7(32'hb81a1580),
	.w8(32'hb90b1a0b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb848c104),
	.w1(32'h38a6fbaf),
	.w2(32'h3914854d),
	.w3(32'hb785d2a8),
	.w4(32'h38feacd9),
	.w5(32'h396f8b6c),
	.w6(32'hb820b700),
	.w7(32'h389ce516),
	.w8(32'h3952cbda),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa725e),
	.w1(32'hb9e34a47),
	.w2(32'hb9b36c40),
	.w3(32'hb9b93af4),
	.w4(32'hb90aadcc),
	.w5(32'hba220b11),
	.w6(32'hba28e260),
	.w7(32'hba700872),
	.w8(32'hbaba35a1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3685b937),
	.w1(32'h35ba9537),
	.w2(32'hb6e2059b),
	.w3(32'hb70cccdd),
	.w4(32'hb7870707),
	.w5(32'h36ef80bd),
	.w6(32'h36f8bb69),
	.w7(32'hb7a4fcd9),
	.w8(32'h37168745),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8965d12),
	.w1(32'hb86bbbe7),
	.w2(32'hb88a679c),
	.w3(32'h37fe7505),
	.w4(32'h37e033eb),
	.w5(32'hb788d89c),
	.w6(32'h3821bd2b),
	.w7(32'h38476fe6),
	.w8(32'hb881b58b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9987912),
	.w1(32'hb9df6177),
	.w2(32'h39e7aaff),
	.w3(32'hb95c6776),
	.w4(32'h37168da5),
	.w5(32'h3a1d7b82),
	.w6(32'hba63f274),
	.w7(32'hb9e92d9f),
	.w8(32'h39e0121a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a767fda),
	.w1(32'h3915d6b5),
	.w2(32'h3a82c28d),
	.w3(32'h3b1679af),
	.w4(32'h3ab09b33),
	.w5(32'h3a7e1131),
	.w6(32'h3a3cc395),
	.w7(32'hb930b7f4),
	.w8(32'h394a1f37),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb823cc80),
	.w1(32'hb8c56be8),
	.w2(32'hb7ab2af2),
	.w3(32'hb9895800),
	.w4(32'h392b2584),
	.w5(32'h39fe1c99),
	.w6(32'hba6944df),
	.w7(32'h3941b85d),
	.w8(32'hb955fd02),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4929e9),
	.w1(32'hba9dcd8d),
	.w2(32'hba2fcde8),
	.w3(32'hba4ae9d4),
	.w4(32'hba019583),
	.w5(32'hba8b2f33),
	.w6(32'hba4fca1a),
	.w7(32'hba57ef5a),
	.w8(32'hb99b1b6b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb61c2),
	.w1(32'hbbc1b6ef),
	.w2(32'hbb7f8d74),
	.w3(32'hbbef3826),
	.w4(32'hbbfa2daf),
	.w5(32'hbbbe18de),
	.w6(32'hbbaded8b),
	.w7(32'hbba29b9d),
	.w8(32'hbb7664e6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00751f),
	.w1(32'h3b7d9d0c),
	.w2(32'h3b224244),
	.w3(32'h3b940251),
	.w4(32'h3bc7fe75),
	.w5(32'h3af69259),
	.w6(32'h3baea71a),
	.w7(32'h3b95e226),
	.w8(32'h3a070688),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393692e6),
	.w1(32'hb8d786dd),
	.w2(32'hb967c393),
	.w3(32'h3912bca8),
	.w4(32'hb8a17683),
	.w5(32'hb8cf8ee1),
	.w6(32'h380061cc),
	.w7(32'hb84fab80),
	.w8(32'hb99e71b8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fbb0bc),
	.w1(32'hb76cc469),
	.w2(32'hb67b8abe),
	.w3(32'hb6c342fd),
	.w4(32'hb6c8de4d),
	.w5(32'hb7f1118b),
	.w6(32'hb86d1e79),
	.w7(32'hb889c163),
	.w8(32'hb7fcc514),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9145842),
	.w1(32'hb86d2eb9),
	.w2(32'hb978c292),
	.w3(32'hb6067c22),
	.w4(32'h38dc8432),
	.w5(32'hb98777c8),
	.w6(32'h37da36d8),
	.w7(32'h3724693d),
	.w8(32'hb9a14f88),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c02291),
	.w1(32'hb7765871),
	.w2(32'h375f5e60),
	.w3(32'h37721135),
	.w4(32'h37182cf4),
	.w5(32'h37946a67),
	.w6(32'hb5f999d5),
	.w7(32'h358cf2bd),
	.w8(32'h37000a87),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a090b33),
	.w1(32'h3a301194),
	.w2(32'h39e71458),
	.w3(32'h39fad7ac),
	.w4(32'h3a4cf104),
	.w5(32'h39bce892),
	.w6(32'h39c84f61),
	.w7(32'h3a2244c4),
	.w8(32'h398a0236),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18026e),
	.w1(32'h3b0e09e0),
	.w2(32'h3a8e0e66),
	.w3(32'h3b1201c4),
	.w4(32'h3b045fb4),
	.w5(32'h3a7ddb48),
	.w6(32'h3ac60dd9),
	.w7(32'h3a7a0b2e),
	.w8(32'h3a18b274),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886ea79),
	.w1(32'h3a9d285c),
	.w2(32'h3abcb6b6),
	.w3(32'h3a87e4ff),
	.w4(32'h3aca0c20),
	.w5(32'h3a609ea5),
	.w6(32'h3afc8afd),
	.w7(32'h3a8ffc15),
	.w8(32'h3aa11a29),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2c3cd),
	.w1(32'hb9c9411f),
	.w2(32'h39056eae),
	.w3(32'hb9aecc68),
	.w4(32'hb8369101),
	.w5(32'h39af527c),
	.w6(32'hb9a5dd19),
	.w7(32'h383cf819),
	.w8(32'h39ee07d0),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf33bd),
	.w1(32'hba5b1ef3),
	.w2(32'hbae1caa4),
	.w3(32'hbab5b4cb),
	.w4(32'hba4e2515),
	.w5(32'hbb2b6ce2),
	.w6(32'hbab64b75),
	.w7(32'hbac7b873),
	.w8(32'hbb03e720),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3532de),
	.w1(32'hba314aaa),
	.w2(32'h39004380),
	.w3(32'hb8e08ea6),
	.w4(32'hb9cd21e1),
	.w5(32'hb8a3676c),
	.w6(32'hb8a62908),
	.w7(32'hb9405866),
	.w8(32'h38a32c54),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3782586c),
	.w1(32'h37ab58c0),
	.w2(32'h38539f3b),
	.w3(32'h3629217e),
	.w4(32'h37810a28),
	.w5(32'h3822e31b),
	.w6(32'h36e1e266),
	.w7(32'h37bcc4cb),
	.w8(32'h382a15e9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b2a733),
	.w1(32'hba3b84cb),
	.w2(32'hba15a369),
	.w3(32'hba12b647),
	.w4(32'hba837c9f),
	.w5(32'hb9aa921d),
	.w6(32'hba4d946a),
	.w7(32'hba08e8b0),
	.w8(32'h3844a300),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e20014),
	.w1(32'h375f34c2),
	.w2(32'h38a2dcb9),
	.w3(32'h37d60536),
	.w4(32'h37cb895e),
	.w5(32'h38a9b30f),
	.w6(32'h38117f32),
	.w7(32'h37b26f6d),
	.w8(32'h38bc6093),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d46c16),
	.w1(32'hb938a73d),
	.w2(32'hb9a960bd),
	.w3(32'hba0bbbd2),
	.w4(32'hb7e28d5f),
	.w5(32'hb9801556),
	.w6(32'hba2fec2d),
	.w7(32'hb96b8b07),
	.w8(32'hb9e84e95),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15cc1e),
	.w1(32'h3b467a9e),
	.w2(32'h3b20845c),
	.w3(32'h3b6a5c0d),
	.w4(32'h3b8e47dc),
	.w5(32'h3b561f50),
	.w6(32'h3b63bc6b),
	.w7(32'h3b59b893),
	.w8(32'h3b13479e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a299630),
	.w1(32'h3a85bc56),
	.w2(32'h39ff1d33),
	.w3(32'h3a9c132e),
	.w4(32'h3acca85b),
	.w5(32'h37a214c7),
	.w6(32'h3ab909c7),
	.w7(32'h3a5c5e0f),
	.w8(32'hb9e29696),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373c4353),
	.w1(32'h3951a3f4),
	.w2(32'h399355da),
	.w3(32'h39c6438c),
	.w4(32'h3a0c99ae),
	.w5(32'h39cbacbd),
	.w6(32'h395e6e93),
	.w7(32'h399f3bfd),
	.w8(32'h39189ba6),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a769378),
	.w1(32'h3aed1fec),
	.w2(32'h3abc0a57),
	.w3(32'h3b288f09),
	.w4(32'h3b1723f0),
	.w5(32'h3a2dbca4),
	.w6(32'h3b47f733),
	.w7(32'h3ae0b3ce),
	.w8(32'h3a05e1f4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9a74e),
	.w1(32'h38ab3355),
	.w2(32'h3a03e4c0),
	.w3(32'hba8e7a14),
	.w4(32'hb99f33b1),
	.w5(32'hb98df057),
	.w6(32'hba0d93c3),
	.w7(32'h385d6e33),
	.w8(32'hb9555de0),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0eb475),
	.w1(32'hba5d026d),
	.w2(32'h3a95c323),
	.w3(32'hbb335255),
	.w4(32'hbabc4acb),
	.w5(32'h39001b2c),
	.w6(32'hbae6fa03),
	.w7(32'hbb067229),
	.w8(32'hba56328f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3792c615),
	.w1(32'h37ac24d8),
	.w2(32'hb759ae27),
	.w3(32'h380d53ad),
	.w4(32'h38116951),
	.w5(32'hb779e6ce),
	.w6(32'hb60f059b),
	.w7(32'h3635d390),
	.w8(32'hb7c9ed49),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7506765),
	.w1(32'hb691adb7),
	.w2(32'h382b46e0),
	.w3(32'hb83dfb39),
	.w4(32'hb74abdde),
	.w5(32'h382009ca),
	.w6(32'hb73afe82),
	.w7(32'hb6ff76d5),
	.w8(32'h3898132d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b71c8),
	.w1(32'h3a6d3b50),
	.w2(32'h3aae0de0),
	.w3(32'h3ad86898),
	.w4(32'h3a856812),
	.w5(32'h39ea99de),
	.w6(32'h39ddf5e2),
	.w7(32'h3966b4d8),
	.w8(32'h398b6f17),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45da4e),
	.w1(32'hba9871ab),
	.w2(32'hba1182f8),
	.w3(32'hbad66bdb),
	.w4(32'hbacc53bf),
	.w5(32'hbac4512f),
	.w6(32'hbb94ecca),
	.w7(32'hbb2a54ce),
	.w8(32'hbb10f366),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a2b9b),
	.w1(32'h3a70d0ed),
	.w2(32'h3b1742bd),
	.w3(32'h3a1f108e),
	.w4(32'h3aa7636e),
	.w5(32'h3ab151b2),
	.w6(32'h3a056154),
	.w7(32'h3a9bc8a8),
	.w8(32'h3a073f0f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff6b3b),
	.w1(32'hba0fd2ac),
	.w2(32'h382873a2),
	.w3(32'hb82a30de),
	.w4(32'h399c930c),
	.w5(32'h3a4f8817),
	.w6(32'hb7940d42),
	.w7(32'hb8cee096),
	.w8(32'hb7913ab4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bedf20),
	.w1(32'h37a2ce99),
	.w2(32'h3890ad24),
	.w3(32'hb80cf30f),
	.w4(32'h3751b381),
	.w5(32'hb5c4a29f),
	.w6(32'hb81188f2),
	.w7(32'hb76ceaa5),
	.w8(32'h37bda6e7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb740682f),
	.w1(32'hb8ac724d),
	.w2(32'h3949317d),
	.w3(32'hb984b3a0),
	.w4(32'hb923805c),
	.w5(32'h39356c8b),
	.w6(32'hb99079e0),
	.w7(32'hb94a7265),
	.w8(32'h38457e92),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ad49b),
	.w1(32'h38e91feb),
	.w2(32'hb9e59e88),
	.w3(32'hb9e00022),
	.w4(32'hba180f1e),
	.w5(32'hba308d1d),
	.w6(32'hbaa7b4ff),
	.w7(32'hb9dde78a),
	.w8(32'hba73b333),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9137c1),
	.w1(32'hbba21314),
	.w2(32'hbb5b0829),
	.w3(32'hbbb45396),
	.w4(32'hbba4a56d),
	.w5(32'hbb4902e2),
	.w6(32'hbba989ab),
	.w7(32'hbb96f620),
	.w8(32'hbaff22a8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3456b),
	.w1(32'hba3963cc),
	.w2(32'hbb2477bc),
	.w3(32'h3a9213f6),
	.w4(32'hbb0bf51e),
	.w5(32'hbb0d8df5),
	.w6(32'hbae2cca0),
	.w7(32'hbb149f86),
	.w8(32'hbb563bf5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31e5c1),
	.w1(32'h3a98347c),
	.w2(32'h3a507a83),
	.w3(32'h3acbef85),
	.w4(32'h3af4ff50),
	.w5(32'h3aac0c9e),
	.w6(32'h3ae3a4f5),
	.w7(32'h3adb5c78),
	.w8(32'h3a7255ec),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0356b),
	.w1(32'h3a25be14),
	.w2(32'h3ab26260),
	.w3(32'hb9229d61),
	.w4(32'h3aec579a),
	.w5(32'h3acddb4a),
	.w6(32'h39be8a0b),
	.w7(32'h3a651194),
	.w8(32'h3a30c06e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376b6d3e),
	.w1(32'h378aef15),
	.w2(32'h37e70272),
	.w3(32'h37912390),
	.w4(32'h3770c18c),
	.w5(32'h37bfc2d5),
	.w6(32'h37dbe7aa),
	.w7(32'h378eebb6),
	.w8(32'h37ad7726),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c60e60),
	.w1(32'hb7de3d63),
	.w2(32'h35be6546),
	.w3(32'h3602b282),
	.w4(32'hb6c0bad4),
	.w5(32'h3611cdad),
	.w6(32'hb5ab3e69),
	.w7(32'hb633c5b4),
	.w8(32'h36e2497d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92666d2),
	.w1(32'h3715e9c2),
	.w2(32'h38ed8f3d),
	.w3(32'h384443d6),
	.w4(32'h392b42b6),
	.w5(32'h38b37cc6),
	.w6(32'h382f1965),
	.w7(32'h38878a8d),
	.w8(32'hb8b69827),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37106d12),
	.w1(32'h36eb9810),
	.w2(32'h380ca888),
	.w3(32'hb7a72d93),
	.w4(32'h3678924a),
	.w5(32'hba90d402),
	.w6(32'hb76355cd),
	.w7(32'h3721e607),
	.w8(32'hba69e3c1),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f72d7),
	.w1(32'hba8e80dd),
	.w2(32'hba4d6216),
	.w3(32'hbaa23af4),
	.w4(32'hba33191f),
	.w5(32'hbb02d379),
	.w6(32'hba6ad4b8),
	.w7(32'hba944679),
	.w8(32'hbaa2360d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbe09f),
	.w1(32'hb91724ee),
	.w2(32'hba3c4054),
	.w3(32'hbb859b56),
	.w4(32'hbad7295a),
	.w5(32'h3ac1b43e),
	.w6(32'hbaeb5798),
	.w7(32'hbae2bd16),
	.w8(32'hba08f460),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7bac2),
	.w1(32'h3a29ae0e),
	.w2(32'h3ab9689a),
	.w3(32'h3b1bac4d),
	.w4(32'h3b42dd32),
	.w5(32'h3a6de091),
	.w6(32'h3add1364),
	.w7(32'h3b0d1d8d),
	.w8(32'hbaa5dc2d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b699e),
	.w1(32'h3a813376),
	.w2(32'h3ac882bb),
	.w3(32'h3a772700),
	.w4(32'h3ad389a1),
	.w5(32'h3a2ee729),
	.w6(32'h3a726434),
	.w7(32'h3ad4f849),
	.w8(32'h3a58124a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad13887),
	.w1(32'hbb652026),
	.w2(32'hbb6ac43c),
	.w3(32'hbb2f5271),
	.w4(32'hbb939740),
	.w5(32'hbaab4a4c),
	.w6(32'hbba86b1e),
	.w7(32'hbb973da5),
	.w8(32'hbaa99926),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1f435),
	.w1(32'h3b16f939),
	.w2(32'h3b10a92d),
	.w3(32'h3a265d14),
	.w4(32'h3878d894),
	.w5(32'hb71a5c47),
	.w6(32'h3ab13040),
	.w7(32'h39c64ebb),
	.w8(32'hbb0bef95),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73d63a9),
	.w1(32'hba8f9e6c),
	.w2(32'hb95d8ba9),
	.w3(32'h3a16c205),
	.w4(32'h3ac1c60e),
	.w5(32'hba90f2f1),
	.w6(32'hbada7b1c),
	.w7(32'hbacfc039),
	.w8(32'hbaabfe61),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2546e9),
	.w1(32'hbb1eba4c),
	.w2(32'hbb257b44),
	.w3(32'hbb5a3aeb),
	.w4(32'hbb097037),
	.w5(32'hbb433d4b),
	.w6(32'hbb581485),
	.w7(32'hbb129324),
	.w8(32'hbb63af73),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46fc79),
	.w1(32'hba75a196),
	.w2(32'hb8a44299),
	.w3(32'hbb2df70e),
	.w4(32'hbb0085ed),
	.w5(32'h3abb348c),
	.w6(32'hbb0d5a33),
	.w7(32'hbb0a1b80),
	.w8(32'h3a99cc61),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d0b19),
	.w1(32'h3aa4a65b),
	.w2(32'h39ac724b),
	.w3(32'h3a9f1f64),
	.w4(32'h3a068e18),
	.w5(32'hbb08649a),
	.w6(32'h3aadd5ad),
	.w7(32'h3a47defc),
	.w8(32'hbb002bc9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d6d32),
	.w1(32'hbb3acaaa),
	.w2(32'hbaf58ed3),
	.w3(32'hbb4a354e),
	.w4(32'hbaf58173),
	.w5(32'h3a30fe5c),
	.w6(32'hbb1eef65),
	.w7(32'hbb043394),
	.w8(32'hb949ea27),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b7b93),
	.w1(32'hb9951bca),
	.w2(32'hb98df36b),
	.w3(32'h39d949b7),
	.w4(32'h3997b5bb),
	.w5(32'hba767fa7),
	.w6(32'hb9455c7e),
	.w7(32'h3625438f),
	.w8(32'hba981a8a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a00a5),
	.w1(32'hba2d93c2),
	.w2(32'h38e922ce),
	.w3(32'hba84f27b),
	.w4(32'h39842d6d),
	.w5(32'h3aec6296),
	.w6(32'h39567a57),
	.w7(32'h3a1441fc),
	.w8(32'h3a91b1ca),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38e8d7),
	.w1(32'h3aade37a),
	.w2(32'h3a547c13),
	.w3(32'h3937ddd6),
	.w4(32'h3afe34af),
	.w5(32'hba608b28),
	.w6(32'hb9c7e12d),
	.w7(32'h39093dff),
	.w8(32'hbb07b4f4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34963f),
	.w1(32'hbb18094a),
	.w2(32'hbabc35e3),
	.w3(32'hbad49ae2),
	.w4(32'hbaaaed49),
	.w5(32'h3a1f65df),
	.w6(32'hbae430f2),
	.w7(32'hbae7b921),
	.w8(32'h3a5b9f35),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b79ba1),
	.w1(32'hb7892e58),
	.w2(32'h3a4796b0),
	.w3(32'hbaa5ae05),
	.w4(32'hbab15b91),
	.w5(32'hbb5c85f9),
	.w6(32'hb9a379d4),
	.w7(32'hb9fbc7c2),
	.w8(32'hbb4abd73),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84ae01),
	.w1(32'h3a4327b0),
	.w2(32'h38dd0453),
	.w3(32'hba0abb1b),
	.w4(32'h3a969023),
	.w5(32'hb7fd0344),
	.w6(32'hba77cdb6),
	.w7(32'hb7f8e7bd),
	.w8(32'hb9000a9d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5b559),
	.w1(32'h38e6157f),
	.w2(32'hb8c97ee7),
	.w3(32'hb8fc9d86),
	.w4(32'h3a6e7dfa),
	.w5(32'h3a6721e2),
	.w6(32'h3a130bd1),
	.w7(32'h39e4ec66),
	.w8(32'h3a5062ec),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e31e8b),
	.w1(32'h3a6fac87),
	.w2(32'h3a342d69),
	.w3(32'h3aab07ff),
	.w4(32'h3a93e28d),
	.w5(32'hb9e3f434),
	.w6(32'h3adb9eb5),
	.w7(32'h3aa26476),
	.w8(32'hba62a558),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba458afe),
	.w1(32'hba830dbb),
	.w2(32'h3600e36b),
	.w3(32'hbad4e267),
	.w4(32'hb949d6ff),
	.w5(32'h3a0f5c46),
	.w6(32'h3594c167),
	.w7(32'hba986440),
	.w8(32'hb8cc955a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ccc2d),
	.w1(32'hba352b96),
	.w2(32'hba3f2b46),
	.w3(32'h3966f78c),
	.w4(32'hb7dcc57d),
	.w5(32'hbb8b7320),
	.w6(32'hb98e9c77),
	.w7(32'hba28e1c3),
	.w8(32'hbb9e74db),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb673317),
	.w1(32'hbba09dda),
	.w2(32'hbb5fbdc0),
	.w3(32'hbba2bb59),
	.w4(32'hbb806de4),
	.w5(32'hb91d1a75),
	.w6(32'hbbb778e0),
	.w7(32'hbb886e5c),
	.w8(32'h3a0ca586),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6eb4ba),
	.w1(32'h3a5eceab),
	.w2(32'hb970cf2a),
	.w3(32'h3abb4dcd),
	.w4(32'h3ac3a856),
	.w5(32'h3a4181f3),
	.w6(32'h3b0606d4),
	.w7(32'h3ac1e175),
	.w8(32'h3a6f789f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a253050),
	.w1(32'h3a36edf6),
	.w2(32'h39e0b6c5),
	.w3(32'h3a83dd73),
	.w4(32'h3ac5b193),
	.w5(32'hb9ef791d),
	.w6(32'hb8e5f482),
	.w7(32'h3a6ba4ee),
	.w8(32'hb8bccad1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d929a0),
	.w1(32'hba26167c),
	.w2(32'hba4065df),
	.w3(32'hbab85044),
	.w4(32'hba773ce3),
	.w5(32'hba389d7f),
	.w6(32'hbaae2b1a),
	.w7(32'hb8433fb3),
	.w8(32'hb9f616fa),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34a05f),
	.w1(32'hba6e0a84),
	.w2(32'hba806700),
	.w3(32'hbac1f5af),
	.w4(32'hbadc1998),
	.w5(32'hbaf343aa),
	.w6(32'hbaa2b8ec),
	.w7(32'hba9fba2b),
	.w8(32'hba6844a5),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f61c1c),
	.w1(32'hb93ceb4c),
	.w2(32'hb9f3880b),
	.w3(32'hbabbdaa5),
	.w4(32'hba988f2c),
	.w5(32'h3a9b62da),
	.w6(32'hba17b3cf),
	.w7(32'hb9d26e01),
	.w8(32'h39e00735),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391937c5),
	.w1(32'h3a0728bd),
	.w2(32'h3a269771),
	.w3(32'h3a8d2a8e),
	.w4(32'h3919bbf2),
	.w5(32'hb8df012e),
	.w6(32'h3988de39),
	.w7(32'hba4f8ef0),
	.w8(32'h39f37cea),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84caba),
	.w1(32'h3aa1b8a6),
	.w2(32'h3a2b3f2a),
	.w3(32'h3a1c9e89),
	.w4(32'h38c605fb),
	.w5(32'hba5d3c85),
	.w6(32'h3add3975),
	.w7(32'h39f406e0),
	.w8(32'hba2b2e45),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41b380),
	.w1(32'hba83f2ad),
	.w2(32'h3adc9ecf),
	.w3(32'h3a28ed70),
	.w4(32'hb7d4e64e),
	.w5(32'h3ae09d9f),
	.w6(32'hbaae6a9a),
	.w7(32'h39691be1),
	.w8(32'h39d8b195),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule