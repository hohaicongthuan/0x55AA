module layer_10_featuremap_96(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3967e5bb),
	.w1(32'h3c071605),
	.w2(32'hbbd804cb),
	.w3(32'hba5f0a3a),
	.w4(32'hbb4b3311),
	.w5(32'hbb18c945),
	.w6(32'h39ec76e6),
	.w7(32'h3b1e43f3),
	.w8(32'h3ba8dbdf),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6736c),
	.w1(32'hb9ab473c),
	.w2(32'h3afaaf60),
	.w3(32'hbb54b2c1),
	.w4(32'hba05da80),
	.w5(32'hb7f4d03e),
	.w6(32'hba9f5fd1),
	.w7(32'h3a0791c4),
	.w8(32'h3af23397),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64ab1b),
	.w1(32'h3a16bc9e),
	.w2(32'h3b6532b6),
	.w3(32'h3a288fc6),
	.w4(32'hba751a39),
	.w5(32'hba895239),
	.w6(32'hb91448e8),
	.w7(32'hba9b60b6),
	.w8(32'h3aff19dc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab54ab8),
	.w1(32'h3b1597ef),
	.w2(32'hbb04d213),
	.w3(32'hbb091cde),
	.w4(32'h3a7b6aa5),
	.w5(32'hbb3670c2),
	.w6(32'h3b108053),
	.w7(32'h3b960e8a),
	.w8(32'hbb4dc82d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba486d13),
	.w1(32'hbb55f2d1),
	.w2(32'h3c7d8559),
	.w3(32'hbae7e2c2),
	.w4(32'h3bfcfa68),
	.w5(32'h3ae501e6),
	.w6(32'hbb0f2576),
	.w7(32'h3c144fa6),
	.w8(32'hb9a4e8aa),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1561bb),
	.w1(32'h399f2f51),
	.w2(32'h3b8acc43),
	.w3(32'hbbdcb550),
	.w4(32'h3ac1b31e),
	.w5(32'h39e3a397),
	.w6(32'h39acdfc8),
	.w7(32'h3b5ca6b6),
	.w8(32'h3b5055d4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40a1c0),
	.w1(32'hb9dd48b9),
	.w2(32'h3bc04494),
	.w3(32'h3adf0e11),
	.w4(32'h3ace47b8),
	.w5(32'h39a4456d),
	.w6(32'hbafbcc62),
	.w7(32'h3a711a7c),
	.w8(32'h3aa4d595),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399acfc9),
	.w1(32'h3a9c3e48),
	.w2(32'h39984962),
	.w3(32'hbb334609),
	.w4(32'h3a896b12),
	.w5(32'hba37a3b0),
	.w6(32'h3ad1db00),
	.w7(32'h3a83b291),
	.w8(32'h3a333c8d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9683677),
	.w1(32'hb6809047),
	.w2(32'hbaa35e10),
	.w3(32'hba1ea886),
	.w4(32'hb6adfe28),
	.w5(32'h3a03440a),
	.w6(32'hb9d3d385),
	.w7(32'hba8ad4f9),
	.w8(32'hb8c1c8b3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39428bc7),
	.w1(32'h3a3d0f99),
	.w2(32'h39a3bb87),
	.w3(32'h3a9fd3e6),
	.w4(32'h3a7db139),
	.w5(32'hb9705173),
	.w6(32'h390fc2ab),
	.w7(32'hbaaef0d5),
	.w8(32'hb9c99f00),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2e58d),
	.w1(32'h3a594ac8),
	.w2(32'hb8c1ef23),
	.w3(32'h3b0c25b5),
	.w4(32'hbadbf2d8),
	.w5(32'hba4bc5fd),
	.w6(32'h3a953962),
	.w7(32'h3b2ebffe),
	.w8(32'hb9e66458),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1adf01),
	.w1(32'hbabdf4bb),
	.w2(32'hbb3a1bf4),
	.w3(32'hba19cea4),
	.w4(32'hba0a2c51),
	.w5(32'hbbc41c00),
	.w6(32'h3b978ae3),
	.w7(32'h3b73bd1a),
	.w8(32'hbb4b07db),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e2f75),
	.w1(32'hbb007543),
	.w2(32'hb9c640bd),
	.w3(32'h390cb75f),
	.w4(32'hba0509d8),
	.w5(32'hba9d1508),
	.w6(32'hbb0f2f48),
	.w7(32'hbb2ba3f7),
	.w8(32'hba574bc7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdc265),
	.w1(32'h3ba785fd),
	.w2(32'hb98df38b),
	.w3(32'hbaede7e0),
	.w4(32'h3b9f8289),
	.w5(32'h3ba1ce24),
	.w6(32'h3be12713),
	.w7(32'h3b61d14f),
	.w8(32'h3ba52356),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50a37f),
	.w1(32'hbb96d4e2),
	.w2(32'hbbb995bc),
	.w3(32'h3b2c1bfe),
	.w4(32'h3bb89131),
	.w5(32'hbba1d41c),
	.w6(32'h39fcf341),
	.w7(32'h3c0d8815),
	.w8(32'hbbfd80d8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02d248),
	.w1(32'hba1dce51),
	.w2(32'hbaa93e26),
	.w3(32'hbbebfa5c),
	.w4(32'hba1e44bb),
	.w5(32'hba5aff1a),
	.w6(32'hba4ced06),
	.w7(32'hba33b82f),
	.w8(32'hba2d08b5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31f7da),
	.w1(32'h3b02bdbb),
	.w2(32'h3bb2699a),
	.w3(32'h39dfe0cb),
	.w4(32'h3af408cc),
	.w5(32'h3b507729),
	.w6(32'h39efcbe0),
	.w7(32'h3b3d5fa6),
	.w8(32'h3b8873d1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7079ff),
	.w1(32'h3a86b48e),
	.w2(32'h3ab2139b),
	.w3(32'h3a81f987),
	.w4(32'h3ae49b3c),
	.w5(32'hb9cc1b4c),
	.w6(32'hbabc7021),
	.w7(32'h3a573ab3),
	.w8(32'h3a8639cb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0213c2),
	.w1(32'hba492ae6),
	.w2(32'hba87fbdb),
	.w3(32'h3a8a76ec),
	.w4(32'h39ec54ce),
	.w5(32'hbacc291f),
	.w6(32'hba9c1325),
	.w7(32'hba87bdb2),
	.w8(32'hba004585),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70791e),
	.w1(32'hba64d1eb),
	.w2(32'hbab64d4e),
	.w3(32'hba0bdea9),
	.w4(32'hba71138b),
	.w5(32'hba851fab),
	.w6(32'hb8e195e9),
	.w7(32'hba3d7bcd),
	.w8(32'h399eedff),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34ddcd),
	.w1(32'hbaad02a7),
	.w2(32'hbb518e0d),
	.w3(32'h3a987964),
	.w4(32'hba66265a),
	.w5(32'hba4c6495),
	.w6(32'h3ab8958d),
	.w7(32'h39938081),
	.w8(32'h3b5bbbc1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04ce17),
	.w1(32'hbaf22092),
	.w2(32'h3b85d4ab),
	.w3(32'h3ae7e207),
	.w4(32'hbbcfb6e1),
	.w5(32'hbbed74a3),
	.w6(32'hbc02a07c),
	.w7(32'hbc2b180a),
	.w8(32'h3b5b67e3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b1131),
	.w1(32'h391c0a88),
	.w2(32'hb9e953f7),
	.w3(32'hbc3e25e9),
	.w4(32'h3af23906),
	.w5(32'h3a949fc1),
	.w6(32'hbaecb47c),
	.w7(32'hb7cdf418),
	.w8(32'hbab1b500),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b084ae8),
	.w1(32'h3a4b1fe2),
	.w2(32'hb9e9116d),
	.w3(32'h3ad182cb),
	.w4(32'h39e37721),
	.w5(32'hb94b8069),
	.w6(32'h3a5488df),
	.w7(32'h393c194f),
	.w8(32'h3a179d75),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33a08d),
	.w1(32'hbab04d6b),
	.w2(32'hb98450ba),
	.w3(32'hba44d310),
	.w4(32'hba299a94),
	.w5(32'hb9be0051),
	.w6(32'hbab5f893),
	.w7(32'h3ab3a5a9),
	.w8(32'h3988d00c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa288d),
	.w1(32'hbb22a12a),
	.w2(32'hbaa13796),
	.w3(32'h3a3a8b01),
	.w4(32'hbad0fb9f),
	.w5(32'hba0591d1),
	.w6(32'hbbc1956e),
	.w7(32'hbb8ee586),
	.w8(32'hbb30e1e1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae90c3e),
	.w1(32'hbad7447e),
	.w2(32'hbaecc1a6),
	.w3(32'h3a3b48cb),
	.w4(32'hbaad7b34),
	.w5(32'hbaa1051f),
	.w6(32'hba103af2),
	.w7(32'hba35d2eb),
	.w8(32'h3925f8ae),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89a3915),
	.w1(32'hbaa414aa),
	.w2(32'hbb29431c),
	.w3(32'hb97e5add),
	.w4(32'hbb3b0a54),
	.w5(32'hbb5f7e03),
	.w6(32'hbb838a27),
	.w7(32'hba138d6e),
	.w8(32'hbb2cbc25),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8faf97),
	.w1(32'h3a673421),
	.w2(32'hbb943c5f),
	.w3(32'hbb3224f0),
	.w4(32'h3b140e40),
	.w5(32'hbb848c96),
	.w6(32'h3b08dbf4),
	.w7(32'hbaeda056),
	.w8(32'h3af384b3),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eab800),
	.w1(32'h3b4c4ab5),
	.w2(32'h3b187eed),
	.w3(32'h3929aaa7),
	.w4(32'h3b3abc4d),
	.w5(32'h3b8fe1c1),
	.w6(32'h3ac18995),
	.w7(32'h3b24af22),
	.w8(32'h3b73294a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a8ed9),
	.w1(32'hba13d247),
	.w2(32'hbab8477c),
	.w3(32'h3b2af66a),
	.w4(32'h367240d1),
	.w5(32'h360e1de8),
	.w6(32'h39dcc539),
	.w7(32'hb9db1661),
	.w8(32'h3aafe674),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f93608),
	.w1(32'hbac314f6),
	.w2(32'hba9f5240),
	.w3(32'h3ab116b1),
	.w4(32'hba89a728),
	.w5(32'hbaff71c4),
	.w6(32'hba6a1b75),
	.w7(32'hba02be1e),
	.w8(32'hb98e1120),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62047b),
	.w1(32'hbb596db8),
	.w2(32'hbb4523ab),
	.w3(32'hbab21839),
	.w4(32'hbb790243),
	.w5(32'hb92035e1),
	.w6(32'hbbe10398),
	.w7(32'hbb8af32d),
	.w8(32'h3aa9f325),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cb4d1),
	.w1(32'h3996a22b),
	.w2(32'hbb8ed0b1),
	.w3(32'h3b53f932),
	.w4(32'hbab8bc4b),
	.w5(32'hbbc4da05),
	.w6(32'h3b9028f7),
	.w7(32'hbbcd02ba),
	.w8(32'hbbedd20c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82cd8c),
	.w1(32'h3ace3b61),
	.w2(32'hbabbf3ca),
	.w3(32'hbb28cdf2),
	.w4(32'hba3bd099),
	.w5(32'hbb4beeaf),
	.w6(32'h3a32d59a),
	.w7(32'hb93fd568),
	.w8(32'h3a99141b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1f788),
	.w1(32'hbada380b),
	.w2(32'hbb64166b),
	.w3(32'h3ac77259),
	.w4(32'hbae21683),
	.w5(32'hbb5a8b3f),
	.w6(32'hba648e32),
	.w7(32'h38cf440e),
	.w8(32'h39ceb888),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3c669),
	.w1(32'hbad6f031),
	.w2(32'h3b05f6d7),
	.w3(32'hbb06b4b5),
	.w4(32'h39fea45e),
	.w5(32'hbaaa723c),
	.w6(32'hbb68bc8e),
	.w7(32'h3a72a28e),
	.w8(32'h39c66c48),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898895a),
	.w1(32'h3a16c50b),
	.w2(32'h3b20e136),
	.w3(32'h386b6a77),
	.w4(32'h3a669a41),
	.w5(32'h3a08aec3),
	.w6(32'hbaf0e181),
	.w7(32'hba0296d5),
	.w8(32'h3a54a498),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2309ba),
	.w1(32'h3a087d65),
	.w2(32'h385d908b),
	.w3(32'h38864499),
	.w4(32'hb73ab7a4),
	.w5(32'h39bc0202),
	.w6(32'hb887664a),
	.w7(32'h3a127871),
	.w8(32'h3a461e58),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ae508),
	.w1(32'h3a3c0457),
	.w2(32'h3ad45e6c),
	.w3(32'hb7ab47db),
	.w4(32'h3a712655),
	.w5(32'h39062032),
	.w6(32'hb9ac3ec7),
	.w7(32'h395fe2fe),
	.w8(32'h3987ae6e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39105124),
	.w1(32'h3aefa3fe),
	.w2(32'h3af82431),
	.w3(32'hba863cb2),
	.w4(32'h3b10325f),
	.w5(32'h3b59bebd),
	.w6(32'h3a347cb7),
	.w7(32'h3b6215f9),
	.w8(32'h3acc6343),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c09ea),
	.w1(32'h3b06f89b),
	.w2(32'hba79b023),
	.w3(32'h38c27d2c),
	.w4(32'h3aae0e7c),
	.w5(32'h398e297c),
	.w6(32'h39a35dec),
	.w7(32'h3b37c946),
	.w8(32'h3a898a11),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a134606),
	.w1(32'hbb20d044),
	.w2(32'hbacb05de),
	.w3(32'h3a7fb6d4),
	.w4(32'hba961040),
	.w5(32'hbad3f8fd),
	.w6(32'hbb14c126),
	.w7(32'hbb2ae12e),
	.w8(32'hbac0cf62),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacab0af),
	.w1(32'h3b690a1a),
	.w2(32'h3b3faf9d),
	.w3(32'hba9a1cb6),
	.w4(32'h3b8e4174),
	.w5(32'h3b1e1eb8),
	.w6(32'h3b44a508),
	.w7(32'hb9ece422),
	.w8(32'h3a1d9ae8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad918dc),
	.w1(32'h3b979346),
	.w2(32'hbb35a3f7),
	.w3(32'h39ffc146),
	.w4(32'h3b94d713),
	.w5(32'h3b687c1d),
	.w6(32'h3b1026bd),
	.w7(32'hbb71744b),
	.w8(32'h3aadac6b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954a1d3),
	.w1(32'hb98454eb),
	.w2(32'h3c035879),
	.w3(32'hbb2a4658),
	.w4(32'h3ab42fe6),
	.w5(32'h3a73db3c),
	.w6(32'hbb4998da),
	.w7(32'hbb5afdc8),
	.w8(32'h3aed8f1f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e36ad),
	.w1(32'hbb6689b3),
	.w2(32'hbbaff3e6),
	.w3(32'hbbfdaec0),
	.w4(32'h3b20a2ad),
	.w5(32'hbb824a72),
	.w6(32'h3b8a7a67),
	.w7(32'h3bbb660d),
	.w8(32'hbbba70ad),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d2ece),
	.w1(32'h3b8b81e4),
	.w2(32'hb95e4756),
	.w3(32'hbaa06c36),
	.w4(32'h3b6722c2),
	.w5(32'h39c6c287),
	.w6(32'h3b22993d),
	.w7(32'h3b610263),
	.w8(32'h3b332647),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4684e8),
	.w1(32'hbac2e481),
	.w2(32'hbae3aed2),
	.w3(32'h3b635c27),
	.w4(32'hba5bb62d),
	.w5(32'hbb019dbe),
	.w6(32'hba89b916),
	.w7(32'hbad24abc),
	.w8(32'hba22f0b8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba763f8e),
	.w1(32'h38ff5564),
	.w2(32'hb991febc),
	.w3(32'hbaa71ca1),
	.w4(32'h399274d4),
	.w5(32'h396a47ce),
	.w6(32'h3ab30ff7),
	.w7(32'h3a03935b),
	.w8(32'hb8a74e42),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba728e8e),
	.w1(32'hbaec16b8),
	.w2(32'hb85feec1),
	.w3(32'hba912b65),
	.w4(32'h3abdf33b),
	.w5(32'h3ab20604),
	.w6(32'hb8ae92a4),
	.w7(32'hba7edb08),
	.w8(32'hbacd430f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a62bb),
	.w1(32'hbb4c9bad),
	.w2(32'h3b11f98d),
	.w3(32'hba5e5b4f),
	.w4(32'hbc262f16),
	.w5(32'hbb72cbdc),
	.w6(32'h3a7525c6),
	.w7(32'hbad7e2cb),
	.w8(32'hbba10c1a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84a261),
	.w1(32'hba118840),
	.w2(32'h3ab946d5),
	.w3(32'h3bbc8248),
	.w4(32'hba9f7d67),
	.w5(32'hbaa6d1b4),
	.w6(32'hba703b44),
	.w7(32'h3b055786),
	.w8(32'h3b1736ec),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9d441),
	.w1(32'hba4661d1),
	.w2(32'h3c585166),
	.w3(32'h3a8ba404),
	.w4(32'h3bc8b330),
	.w5(32'hbb695186),
	.w6(32'hbb23156b),
	.w7(32'h3bedce59),
	.w8(32'h3b443e2a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc0d45),
	.w1(32'hbb6a708d),
	.w2(32'hba9ddea6),
	.w3(32'hbbb54c66),
	.w4(32'hbb215f07),
	.w5(32'hbafd8d90),
	.w6(32'hbb68f90d),
	.w7(32'hbb081038),
	.w8(32'hbabd1c2b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01efef),
	.w1(32'hba6ab16f),
	.w2(32'hba66fb56),
	.w3(32'hba88d7a1),
	.w4(32'hba6daedf),
	.w5(32'hbac5189b),
	.w6(32'hbb950b2e),
	.w7(32'hb6d4cce4),
	.w8(32'hba6700b9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14a642),
	.w1(32'hbb824b61),
	.w2(32'hbacdfec8),
	.w3(32'hbb04f7d4),
	.w4(32'hbaf253c0),
	.w5(32'h3b370c22),
	.w6(32'hbb6da886),
	.w7(32'hbb9f16c5),
	.w8(32'h3b2a9dec),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8930c6),
	.w1(32'hbbbbfeab),
	.w2(32'h3ca172f7),
	.w3(32'h3af5b524),
	.w4(32'h3c051d0e),
	.w5(32'h3b28537b),
	.w6(32'hbb57bd6d),
	.w7(32'h3c1f58f5),
	.w8(32'h3be85f8e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c58c4),
	.w1(32'h3acc07bb),
	.w2(32'h3aa1237f),
	.w3(32'hbba920cb),
	.w4(32'hb93c0359),
	.w5(32'h39d1c270),
	.w6(32'h3acf5253),
	.w7(32'h3ade5767),
	.w8(32'h3a10dffc),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7cda2),
	.w1(32'h3a37835d),
	.w2(32'hba530fe8),
	.w3(32'hbabd26e7),
	.w4(32'hb97a01f6),
	.w5(32'hb5e32d9a),
	.w6(32'h397b0abb),
	.w7(32'hb8bdac6c),
	.w8(32'h3a440898),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952b15a),
	.w1(32'hb92403da),
	.w2(32'h3a3a696e),
	.w3(32'hb9c1cdf6),
	.w4(32'h39377ab2),
	.w5(32'hba23ba1e),
	.w6(32'hba82ada0),
	.w7(32'hb9c79a99),
	.w8(32'hb8485f54),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fed0f),
	.w1(32'h3a32e49e),
	.w2(32'hbb11efef),
	.w3(32'hba8f9680),
	.w4(32'hb9e43ef1),
	.w5(32'h3a11b512),
	.w6(32'h384fa511),
	.w7(32'hbac0aceb),
	.w8(32'h3a8cfac0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bf3a1),
	.w1(32'h3b659ab9),
	.w2(32'h396f7e43),
	.w3(32'hba07f077),
	.w4(32'hbb18677c),
	.w5(32'h3b2257b7),
	.w6(32'hba769a51),
	.w7(32'h390e2dba),
	.w8(32'h3b665900),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5ca03),
	.w1(32'h3b10d190),
	.w2(32'h3adc7f79),
	.w3(32'h3bf85f8e),
	.w4(32'h3b217e6f),
	.w5(32'h3a5cab41),
	.w6(32'h3af97e7d),
	.w7(32'hb90f07d2),
	.w8(32'h398ffa25),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a298c65),
	.w1(32'hbb5b8c7e),
	.w2(32'h3a332d6d),
	.w3(32'hb8e70da4),
	.w4(32'hbadeb79a),
	.w5(32'h39203bcf),
	.w6(32'hbb1e6101),
	.w7(32'hba0df9c7),
	.w8(32'h3b1d77aa),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadeb50),
	.w1(32'hbac48aab),
	.w2(32'h3c7f79c5),
	.w3(32'hb98ae432),
	.w4(32'h3bb47685),
	.w5(32'h39690a01),
	.w6(32'hbadd6849),
	.w7(32'h3ae20e65),
	.w8(32'h3b4dfaa9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab6030),
	.w1(32'hb9db9c58),
	.w2(32'h3b990a81),
	.w3(32'hbc0f4514),
	.w4(32'h3a731628),
	.w5(32'h3b67ff86),
	.w6(32'hbb4436a7),
	.w7(32'h3aa53c05),
	.w8(32'h3a09f673),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab450d6),
	.w1(32'h3a7942a3),
	.w2(32'h3a2e32ba),
	.w3(32'h3a59627d),
	.w4(32'h3b53f463),
	.w5(32'h3af648db),
	.w6(32'h3984a9d4),
	.w7(32'h3b25ffb3),
	.w8(32'hb994498e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e33aa),
	.w1(32'hbad76784),
	.w2(32'hb9963f92),
	.w3(32'h3997b69e),
	.w4(32'hb9a7af3b),
	.w5(32'h398a9a5b),
	.w6(32'hbaa7893d),
	.w7(32'hb90c73c9),
	.w8(32'h3a73b84d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904d948),
	.w1(32'h39fd14a3),
	.w2(32'h3c2b4893),
	.w3(32'h3a123259),
	.w4(32'h3c2a5fbf),
	.w5(32'h3b8a4fd6),
	.w6(32'h3b090019),
	.w7(32'h3b979b0b),
	.w8(32'h3b96fcc8),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63a0c2),
	.w1(32'h3b098d55),
	.w2(32'h39f78b91),
	.w3(32'hbb990355),
	.w4(32'h3a9f5345),
	.w5(32'hba10628d),
	.w6(32'h3a4425de),
	.w7(32'h3a3c92e8),
	.w8(32'h3a0fba7b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92e3f5),
	.w1(32'hb9eefeb9),
	.w2(32'h3a7b6979),
	.w3(32'h3a09b35c),
	.w4(32'h3a928549),
	.w5(32'h3aa9d1f6),
	.w6(32'hba968744),
	.w7(32'h3a31ceeb),
	.w8(32'h3afdc253),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b9134),
	.w1(32'h3a0964dc),
	.w2(32'hb9a440cd),
	.w3(32'hba794786),
	.w4(32'h38ef8adf),
	.w5(32'h39873756),
	.w6(32'hb9a708b8),
	.w7(32'h39936330),
	.w8(32'h3a3a6603),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3975e35b),
	.w1(32'hbad6b830),
	.w2(32'hbb09ce9d),
	.w3(32'hb8a0427c),
	.w4(32'hbacbd140),
	.w5(32'hbad29845),
	.w6(32'hb9111f56),
	.w7(32'hb9b1c8fe),
	.w8(32'h3a86d481),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a15093),
	.w1(32'h3a0b56f4),
	.w2(32'h3a7820b6),
	.w3(32'hba7c24ac),
	.w4(32'hba3e43e1),
	.w5(32'hb99f73e2),
	.w6(32'h3a242ceb),
	.w7(32'h3b516d22),
	.w8(32'h3a801cde),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb794ecbd),
	.w1(32'hbb7b5b2f),
	.w2(32'h3b1e3957),
	.w3(32'h3a7e778d),
	.w4(32'hbab1ecba),
	.w5(32'h3a275355),
	.w6(32'hbb9a7c59),
	.w7(32'hb9a3eee4),
	.w8(32'hbbb4245c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65c2fd),
	.w1(32'h3aeb676d),
	.w2(32'h354e7851),
	.w3(32'h3b0edba9),
	.w4(32'h3b239854),
	.w5(32'h3a91930e),
	.w6(32'h3b2a094c),
	.w7(32'h3a35a5df),
	.w8(32'h3aacb109),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a181bab),
	.w1(32'h3b092725),
	.w2(32'hba855cd2),
	.w3(32'h3a629f9f),
	.w4(32'h3aaaec89),
	.w5(32'h3a97aca2),
	.w6(32'hba7ded8a),
	.w7(32'hb9ca05a4),
	.w8(32'hba9bcb3e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed7c2d),
	.w1(32'hbbc81bf5),
	.w2(32'hba268156),
	.w3(32'h3b424ea5),
	.w4(32'hbb72fd9f),
	.w5(32'hbac6275d),
	.w6(32'hbbd937c1),
	.w7(32'hbbbb66e4),
	.w8(32'hbb1f5b2b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9430edb),
	.w1(32'hba5dca04),
	.w2(32'hbb2803c7),
	.w3(32'hb9935c3c),
	.w4(32'h3a82a614),
	.w5(32'h399e125b),
	.w6(32'h3a7a9e6f),
	.w7(32'hba924a56),
	.w8(32'h3a0a5803),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9381b09),
	.w1(32'h3a96d603),
	.w2(32'h3a302d3b),
	.w3(32'h3a9c8647),
	.w4(32'h3b0ccd2d),
	.w5(32'h3a49113a),
	.w6(32'h3a334b8f),
	.w7(32'h3b18839d),
	.w8(32'h3a1f5e7c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3929acab),
	.w1(32'hb97726a7),
	.w2(32'h3b260a21),
	.w3(32'hb9439dd3),
	.w4(32'hba592f50),
	.w5(32'h3b1a2ba3),
	.w6(32'h3b09ea51),
	.w7(32'h3b203ebd),
	.w8(32'h3aef24ca),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54dd6f),
	.w1(32'h39a6a3d5),
	.w2(32'hb8973786),
	.w3(32'h3a18264d),
	.w4(32'hb87fdb7c),
	.w5(32'hb80f5133),
	.w6(32'hba9c61fa),
	.w7(32'h3add6a1b),
	.w8(32'h3ae874f8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f5f525),
	.w1(32'h3b1ab8e9),
	.w2(32'h3b36002d),
	.w3(32'h3a74c167),
	.w4(32'hba28a7f9),
	.w5(32'hba3cab6b),
	.w6(32'h3a6d9990),
	.w7(32'h3ac61cfa),
	.w8(32'h3a83c799),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6f58a),
	.w1(32'h3b117848),
	.w2(32'hbb3f81d4),
	.w3(32'hbb008a5e),
	.w4(32'hb9d76292),
	.w5(32'hb9bfd990),
	.w6(32'h3b368604),
	.w7(32'h3a5289a6),
	.w8(32'hbb27007f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4471e3),
	.w1(32'hbab1f84e),
	.w2(32'h3b7bfaeb),
	.w3(32'h3a3041b9),
	.w4(32'hba256f19),
	.w5(32'h3b0ddd8d),
	.w6(32'hbb3197b9),
	.w7(32'hb9b843ef),
	.w8(32'h3ae7a256),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35405b),
	.w1(32'h3a6da1f8),
	.w2(32'hb9888d91),
	.w3(32'h3a4f6658),
	.w4(32'h3b2f4f4b),
	.w5(32'h3ae32871),
	.w6(32'h3b1d4407),
	.w7(32'h3b378684),
	.w8(32'h3a8d9c68),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9b372),
	.w1(32'hba85430d),
	.w2(32'hbabc60c8),
	.w3(32'h3b4367f6),
	.w4(32'hb9d2a6cd),
	.w5(32'h398cd0d6),
	.w6(32'h39b65c11),
	.w7(32'hb9a12561),
	.w8(32'h3ac08cb0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a881d10),
	.w1(32'hbb07573c),
	.w2(32'hbaab8539),
	.w3(32'h3a963a72),
	.w4(32'hbabcff2f),
	.w5(32'hbac7801e),
	.w6(32'hbadf53da),
	.w7(32'hbabbabc3),
	.w8(32'hba21fc2b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdfd6f),
	.w1(32'hbabe6eec),
	.w2(32'hbb34411c),
	.w3(32'hba2eb4db),
	.w4(32'hba74fb15),
	.w5(32'hbabcad86),
	.w6(32'hb8d2e12f),
	.w7(32'hba180aa5),
	.w8(32'h3a842c19),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954a64c),
	.w1(32'hba28c60f),
	.w2(32'hba1b86aa),
	.w3(32'h3a13f1c8),
	.w4(32'hba9924a1),
	.w5(32'hb923beb5),
	.w6(32'h39029050),
	.w7(32'h397e2a4b),
	.w8(32'h3adb0247),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d72b8c),
	.w1(32'h397c63c0),
	.w2(32'h3aa793dd),
	.w3(32'h3a6cb01f),
	.w4(32'h3b3c97f9),
	.w5(32'h3afdd9c3),
	.w6(32'hba0f0350),
	.w7(32'hbaa9bcc7),
	.w8(32'h3accf9a2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ca0eb),
	.w1(32'h39936c55),
	.w2(32'h3ace3678),
	.w3(32'h3b13b355),
	.w4(32'hbb08c11b),
	.w5(32'hb9bc7ee4),
	.w6(32'hb9061842),
	.w7(32'h3b0e57b8),
	.w8(32'h3b1d7b93),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb851f1b4),
	.w1(32'h395907de),
	.w2(32'hbadaddb4),
	.w3(32'h3a3042ea),
	.w4(32'h3adfac35),
	.w5(32'hbaac1f7a),
	.w6(32'h3a6ae9e3),
	.w7(32'h3964daf7),
	.w8(32'hb9365aa6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4d88f),
	.w1(32'h3b11b52a),
	.w2(32'h3b29dbe4),
	.w3(32'hbaded0be),
	.w4(32'hba102969),
	.w5(32'hbac49fd0),
	.w6(32'hba290de1),
	.w7(32'hb946a5bc),
	.w8(32'h3ac93021),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33730b),
	.w1(32'hba840ea0),
	.w2(32'h3c4132a6),
	.w3(32'hba8bd8e3),
	.w4(32'hb8b2a9ce),
	.w5(32'h3afc68c0),
	.w6(32'hbb1389c3),
	.w7(32'h3b2d5827),
	.w8(32'h3b17f7fb),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8ec1d),
	.w1(32'hbb337bfc),
	.w2(32'hba465d50),
	.w3(32'hbb0e44cc),
	.w4(32'hba8dcc58),
	.w5(32'h3ad13aff),
	.w6(32'hbb780abe),
	.w7(32'hba424ee9),
	.w8(32'hba9da7c7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a994532),
	.w1(32'hbafebdd5),
	.w2(32'hbb3a44f4),
	.w3(32'h3afeb03b),
	.w4(32'hbb8e843b),
	.w5(32'hbb07728c),
	.w6(32'hbb5dad96),
	.w7(32'hba4e0411),
	.w8(32'hbb8a4648),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcee63),
	.w1(32'h3a92e139),
	.w2(32'h3b6125f8),
	.w3(32'hbb563199),
	.w4(32'h3978fe97),
	.w5(32'h3a872d6d),
	.w6(32'h3ae59dae),
	.w7(32'h3b086301),
	.w8(32'h3b16c659),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44ef95),
	.w1(32'h3a5e2c91),
	.w2(32'h39b9a9d9),
	.w3(32'hb9d68b51),
	.w4(32'hba2c3007),
	.w5(32'hba956ec5),
	.w6(32'hbad02013),
	.w7(32'h3ace44fc),
	.w8(32'h3a9bdca7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce0d5a),
	.w1(32'hbc6665cc),
	.w2(32'h3bf5e027),
	.w3(32'h3ada9e1e),
	.w4(32'h3a05ea8b),
	.w5(32'hbbc6ac29),
	.w6(32'hbc1a0197),
	.w7(32'hbc00dc9d),
	.w8(32'hba9a6b70),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb783432),
	.w1(32'hbb1f3dee),
	.w2(32'h3d2a5e9e),
	.w3(32'hbba9b17a),
	.w4(32'hbb5fe378),
	.w5(32'h3ba3914a),
	.w6(32'hbbfa422a),
	.w7(32'h3856153d),
	.w8(32'h3a65b160),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eda19),
	.w1(32'h3b3a9a35),
	.w2(32'h3a04eaa4),
	.w3(32'hbc524cc3),
	.w4(32'h3b866bf6),
	.w5(32'h3b02d8a0),
	.w6(32'h3b82d169),
	.w7(32'h3aa34a51),
	.w8(32'h3b0d0033),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78c918),
	.w1(32'hbb0bf676),
	.w2(32'h3a0b23d9),
	.w3(32'h3aa2f1f4),
	.w4(32'h39eba261),
	.w5(32'h394ae826),
	.w6(32'hbaa14b8b),
	.w7(32'h3a1f7e5a),
	.w8(32'h3a85e742),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a199efd),
	.w1(32'h3ac62c74),
	.w2(32'h38ccb09c),
	.w3(32'hba0ebad9),
	.w4(32'h3ac899e5),
	.w5(32'h3a734db0),
	.w6(32'h3b1775ba),
	.w7(32'h39f0d80f),
	.w8(32'h3a5eb634),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c56cd6),
	.w1(32'hba9afd15),
	.w2(32'hbb0b7ef3),
	.w3(32'h3a2743ef),
	.w4(32'hba7ff41c),
	.w5(32'hba2c95c1),
	.w6(32'hbaa0cbe3),
	.w7(32'hbaa72e43),
	.w8(32'hb7ee7bcd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39591853),
	.w1(32'h3b166d15),
	.w2(32'h3b19649c),
	.w3(32'h3a8fdd00),
	.w4(32'hbae75b41),
	.w5(32'hbab4c35b),
	.w6(32'h3ac9b036),
	.w7(32'h39af6c1e),
	.w8(32'h3a93a8a4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad1a12),
	.w1(32'hbab2461b),
	.w2(32'hbafd6639),
	.w3(32'hbacb9de5),
	.w4(32'hbaca124f),
	.w5(32'h3a47bf6c),
	.w6(32'h3a47cbaf),
	.w7(32'h3936df67),
	.w8(32'h3b5adc90),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e868b),
	.w1(32'h3ac53ffb),
	.w2(32'h3a1aaa58),
	.w3(32'h3b38f4b2),
	.w4(32'h3b0bceee),
	.w5(32'h3aa4e090),
	.w6(32'h3b0a8e6b),
	.w7(32'h3a399f55),
	.w8(32'h3aaa5c9b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c9e92),
	.w1(32'h3b4bbf9d),
	.w2(32'h3b0721a7),
	.w3(32'h3a363114),
	.w4(32'h3b7eec34),
	.w5(32'h3b72c64a),
	.w6(32'h3a1d78f5),
	.w7(32'hbaaad6b5),
	.w8(32'h3b22fa50),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19c75a),
	.w1(32'hbaca68a7),
	.w2(32'hbb14673a),
	.w3(32'h3b26740e),
	.w4(32'hbb51a9b0),
	.w5(32'hbb1aacd5),
	.w6(32'hba105315),
	.w7(32'hba9b3b04),
	.w8(32'hba2d4ad6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab04db),
	.w1(32'h3afb9364),
	.w2(32'hbbcca1d4),
	.w3(32'h3a2d8809),
	.w4(32'hbb49fdeb),
	.w5(32'hb992408d),
	.w6(32'hbb4930ff),
	.w7(32'hbb9517b6),
	.w8(32'h3a5a990e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a42f5),
	.w1(32'hba88ab81),
	.w2(32'hbad69d8c),
	.w3(32'h3b80a241),
	.w4(32'hbad32cc1),
	.w5(32'hbadee6cc),
	.w6(32'hba481259),
	.w7(32'h3a36efae),
	.w8(32'hb7fb9ff9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58c215),
	.w1(32'h3af4b47b),
	.w2(32'h3836893f),
	.w3(32'h3a3af2d8),
	.w4(32'h398dba3d),
	.w5(32'h3a4f5b63),
	.w6(32'h3af452e7),
	.w7(32'h39c88c5f),
	.w8(32'hb974c367),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0324ab),
	.w1(32'hbb813a26),
	.w2(32'hbbcbe3b7),
	.w3(32'hba480df5),
	.w4(32'hbb9a0d69),
	.w5(32'hbb88baec),
	.w6(32'hbb7d7082),
	.w7(32'hbb71d28c),
	.w8(32'hba8b570d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cabe2),
	.w1(32'h3b038bf0),
	.w2(32'h39c9600d),
	.w3(32'hbaeb0169),
	.w4(32'h3b3ae101),
	.w5(32'h3aca647e),
	.w6(32'h3b3f955e),
	.w7(32'h3a5f9fe6),
	.w8(32'h3ad7e707),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30b2fa),
	.w1(32'h3a9e6959),
	.w2(32'h3a8faa58),
	.w3(32'h3a81ad4d),
	.w4(32'h3ac6b389),
	.w5(32'h3a3664bf),
	.w6(32'h3a4c8b1e),
	.w7(32'h3ab43916),
	.w8(32'h3abad54d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a285c7c),
	.w1(32'h3abe1337),
	.w2(32'h3a95615d),
	.w3(32'h39cd161c),
	.w4(32'h3ab39a2e),
	.w5(32'h39dffca1),
	.w6(32'h3ab438e1),
	.w7(32'h3b085856),
	.w8(32'h3ab9303e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a328b60),
	.w1(32'h3be73bc6),
	.w2(32'h3c15ae79),
	.w3(32'h3a8acb1c),
	.w4(32'h3b6831be),
	.w5(32'h3b2b355a),
	.w6(32'hbaee3330),
	.w7(32'hbb3a849f),
	.w8(32'h3c0a3820),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba015f9),
	.w1(32'hbb88adac),
	.w2(32'hb9b936fd),
	.w3(32'hbbd47ae3),
	.w4(32'hbb0105a4),
	.w5(32'hbc036ab6),
	.w6(32'hbb62575a),
	.w7(32'hbbc2fb03),
	.w8(32'hbb4b995b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b76b7),
	.w1(32'hb9b5d464),
	.w2(32'hbaf64b86),
	.w3(32'hbb82b8c7),
	.w4(32'hba826257),
	.w5(32'hbb5513fd),
	.w6(32'hb9866991),
	.w7(32'h3ab9d249),
	.w8(32'h3a2f7067),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edb95d),
	.w1(32'h3ae6695c),
	.w2(32'hba9e1bdf),
	.w3(32'h379637c6),
	.w4(32'hbacad109),
	.w5(32'hba9e4003),
	.w6(32'h3a88c04c),
	.w7(32'h3a04b72e),
	.w8(32'h3a1c71bf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a377031),
	.w1(32'h39db3acc),
	.w2(32'hb9a99b91),
	.w3(32'h3a658465),
	.w4(32'hb8bff525),
	.w5(32'h38eb9680),
	.w6(32'h3a009743),
	.w7(32'hb8ff9d87),
	.w8(32'h3a0af5e7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38e24f),
	.w1(32'h3bc62a79),
	.w2(32'h3ce4837f),
	.w3(32'hba561a16),
	.w4(32'h3bd5f516),
	.w5(32'h3c468bab),
	.w6(32'hbbe4ebe8),
	.w7(32'hba2e6ff3),
	.w8(32'h3c1aacf8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13601f),
	.w1(32'hba2fb3b3),
	.w2(32'h3ba807bb),
	.w3(32'hbbf93453),
	.w4(32'hba4c8b74),
	.w5(32'h3a4356a6),
	.w6(32'hb83b70d9),
	.w7(32'h3b0eb2ca),
	.w8(32'h3b13eb9b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bf6da),
	.w1(32'hba58d780),
	.w2(32'hbb0580ff),
	.w3(32'h3a041cec),
	.w4(32'hba2dd8e4),
	.w5(32'h399ef43e),
	.w6(32'h3a189a6c),
	.w7(32'hb9c5a44d),
	.w8(32'h3abaf541),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e8515),
	.w1(32'h374c0600),
	.w2(32'h36f7bef4),
	.w3(32'h3ae0553c),
	.w4(32'h36989d99),
	.w5(32'hb6337bd0),
	.w6(32'h36db91a6),
	.w7(32'h3603f53b),
	.w8(32'h371b6b5f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a9ea5e),
	.w1(32'hb8b0a5c4),
	.w2(32'hb907ee77),
	.w3(32'h384c312a),
	.w4(32'hb6b86086),
	.w5(32'hb950c9ce),
	.w6(32'hb6f8bd0c),
	.w7(32'hb7fcd1c5),
	.w8(32'hb7be7527),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38219d0b),
	.w1(32'hb80dd0a1),
	.w2(32'hb8a9f365),
	.w3(32'hb82295c8),
	.w4(32'hb888f182),
	.w5(32'hb9136109),
	.w6(32'hb8564aee),
	.w7(32'hb7b800eb),
	.w8(32'hb8bace76),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ac9033),
	.w1(32'hb748b555),
	.w2(32'hb7b486f8),
	.w3(32'hb5d38c4c),
	.w4(32'h36b7a42a),
	.w5(32'hb7adbe74),
	.w6(32'h36e08926),
	.w7(32'hb6c6c5cc),
	.w8(32'hb7423cb1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86451f5),
	.w1(32'hb78df193),
	.w2(32'hb58dc24e),
	.w3(32'h36cf2ef7),
	.w4(32'hb64f117d),
	.w5(32'hb7bfe101),
	.w6(32'h3620c7ef),
	.w7(32'h37878a2b),
	.w8(32'hb71d599e),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d6e11d),
	.w1(32'h3746e7b4),
	.w2(32'h37e85bff),
	.w3(32'hb76c492e),
	.w4(32'h37eb5298),
	.w5(32'h37899d54),
	.w6(32'hb771b709),
	.w7(32'hb77c5572),
	.w8(32'hb7e92d35),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e333a8),
	.w1(32'hb7043c5b),
	.w2(32'hb8248424),
	.w3(32'hb7d7af5d),
	.w4(32'hb80d785d),
	.w5(32'hb827c12d),
	.w6(32'h377d381b),
	.w7(32'hb7b41839),
	.w8(32'hb84e08fa),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d1534f),
	.w1(32'h379bb10a),
	.w2(32'h37843cbb),
	.w3(32'h37ee3e44),
	.w4(32'h37816431),
	.w5(32'h37d4b42e),
	.w6(32'h36ca050a),
	.w7(32'hb73df33d),
	.w8(32'hb7b1ddca),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394307b9),
	.w1(32'hb8fd1403),
	.w2(32'hb9850584),
	.w3(32'hb8f9d15a),
	.w4(32'h37aa3ad3),
	.w5(32'hb99695f9),
	.w6(32'hb8009812),
	.w7(32'h389dbb00),
	.w8(32'hb964439d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80f14ec),
	.w1(32'h37a37fa4),
	.w2(32'h36a088cc),
	.w3(32'hb638f8db),
	.w4(32'hb7b2c09d),
	.w5(32'h37036a1a),
	.w6(32'hb8550af7),
	.w7(32'hb82308c3),
	.w8(32'hb7ea74f4),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb874a02a),
	.w1(32'hb6b130c2),
	.w2(32'h37e90975),
	.w3(32'hb854e0ef),
	.w4(32'hb61e0b4f),
	.w5(32'hb813d3ae),
	.w6(32'h36f310c2),
	.w7(32'hb8027146),
	.w8(32'hb7634f8c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d89b4),
	.w1(32'h3869c88d),
	.w2(32'hb9cc16f7),
	.w3(32'hb88ad5ae),
	.w4(32'hb85f7f9f),
	.w5(32'hb9acbe83),
	.w6(32'h37bf92da),
	.w7(32'h389dc878),
	.w8(32'hb982c1fe),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e87617),
	.w1(32'h37d915ca),
	.w2(32'hb79d480a),
	.w3(32'h379ca8a6),
	.w4(32'h377163b8),
	.w5(32'h38229c82),
	.w6(32'hb6b72f79),
	.w7(32'hb82e1609),
	.w8(32'hb75e8a86),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37459264),
	.w1(32'hb7fc2685),
	.w2(32'hb8a31b4d),
	.w3(32'hb85b8c34),
	.w4(32'hb72968df),
	.w5(32'hb8a46c5f),
	.w6(32'hb846fdb6),
	.w7(32'hb8559a90),
	.w8(32'hb89c68bd),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6be6bc0),
	.w1(32'hb681e6e5),
	.w2(32'hb73bd2ee),
	.w3(32'hb6ec0c08),
	.w4(32'hb7a074d7),
	.w5(32'hb799036b),
	.w6(32'hb6ced0c6),
	.w7(32'hb7061597),
	.w8(32'hb78fe032),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b1188d),
	.w1(32'h3698faac),
	.w2(32'h3744faee),
	.w3(32'hb88f9e6c),
	.w4(32'h38196042),
	.w5(32'h37bf97a6),
	.w6(32'hb86bc0cc),
	.w7(32'hb6d6d6b9),
	.w8(32'hb7aed8a3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83b809a),
	.w1(32'hb7f137e3),
	.w2(32'hb7bd8a31),
	.w3(32'hb8340e0c),
	.w4(32'h373342b8),
	.w5(32'hb6a4ac40),
	.w6(32'hb82a6639),
	.w7(32'hb8190549),
	.w8(32'h361817ea),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37770d9f),
	.w1(32'h36740f9c),
	.w2(32'h36bb0312),
	.w3(32'hb681811a),
	.w4(32'hb58c83ba),
	.w5(32'h361a8465),
	.w6(32'hb5f3cf5a),
	.w7(32'hb71092d5),
	.w8(32'hb6e9a188),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365fa868),
	.w1(32'h3757b8d3),
	.w2(32'h35cb79d7),
	.w3(32'h369bea40),
	.w4(32'h36ce6b8f),
	.w5(32'hb7902e19),
	.w6(32'h374a0ad4),
	.w7(32'h375e7e14),
	.w8(32'hb535eb55),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76dd219),
	.w1(32'h387f13a9),
	.w2(32'h38325e97),
	.w3(32'hb6b71205),
	.w4(32'h3690f7b1),
	.w5(32'h380d1dea),
	.w6(32'h36f8701b),
	.w7(32'hb7eddcd6),
	.w8(32'h380c6e5d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7feca7b),
	.w1(32'h384e7e2b),
	.w2(32'hb842ebe2),
	.w3(32'hb890eeb4),
	.w4(32'h37aadc90),
	.w5(32'h34f579a3),
	.w6(32'hb72c7364),
	.w7(32'hb809bfd9),
	.w8(32'hb846768a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ecab00),
	.w1(32'hb84a267d),
	.w2(32'hb8c3e46c),
	.w3(32'hb6849d60),
	.w4(32'hb7972dfe),
	.w5(32'hb8ac41f9),
	.w6(32'hb7a2a66d),
	.w7(32'hb8220aa0),
	.w8(32'hb8f545fa),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb604844c),
	.w1(32'h37cf7f90),
	.w2(32'h379bdfba),
	.w3(32'h35f1c0c1),
	.w4(32'h370aca9d),
	.w5(32'h35ed384c),
	.w6(32'h37d88088),
	.w7(32'h3781c857),
	.w8(32'h37a60cab),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ab42c4),
	.w1(32'hb5ce94f1),
	.w2(32'hb88d5c4b),
	.w3(32'hb809ce4b),
	.w4(32'hb8e7c546),
	.w5(32'hb8f4f1ca),
	.w6(32'hb7a8040b),
	.w7(32'hb80a88e2),
	.w8(32'hb83c467c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb897a0aa),
	.w1(32'h3834694c),
	.w2(32'hb6b90fbb),
	.w3(32'hb7f80d34),
	.w4(32'hb6cf3d22),
	.w5(32'hb8006489),
	.w6(32'h3768aeb1),
	.w7(32'hb7873705),
	.w8(32'hb828a6af),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383c2276),
	.w1(32'hb912f47f),
	.w2(32'hb901452d),
	.w3(32'hb94db062),
	.w4(32'h38334d7b),
	.w5(32'hb983fbae),
	.w6(32'h377ee2d0),
	.w7(32'h39425982),
	.w8(32'hb8377ed1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80b02eb),
	.w1(32'hb689eb0b),
	.w2(32'h3810f5bc),
	.w3(32'hb7cb9f20),
	.w4(32'h38284583),
	.w5(32'h3825d740),
	.w6(32'hb82504ee),
	.w7(32'h36b2babf),
	.w8(32'hb89b377d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d95fb8),
	.w1(32'h381d3052),
	.w2(32'h38335917),
	.w3(32'hb73b9ad4),
	.w4(32'h37f694ce),
	.w5(32'h378e8f7e),
	.w6(32'h38514214),
	.w7(32'h38414471),
	.w8(32'h386b10d4),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3746f6c9),
	.w1(32'hb60ebf29),
	.w2(32'hb6cd3551),
	.w3(32'hb805bf1a),
	.w4(32'hb713d468),
	.w5(32'hb72eea50),
	.w6(32'hb6ae9410),
	.w7(32'hb76b8ca8),
	.w8(32'hb615227a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88a60d6),
	.w1(32'h375f9a32),
	.w2(32'hb827445b),
	.w3(32'hb667a30b),
	.w4(32'h37d1b5d2),
	.w5(32'hb6c1d816),
	.w6(32'hb8209825),
	.w7(32'h357b57e8),
	.w8(32'hb7e182ac),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cc0343),
	.w1(32'h38726183),
	.w2(32'h38c37349),
	.w3(32'hb6bd4218),
	.w4(32'h38192154),
	.w5(32'h3848dd90),
	.w6(32'h37e95ae8),
	.w7(32'h3802d593),
	.w8(32'h38324f88),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84cdb31),
	.w1(32'h35ca626f),
	.w2(32'hb5e43b40),
	.w3(32'hb884e5ec),
	.w4(32'h3735b86e),
	.w5(32'h37835113),
	.w6(32'hb78eea4e),
	.w7(32'hb6db0582),
	.w8(32'hb62f720d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b92ef8),
	.w1(32'h38160b20),
	.w2(32'hb7d5b676),
	.w3(32'hb856d446),
	.w4(32'h37b6b594),
	.w5(32'hb8267713),
	.w6(32'h36fb383d),
	.w7(32'h37ef573a),
	.w8(32'hb6a05514),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f14703),
	.w1(32'hb586169c),
	.w2(32'h373f5c3b),
	.w3(32'h37af8c2e),
	.w4(32'h36eefd2e),
	.w5(32'hb78d8049),
	.w6(32'h37f34895),
	.w7(32'h3790f182),
	.w8(32'hb792db37),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c0e1c1),
	.w1(32'hb76ca4db),
	.w2(32'hb7801cf0),
	.w3(32'hb8fad5bb),
	.w4(32'h382a72ce),
	.w5(32'hb8e4c248),
	.w6(32'h385065b8),
	.w7(32'h37788fb9),
	.w8(32'hb8abf2a6),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb791d088),
	.w1(32'hb7e66a2f),
	.w2(32'h36008320),
	.w3(32'hb70dde62),
	.w4(32'hb7ba1a55),
	.w5(32'hb4a2c922),
	.w6(32'hb74e341f),
	.w7(32'h37d0d8c7),
	.w8(32'hb765212a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e6f2d9),
	.w1(32'hb70bf4dc),
	.w2(32'h37828141),
	.w3(32'h384b7590),
	.w4(32'hb7b5c2f6),
	.w5(32'hb6dfa949),
	.w6(32'h37db1d0a),
	.w7(32'hb7b21c4c),
	.w8(32'hb7dd7896),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b3b0ee),
	.w1(32'hb6bac355),
	.w2(32'hb675dd76),
	.w3(32'hb6f2885b),
	.w4(32'h34ac9075),
	.w5(32'hb6c073da),
	.w6(32'hb3daa0d6),
	.w7(32'hb771718f),
	.w8(32'h35bdabeb),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73e3bed),
	.w1(32'h3777b8f7),
	.w2(32'h37b6ca54),
	.w3(32'hb71c81ef),
	.w4(32'h37cd465d),
	.w5(32'h38138dfa),
	.w6(32'h37450d37),
	.w7(32'h3811265a),
	.w8(32'h382577a6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37836fd3),
	.w1(32'h3685a3be),
	.w2(32'hb55649d5),
	.w3(32'h37443fb3),
	.w4(32'h360110a1),
	.w5(32'hb5f43df4),
	.w6(32'h372fd2b2),
	.w7(32'h361f0fa5),
	.w8(32'h36f0811a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375840aa),
	.w1(32'hb6d5e4af),
	.w2(32'hb78f2fd9),
	.w3(32'h3627986b),
	.w4(32'hb6a4aa34),
	.w5(32'hb7b80c59),
	.w6(32'h361f1960),
	.w7(32'h36c7e97e),
	.w8(32'hb7176daa),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3722b9cc),
	.w1(32'hb746b553),
	.w2(32'hb6250177),
	.w3(32'hb73802f4),
	.w4(32'hb758e956),
	.w5(32'hb59c999f),
	.w6(32'hb7e6f9cb),
	.w7(32'hb79dfcad),
	.w8(32'hb81b05a5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82fbbf3),
	.w1(32'h3782401f),
	.w2(32'hb9690b3b),
	.w3(32'hb90f009d),
	.w4(32'hb88046a8),
	.w5(32'hb94e5eeb),
	.w6(32'hb8705941),
	.w7(32'hb89715a1),
	.w8(32'hb9005db8),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8904e47),
	.w1(32'hb772fa85),
	.w2(32'hb7a6e46a),
	.w3(32'hb891aa13),
	.w4(32'h377ce167),
	.w5(32'h36f627df),
	.w6(32'hb7782079),
	.w7(32'hb7c887af),
	.w8(32'hb7511e65),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b63e40),
	.w1(32'hb7ffd1f4),
	.w2(32'h34c6b7a7),
	.w3(32'hb85db5a4),
	.w4(32'hb80fb1c4),
	.w5(32'hb8392b68),
	.w6(32'hb7b0f5ec),
	.w7(32'hb7dbd3e7),
	.w8(32'hb87572dd),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3527872c),
	.w1(32'h37438d6d),
	.w2(32'h3702c215),
	.w3(32'h354636e2),
	.w4(32'h37c7b9dc),
	.w5(32'h37adfac8),
	.w6(32'hb7de41dd),
	.w7(32'hb7aa8297),
	.w8(32'hb7bf5465),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8973f85),
	.w1(32'hb8c37a26),
	.w2(32'hb8c4cd0a),
	.w3(32'hb8d9cb5e),
	.w4(32'hb8bc92d9),
	.w5(32'hb9083795),
	.w6(32'hb80f6154),
	.w7(32'hb805bb09),
	.w8(32'hb89fee2f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7585e80),
	.w1(32'h37970876),
	.w2(32'hb8818234),
	.w3(32'hb7f8c1fc),
	.w4(32'hb517994d),
	.w5(32'hb8926d86),
	.w6(32'hb84f527c),
	.w7(32'h36f82edb),
	.w8(32'hb7df53cb),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385ee3ef),
	.w1(32'hb8a88cde),
	.w2(32'hb90c46dc),
	.w3(32'hb7ce3b6c),
	.w4(32'hb7ba8552),
	.w5(32'hb918002e),
	.w6(32'hb83aaa4c),
	.w7(32'hb78997a6),
	.w8(32'hb8c2b308),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376efe08),
	.w1(32'h37d3c9f8),
	.w2(32'h3732dbd4),
	.w3(32'hb78c5fd6),
	.w4(32'h374330bf),
	.w5(32'hb78e4397),
	.w6(32'h37ac1f31),
	.w7(32'hb6b36abd),
	.w8(32'hb7f10295),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h350d32dd),
	.w1(32'hb903fa38),
	.w2(32'hb86b9e8d),
	.w3(32'hb82e3478),
	.w4(32'hb88d8825),
	.w5(32'hb90aadc1),
	.w6(32'hb7aa00b9),
	.w7(32'hb78db973),
	.w8(32'hb8c6d233),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35caefa3),
	.w1(32'hb543a820),
	.w2(32'h362a40f9),
	.w3(32'hb73461ce),
	.w4(32'hb725d428),
	.w5(32'hb561f589),
	.w6(32'hb62471c4),
	.w7(32'hb60d5725),
	.w8(32'hb6cf0e9b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375fcacd),
	.w1(32'hb65cc13c),
	.w2(32'hb7a59b0b),
	.w3(32'h37a6f7a1),
	.w4(32'hb7b74832),
	.w5(32'hb803ae7a),
	.w6(32'h36aed9b7),
	.w7(32'hb7c0da44),
	.w8(32'hb7e208f8),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eb5ee2),
	.w1(32'hb84f1b9a),
	.w2(32'hb82c45a2),
	.w3(32'h37e61256),
	.w4(32'h3761575b),
	.w5(32'hb7913a30),
	.w6(32'hb846370d),
	.w7(32'h350294a2),
	.w8(32'hb842bfa8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb678d3e8),
	.w1(32'h379efc53),
	.w2(32'hb806280c),
	.w3(32'hb792bed6),
	.w4(32'hb68be620),
	.w5(32'hb7f01210),
	.w6(32'hb761e391),
	.w7(32'hb7faf533),
	.w8(32'hb885c48c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370e8ad6),
	.w1(32'hb679e931),
	.w2(32'hb7c03910),
	.w3(32'hb62e37b5),
	.w4(32'hb78ee882),
	.w5(32'hb72309a5),
	.w6(32'h3759f34a),
	.w7(32'hb6e6536d),
	.w8(32'h3697ce5f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d28c24),
	.w1(32'h36983a54),
	.w2(32'h3693193e),
	.w3(32'hb64e3625),
	.w4(32'h37534083),
	.w5(32'h3711c6b9),
	.w6(32'hb5b0c52c),
	.w7(32'hb4c3d312),
	.w8(32'hb78f0d26),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9101400),
	.w1(32'h35f13880),
	.w2(32'hb8916970),
	.w3(32'h38486f97),
	.w4(32'h378b6d0a),
	.w5(32'hb8b4464c),
	.w6(32'h379a0061),
	.w7(32'hb7303ceb),
	.w8(32'hb7d7ae04),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88a79ea),
	.w1(32'hb702a374),
	.w2(32'hb8b474cf),
	.w3(32'hb8e38071),
	.w4(32'h3865e89a),
	.w5(32'hb8c78404),
	.w6(32'hb77c9bae),
	.w7(32'h37e31496),
	.w8(32'h37cc1b9a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb72cf),
	.w1(32'h3892e1fa),
	.w2(32'hb703f6d0),
	.w3(32'hb8a3e981),
	.w4(32'h3882f787),
	.w5(32'h376f21ba),
	.w6(32'h377e6769),
	.w7(32'hb73a550a),
	.w8(32'h38eacfd3),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3806e6b7),
	.w1(32'hb5a05a4b),
	.w2(32'hb73084db),
	.w3(32'h3843e985),
	.w4(32'hb607830b),
	.w5(32'hb5c17a44),
	.w6(32'h37e9d900),
	.w7(32'h378f59ad),
	.w8(32'h37253e4e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381a9e0f),
	.w1(32'hb98aa8f7),
	.w2(32'hb985fdf7),
	.w3(32'hb8eda9a6),
	.w4(32'hb82b3ad0),
	.w5(32'hb9aaa69b),
	.w6(32'hb6e58eed),
	.w7(32'hb7bde742),
	.w8(32'hb8bc4548),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3860073f),
	.w1(32'h37e3ae19),
	.w2(32'h38baf59c),
	.w3(32'h382fda8b),
	.w4(32'hb812e0e7),
	.w5(32'h38c35cd5),
	.w6(32'hb82acdc2),
	.w7(32'hb8a8574e),
	.w8(32'h3605004f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37afa78a),
	.w1(32'h37c37f44),
	.w2(32'hb578e802),
	.w3(32'hb7da11fc),
	.w4(32'hb7a9b472),
	.w5(32'hb7b352a3),
	.w6(32'h36053940),
	.w7(32'h3627a9bd),
	.w8(32'hb74ff832),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36db1fd3),
	.w1(32'hb764c425),
	.w2(32'h36813c62),
	.w3(32'h3619dde7),
	.w4(32'hb7c0d32b),
	.w5(32'h369b2a2c),
	.w6(32'h3701bbdb),
	.w7(32'h37a3cad0),
	.w8(32'h36226484),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb526dd13),
	.w1(32'h303ad616),
	.w2(32'hb690dc46),
	.w3(32'h38080457),
	.w4(32'h377ba01a),
	.w5(32'h36be11e8),
	.w6(32'hb6ce9986),
	.w7(32'hb7348242),
	.w8(32'hb75884bf),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7186367),
	.w1(32'hb7483f3e),
	.w2(32'hb77755a2),
	.w3(32'hb68bc756),
	.w4(32'hb728fdcc),
	.w5(32'hb77055de),
	.w6(32'hb70e6298),
	.w7(32'hb76dd60b),
	.w8(32'hb776934b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f9f9ce),
	.w1(32'h3819dc14),
	.w2(32'hb8819f8b),
	.w3(32'hb80fc9c2),
	.w4(32'h3813ec87),
	.w5(32'hb84cf942),
	.w6(32'h378a520b),
	.w7(32'h3772cbb4),
	.w8(32'h37e6dad0),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7898332),
	.w1(32'h36486cdb),
	.w2(32'hb734f773),
	.w3(32'hb74aaab9),
	.w4(32'hb87deb53),
	.w5(32'hb7def25d),
	.w6(32'hb816d9fc),
	.w7(32'hb777f413),
	.w8(32'h36dbba42),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f023fe),
	.w1(32'h38677ead),
	.w2(32'h36bd452a),
	.w3(32'hb87a3b49),
	.w4(32'hb6a5a161),
	.w5(32'hb798643a),
	.w6(32'h36c0027c),
	.w7(32'hb8046aa2),
	.w8(32'hb8b8d85a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87d7c32),
	.w1(32'h365129b5),
	.w2(32'hb57e3498),
	.w3(32'hb858c6d4),
	.w4(32'h3774fffa),
	.w5(32'hb579c8e5),
	.w6(32'hb5d16fd3),
	.w7(32'hb43cd428),
	.w8(32'hb6d42fee),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71f36ad),
	.w1(32'hb886e179),
	.w2(32'hb920351c),
	.w3(32'hb8c35827),
	.w4(32'hb813b2ae),
	.w5(32'hb92771ae),
	.w6(32'hb85156cf),
	.w7(32'hb7b1f50d),
	.w8(32'hb8cc8428),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82b1776),
	.w1(32'h37622f96),
	.w2(32'hb7ed5111),
	.w3(32'hb83bcdeb),
	.w4(32'h37c6d850),
	.w5(32'h37e48585),
	.w6(32'h37b12cd2),
	.w7(32'h378035cb),
	.w8(32'h388e5ef1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367a7d73),
	.w1(32'h369f7185),
	.w2(32'h358da020),
	.w3(32'h36a02af8),
	.w4(32'hb708e1fc),
	.w5(32'hb6d455de),
	.w6(32'h3624b1c4),
	.w7(32'hb6f0fd53),
	.w8(32'hb5058b32),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d8b5a1),
	.w1(32'h39017164),
	.w2(32'hb807a41d),
	.w3(32'hb8844a70),
	.w4(32'hb6c80d89),
	.w5(32'hb819caec),
	.w6(32'h38a5c86d),
	.w7(32'hb7e5504a),
	.w8(32'h37dac756),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c3d36d),
	.w1(32'h374e8a6e),
	.w2(32'h371f31f5),
	.w3(32'h364138d9),
	.w4(32'h36d115e0),
	.w5(32'hb6f3e1ca),
	.w6(32'h37494828),
	.w7(32'h36612457),
	.w8(32'h36e52ed5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ac1644),
	.w1(32'hb8156623),
	.w2(32'hb8ae4953),
	.w3(32'hb85ff566),
	.w4(32'hb7ee706b),
	.w5(32'hb88f121d),
	.w6(32'hb80d4e62),
	.w7(32'hb8318eb6),
	.w8(32'hb8ba67cb),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85209d9),
	.w1(32'h37ecf92e),
	.w2(32'h38a67d19),
	.w3(32'hb7c72992),
	.w4(32'h3847de9b),
	.w5(32'h389839cc),
	.w6(32'hb7ba5742),
	.w7(32'h36cc67ac),
	.w8(32'h385503b2),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7feb32f),
	.w1(32'h37a7c851),
	.w2(32'h381c15d9),
	.w3(32'hb8204f29),
	.w4(32'hb7c0b6d2),
	.w5(32'hb58b44ab),
	.w6(32'hb85c0cbb),
	.w7(32'hb78e1bb7),
	.w8(32'hb823aa02),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7058274),
	.w1(32'h36be7c65),
	.w2(32'hb6140e83),
	.w3(32'hb7321786),
	.w4(32'h36baa264),
	.w5(32'h3620da2a),
	.w6(32'h37b14a1f),
	.w7(32'h37669c1f),
	.w8(32'h36edfd95),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ce14ac),
	.w1(32'h37b36eab),
	.w2(32'hb6c80437),
	.w3(32'hb81c3191),
	.w4(32'h3872cef4),
	.w5(32'h37998972),
	.w6(32'hb82912da),
	.w7(32'hb7cfa4d1),
	.w8(32'hb782d57d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb814a109),
	.w1(32'h378bb996),
	.w2(32'hb72e7221),
	.w3(32'hb8739769),
	.w4(32'hb759643e),
	.w5(32'hb82a7d58),
	.w6(32'h36a503aa),
	.w7(32'hb78fe647),
	.w8(32'hb82d7f40),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5cc0796),
	.w1(32'hb6c3959b),
	.w2(32'hb8a378f6),
	.w3(32'hb80155f3),
	.w4(32'hb7a22061),
	.w5(32'hb901eff9),
	.w6(32'hb6ee7447),
	.w7(32'hb812e6e3),
	.w8(32'hb8c82684),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8335a98),
	.w1(32'h35bed84b),
	.w2(32'hb71dc889),
	.w3(32'hb86a0c28),
	.w4(32'hb6d1acb0),
	.w5(32'h3393c8c4),
	.w6(32'h371435f7),
	.w7(32'hb68d2c54),
	.w8(32'hb6ee6505),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e15b26),
	.w1(32'h3707230b),
	.w2(32'hb3894c69),
	.w3(32'hb62858a5),
	.w4(32'h37525643),
	.w5(32'hb6c54571),
	.w6(32'h3694ddca),
	.w7(32'hb6f055b5),
	.w8(32'hb75b3c59),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc4f72),
	.w1(32'hb78f1dbd),
	.w2(32'hb7229c6a),
	.w3(32'hb8675dbf),
	.w4(32'h36ac1e0e),
	.w5(32'hb7c852c1),
	.w6(32'hb7cd5e90),
	.w7(32'h37ca8aad),
	.w8(32'h379158c7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b4d8a4),
	.w1(32'hb792fa8b),
	.w2(32'hb90e18a8),
	.w3(32'hb919d04d),
	.w4(32'hb76c4bb9),
	.w5(32'hb91d9b16),
	.w6(32'hb818d516),
	.w7(32'hb828fdeb),
	.w8(32'hb871837d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ef709),
	.w1(32'h3735f7c3),
	.w2(32'hb81002f5),
	.w3(32'h38bab73f),
	.w4(32'h382387ac),
	.w5(32'hb82b41fd),
	.w6(32'hb83d7147),
	.w7(32'h38535ac4),
	.w8(32'hb8ce76b2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d6803),
	.w1(32'h381bf96c),
	.w2(32'hb8c2a0e8),
	.w3(32'hb7f5495e),
	.w4(32'h37f058db),
	.w5(32'hb8f86e95),
	.w6(32'h379f72f3),
	.w7(32'h38040d0a),
	.w8(32'hb7e2db36),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361dfb49),
	.w1(32'h37410c52),
	.w2(32'h3748cd68),
	.w3(32'hb6626b1c),
	.w4(32'h36a389fb),
	.w5(32'h360cabd4),
	.w6(32'h375168a3),
	.w7(32'h36b91983),
	.w8(32'h370075ee),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37826d70),
	.w1(32'h33a47dd7),
	.w2(32'hb58a2491),
	.w3(32'h36bb0f48),
	.w4(32'h368bfaf6),
	.w5(32'hb66345be),
	.w6(32'h366b1b5f),
	.w7(32'hb730296c),
	.w8(32'hb7f53366),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d6efa),
	.w1(32'h399acd24),
	.w2(32'hb93e2d63),
	.w3(32'hb891ea76),
	.w4(32'h391669e7),
	.w5(32'hb8da5c10),
	.w6(32'h388d9bf9),
	.w7(32'h38999be3),
	.w8(32'h376c187b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e38497),
	.w1(32'hb8f49bcc),
	.w2(32'hb996f79c),
	.w3(32'hb8db9b4e),
	.w4(32'hb7af71c2),
	.w5(32'hb9a80476),
	.w6(32'h37828887),
	.w7(32'h380f043a),
	.w8(32'hb70dcb26),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901eec6),
	.w1(32'h387a89a8),
	.w2(32'hb97400b8),
	.w3(32'hb893c893),
	.w4(32'h37942aa8),
	.w5(32'hb9458713),
	.w6(32'h3789442c),
	.w7(32'h37e04627),
	.w8(32'hb845f770),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898178b),
	.w1(32'h37d584f1),
	.w2(32'h383f4e0d),
	.w3(32'hb7e0d051),
	.w4(32'h38506dfd),
	.w5(32'h38b62eb2),
	.w6(32'h379ac4d7),
	.w7(32'h381371ad),
	.w8(32'h387ab2d1),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77947ae),
	.w1(32'h37e2141a),
	.w2(32'h37ae8506),
	.w3(32'hb77af423),
	.w4(32'h37aacc22),
	.w5(32'hb62888f2),
	.w6(32'h368dfe74),
	.w7(32'hb7e4235b),
	.w8(32'hb7bccfb3),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8131a0c),
	.w1(32'h32f981a1),
	.w2(32'hb65327b3),
	.w3(32'hb84b0627),
	.w4(32'h360c9199),
	.w5(32'hb6aa4875),
	.w6(32'hb4aaa5df),
	.w7(32'hb652d9b5),
	.w8(32'h36b07afe),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb650dc9a),
	.w1(32'hb3b5534b),
	.w2(32'hb7a2e2c5),
	.w3(32'hb7706be2),
	.w4(32'hb8077229),
	.w5(32'hb7bf6020),
	.w6(32'hb571c200),
	.w7(32'hb6b1f9ce),
	.w8(32'h368e8b41),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78fcf09),
	.w1(32'h379e18fe),
	.w2(32'hb3b7406c),
	.w3(32'hb7bbae78),
	.w4(32'hb60b3a62),
	.w5(32'hb60d73f8),
	.w6(32'h379bb791),
	.w7(32'hb66ee3c4),
	.w8(32'hb7da2369),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83aeb57),
	.w1(32'hb7ca1ad9),
	.w2(32'h35004fac),
	.w3(32'hb848b352),
	.w4(32'hb7a2d2dd),
	.w5(32'h36e5887b),
	.w6(32'hb76e4e74),
	.w7(32'hb733e465),
	.w8(32'hb7562d4d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35538845),
	.w1(32'hb6695c3f),
	.w2(32'hb77e890a),
	.w3(32'hb64ee744),
	.w4(32'h358d75e3),
	.w5(32'hb6c7328e),
	.w6(32'h3708c209),
	.w7(32'hb72230ae),
	.w8(32'h36fa1710),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec897c),
	.w1(32'hb8c78610),
	.w2(32'hb9027d65),
	.w3(32'hb6652e84),
	.w4(32'h362d62f0),
	.w5(32'hb91e17c9),
	.w6(32'h3700af4a),
	.w7(32'h35af1c57),
	.w8(32'hb8b17bb3),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82347ca),
	.w1(32'hb525639c),
	.w2(32'hb851d8d6),
	.w3(32'hb7aed61d),
	.w4(32'hb7f42fba),
	.w5(32'hb80d7ba2),
	.w6(32'hb7232818),
	.w7(32'hb7c08223),
	.w8(32'hb7875006),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c67740),
	.w1(32'h37e8c059),
	.w2(32'hb77f735b),
	.w3(32'h37bc2d77),
	.w4(32'hb78c25bc),
	.w5(32'hb7a8571c),
	.w6(32'h38649fbe),
	.w7(32'h37e1ead6),
	.w8(32'h37adcbba),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f79fc),
	.w1(32'h38d1f320),
	.w2(32'hb9f312be),
	.w3(32'hb9887fc1),
	.w4(32'h38bea858),
	.w5(32'hb9d097e9),
	.w6(32'hb82bb71e),
	.w7(32'h3921a618),
	.w8(32'hb9158038),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aba921),
	.w1(32'hb82c2c8d),
	.w2(32'hb879101c),
	.w3(32'hb831a52c),
	.w4(32'hb7e9517e),
	.w5(32'hb8ac991c),
	.w6(32'hb68b7f5b),
	.w7(32'hb6855ac3),
	.w8(32'hb86e1fa1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36eba686),
	.w1(32'h36059ab8),
	.w2(32'h36ff9f97),
	.w3(32'h353f4c4e),
	.w4(32'hb6c93e02),
	.w5(32'h36779d9c),
	.w6(32'hb70ff3b7),
	.w7(32'hb6f33511),
	.w8(32'hb7048291),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3842f56d),
	.w1(32'hb6d7b52f),
	.w2(32'hb8977cd5),
	.w3(32'hb85764db),
	.w4(32'h37d35d8e),
	.w5(32'hb8b9ee6d),
	.w6(32'hb6f64a4c),
	.w7(32'h3783def9),
	.w8(32'hb80f58af),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363cedb1),
	.w1(32'hb3f26f46),
	.w2(32'h35207897),
	.w3(32'hb4e92ecd),
	.w4(32'hb636eb5c),
	.w5(32'hb6bc01b3),
	.w6(32'h356ada34),
	.w7(32'hb6a77ff1),
	.w8(32'hb6ddcbde),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f10add),
	.w1(32'h37c6530a),
	.w2(32'h37fb0e96),
	.w3(32'hb72bc4f8),
	.w4(32'h36efa012),
	.w5(32'h37164294),
	.w6(32'h37e4136d),
	.w7(32'h3798c6a7),
	.w8(32'h37d09880),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3809fe34),
	.w1(32'h36860cd7),
	.w2(32'h36ee2539),
	.w3(32'h370a734d),
	.w4(32'hb72685cc),
	.w5(32'hb2de3e50),
	.w6(32'hb72cf01f),
	.w7(32'hb7036b15),
	.w8(32'hb72d5697),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3640ab26),
	.w1(32'h370913cd),
	.w2(32'h35bcbab0),
	.w3(32'hb64099a3),
	.w4(32'h36df400c),
	.w5(32'hb703e67b),
	.w6(32'h3776ced7),
	.w7(32'hb71c4920),
	.w8(32'hb7d32dff),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b19ffc),
	.w1(32'h376c58ff),
	.w2(32'hb79d729c),
	.w3(32'h36dec6b2),
	.w4(32'h357fb2de),
	.w5(32'h35e52078),
	.w6(32'h36a2054f),
	.w7(32'h36d39db2),
	.w8(32'h3742a39c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3768dc9a),
	.w1(32'hb866eb38),
	.w2(32'hb8792d8a),
	.w3(32'hb8078668),
	.w4(32'hb8397c0d),
	.w5(32'hb894ffbe),
	.w6(32'hb8802e95),
	.w7(32'hb803974e),
	.w8(32'hb908b504),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a32f67),
	.w1(32'hb837dd2c),
	.w2(32'hb8f7902a),
	.w3(32'hb8136370),
	.w4(32'hb7f76d62),
	.w5(32'hb91f8440),
	.w6(32'hb8328140),
	.w7(32'hb738cd7a),
	.w8(32'hb8d1f044),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382a05d3),
	.w1(32'hb84b8c53),
	.w2(32'hb8c0ecaf),
	.w3(32'hb7d68461),
	.w4(32'hb7a4534a),
	.w5(32'hb8f93785),
	.w6(32'hb7a067e9),
	.w7(32'hb7e1181e),
	.w8(32'hb8c77737),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79a7937),
	.w1(32'hb6a2e51b),
	.w2(32'h379cae0d),
	.w3(32'hb75c09a2),
	.w4(32'hb57a070c),
	.w5(32'h37ad5ddd),
	.w6(32'hb58b3db4),
	.w7(32'h3739de8d),
	.w8(32'h36d709e5),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37155752),
	.w1(32'h367f56d2),
	.w2(32'h37255a2c),
	.w3(32'h36cc11ea),
	.w4(32'hb77a932e),
	.w5(32'hb542952e),
	.w6(32'hb77a5299),
	.w7(32'hb76a57c0),
	.w8(32'hb79ffbda),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363e2ea5),
	.w1(32'h351c15af),
	.w2(32'hb5100763),
	.w3(32'hb67d2268),
	.w4(32'hb73db790),
	.w5(32'hb6641491),
	.w6(32'hb6ae7a21),
	.w7(32'hb707ed20),
	.w8(32'hb7162e45),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb53574f9),
	.w1(32'h354cfc48),
	.w2(32'hb28e55aa),
	.w3(32'hb595d751),
	.w4(32'hb72bd2a5),
	.w5(32'hb65c56a0),
	.w6(32'hb6a685bc),
	.w7(32'hb734f37e),
	.w8(32'hb725a3aa),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37817e16),
	.w1(32'hb8b4c32a),
	.w2(32'hb9239298),
	.w3(32'hb846aa19),
	.w4(32'hb8dc4e51),
	.w5(32'hb945a9d9),
	.w6(32'hb7790106),
	.w7(32'hb7cd3325),
	.w8(32'hb9096b03),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77e3549),
	.w1(32'hb75b496d),
	.w2(32'hb668ca56),
	.w3(32'hb778af2e),
	.w4(32'hb6bf95f9),
	.w5(32'h3771732c),
	.w6(32'hb6e9b8a7),
	.w7(32'hb6370609),
	.w8(32'h37cd7f06),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369a4034),
	.w1(32'hb6fbed89),
	.w2(32'hb74d85b5),
	.w3(32'h36e554fa),
	.w4(32'hb60f48ca),
	.w5(32'hb710abba),
	.w6(32'hb6cf0162),
	.w7(32'hb7620feb),
	.w8(32'hb2cc6535),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364b176e),
	.w1(32'hb774d2c2),
	.w2(32'hb33c8ea9),
	.w3(32'hb74b4f8a),
	.w4(32'hb697c350),
	.w5(32'hb5dedab0),
	.w6(32'hb7e05cc1),
	.w7(32'hb7fc2f47),
	.w8(32'hb76bd239),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb730dc39),
	.w1(32'h35441b31),
	.w2(32'h3648a1d2),
	.w3(32'h34f0b1e1),
	.w4(32'hb7523436),
	.w5(32'hb65de22d),
	.w6(32'hb6815119),
	.w7(32'hb6be6fcc),
	.w8(32'hb70d2e60),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bd2729),
	.w1(32'hb75feb14),
	.w2(32'hb892f586),
	.w3(32'hb6b7b18b),
	.w4(32'hb8354ee1),
	.w5(32'hb8d013ef),
	.w6(32'hb74410fc),
	.w7(32'h382006c4),
	.w8(32'hb710afd6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86b57e3),
	.w1(32'h37ae4cf9),
	.w2(32'h35d38614),
	.w3(32'hb80f0fd5),
	.w4(32'h36080d4c),
	.w5(32'hb6e6f753),
	.w6(32'h375c157d),
	.w7(32'hb6c9e13a),
	.w8(32'hb6a73ae4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b8ee45),
	.w1(32'hb85a3d36),
	.w2(32'hb75d751c),
	.w3(32'hb7bc9bab),
	.w4(32'h37240269),
	.w5(32'hb83bef29),
	.w6(32'h39312707),
	.w7(32'hb623b27f),
	.w8(32'hb8e9aa21),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b1b187),
	.w1(32'h3b20e7df),
	.w2(32'h3bcd3205),
	.w3(32'h36f1f85c),
	.w4(32'h3ac199c7),
	.w5(32'h3b96aed8),
	.w6(32'h3a1cf114),
	.w7(32'h3b992906),
	.w8(32'hb9dd3b44),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdd1d5),
	.w1(32'h3b02a648),
	.w2(32'h3b8ae7ea),
	.w3(32'hba3998b4),
	.w4(32'hbb2d6802),
	.w5(32'h3a424ae1),
	.w6(32'hbb345bf4),
	.w7(32'h3a5cf152),
	.w8(32'hbac551d1),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule