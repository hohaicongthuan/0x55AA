module layer_10_featuremap_46(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94dce66),
	.w1(32'h3af40055),
	.w2(32'h3a58aae6),
	.w3(32'hbbcc3265),
	.w4(32'hbb579806),
	.w5(32'h3b709728),
	.w6(32'hbc47eda4),
	.w7(32'hbc6e9dde),
	.w8(32'h3ad5cb95),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb0837),
	.w1(32'h3b906507),
	.w2(32'h3afe4bd9),
	.w3(32'hbc34013c),
	.w4(32'h3955a5c9),
	.w5(32'hbb7e2fc6),
	.w6(32'hbbf0616c),
	.w7(32'h3b1aca54),
	.w8(32'hb8a1252b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d8c5d),
	.w1(32'h37d721bc),
	.w2(32'h3be63ec5),
	.w3(32'h3ab8d4b2),
	.w4(32'h3a6c90fe),
	.w5(32'h3ab911b9),
	.w6(32'hbac494ed),
	.w7(32'h3b6cbcb5),
	.w8(32'h3abb011a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33f651),
	.w1(32'h3a3c03dc),
	.w2(32'hb971bd00),
	.w3(32'h3b0927c7),
	.w4(32'hba1189b6),
	.w5(32'hbaee0d93),
	.w6(32'hbba2ee98),
	.w7(32'hba82b5cd),
	.w8(32'hbbde0771),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb554310),
	.w1(32'h3b92eeb5),
	.w2(32'h38fa6dd2),
	.w3(32'hbbb1f546),
	.w4(32'hba89fc29),
	.w5(32'hbb83bd67),
	.w6(32'hbba8fc5a),
	.w7(32'hbbade141),
	.w8(32'hbadd0b5d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc049f9f),
	.w1(32'hbbd52c94),
	.w2(32'h3d51f3a1),
	.w3(32'h3b097e3c),
	.w4(32'hb8c36ff7),
	.w5(32'h3dbc9621),
	.w6(32'hbb845534),
	.w7(32'h3be72a49),
	.w8(32'h3d8605ac),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d1e5b),
	.w1(32'hbd4cd19d),
	.w2(32'hbbcf5b33),
	.w3(32'h3b6b78e7),
	.w4(32'hbdbfa190),
	.w5(32'hbb80c60b),
	.w6(32'h3c89d31c),
	.w7(32'hbd31ccf9),
	.w8(32'h3b37e653),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09c8f3),
	.w1(32'hbb88b941),
	.w2(32'h3ad97d4e),
	.w3(32'hbb9f2d54),
	.w4(32'hbbbc2899),
	.w5(32'h3c05e9ad),
	.w6(32'hb9cbfb54),
	.w7(32'hbc2917f7),
	.w8(32'h3c03f8db),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06a38f),
	.w1(32'hbbfacecc),
	.w2(32'hbb0ee84b),
	.w3(32'hb9694e5b),
	.w4(32'h39fa225b),
	.w5(32'hbc0685e9),
	.w6(32'h3c00d0ac),
	.w7(32'h3a3e02cd),
	.w8(32'hbb43e496),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53ef9b),
	.w1(32'hba37136c),
	.w2(32'hbd38c071),
	.w3(32'hbbb9a4e3),
	.w4(32'h3c2c522d),
	.w5(32'hbd739a88),
	.w6(32'h3b7182b3),
	.w7(32'h3c883deb),
	.w8(32'hbd261c4a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75da1f),
	.w1(32'h3d19e48a),
	.w2(32'h3bbc49dc),
	.w3(32'h3c112378),
	.w4(32'h3d991eea),
	.w5(32'h3b8acc00),
	.w6(32'hbb255367),
	.w7(32'h3d26f0d5),
	.w8(32'h3b20c7b7),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c135d),
	.w1(32'hbb3e04e3),
	.w2(32'h3b4a68b0),
	.w3(32'h3bc47bc6),
	.w4(32'hbb0b00a4),
	.w5(32'h3c50926a),
	.w6(32'hbb0483b1),
	.w7(32'hbae0d742),
	.w8(32'h3c4177e7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb94fe1),
	.w1(32'hbc5bc440),
	.w2(32'hbba22798),
	.w3(32'h3b9ba5fb),
	.w4(32'hbc4ce1b3),
	.w5(32'h3b560620),
	.w6(32'h3c19a688),
	.w7(32'hba04c7aa),
	.w8(32'h3bab8072),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ad1ff),
	.w1(32'h3b112522),
	.w2(32'h3ba3d0ab),
	.w3(32'h3b828396),
	.w4(32'h3b0d9aea),
	.w5(32'hbafdfa93),
	.w6(32'hb920f0cc),
	.w7(32'hbb591f2c),
	.w8(32'h3a15f92d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f2c84),
	.w1(32'hbab610bd),
	.w2(32'h3a3619a6),
	.w3(32'h3b0cc2b8),
	.w4(32'h3bc154b8),
	.w5(32'hbbc07c6e),
	.w6(32'hb9beff0a),
	.w7(32'h3b9365c0),
	.w8(32'hb9d21038),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5960f0),
	.w1(32'hbb0a3b72),
	.w2(32'hbcf88eb7),
	.w3(32'hbba2394d),
	.w4(32'h3acf5ef2),
	.w5(32'hbd0f44b8),
	.w6(32'hbb46dca5),
	.w7(32'h3b168973),
	.w8(32'hbcd5d56c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a531a4d),
	.w1(32'h3cb07ac1),
	.w2(32'h3b376615),
	.w3(32'h3b8886d8),
	.w4(32'h3d33ee37),
	.w5(32'hbb18f202),
	.w6(32'hbb857097),
	.w7(32'h3cc677e7),
	.w8(32'h38058800),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e6687),
	.w1(32'hbbefba12),
	.w2(32'hbbd8b020),
	.w3(32'hbbfc921f),
	.w4(32'hbaa731a5),
	.w5(32'hba9e4c89),
	.w6(32'hbbe777a0),
	.w7(32'hba952b1e),
	.w8(32'hbba97427),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3a32e),
	.w1(32'hbb4b8637),
	.w2(32'h39c6c963),
	.w3(32'h39abc448),
	.w4(32'h3b8b9448),
	.w5(32'h3ad95fa0),
	.w6(32'hba9eb3be),
	.w7(32'h3bb9d906),
	.w8(32'h3ba42de8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15a5b6),
	.w1(32'hbc35857c),
	.w2(32'h3b39d1d1),
	.w3(32'h3b1a46f6),
	.w4(32'hbc12291e),
	.w5(32'hba9aabdc),
	.w6(32'hbb8c2462),
	.w7(32'hbb9612b4),
	.w8(32'hbb4e2722),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf10d82),
	.w1(32'h3bd7f86b),
	.w2(32'hb94af7ce),
	.w3(32'hbc9ffcd1),
	.w4(32'hbbf76edf),
	.w5(32'h3b81e836),
	.w6(32'hbc165978),
	.w7(32'hbb2f6bd0),
	.w8(32'hbb748624),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d2037),
	.w1(32'h3adcabaa),
	.w2(32'h3b8d693e),
	.w3(32'hba2afe1f),
	.w4(32'h3bc91a0d),
	.w5(32'h3b4f6486),
	.w6(32'h3b4f756e),
	.w7(32'hbae03242),
	.w8(32'h3b244944),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60f80b),
	.w1(32'hbc4a49f5),
	.w2(32'hbd380e44),
	.w3(32'hbc085ea1),
	.w4(32'hbbb5baf7),
	.w5(32'hbd7ef6b2),
	.w6(32'hbbb6bad0),
	.w7(32'hbb7561a3),
	.w8(32'hbd1db3f2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdeb1b7),
	.w1(32'h3d0244dd),
	.w2(32'hbb0d6c39),
	.w3(32'h3c0df0c6),
	.w4(32'h3da68e4d),
	.w5(32'h3b2f2127),
	.w6(32'hbaa309ad),
	.w7(32'h3d4c6d7d),
	.w8(32'hba44e291),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82a127),
	.w1(32'h3a1b861b),
	.w2(32'h3bb965db),
	.w3(32'hbbd73468),
	.w4(32'h3bda3da6),
	.w5(32'h3c11b2ae),
	.w6(32'hbb63f872),
	.w7(32'h3b8fb8bf),
	.w8(32'h3b0405d7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb108091),
	.w1(32'hbc3c7bb1),
	.w2(32'h3bb6ab5a),
	.w3(32'hbc73328c),
	.w4(32'hbc87db60),
	.w5(32'h3be63745),
	.w6(32'hbc0a093b),
	.w7(32'hbbb9b4fe),
	.w8(32'h3a98cbbe),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba440f7),
	.w1(32'hba92c4b1),
	.w2(32'hb81d2544),
	.w3(32'h3b5be680),
	.w4(32'hba1ad0e7),
	.w5(32'h3a05b889),
	.w6(32'h3b263b26),
	.w7(32'hbc35b1de),
	.w8(32'hba7be8f3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52be83),
	.w1(32'hb9d055fc),
	.w2(32'h3b93e574),
	.w3(32'hbb966a7d),
	.w4(32'hbbac3b2e),
	.w5(32'h3c202007),
	.w6(32'hbbf1caa8),
	.w7(32'hbb66f692),
	.w8(32'h3c90e5f1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba024c6),
	.w1(32'h3b7ce03d),
	.w2(32'h3c0dbc53),
	.w3(32'hbb99c408),
	.w4(32'hbafd0410),
	.w5(32'hb9f338d0),
	.w6(32'h3ae47699),
	.w7(32'hbada14c3),
	.w8(32'hbb79b0a7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f296a),
	.w1(32'hbc1ffc56),
	.w2(32'h3a85c53d),
	.w3(32'hbc776daa),
	.w4(32'hbb90b544),
	.w5(32'hba8d9cd6),
	.w6(32'hbb98f5ac),
	.w7(32'h3b5269a7),
	.w8(32'hbb967867),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8d2a0),
	.w1(32'hbacf6cb3),
	.w2(32'hb90cac46),
	.w3(32'h3a8a06e6),
	.w4(32'hba04badf),
	.w5(32'hbc99f56e),
	.w6(32'hbb64e5a0),
	.w7(32'hbb558310),
	.w8(32'hbc949c45),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc59a4),
	.w1(32'hbb84258f),
	.w2(32'hba9055d7),
	.w3(32'hbc0c32bc),
	.w4(32'h3c85906a),
	.w5(32'h3ba7f7be),
	.w6(32'hba67fc67),
	.w7(32'h3cc3c48e),
	.w8(32'h3b9a47dd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc290132),
	.w1(32'hbb8fe851),
	.w2(32'hbbebed72),
	.w3(32'h3b8575de),
	.w4(32'h3c27302f),
	.w5(32'h3ab34e98),
	.w6(32'h3bd8dec8),
	.w7(32'h3cacc452),
	.w8(32'hba72ca57),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6917f),
	.w1(32'h39bc3e82),
	.w2(32'h3b21682b),
	.w3(32'h3b45ba80),
	.w4(32'h3a556506),
	.w5(32'h3bf1f0f3),
	.w6(32'hbabfe674),
	.w7(32'hbb875e3f),
	.w8(32'h3c280857),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a2bf5),
	.w1(32'h3a10d1c9),
	.w2(32'h3a6fae2e),
	.w3(32'h3c16fa1c),
	.w4(32'h3b0b08e8),
	.w5(32'hb9d3e40a),
	.w6(32'h3c4cd4a7),
	.w7(32'h3bba6b6b),
	.w8(32'h3ace8856),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba098206),
	.w1(32'h3a803a98),
	.w2(32'h3bceaa9d),
	.w3(32'hbb030ea2),
	.w4(32'hbb3869ef),
	.w5(32'h3ca7cb1e),
	.w6(32'h3aa9fde4),
	.w7(32'h3a188a42),
	.w8(32'h3b7f36c8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fdc18),
	.w1(32'hbc6c0009),
	.w2(32'hbc5c35ca),
	.w3(32'h3c23be09),
	.w4(32'hbc3e2fa7),
	.w5(32'h3b17ffc4),
	.w6(32'h3c70cad4),
	.w7(32'h3cc82a53),
	.w8(32'h3afee8fb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc536ad0),
	.w1(32'h3bc2c831),
	.w2(32'h3a60040b),
	.w3(32'hbbf4f175),
	.w4(32'h3bfe268a),
	.w5(32'hba845e4c),
	.w6(32'hbc70c330),
	.w7(32'hbb9f11bf),
	.w8(32'h3c4dea1f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6a528),
	.w1(32'h3c134b2d),
	.w2(32'h3bd71ef9),
	.w3(32'hbc464c53),
	.w4(32'h3c04e6fe),
	.w5(32'h3c87652a),
	.w6(32'hbc3221af),
	.w7(32'hbc453f3e),
	.w8(32'h3bff8597),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb655f5),
	.w1(32'h3aa1cdb8),
	.w2(32'hb9a4556e),
	.w3(32'hbbde2192),
	.w4(32'h3b8487b1),
	.w5(32'hbbcb3942),
	.w6(32'hbc83d361),
	.w7(32'hb9af40d2),
	.w8(32'hbbfeb24c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b472726),
	.w1(32'h3b8299b6),
	.w2(32'h3b27fec6),
	.w3(32'hba9e4a38),
	.w4(32'hbbcea959),
	.w5(32'hba815a07),
	.w6(32'hbb9b693a),
	.w7(32'hbbdae43d),
	.w8(32'hba13329d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27fd49),
	.w1(32'h3b10ea07),
	.w2(32'hba90f50e),
	.w3(32'h3abe7f6b),
	.w4(32'h3b3109e8),
	.w5(32'h3c0372f3),
	.w6(32'hbaf3e67c),
	.w7(32'hbc0c57bb),
	.w8(32'h3c09d72e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cdc01),
	.w1(32'h3bacf9b5),
	.w2(32'h3a3a6684),
	.w3(32'h3bc2cde7),
	.w4(32'h3ba7f63f),
	.w5(32'hbadb9340),
	.w6(32'h3c64849c),
	.w7(32'h3c9aeaaf),
	.w8(32'hb6d5649c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d3b05),
	.w1(32'hbc3431dc),
	.w2(32'hbc2d97e6),
	.w3(32'hbc159517),
	.w4(32'hbb85f219),
	.w5(32'hbc8dedc6),
	.w6(32'hbb7a45d7),
	.w7(32'hbb029975),
	.w8(32'hbc5bdc29),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b5115),
	.w1(32'h3bba5fd3),
	.w2(32'h3b8cceab),
	.w3(32'hbd00b471),
	.w4(32'hbbfae720),
	.w5(32'h3c955882),
	.w6(32'hbc8e612b),
	.w7(32'h3b8d34ec),
	.w8(32'h3c85a477),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba00193),
	.w1(32'hbc676ce9),
	.w2(32'hbc781798),
	.w3(32'hbc0fd88d),
	.w4(32'hbc4e7314),
	.w5(32'h39d9b39b),
	.w6(32'hbc0bc74c),
	.w7(32'hbc1eef9b),
	.w8(32'hbb51186a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35f586),
	.w1(32'hbbd3b86f),
	.w2(32'hb9ab9757),
	.w3(32'hba5c9ac8),
	.w4(32'hbbde9eca),
	.w5(32'hbb202668),
	.w6(32'hbbf8a91f),
	.w7(32'hbbd10e9f),
	.w8(32'h3b281b52),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cc543),
	.w1(32'hbbcfcd8f),
	.w2(32'hbc01b66d),
	.w3(32'h3c43d0fe),
	.w4(32'hbb39ea26),
	.w5(32'hba21e10e),
	.w6(32'h3c80c165),
	.w7(32'h3bd33189),
	.w8(32'h3ac5bec7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3e787),
	.w1(32'hbafe2fa0),
	.w2(32'h3a872614),
	.w3(32'hbb491375),
	.w4(32'h3a937aa5),
	.w5(32'hbb6337d1),
	.w6(32'h39da5498),
	.w7(32'h3a8076cd),
	.w8(32'hbb299e9c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4cc66f),
	.w1(32'h3bc50f89),
	.w2(32'h3b506ec7),
	.w3(32'h3c3d2685),
	.w4(32'h3c2904c7),
	.w5(32'h3c05f282),
	.w6(32'hba8c067d),
	.w7(32'hbaafa59c),
	.w8(32'h3cc643e2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb163565),
	.w1(32'hbc213306),
	.w2(32'h3b9ecfd6),
	.w3(32'hbb62aa65),
	.w4(32'hbcbf0366),
	.w5(32'h3c122423),
	.w6(32'h3c604073),
	.w7(32'hbc41bc98),
	.w8(32'h3c0cb75b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa6fa7),
	.w1(32'hbc00ff27),
	.w2(32'hbb4321f9),
	.w3(32'h3b0112e0),
	.w4(32'hba7f43db),
	.w5(32'h3c82bf5e),
	.w6(32'hbb8730b2),
	.w7(32'h3b8794a6),
	.w8(32'h3cc6ec18),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9466c8),
	.w1(32'hbc73dd12),
	.w2(32'hba267c53),
	.w3(32'hbb94ba10),
	.w4(32'hbcc8747c),
	.w5(32'h3bb8ea2f),
	.w6(32'h3c55532f),
	.w7(32'hbc2fe235),
	.w8(32'h3beabd98),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc276f4e),
	.w1(32'hbc155aa4),
	.w2(32'h393f97bb),
	.w3(32'h3bfba862),
	.w4(32'h3b078c8f),
	.w5(32'hbb4cf63f),
	.w6(32'h3b0ef0ae),
	.w7(32'h3b8aef20),
	.w8(32'h3a55d1cd),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa74e05),
	.w1(32'hbc390580),
	.w2(32'h3bace7c3),
	.w3(32'hbb901359),
	.w4(32'hb948f2bb),
	.w5(32'hbb7e2e98),
	.w6(32'h3b360ddc),
	.w7(32'h3b802ed2),
	.w8(32'hbce19e28),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d4b48),
	.w1(32'hbb4a6d30),
	.w2(32'h3ad5cabf),
	.w3(32'hbc03de14),
	.w4(32'h3c04a93c),
	.w5(32'h3b85a09b),
	.w6(32'hbba56c02),
	.w7(32'h3c98edab),
	.w8(32'hba40a3a1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b6373),
	.w1(32'hbad0381b),
	.w2(32'hbb13af36),
	.w3(32'h3a547542),
	.w4(32'h3adc603e),
	.w5(32'h3981b220),
	.w6(32'hbb8724ef),
	.w7(32'hbc11cb5d),
	.w8(32'h39d70dab),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba901449),
	.w1(32'hbb0c9353),
	.w2(32'hbb4c2ee4),
	.w3(32'h39de0012),
	.w4(32'hbb4f0a77),
	.w5(32'hbadfe2dd),
	.w6(32'hbb317903),
	.w7(32'hbaa04486),
	.w8(32'h3b62a37e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18b045),
	.w1(32'h3c83339a),
	.w2(32'h3a628fe1),
	.w3(32'hbbb04a23),
	.w4(32'h3c45ade8),
	.w5(32'h3b584637),
	.w6(32'hbb025d7e),
	.w7(32'h3c86cbfd),
	.w8(32'h3bfd75c9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a6a4e),
	.w1(32'hbc0559e7),
	.w2(32'h3c216ca4),
	.w3(32'h3b35cf36),
	.w4(32'hb8d3f56b),
	.w5(32'h3c284e2d),
	.w6(32'hba1961a8),
	.w7(32'hbb5d174f),
	.w8(32'h3c38bb8a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2609e3),
	.w1(32'hbb784d8e),
	.w2(32'hbb9cbef4),
	.w3(32'hbaecfe0d),
	.w4(32'h3b68e8ab),
	.w5(32'h3bd5f95d),
	.w6(32'h3bb06dd5),
	.w7(32'h3bb9bd37),
	.w8(32'h3b2d9683),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba959b3c),
	.w1(32'hbb914bb1),
	.w2(32'h3c4b9d0c),
	.w3(32'h3bc610f9),
	.w4(32'hbb502d8b),
	.w5(32'h3ca9c906),
	.w6(32'hbbc0c332),
	.w7(32'hbbe302c6),
	.w8(32'h3bc94bdb),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c115e92),
	.w1(32'h3b3b737d),
	.w2(32'hbb95c8b7),
	.w3(32'hbad16bcf),
	.w4(32'hbcb5edde),
	.w5(32'h3c01bc0b),
	.w6(32'hbc61beb4),
	.w7(32'hbd06cecd),
	.w8(32'h398928da),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab02a58),
	.w1(32'h3ab735b1),
	.w2(32'hbb5cacd1),
	.w3(32'h3ad59995),
	.w4(32'h385e5474),
	.w5(32'hbc98328e),
	.w6(32'hbbb38bd0),
	.w7(32'hbb80d202),
	.w8(32'hbd115958),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe83ae6),
	.w1(32'h3a2524a8),
	.w2(32'h3b2409f4),
	.w3(32'h3ac2dfe2),
	.w4(32'h3cb020d1),
	.w5(32'hb9cf844b),
	.w6(32'hbbad3961),
	.w7(32'h3cb748b0),
	.w8(32'hb9d89533),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12d0a0),
	.w1(32'h3b606c29),
	.w2(32'h3bf2fe96),
	.w3(32'hbaa93a6a),
	.w4(32'h3ac256d9),
	.w5(32'h3c456598),
	.w6(32'hbb203b75),
	.w7(32'h3b1b9fe2),
	.w8(32'h3c11811c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd93dc),
	.w1(32'hbc304541),
	.w2(32'hbc9aea22),
	.w3(32'hba7b79bd),
	.w4(32'hbc052e66),
	.w5(32'hbc70f5d3),
	.w6(32'hbb2cd02b),
	.w7(32'hbbb4509b),
	.w8(32'h3b1c3fdf),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc98997),
	.w1(32'hb8ed676f),
	.w2(32'hbc225057),
	.w3(32'hbc1a4fba),
	.w4(32'hbac4f7d8),
	.w5(32'h3ba22c2d),
	.w6(32'h3c265486),
	.w7(32'hb912db4e),
	.w8(32'h3b970692),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36e41e),
	.w1(32'hbba20cf5),
	.w2(32'hbc0e2508),
	.w3(32'hbb2109fc),
	.w4(32'hbc1bd883),
	.w5(32'hbbb24401),
	.w6(32'h3bac0c33),
	.w7(32'hbc64b455),
	.w8(32'hbbbf5f0b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba26618),
	.w1(32'h3bdfa761),
	.w2(32'h3c017cda),
	.w3(32'hbb9c2ead),
	.w4(32'h3bc51569),
	.w5(32'h3c10cfd6),
	.w6(32'hbb9ef91d),
	.w7(32'h3b85482e),
	.w8(32'h3c09a218),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb128fdc),
	.w1(32'h3c1c846c),
	.w2(32'hbb8a2d28),
	.w3(32'h3ab5306e),
	.w4(32'h3c1a6492),
	.w5(32'h3b78c477),
	.w6(32'hbc018125),
	.w7(32'h3bfbc74c),
	.w8(32'h3bcf024d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb49be4),
	.w1(32'h3b1423c1),
	.w2(32'hba2cefa0),
	.w3(32'hbaedd7ef),
	.w4(32'h3b9d9a7a),
	.w5(32'hbb9316d8),
	.w6(32'h3ac308b7),
	.w7(32'h3b87be25),
	.w8(32'hbb480ef3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c2269),
	.w1(32'h3bc388bb),
	.w2(32'hbc2d63b7),
	.w3(32'h3b2aa67d),
	.w4(32'hbc09d723),
	.w5(32'hbcc51a87),
	.w6(32'hbbb7cc68),
	.w7(32'hbb8fd581),
	.w8(32'hbcbd298a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91c5ca),
	.w1(32'h3aa85c6b),
	.w2(32'hbac339af),
	.w3(32'hbbf23eac),
	.w4(32'h3d03e8e9),
	.w5(32'hb9ad2ce4),
	.w6(32'hbc73b16d),
	.w7(32'h3ccaead3),
	.w8(32'h397031e1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ab38c),
	.w1(32'h3b73f3c9),
	.w2(32'h3bf928f7),
	.w3(32'hba979cc3),
	.w4(32'h3b5e8776),
	.w5(32'hb9f2e8d3),
	.w6(32'h3b8b06f1),
	.w7(32'h3be8a221),
	.w8(32'hbaaac1ca),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a983e3e),
	.w1(32'hb995a6f1),
	.w2(32'h3b8b4cfd),
	.w3(32'h3b299239),
	.w4(32'hbb2b06de),
	.w5(32'h3c1bdca0),
	.w6(32'h3af867a0),
	.w7(32'h3aca0988),
	.w8(32'h3b8e7201),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6cf56f),
	.w1(32'hbc25c963),
	.w2(32'h3ab19418),
	.w3(32'h3c53ce32),
	.w4(32'h3c1c2d36),
	.w5(32'h39c58285),
	.w6(32'h3bcc19e7),
	.w7(32'h3ba5113c),
	.w8(32'hbaf88f7b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cd519),
	.w1(32'hbb73adcb),
	.w2(32'hbba1e0a8),
	.w3(32'h3c70a3b3),
	.w4(32'h3c5994d7),
	.w5(32'h3b3ea5b1),
	.w6(32'hba66250f),
	.w7(32'h3c430905),
	.w8(32'hbbcdc6ce),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ba0c2),
	.w1(32'hbc15e75e),
	.w2(32'hbb7362e6),
	.w3(32'hbaed4cfd),
	.w4(32'hbc3fe4df),
	.w5(32'hbba51805),
	.w6(32'hbbd7d08c),
	.w7(32'hbbcbae07),
	.w8(32'hbb7644d4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42a078),
	.w1(32'hbb633fe1),
	.w2(32'hbc546cb0),
	.w3(32'hbaed8e23),
	.w4(32'hbb92e2ba),
	.w5(32'hbbb0deb6),
	.w6(32'h3a990e69),
	.w7(32'hb8fd86cb),
	.w8(32'hbb09a6f1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d2783),
	.w1(32'hbb772f90),
	.w2(32'hbb3bff96),
	.w3(32'hbbe4a7a3),
	.w4(32'h3b0b301a),
	.w5(32'hb93fa4dd),
	.w6(32'hbb8e48ee),
	.w7(32'h3b1f934b),
	.w8(32'hbb6cb4a7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4162f4),
	.w1(32'hbb81a30c),
	.w2(32'hbbc12f7b),
	.w3(32'hbae27ca8),
	.w4(32'hbb66be3c),
	.w5(32'h3c5ebbe1),
	.w6(32'hbb9182f6),
	.w7(32'hbb8fb56f),
	.w8(32'h3cfd037a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23a669),
	.w1(32'h3c1d66fb),
	.w2(32'hbb4761ac),
	.w3(32'h3ca380bf),
	.w4(32'h3c30528d),
	.w5(32'h3c034d1a),
	.w6(32'h3ce96b97),
	.w7(32'h3af368a3),
	.w8(32'h3a5c0dc8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4480bf),
	.w1(32'h3ac951f2),
	.w2(32'h3b5f6d71),
	.w3(32'h3b6ee341),
	.w4(32'hbc539fab),
	.w5(32'h3c37224b),
	.w6(32'hbbb74798),
	.w7(32'hbb185bdd),
	.w8(32'h3c030302),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38ad3a),
	.w1(32'h3b878151),
	.w2(32'hbb2959bf),
	.w3(32'h3c7736e7),
	.w4(32'hbc7f6e86),
	.w5(32'h3c39e6ca),
	.w6(32'hbbd3361c),
	.w7(32'hbc8bdb92),
	.w8(32'h3b88339f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8217a),
	.w1(32'hba453ae5),
	.w2(32'h3b5964eb),
	.w3(32'hbc98b1ff),
	.w4(32'h3b22da79),
	.w5(32'h3b6bda1f),
	.w6(32'h3b11483a),
	.w7(32'h3aeaec5d),
	.w8(32'h3b939222),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb995d8d),
	.w1(32'h3ba5b524),
	.w2(32'hbb0b7b0c),
	.w3(32'hbb200520),
	.w4(32'h3c045c54),
	.w5(32'hbb682f09),
	.w6(32'hbbb0963a),
	.w7(32'h3b058a67),
	.w8(32'hbbc619ff),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdaf0a),
	.w1(32'h3aadc270),
	.w2(32'h3b2440d4),
	.w3(32'hbb112dd2),
	.w4(32'hbb46d81b),
	.w5(32'h3bf1c38f),
	.w6(32'hbbd62c63),
	.w7(32'hbb6d390d),
	.w8(32'h3ca0f132),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb054c7a),
	.w1(32'hbc4947ec),
	.w2(32'h3a50a802),
	.w3(32'hbbbb9d1c),
	.w4(32'hbcac4f56),
	.w5(32'hbaa7372a),
	.w6(32'h3c41da7c),
	.w7(32'hbcb317f3),
	.w8(32'hbbb8d2ca),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d39ef),
	.w1(32'hbbf03aa1),
	.w2(32'h3b274425),
	.w3(32'hbc1ba1a3),
	.w4(32'h38fd13da),
	.w5(32'h3c5cb5e4),
	.w6(32'hbc0a9e1c),
	.w7(32'h3b8d6830),
	.w8(32'h3c88542d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0562b6),
	.w1(32'hba842962),
	.w2(32'h3c13a731),
	.w3(32'hbba21c65),
	.w4(32'hbbe3a894),
	.w5(32'h3cae429e),
	.w6(32'hbbdfc5fe),
	.w7(32'hbc1fb261),
	.w8(32'h3cba0277),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0957c),
	.w1(32'hbb46fb5b),
	.w2(32'hbbcf7663),
	.w3(32'h3c0b1cca),
	.w4(32'h3bbd7a71),
	.w5(32'hbb2638af),
	.w6(32'h3c436b64),
	.w7(32'h3bdc4bcf),
	.w8(32'hbb8afc53),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc6177),
	.w1(32'h3b60197c),
	.w2(32'h3c04dd55),
	.w3(32'hbbaf5f6d),
	.w4(32'hbb7beb02),
	.w5(32'h3bf2ac67),
	.w6(32'hbbf79552),
	.w7(32'hbba662f3),
	.w8(32'h3bd39d5c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa23ca2),
	.w1(32'hbbaf5a53),
	.w2(32'h3a4e55e5),
	.w3(32'hba637e3a),
	.w4(32'hbb390e60),
	.w5(32'h3c5435e0),
	.w6(32'hba88e541),
	.w7(32'hb99d2e02),
	.w8(32'h3c461e63),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78a5f20),
	.w1(32'hbc16675f),
	.w2(32'hbb169020),
	.w3(32'hb9a963d9),
	.w4(32'hbc9887a5),
	.w5(32'hbc2f1281),
	.w6(32'hba0dac66),
	.w7(32'hbc6ccdcf),
	.w8(32'h3b674bd4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39edee67),
	.w1(32'h3ca25028),
	.w2(32'h3bb58227),
	.w3(32'h39cb7c23),
	.w4(32'h3c6142de),
	.w5(32'h3bcf2269),
	.w6(32'hba792d7b),
	.w7(32'hbb9d6b3e),
	.w8(32'hbb7a3469),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bbe50),
	.w1(32'h3a93d9bc),
	.w2(32'h3c8bba0d),
	.w3(32'hb98aa5fa),
	.w4(32'hbc2d7e72),
	.w5(32'h3cc0974e),
	.w6(32'h3977ec2e),
	.w7(32'hbb6c390b),
	.w8(32'h3c795c66),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0741e),
	.w1(32'hbbdb99bd),
	.w2(32'hbbb2d75d),
	.w3(32'h3b65adb5),
	.w4(32'hbcb6b355),
	.w5(32'h3a4b87e2),
	.w6(32'hbc156f2c),
	.w7(32'hbcb23276),
	.w8(32'hbc20165e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ef7f9),
	.w1(32'hbc9585da),
	.w2(32'hbbb50edc),
	.w3(32'h3b9b75d4),
	.w4(32'hbc0ee876),
	.w5(32'h3bd6c172),
	.w6(32'h3bb19efa),
	.w7(32'h3be315b2),
	.w8(32'h3c128c2f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab423b0),
	.w1(32'h3aabbe75),
	.w2(32'hbccaf536),
	.w3(32'h3af8f6df),
	.w4(32'hbb8120cf),
	.w5(32'hbd3889ad),
	.w6(32'h3ba46a74),
	.w7(32'h3b126ed7),
	.w8(32'hbcc9e2c1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c2f53),
	.w1(32'h3c9213a1),
	.w2(32'h3ac5ad11),
	.w3(32'hbc01924e),
	.w4(32'h3d228b1a),
	.w5(32'hbd1a2c91),
	.w6(32'hbbc1726b),
	.w7(32'h3d2522ab),
	.w8(32'hbd08cb77),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3810690a),
	.w1(32'h3c20b2f0),
	.w2(32'hbbefeef9),
	.w3(32'hbb3c8a54),
	.w4(32'h3d43f9f9),
	.w5(32'hbb896fb9),
	.w6(32'h3b2f617a),
	.w7(32'h3d3f3e0f),
	.w8(32'hba555b25),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabfa1c),
	.w1(32'h3ba564da),
	.w2(32'hbc4b36e7),
	.w3(32'h3bd10798),
	.w4(32'h3b9e66c1),
	.w5(32'hbbb84c33),
	.w6(32'h3b4d9726),
	.w7(32'h3c1cbb4a),
	.w8(32'hb7bdd855),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdefca),
	.w1(32'hbac68af0),
	.w2(32'hbbaa7d24),
	.w3(32'hbb8ca108),
	.w4(32'hbb4d05b5),
	.w5(32'hbab13856),
	.w6(32'hbb80a462),
	.w7(32'h39b523ed),
	.w8(32'h3bf7f890),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3751e),
	.w1(32'hbc05c00d),
	.w2(32'hbc2bc6b1),
	.w3(32'hbb24ccc3),
	.w4(32'hbb65e5fb),
	.w5(32'hb5eeff58),
	.w6(32'h3b252bc4),
	.w7(32'h3b8912fa),
	.w8(32'h3b898de7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb7482),
	.w1(32'h3b4bbd24),
	.w2(32'hbbb3381e),
	.w3(32'h3a5ac140),
	.w4(32'h399013ee),
	.w5(32'hbab79026),
	.w6(32'hbadca8c5),
	.w7(32'hba52794a),
	.w8(32'hba40e668),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2da51c),
	.w1(32'h3bac2315),
	.w2(32'hbaebba12),
	.w3(32'hbad55323),
	.w4(32'h3b84f0f1),
	.w5(32'hbbe87c5a),
	.w6(32'hbb952d51),
	.w7(32'h3b8939ef),
	.w8(32'h3848690f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24ed8e),
	.w1(32'hbb698157),
	.w2(32'h3c09fd69),
	.w3(32'hbbfd1917),
	.w4(32'hbbd83d1b),
	.w5(32'h3c103eea),
	.w6(32'hbc09ca0f),
	.w7(32'hbbb3d865),
	.w8(32'hbbe05ad4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c834c),
	.w1(32'hbb8e23ce),
	.w2(32'hbbb624fc),
	.w3(32'h3c05dbf7),
	.w4(32'hbbb75292),
	.w5(32'hbc8a1a45),
	.w6(32'hbbf57522),
	.w7(32'hbc4364b6),
	.w8(32'hbc5d68e5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a2fdd),
	.w1(32'hb877899b),
	.w2(32'h3c8391c9),
	.w3(32'hbb403550),
	.w4(32'h3ca146a0),
	.w5(32'h3ccd3794),
	.w6(32'h394415fe),
	.w7(32'h3cf57d29),
	.w8(32'h3cbbaaad),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba47bfd),
	.w1(32'hbad64b87),
	.w2(32'hbc0e2581),
	.w3(32'hba8cfc3b),
	.w4(32'hbc360f87),
	.w5(32'hbbc96091),
	.w6(32'hbb3573c1),
	.w7(32'hbc9ae36a),
	.w8(32'hbb2552b2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55821e),
	.w1(32'h3b00c4ea),
	.w2(32'hbac1973c),
	.w3(32'hbc1d7fd3),
	.w4(32'h3aff0795),
	.w5(32'h3c23747f),
	.w6(32'hbbaab59c),
	.w7(32'hbacf4c1b),
	.w8(32'h3c8934dc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03c196),
	.w1(32'h3a4be72f),
	.w2(32'hbb96844c),
	.w3(32'h3b8720ae),
	.w4(32'hbb096116),
	.w5(32'hbb46c3f3),
	.w6(32'h3ca17731),
	.w7(32'hbb8bbe0d),
	.w8(32'h3a9dfe51),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8ed35),
	.w1(32'hbc8eec99),
	.w2(32'hbbcb6542),
	.w3(32'hbb492c36),
	.w4(32'h3c1726d6),
	.w5(32'hbc0af893),
	.w6(32'h3b43964f),
	.w7(32'h3c94182b),
	.w8(32'hbc1a025b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc001f12),
	.w1(32'hbc249a52),
	.w2(32'h3b858ce2),
	.w3(32'hbbcfd420),
	.w4(32'hbc1ae743),
	.w5(32'h3b4c60c6),
	.w6(32'hbbf93012),
	.w7(32'hb80965d6),
	.w8(32'h3b12d998),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f2991),
	.w1(32'h3b9c84e8),
	.w2(32'h3b2d8686),
	.w3(32'hba4ac9f5),
	.w4(32'hbbbd7bf2),
	.w5(32'h3b5beb97),
	.w6(32'hbb6f4b49),
	.w7(32'hbc02bab0),
	.w8(32'h3be7064b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb092cf5),
	.w1(32'hbbc47505),
	.w2(32'hb9c8279a),
	.w3(32'hbb94b88b),
	.w4(32'hbc76b04d),
	.w5(32'h3a52af0b),
	.w6(32'hbb4da7a7),
	.w7(32'hb88442e8),
	.w8(32'h3b70c18a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9da2b8),
	.w1(32'h3b571941),
	.w2(32'h3b158271),
	.w3(32'h3a8f4e11),
	.w4(32'h3a93070f),
	.w5(32'hbbf3619d),
	.w6(32'h39bb3d19),
	.w7(32'h3ae1cd22),
	.w8(32'hbc2b2d01),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a45371),
	.w1(32'h3b4ca975),
	.w2(32'hbb2bf34d),
	.w3(32'h3b199753),
	.w4(32'h3c6852fe),
	.w5(32'hbd0f8f79),
	.w6(32'hbb965f98),
	.w7(32'h3c6efa1d),
	.w8(32'hbd1c80ba),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395e4758),
	.w1(32'h3c06abcc),
	.w2(32'h3a2a6424),
	.w3(32'hbb9b0033),
	.w4(32'h3d4205e7),
	.w5(32'h3c848588),
	.w6(32'h3a82ab4e),
	.w7(32'h3d49ec81),
	.w8(32'h3ca43438),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0ec4a),
	.w1(32'hbbaf7090),
	.w2(32'hba24ecbb),
	.w3(32'h3bac4280),
	.w4(32'hbc9bf66c),
	.w5(32'hbb92c36d),
	.w6(32'h3baa9293),
	.w7(32'hbc938a50),
	.w8(32'hbb7aca3a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d54741),
	.w1(32'h38696fc4),
	.w2(32'hbb4457c6),
	.w3(32'h3a9f140e),
	.w4(32'hba929090),
	.w5(32'hbaf77cdd),
	.w6(32'h3a789e42),
	.w7(32'hbae2cad1),
	.w8(32'hbb53a84d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e601a),
	.w1(32'h3b477ea0),
	.w2(32'hbba48126),
	.w3(32'hbb37e905),
	.w4(32'h3b390bb8),
	.w5(32'h3a46cffb),
	.w6(32'hbbe307bb),
	.w7(32'hbb139528),
	.w8(32'hba980f9b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b405061),
	.w1(32'hbb638e9c),
	.w2(32'h39446d72),
	.w3(32'h3a122c18),
	.w4(32'hbbdb1875),
	.w5(32'hbb31acbf),
	.w6(32'h3ad12ff8),
	.w7(32'hbbaf1d3b),
	.w8(32'hbab655ce),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80303d),
	.w1(32'h3afd67e4),
	.w2(32'hbb881e30),
	.w3(32'hbb8bc87e),
	.w4(32'h3aace9c8),
	.w5(32'hba82230d),
	.w6(32'hbae8cdd4),
	.w7(32'hb8fd08b2),
	.w8(32'h3bca40be),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50ac98),
	.w1(32'hbc2d9c09),
	.w2(32'hbb9fad25),
	.w3(32'h3b198b47),
	.w4(32'hbc567265),
	.w5(32'hbbef03e5),
	.w6(32'h3bdd5d0b),
	.w7(32'hbbcd9c58),
	.w8(32'hbb02528f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbea369),
	.w1(32'h3b7d891d),
	.w2(32'hbc60281e),
	.w3(32'hbbe40a13),
	.w4(32'h3a0cb8f5),
	.w5(32'hbc2ebba5),
	.w6(32'h3b908703),
	.w7(32'hbb82ab4a),
	.w8(32'hbac2ee1c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a368883),
	.w1(32'h3a02f572),
	.w2(32'hbb3a9cc8),
	.w3(32'h3bd7a1bf),
	.w4(32'hbbdbda98),
	.w5(32'hb84e7f5e),
	.w6(32'h3c418f52),
	.w7(32'h3a95258b),
	.w8(32'hbb000b87),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a7f47),
	.w1(32'hbbe29078),
	.w2(32'hbba444f8),
	.w3(32'h3b39c249),
	.w4(32'hbb425611),
	.w5(32'h3b9dc2d8),
	.w6(32'hbb010cdb),
	.w7(32'h3baf3b79),
	.w8(32'h3c0898ee),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdc1d5),
	.w1(32'hbb0ce70c),
	.w2(32'hbb17584b),
	.w3(32'hbb60deef),
	.w4(32'hbbea1b29),
	.w5(32'hbc36a4de),
	.w6(32'h3b0fc01c),
	.w7(32'hbc5a50a8),
	.w8(32'hbc523246),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aadcf),
	.w1(32'h3be4d285),
	.w2(32'hba68d786),
	.w3(32'hbbc6d408),
	.w4(32'h3cc198b8),
	.w5(32'h3ab27465),
	.w6(32'hbb4aad19),
	.w7(32'h3c6d9ee2),
	.w8(32'h3c957fe8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc380411),
	.w1(32'hbc09d3dc),
	.w2(32'h3bc4c8bf),
	.w3(32'h3bc04197),
	.w4(32'hbb00b86f),
	.w5(32'h3b153c1e),
	.w6(32'h3c8e0f3e),
	.w7(32'h3bc32974),
	.w8(32'h3b7861cd),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfe285),
	.w1(32'h3a8a3227),
	.w2(32'hbc2f09c9),
	.w3(32'h3c8a545d),
	.w4(32'h3c1496ad),
	.w5(32'hbc3a3e8f),
	.w6(32'hbb9824b6),
	.w7(32'hbab9b625),
	.w8(32'h3b85bc1f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd06721),
	.w1(32'h3c6985ea),
	.w2(32'hbbe817d2),
	.w3(32'hbb11caab),
	.w4(32'h3cf7fc77),
	.w5(32'hbb936933),
	.w6(32'h3c2873d9),
	.w7(32'h3cf665f5),
	.w8(32'hbbc81cbb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3ee91),
	.w1(32'hbc204d36),
	.w2(32'hbc6c4a7e),
	.w3(32'hbb7074ad),
	.w4(32'hbb89f5c4),
	.w5(32'hbba20e7c),
	.w6(32'hb98a7f8e),
	.w7(32'h3ae3c286),
	.w8(32'h3a47e1ed),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af07227),
	.w1(32'h3be91f8a),
	.w2(32'h3b29c6ad),
	.w3(32'h3ba1d70b),
	.w4(32'hbaac271d),
	.w5(32'hb817b5c0),
	.w6(32'h3b65af45),
	.w7(32'hbb3e9ee7),
	.w8(32'hbb20a1c7),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c34c1),
	.w1(32'hbb5e0889),
	.w2(32'hbc520e5e),
	.w3(32'h3b0622ac),
	.w4(32'h3b541934),
	.w5(32'hbb850ef5),
	.w6(32'hbb8773bc),
	.w7(32'h3b650045),
	.w8(32'hbb0668d5),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ce79d),
	.w1(32'hbbe03d62),
	.w2(32'hbb30610d),
	.w3(32'hbc4ded74),
	.w4(32'hbc1db3e0),
	.w5(32'h3af947ae),
	.w6(32'hbbb3ee0d),
	.w7(32'hbb906fcf),
	.w8(32'h3b6dd8fa),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3c45d),
	.w1(32'h3baabb23),
	.w2(32'h3a510535),
	.w3(32'h3b85da14),
	.w4(32'h3ba2a2ab),
	.w5(32'hbb620aa9),
	.w6(32'h3b38a3ef),
	.w7(32'h3b8c03a8),
	.w8(32'h3bd612fe),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02ea6a),
	.w1(32'h3b0a38fa),
	.w2(32'hbba034b0),
	.w3(32'hba98eed5),
	.w4(32'h3b847c26),
	.w5(32'hbaa9f6a1),
	.w6(32'h3cb18005),
	.w7(32'h3cd5eb98),
	.w8(32'h38539cf3),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ebca9),
	.w1(32'h3a20a0ef),
	.w2(32'h3b736fcd),
	.w3(32'h38f8a6ab),
	.w4(32'h3a793a25),
	.w5(32'h3c0d0334),
	.w6(32'h3b5261ed),
	.w7(32'h3b8eb90f),
	.w8(32'h3bc29f37),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6dfaa),
	.w1(32'h3c2c5c29),
	.w2(32'h3c0aa4f7),
	.w3(32'hbbeee066),
	.w4(32'hba84b47d),
	.w5(32'hbc84b561),
	.w6(32'hbc3b759e),
	.w7(32'hba4f765d),
	.w8(32'hbbc9979a),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60ab4b),
	.w1(32'h3cdbb277),
	.w2(32'hb9b02818),
	.w3(32'h3bf14e9d),
	.w4(32'h3ced9e7c),
	.w5(32'hbb4199ed),
	.w6(32'hbc5cdecb),
	.w7(32'h3ac27b32),
	.w8(32'hbabe5041),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e04603),
	.w1(32'h3a956903),
	.w2(32'h3bc7a106),
	.w3(32'hbb17cd75),
	.w4(32'h39dbc30f),
	.w5(32'h3bc6cbbe),
	.w6(32'hbbaa2678),
	.w7(32'hbb86b96f),
	.w8(32'h3bbfe691),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e3227),
	.w1(32'h3b2dad1e),
	.w2(32'hbae64d56),
	.w3(32'h3b5559c7),
	.w4(32'h3a8d6556),
	.w5(32'hbaf83ebe),
	.w6(32'h3b29bc99),
	.w7(32'h3ac31683),
	.w8(32'h393916b5),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8dbe0),
	.w1(32'h3b3af907),
	.w2(32'h3b7f3a63),
	.w3(32'hbb7fc6c9),
	.w4(32'h3be4e5ac),
	.w5(32'h3c8313b2),
	.w6(32'hba9f6bac),
	.w7(32'h3c183ed8),
	.w8(32'h3c3d0373),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbede82f),
	.w1(32'h3bec8da2),
	.w2(32'h3c80bd09),
	.w3(32'h39c8a6ed),
	.w4(32'hba84f836),
	.w5(32'h3c75e806),
	.w6(32'hbb9228c1),
	.w7(32'h3bb6d7f6),
	.w8(32'h3c340ca4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c287bfd),
	.w1(32'hbb71a766),
	.w2(32'hbbcd7eb8),
	.w3(32'h3c2097a1),
	.w4(32'h3987f7c5),
	.w5(32'h3a2eb931),
	.w6(32'h3c01d617),
	.w7(32'hbb358766),
	.w8(32'hbaa9f90c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c780a),
	.w1(32'h3c07251f),
	.w2(32'h3c80c5c6),
	.w3(32'h3b101bf0),
	.w4(32'h3bd1a604),
	.w5(32'h3cd4fdfc),
	.w6(32'h3a9dacca),
	.w7(32'h3c2837ba),
	.w8(32'h3bf5e26b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a8c0c),
	.w1(32'hbc17634b),
	.w2(32'hbbc7fa8d),
	.w3(32'h3c25dd3f),
	.w4(32'hbc9d53e0),
	.w5(32'hb9fe7020),
	.w6(32'h3b83b838),
	.w7(32'hbcd311a2),
	.w8(32'hbb9daaa6),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf095e8),
	.w1(32'hbb643782),
	.w2(32'hbc00debe),
	.w3(32'hbb9c5fa8),
	.w4(32'hbc2ed845),
	.w5(32'hbbf27036),
	.w6(32'h3b52a451),
	.w7(32'h399621b8),
	.w8(32'hbc0240c2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf32bf2),
	.w1(32'hbb589e45),
	.w2(32'hbc3cc5b7),
	.w3(32'hba54aa0f),
	.w4(32'hbb516836),
	.w5(32'h3c148332),
	.w6(32'hba412a96),
	.w7(32'hb9062996),
	.w8(32'h3c2ecf83),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e837c),
	.w1(32'h3aee1b3d),
	.w2(32'hbc38e1bc),
	.w3(32'hbb1f65e7),
	.w4(32'hba6abfe9),
	.w5(32'hbbadd63a),
	.w6(32'hbc1d9675),
	.w7(32'h3af45f7e),
	.w8(32'h3bf17a07),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c2c47),
	.w1(32'h3bb60ec4),
	.w2(32'h3be8df0d),
	.w3(32'hbabd2037),
	.w4(32'h3c478b60),
	.w5(32'h3c4e9c44),
	.w6(32'hbb8f8369),
	.w7(32'hbc0d68ec),
	.w8(32'h3c58fca2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafa507),
	.w1(32'hbbbd06c6),
	.w2(32'h3a660fa1),
	.w3(32'h3c922df7),
	.w4(32'hbbcff5ff),
	.w5(32'h3ae77de0),
	.w6(32'h3c45d792),
	.w7(32'hbb23bf5c),
	.w8(32'h38fb4ae4),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d016c),
	.w1(32'h3b0ae87a),
	.w2(32'h3b65a7dc),
	.w3(32'hbad38b33),
	.w4(32'h3b840e85),
	.w5(32'h3b14b21a),
	.w6(32'hbb6fd43c),
	.w7(32'h3b27bbc4),
	.w8(32'h3b297b81),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39806e6e),
	.w1(32'h3a58240f),
	.w2(32'hbbe53ee3),
	.w3(32'h3ba06399),
	.w4(32'h3b837fb8),
	.w5(32'h385e06d9),
	.w6(32'h3b68192b),
	.w7(32'h3b84daff),
	.w8(32'h3aa1d1cd),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17ec49),
	.w1(32'hbc0fb9c5),
	.w2(32'h3b4fce54),
	.w3(32'hbc0c12e6),
	.w4(32'h39446dbc),
	.w5(32'hb9eb7949),
	.w6(32'hb99ccd82),
	.w7(32'h3b32cab4),
	.w8(32'hbb625b44),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7936ca),
	.w1(32'h3a2d116d),
	.w2(32'hbc24e7ae),
	.w3(32'hbb865416),
	.w4(32'hbaa33f23),
	.w5(32'hbc1dd5ea),
	.w6(32'hbbda1476),
	.w7(32'hbb0f6c0d),
	.w8(32'hbb9d854c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7f001),
	.w1(32'hb794c5c2),
	.w2(32'hbc0c1756),
	.w3(32'hbc81c018),
	.w4(32'hbc40d813),
	.w5(32'hbc93d101),
	.w6(32'hbc112ab7),
	.w7(32'hbc4e2873),
	.w8(32'hbc89d1fb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be23a),
	.w1(32'hbaef46d1),
	.w2(32'hbb737f5b),
	.w3(32'hbc52ca36),
	.w4(32'hbb4bd2a2),
	.w5(32'hba9d25d1),
	.w6(32'hbc900ba8),
	.w7(32'hbc98e8ca),
	.w8(32'hbb0a0296),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a3f93),
	.w1(32'h3b02adaf),
	.w2(32'hbb9c323e),
	.w3(32'h3ac07452),
	.w4(32'h3ad9f7d3),
	.w5(32'hbab9053f),
	.w6(32'h3b3a682a),
	.w7(32'h3b540699),
	.w8(32'h3b270c2a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45fc3a),
	.w1(32'hbb2bf0e0),
	.w2(32'hbb0fd6ef),
	.w3(32'hbb5e0116),
	.w4(32'hbb85c291),
	.w5(32'hbabeed26),
	.w6(32'hbbcdc6b6),
	.w7(32'hbb5069e9),
	.w8(32'hba9fba8d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36962e),
	.w1(32'hba164b1d),
	.w2(32'h3b92225f),
	.w3(32'hbb1d9459),
	.w4(32'hbac244b9),
	.w5(32'h3981006d),
	.w6(32'h3a2e62ed),
	.w7(32'hba3d4d9d),
	.w8(32'hbc163d31),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a719e5),
	.w1(32'hb9d609d2),
	.w2(32'hbbfa600b),
	.w3(32'h3b6f16e8),
	.w4(32'hb94ba83d),
	.w5(32'hbb5237f7),
	.w6(32'h3a61a429),
	.w7(32'h3a61e3ae),
	.w8(32'hbc08f6a5),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb911089),
	.w1(32'hbbedba96),
	.w2(32'hbc496b84),
	.w3(32'h3859a83c),
	.w4(32'hbb54b4bc),
	.w5(32'hbc074c09),
	.w6(32'hba150077),
	.w7(32'hbba5d7e4),
	.w8(32'h39a7ce1a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc754dbb),
	.w1(32'hbaa8bf1e),
	.w2(32'hba8f77a7),
	.w3(32'hbc45f6b7),
	.w4(32'hbbdcafb6),
	.w5(32'h3b801ecb),
	.w6(32'hbc66f24e),
	.w7(32'hbc6eb1e5),
	.w8(32'h3b2ebee2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a948af5),
	.w1(32'h3ba7dd22),
	.w2(32'hbab6115a),
	.w3(32'h3b9acd5c),
	.w4(32'h3bb38afb),
	.w5(32'h3ab9954c),
	.w6(32'h38efdddd),
	.w7(32'h3a564359),
	.w8(32'h3a9d6e5a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbb060),
	.w1(32'hb9f2dc45),
	.w2(32'hbc6ea69e),
	.w3(32'hba8d371d),
	.w4(32'h3b13e817),
	.w5(32'hbc8f88cc),
	.w6(32'h3aaa704b),
	.w7(32'h3a98ce49),
	.w8(32'hbca36fe9),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a1970),
	.w1(32'h3bc458d3),
	.w2(32'hbc30c18f),
	.w3(32'hbc3167a5),
	.w4(32'hbb95250f),
	.w5(32'hbc812254),
	.w6(32'hbc7502db),
	.w7(32'hbc7b5f78),
	.w8(32'hbbc0cdfb),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43ddb5),
	.w1(32'h3b96a127),
	.w2(32'hbbd784eb),
	.w3(32'hbc40eceb),
	.w4(32'hbc24e9dd),
	.w5(32'hbac9fa0d),
	.w6(32'hbc673e12),
	.w7(32'hbbf356ee),
	.w8(32'h3ad582f2),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0c15f),
	.w1(32'hbbd42495),
	.w2(32'hbbe25fcf),
	.w3(32'hbb00f517),
	.w4(32'hbb3837de),
	.w5(32'hbb495e03),
	.w6(32'h3b416228),
	.w7(32'hb986521a),
	.w8(32'hba8a9fdf),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4871ab),
	.w1(32'hbba5d974),
	.w2(32'hbbb8f477),
	.w3(32'hbbb2661f),
	.w4(32'h3aa1ec1e),
	.w5(32'h3b8ff608),
	.w6(32'hbb362ccc),
	.w7(32'h3b836d3e),
	.w8(32'h3ada59a1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabe3fd),
	.w1(32'hbb79bc8d),
	.w2(32'hbc63fbd6),
	.w3(32'h3bd37f62),
	.w4(32'h3b52d42e),
	.w5(32'hbbd33ac9),
	.w6(32'h3b2856b2),
	.w7(32'h3bd53283),
	.w8(32'hbc07d669),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3235c6),
	.w1(32'hbc15a31b),
	.w2(32'hbc785ed2),
	.w3(32'hba8fc64a),
	.w4(32'hbc222a0c),
	.w5(32'hbc974856),
	.w6(32'hbb8ae463),
	.w7(32'hbc3a592e),
	.w8(32'hbc34fbbb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3dfd32),
	.w1(32'h3b5b52f3),
	.w2(32'hbb920d18),
	.w3(32'hbc6006fc),
	.w4(32'hbbd1ba8b),
	.w5(32'hbb21ff7c),
	.w6(32'hbc4ee49e),
	.w7(32'hbc7c611b),
	.w8(32'hb9f94fda),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb91917),
	.w1(32'hbb9d3eaf),
	.w2(32'hbb426519),
	.w3(32'hb9e554e2),
	.w4(32'hbafcb6a0),
	.w5(32'hbbd08218),
	.w6(32'h3addec35),
	.w7(32'hba282ada),
	.w8(32'hbb1d22f8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2ae51),
	.w1(32'h3bd6c32b),
	.w2(32'h3b16d817),
	.w3(32'hbbca9be9),
	.w4(32'hb8b469f7),
	.w5(32'h38a9b0f1),
	.w6(32'hbb0a5d63),
	.w7(32'h3b7bc929),
	.w8(32'h3b8de950),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3140c9),
	.w1(32'hbaaeed57),
	.w2(32'h3be62529),
	.w3(32'hbba2c5d5),
	.w4(32'h39faf999),
	.w5(32'h3bc31bf2),
	.w6(32'h3b8e1485),
	.w7(32'h3bf0e4c8),
	.w8(32'hbb1554ca),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ed420),
	.w1(32'h3b17746e),
	.w2(32'h3ac437c8),
	.w3(32'h3b363ea0),
	.w4(32'hb8d4451c),
	.w5(32'hb878277e),
	.w6(32'hbc253b12),
	.w7(32'hbb1d4568),
	.w8(32'h3bfa4771),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10dbf7),
	.w1(32'hbb2793d0),
	.w2(32'hb8e36daa),
	.w3(32'hbb569933),
	.w4(32'h3ac9ae90),
	.w5(32'h3ba18f63),
	.w6(32'hbade54b4),
	.w7(32'h3ba52391),
	.w8(32'h3a2e8810),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3d0a3),
	.w1(32'h3c2e48dd),
	.w2(32'h3aba2b2d),
	.w3(32'h3bca27ad),
	.w4(32'h3b4fc2ea),
	.w5(32'h3b8bb584),
	.w6(32'h3be86713),
	.w7(32'h3c0cbf5a),
	.w8(32'hbbda1043),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad6d5c),
	.w1(32'h3be10441),
	.w2(32'hbabbdf05),
	.w3(32'h3b81bb8b),
	.w4(32'h3c145410),
	.w5(32'hbb5a47c2),
	.w6(32'hbb1f3c43),
	.w7(32'h3bd4764d),
	.w8(32'h3b8db413),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab21c5e),
	.w1(32'h3b825c73),
	.w2(32'hbc210d18),
	.w3(32'h38051d47),
	.w4(32'h3ba99445),
	.w5(32'h3894f7e1),
	.w6(32'hb9cc2b43),
	.w7(32'h3a369d9a),
	.w8(32'h3a5a7ecf),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98aa9b),
	.w1(32'hb9b1ccae),
	.w2(32'h3a8a2360),
	.w3(32'hbcb5a262),
	.w4(32'hbc269ff8),
	.w5(32'h3a94a0d0),
	.w6(32'hbc19d8ce),
	.w7(32'hbc796d1d),
	.w8(32'hbb4b5d59),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c015344),
	.w1(32'h3bd1eeaa),
	.w2(32'hbb8ba9ee),
	.w3(32'h3bbfac7d),
	.w4(32'h3c002a6a),
	.w5(32'hbb3f2f4f),
	.w6(32'h3b2fe579),
	.w7(32'h3bce2a62),
	.w8(32'h3bf38b03),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e36267),
	.w1(32'hbbb1da06),
	.w2(32'hbc022530),
	.w3(32'h3a971dda),
	.w4(32'hbbb67d48),
	.w5(32'hbc59ca94),
	.w6(32'h3c094510),
	.w7(32'h3a22273c),
	.w8(32'hbb5ec39c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc068ba6),
	.w1(32'hbba71bc1),
	.w2(32'hbc0de5c9),
	.w3(32'hbba4c8a6),
	.w4(32'hbb6cce06),
	.w5(32'hbbf87c02),
	.w6(32'h3b066527),
	.w7(32'h3b3d1129),
	.w8(32'hbc1b35e4),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31294d),
	.w1(32'h3c5cd462),
	.w2(32'hbc82056b),
	.w3(32'h3bd92dd8),
	.w4(32'h3ca16f1c),
	.w5(32'hbc4559e8),
	.w6(32'hbc33f104),
	.w7(32'h3c67f51f),
	.w8(32'hbbb45a23),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf3e07),
	.w1(32'hbb7e0b40),
	.w2(32'h3b80229f),
	.w3(32'hbb1cb539),
	.w4(32'hbb8ce9aa),
	.w5(32'hbb0dac63),
	.w6(32'h3aa423d9),
	.w7(32'hbbf00370),
	.w8(32'hbb493ee8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcde6d5),
	.w1(32'hb9b007d9),
	.w2(32'h3baa68d5),
	.w3(32'h3c069fa4),
	.w4(32'h3a71f6d6),
	.w5(32'h3c1382d0),
	.w6(32'h3ba3e578),
	.w7(32'h3b4861f4),
	.w8(32'h3b4ee733),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c354dc5),
	.w1(32'h3c0285fb),
	.w2(32'h3b9dc384),
	.w3(32'h3c7ffeb8),
	.w4(32'h3c2b38b0),
	.w5(32'h3baa8b03),
	.w6(32'h3c1c3e8e),
	.w7(32'h3ba4bf5a),
	.w8(32'h3a03d94f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f44c71),
	.w1(32'h3acb1331),
	.w2(32'h3c6062ec),
	.w3(32'hba62a5ad),
	.w4(32'hbb49dae0),
	.w5(32'h3c416481),
	.w6(32'hbbb996dd),
	.w7(32'hbbe2b304),
	.w8(32'h3bee436c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c931b9f),
	.w1(32'h3c4929e6),
	.w2(32'hbbc8c601),
	.w3(32'h3c9df86e),
	.w4(32'h3c5decb5),
	.w5(32'h3997dc4f),
	.w6(32'h3c4ad0fd),
	.w7(32'h3c4db260),
	.w8(32'h3a576975),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e51d5),
	.w1(32'hbbab494c),
	.w2(32'hbbdf4eab),
	.w3(32'h3b81bf58),
	.w4(32'h39bafb77),
	.w5(32'hbbde3351),
	.w6(32'h3b9f12a9),
	.w7(32'h3b0201f1),
	.w8(32'hbc097f04),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e117b),
	.w1(32'hbb88d3c9),
	.w2(32'hb9c8f0a7),
	.w3(32'hbc1c35bf),
	.w4(32'hb8532c59),
	.w5(32'hbb0fbfb1),
	.w6(32'hbc02b872),
	.w7(32'hba969922),
	.w8(32'h3b832bf0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc18d99),
	.w1(32'h3af775f1),
	.w2(32'h3c010092),
	.w3(32'h3b05b9ec),
	.w4(32'h371a6cba),
	.w5(32'h3c09f4b2),
	.w6(32'h3b85ea91),
	.w7(32'h3b80db01),
	.w8(32'h3bd6ef8a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01f75d),
	.w1(32'h3b4a8460),
	.w2(32'hbcbf6c8e),
	.w3(32'h3c65fe76),
	.w4(32'h3c31ee4e),
	.w5(32'hbc682878),
	.w6(32'h3c4a15d8),
	.w7(32'h3c35fc89),
	.w8(32'hbb6eb2ab),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7eefa9),
	.w1(32'hbc6a34fd),
	.w2(32'h3a0692e9),
	.w3(32'hbc839b06),
	.w4(32'hbc7fbf0b),
	.w5(32'hbaa371ac),
	.w6(32'hbc2c9afb),
	.w7(32'hbc65ed2f),
	.w8(32'hb99675c1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a6b5b),
	.w1(32'h3c15b7ec),
	.w2(32'hbb8a1df4),
	.w3(32'h3bf2a164),
	.w4(32'h3c01b3fb),
	.w5(32'hbc232e72),
	.w6(32'h3ba07c17),
	.w7(32'h3be86666),
	.w8(32'hbbf58605),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e3b4d),
	.w1(32'hbbb40761),
	.w2(32'hbbbfc402),
	.w3(32'hbc88a70a),
	.w4(32'hbc23e3a6),
	.w5(32'hbb6a3261),
	.w6(32'hbc97b2ce),
	.w7(32'hbc58bfb6),
	.w8(32'hbb0c580c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcff4bf),
	.w1(32'hbbca5bb9),
	.w2(32'hba72a040),
	.w3(32'hbbe5aaba),
	.w4(32'h3a9ab677),
	.w5(32'hba72ee2b),
	.w6(32'hbc224c56),
	.w7(32'hbbc5c00d),
	.w8(32'hba2dc93c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20f882),
	.w1(32'hbaef33f9),
	.w2(32'hbc28adb4),
	.w3(32'hbb751a88),
	.w4(32'h3b02405c),
	.w5(32'hbba5f74a),
	.w6(32'hbb951ada),
	.w7(32'h39c03a39),
	.w8(32'hbbf6b000),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42b621),
	.w1(32'hbb3ffb19),
	.w2(32'h3b6df111),
	.w3(32'hbc292195),
	.w4(32'hba2798ef),
	.w5(32'h3a24a187),
	.w6(32'hbc3b5ef0),
	.w7(32'hba83c3e3),
	.w8(32'hbab60ed3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd75221),
	.w1(32'h3b1ef99a),
	.w2(32'hbaeac2e5),
	.w3(32'hbb2dc7a8),
	.w4(32'hbb42d259),
	.w5(32'hbc0945bf),
	.w6(32'hbc2b03cc),
	.w7(32'hbbde50b5),
	.w8(32'hbc20fd44),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb216df7),
	.w1(32'hbbcde64a),
	.w2(32'hbc5b145a),
	.w3(32'hbc3db249),
	.w4(32'hbbea445e),
	.w5(32'hbbfcb6f7),
	.w6(32'hbc04a88f),
	.w7(32'hbc015464),
	.w8(32'hbbc8ef6b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66592d),
	.w1(32'h39603d03),
	.w2(32'hba389fe8),
	.w3(32'hbc70f7c9),
	.w4(32'hbc1f69a8),
	.w5(32'h3a4e1dbe),
	.w6(32'hbc6d2980),
	.w7(32'hbc4eeff8),
	.w8(32'hba72a0cc),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ee955f),
	.w1(32'hbb0b06ac),
	.w2(32'hbc103766),
	.w3(32'h3b2b3d63),
	.w4(32'h3acc7848),
	.w5(32'hbbeb7137),
	.w6(32'h3b1d9c67),
	.w7(32'h3b008b95),
	.w8(32'hbba061ef),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b02d8),
	.w1(32'hbc2fa72b),
	.w2(32'hbbf176b6),
	.w3(32'hbba08de7),
	.w4(32'hbbde240f),
	.w5(32'hbb2b8192),
	.w6(32'hbb7f1cfb),
	.w7(32'hbb50f9d3),
	.w8(32'hba9b164e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02a8cb),
	.w1(32'hb9bb9aaa),
	.w2(32'h3ad699f8),
	.w3(32'hbafb8153),
	.w4(32'h38958fac),
	.w5(32'h3b47126b),
	.w6(32'hbb4ab814),
	.w7(32'h39f31dfa),
	.w8(32'hbb12ddd7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c9c52),
	.w1(32'h39e5e5c7),
	.w2(32'h3b3bd8a1),
	.w3(32'hbb08a68c),
	.w4(32'hbbaeb7af),
	.w5(32'h3b6f5dfb),
	.w6(32'hba650ab3),
	.w7(32'hbbe66de8),
	.w8(32'h3bc9b896),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c485ddf),
	.w1(32'hbabeb198),
	.w2(32'hbca63faf),
	.w3(32'h3c83e3b9),
	.w4(32'h3c68c199),
	.w5(32'hbb72439f),
	.w6(32'h3c30237e),
	.w7(32'h3bc894cf),
	.w8(32'hbb5f7dc8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc312378),
	.w1(32'hbbd2acaf),
	.w2(32'hbafcb4d4),
	.w3(32'hbc3577c4),
	.w4(32'hbbb5e6b6),
	.w5(32'h38a74745),
	.w6(32'hbaaf9ad0),
	.w7(32'hbb730f8b),
	.w8(32'hbba42736),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e63237),
	.w1(32'h3b078f9f),
	.w2(32'h3b45c715),
	.w3(32'hbb1b9355),
	.w4(32'h3bea82fa),
	.w5(32'h3bedb374),
	.w6(32'hbb9e3af6),
	.w7(32'h3bcce381),
	.w8(32'h3beb0493),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be82ea8),
	.w1(32'h3b13d289),
	.w2(32'hbbb412bf),
	.w3(32'h3c550834),
	.w4(32'h3b22f693),
	.w5(32'hbb548e64),
	.w6(32'h3c2675c7),
	.w7(32'h3b9a36e9),
	.w8(32'hba769893),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac59cb9),
	.w1(32'hbafe3124),
	.w2(32'h3b083e97),
	.w3(32'hbb6b46ed),
	.w4(32'hbb05429e),
	.w5(32'h3ab36cfd),
	.w6(32'hbb064243),
	.w7(32'h39292321),
	.w8(32'h3c02878c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a289d),
	.w1(32'h3aa25a44),
	.w2(32'h3bab40d3),
	.w3(32'h3ab79893),
	.w4(32'hbaaeb26e),
	.w5(32'h3c201b69),
	.w6(32'h3ba1763f),
	.w7(32'h3bda1e57),
	.w8(32'h3c1821db),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0537f1),
	.w1(32'h3bd04b40),
	.w2(32'h3b13a5f5),
	.w3(32'h3c75d9e4),
	.w4(32'h3c4ca9a1),
	.w5(32'h3c22255f),
	.w6(32'h3c9cac9d),
	.w7(32'h3ca57519),
	.w8(32'h3c223657),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc60c69),
	.w1(32'h3bc2a457),
	.w2(32'hbc0fd82f),
	.w3(32'h3cd3ba8f),
	.w4(32'h3c79a2d1),
	.w5(32'h3a548a3a),
	.w6(32'h3caa2b9c),
	.w7(32'h3ca4d0e7),
	.w8(32'h3ae714cf),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1d391),
	.w1(32'h3a8c312e),
	.w2(32'hba6d709d),
	.w3(32'h3c698e9b),
	.w4(32'h3c1e5264),
	.w5(32'hb9761f8e),
	.w6(32'h3c81066b),
	.w7(32'h3c1e44a9),
	.w8(32'h3944a468),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d03fa),
	.w1(32'h3bc02f23),
	.w2(32'h3b53ac48),
	.w3(32'hbae5cc30),
	.w4(32'h3b0aef0b),
	.w5(32'h3a9dfab8),
	.w6(32'hbadf224f),
	.w7(32'h3b31e24f),
	.w8(32'h3a28aacf),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc0f2c),
	.w1(32'h3b6e64a1),
	.w2(32'hbb3228a9),
	.w3(32'hbafd6f4d),
	.w4(32'h3b9b9705),
	.w5(32'h3b9e5785),
	.w6(32'hbb44fcc0),
	.w7(32'h3b6b41d9),
	.w8(32'h3b15ec39),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17b3fd),
	.w1(32'h38dcbf17),
	.w2(32'hbb694a6b),
	.w3(32'hba0ee294),
	.w4(32'hbb409bd2),
	.w5(32'hbb6eabfa),
	.w6(32'hb9c39257),
	.w7(32'h39befc0c),
	.w8(32'hb883acbc),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b79b0),
	.w1(32'hbacfb3a4),
	.w2(32'h3b2d4491),
	.w3(32'hbbf2176b),
	.w4(32'hbbf827dc),
	.w5(32'h3b72f83e),
	.w6(32'hbbd9acf7),
	.w7(32'hbb6c78ff),
	.w8(32'h3b21b443),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0b920),
	.w1(32'h3bf5548a),
	.w2(32'h363f33a4),
	.w3(32'h38d3f840),
	.w4(32'h3a958b99),
	.w5(32'hbacfe862),
	.w6(32'h3b6e7bc3),
	.w7(32'h3bcd1e73),
	.w8(32'h3b40b1cc),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb920f0d),
	.w1(32'h3bcba31b),
	.w2(32'hba9fe40a),
	.w3(32'hbb54d746),
	.w4(32'hbb88a147),
	.w5(32'hbafbbb67),
	.w6(32'h3b11e7d4),
	.w7(32'h3b83fc32),
	.w8(32'hbb9d30d8),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a07e9),
	.w1(32'hbb7ddc0d),
	.w2(32'hbbbc00e8),
	.w3(32'hb893e7aa),
	.w4(32'hb8e8dd21),
	.w5(32'hbb63b62f),
	.w6(32'h3b154436),
	.w7(32'h3b0be543),
	.w8(32'hbbb245f1),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99514b),
	.w1(32'hbb1d08fb),
	.w2(32'hbbe1de9d),
	.w3(32'h3b6f693c),
	.w4(32'h3a92ad49),
	.w5(32'hbc01ceb4),
	.w6(32'h3b07df42),
	.w7(32'hba7c0e99),
	.w8(32'hbbb2392b),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67bbda),
	.w1(32'hba9fa030),
	.w2(32'hbbdeac49),
	.w3(32'hbc59acca),
	.w4(32'h3a8e8e71),
	.w5(32'hbaf38f5e),
	.w6(32'hbbbf31b7),
	.w7(32'hbbd69535),
	.w8(32'hbb96e531),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc071795),
	.w1(32'hbbb02d20),
	.w2(32'hbb95daa6),
	.w3(32'hbc289442),
	.w4(32'hbbdf9f5b),
	.w5(32'hbb70c0d1),
	.w6(32'hbc23dc88),
	.w7(32'hbba5f60b),
	.w8(32'hbae44072),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc27bd1),
	.w1(32'hba8f9960),
	.w2(32'hbc07d360),
	.w3(32'hba647a3d),
	.w4(32'hbaa75732),
	.w5(32'hb8061eef),
	.w6(32'h3b586af1),
	.w7(32'h3b8af788),
	.w8(32'hbb1d6f97),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b21467),
	.w1(32'h3aca3248),
	.w2(32'hbc357559),
	.w3(32'h3b90a092),
	.w4(32'h3acbd83f),
	.w5(32'hbbef1888),
	.w6(32'h3bb15214),
	.w7(32'h3b993952),
	.w8(32'hbb0c9dc8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d6056),
	.w1(32'hb9a40a89),
	.w2(32'h3bd6a7bc),
	.w3(32'hbbcc2336),
	.w4(32'h3b9f5e8c),
	.w5(32'h3b9b916e),
	.w6(32'hbb0ca3dc),
	.w7(32'h3a8ec77f),
	.w8(32'h3b9050e3),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b839b18),
	.w1(32'h3b9d700c),
	.w2(32'h3958d236),
	.w3(32'h3bbdb398),
	.w4(32'h3b750d2a),
	.w5(32'h3a907862),
	.w6(32'h3b8bb0a6),
	.w7(32'h3b919a97),
	.w8(32'h3b00f6fe),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29967e),
	.w1(32'h3bc9da52),
	.w2(32'hbc3aa4fb),
	.w3(32'h3c0998dc),
	.w4(32'h3bd0e4dc),
	.w5(32'hbb92a012),
	.w6(32'h3bd16f7f),
	.w7(32'h3ba9a229),
	.w8(32'hbb4ff963),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe82c64),
	.w1(32'hbbc0ffb6),
	.w2(32'hbc190211),
	.w3(32'hbc11d716),
	.w4(32'hbbef1063),
	.w5(32'hbbd18ed7),
	.w6(32'hbb3c9514),
	.w7(32'hbbd93f2b),
	.w8(32'hbb889bd1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3403ea),
	.w1(32'h3a9f7434),
	.w2(32'hbc01f371),
	.w3(32'hbc84d5fd),
	.w4(32'hbbaf6c68),
	.w5(32'hbc3dcced),
	.w6(32'hbc81a9b0),
	.w7(32'hbbb1aad7),
	.w8(32'hbc129efe),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99bcca),
	.w1(32'h3b5e12f0),
	.w2(32'h3b4d633e),
	.w3(32'hbbd6e1ae),
	.w4(32'hbb388039),
	.w5(32'h3a4b8c3d),
	.w6(32'hbb0ed1b0),
	.w7(32'hbb6b7bdb),
	.w8(32'h3ae8dbd1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10898d),
	.w1(32'h3bca4505),
	.w2(32'hbb358550),
	.w3(32'hbbbe9d19),
	.w4(32'hbb337b6b),
	.w5(32'hbb345460),
	.w6(32'h385ca351),
	.w7(32'h3aa61352),
	.w8(32'hbb667406),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca76992),
	.w1(32'hbc0c429c),
	.w2(32'hbc7b58a9),
	.w3(32'hbc699c97),
	.w4(32'hbc42e4d1),
	.w5(32'hbc51ae04),
	.w6(32'hbc31a88e),
	.w7(32'hbc330fef),
	.w8(32'hbbb4bcbe),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d6dec),
	.w1(32'h3b03a05b),
	.w2(32'hbcb64ec8),
	.w3(32'h3c1a6a62),
	.w4(32'h3bd4449f),
	.w5(32'hbc202798),
	.w6(32'h3c0590c2),
	.w7(32'h3b60c72f),
	.w8(32'hbc0d73d9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cee35),
	.w1(32'hbc267742),
	.w2(32'hbbfad520),
	.w3(32'hbc766214),
	.w4(32'hbc06935d),
	.w5(32'hbb5509c6),
	.w6(32'hbb087b51),
	.w7(32'hbb871bcd),
	.w8(32'hbbe2506f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d2c3e),
	.w1(32'hb9cd07f9),
	.w2(32'hbc06d161),
	.w3(32'h3b3fcdaf),
	.w4(32'h3b1734d2),
	.w5(32'hbc339901),
	.w6(32'hbb257fde),
	.w7(32'hba9f4f1d),
	.w8(32'hbc1667c0),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc153ce8),
	.w1(32'hbc16a79c),
	.w2(32'h3bf59425),
	.w3(32'hbc3b28ec),
	.w4(32'hbc43b116),
	.w5(32'h3c093a66),
	.w6(32'hbc50534e),
	.w7(32'hbc6cb05f),
	.w8(32'hb93cf3eb),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12f77d),
	.w1(32'h3c15b9a7),
	.w2(32'hbb36a51b),
	.w3(32'h3c4e9ce7),
	.w4(32'h3c36e172),
	.w5(32'hbc12a35e),
	.w6(32'h3c0c3465),
	.w7(32'h3c5389ba),
	.w8(32'hbc1438aa),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb389217),
	.w1(32'hba8790e6),
	.w2(32'hbbe53318),
	.w3(32'hbc1c85d0),
	.w4(32'hbbbb81bd),
	.w5(32'hbc228483),
	.w6(32'hbc56602a),
	.w7(32'hbc46df4d),
	.w8(32'hbb233c57),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd23cef),
	.w1(32'hbbaf1899),
	.w2(32'hbc457664),
	.w3(32'hbc1d5ffe),
	.w4(32'hbc26353b),
	.w5(32'hbc1a0933),
	.w6(32'hbc2398e2),
	.w7(32'hbc585636),
	.w8(32'hbba7ab5a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2464d),
	.w1(32'h3b1c80af),
	.w2(32'h3bc28357),
	.w3(32'hbc7653ae),
	.w4(32'hbb2d66df),
	.w5(32'h3baff112),
	.w6(32'hbc2cd6c1),
	.w7(32'hbc30c1c3),
	.w8(32'hbaf1ef8e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78e91c),
	.w1(32'hbb82b089),
	.w2(32'hbb57875a),
	.w3(32'h3bde2d3c),
	.w4(32'h3b44cd89),
	.w5(32'hbbc25198),
	.w6(32'h3a489f81),
	.w7(32'h3bb67c8c),
	.w8(32'hbbe3fa55),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89fc70),
	.w1(32'hba3cb6fa),
	.w2(32'hbb7f6137),
	.w3(32'hbbd8a761),
	.w4(32'hbb74651c),
	.w5(32'hbbcc181f),
	.w6(32'hbbd4f662),
	.w7(32'hbbb8e91a),
	.w8(32'hbbad8d97),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb578602),
	.w1(32'hb96feede),
	.w2(32'h3bdde41e),
	.w3(32'hbbe08116),
	.w4(32'hbb2c016a),
	.w5(32'h3b84cb18),
	.w6(32'hbbd58fba),
	.w7(32'hbb310891),
	.w8(32'hbb6d88b1),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd7752),
	.w1(32'h3c1b1835),
	.w2(32'h3b9f431c),
	.w3(32'h3c681038),
	.w4(32'h3c8814f9),
	.w5(32'h3b210dc8),
	.w6(32'h3c723275),
	.w7(32'h3bc036dc),
	.w8(32'h3adaf22b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8148e),
	.w1(32'h3be949bb),
	.w2(32'hbb5a8b5a),
	.w3(32'h3b9b6806),
	.w4(32'h3bddb8ef),
	.w5(32'hbbac66d5),
	.w6(32'h39ff6850),
	.w7(32'h3b053f99),
	.w8(32'hbb58d772),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02c9da),
	.w1(32'hbb10eb0b),
	.w2(32'hbc436c4b),
	.w3(32'h39bc9ed4),
	.w4(32'hbaad8464),
	.w5(32'h3a01c923),
	.w6(32'hbb4414ef),
	.w7(32'hbb0f7b48),
	.w8(32'hbb0890b2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc272295),
	.w1(32'h3af8dcde),
	.w2(32'hbbfbdfca),
	.w3(32'hbbabc7f2),
	.w4(32'h3b9822ea),
	.w5(32'hbc24e06f),
	.w6(32'hbc3e3e54),
	.w7(32'hbbbb31c9),
	.w8(32'hbb196ebb),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc392c52),
	.w1(32'h3a81fd11),
	.w2(32'h3bcfca79),
	.w3(32'hbc6a0d36),
	.w4(32'hbaaf0611),
	.w5(32'h3c202563),
	.w6(32'hbc7089c0),
	.w7(32'hbb45632a),
	.w8(32'h3bd11fbf),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule