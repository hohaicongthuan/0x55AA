module layer_6_featuremap_29(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d01cc),
	.w1(32'hbb6a4447),
	.w2(32'h3b88e4eb),
	.w3(32'hbc0c4122),
	.w4(32'hbb92faf7),
	.w5(32'hbbd406f4),
	.w6(32'hbb820f7f),
	.w7(32'h3bf1187f),
	.w8(32'h3bc7e448),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01b64a),
	.w1(32'h3a28df6a),
	.w2(32'h3b341c81),
	.w3(32'hb9e7c2b6),
	.w4(32'h3a821ce1),
	.w5(32'h39f1d4b7),
	.w6(32'hbc36778b),
	.w7(32'hbc062e6d),
	.w8(32'h3a59a0e3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b863276),
	.w1(32'h3ba61e21),
	.w2(32'h3a5cc9ac),
	.w3(32'h3c0e3258),
	.w4(32'hb9e863cd),
	.w5(32'h3c14e2df),
	.w6(32'h3bd049d9),
	.w7(32'h3b94160f),
	.w8(32'h3be8f358),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff70c7),
	.w1(32'h3b25636c),
	.w2(32'h3aaf79fc),
	.w3(32'h3b356aa9),
	.w4(32'h3a838b0c),
	.w5(32'h3b6db8bf),
	.w6(32'h3ae722be),
	.w7(32'h3ab89f26),
	.w8(32'h3b1d6068),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e659c),
	.w1(32'hbbe399cb),
	.w2(32'h39cf144c),
	.w3(32'hbb328458),
	.w4(32'hbc21895d),
	.w5(32'hbabff135),
	.w6(32'hbc16c4be),
	.w7(32'hbb427d6b),
	.w8(32'h3c78320f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c302ccf),
	.w1(32'hbc268e6b),
	.w2(32'hbc3d938c),
	.w3(32'hbbb23f68),
	.w4(32'hbc3f198f),
	.w5(32'hbc0f18c7),
	.w6(32'hbc2a085d),
	.w7(32'hbc77a4b7),
	.w8(32'hbbefd449),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb016eb1),
	.w1(32'h3c13576c),
	.w2(32'h3c99e11c),
	.w3(32'hb9819fe3),
	.w4(32'h3ac2516d),
	.w5(32'h3b4ba7ca),
	.w6(32'h3bdd6340),
	.w7(32'h3caf73ab),
	.w8(32'h3c974db4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64b289),
	.w1(32'hbba3b074),
	.w2(32'h3a13aca7),
	.w3(32'hbbca6fbe),
	.w4(32'hbc00d4b8),
	.w5(32'h3b5a5a9f),
	.w6(32'hbc620678),
	.w7(32'hbb1c7e86),
	.w8(32'hbb0f3771),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b4e7a),
	.w1(32'hbc707fd3),
	.w2(32'hbb6b4afe),
	.w3(32'hbbc9ca6a),
	.w4(32'hbc4aca11),
	.w5(32'hbaf20ed8),
	.w6(32'hbc0638ee),
	.w7(32'hbb685e98),
	.w8(32'h3b0c93ff),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2a0fa),
	.w1(32'hbbbf3845),
	.w2(32'hbad64a42),
	.w3(32'hba29b60f),
	.w4(32'hbbd6a214),
	.w5(32'hbbf78c20),
	.w6(32'hbb7ffdd4),
	.w7(32'hba1a2807),
	.w8(32'hbad9e881),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb504d3d),
	.w1(32'hbbc2e056),
	.w2(32'hbbced9b5),
	.w3(32'hbb18ec00),
	.w4(32'hbb8c365c),
	.w5(32'hbb943940),
	.w6(32'hbbe21e8e),
	.w7(32'hbb65a80d),
	.w8(32'hbbd14c4b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3524f626),
	.w1(32'hbaf01bdf),
	.w2(32'hbba27199),
	.w3(32'hb8a059de),
	.w4(32'hbbac565b),
	.w5(32'hbb2f9e39),
	.w6(32'h394b151b),
	.w7(32'hbaa25ce5),
	.w8(32'hbb17fad8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3fd95),
	.w1(32'hbcc4d8df),
	.w2(32'h3d0c7ff2),
	.w3(32'hbcfc4113),
	.w4(32'hbb59ac49),
	.w5(32'hbce08c9d),
	.w6(32'hbc659484),
	.w7(32'h3d725ccb),
	.w8(32'hba641204),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbbbc91),
	.w1(32'hba2e93cc),
	.w2(32'hbb12f8b6),
	.w3(32'h35b8b043),
	.w4(32'hba77e815),
	.w5(32'hbb6889b3),
	.w6(32'h3b8e7dd0),
	.w7(32'hbb4a5625),
	.w8(32'h3b0d9054),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e1906),
	.w1(32'h3bae19aa),
	.w2(32'hbacd448e),
	.w3(32'hba98a276),
	.w4(32'hbbf85d09),
	.w5(32'hb9997a57),
	.w6(32'h3c00f85c),
	.w7(32'h3a6bd56c),
	.w8(32'h3bf7c39b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0367cc),
	.w1(32'hbb362973),
	.w2(32'hbb2f4192),
	.w3(32'hbb829f99),
	.w4(32'hbbb77dd7),
	.w5(32'hbb349429),
	.w6(32'hbbad2856),
	.w7(32'hbba0ed93),
	.w8(32'h3b244241),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba505f29),
	.w1(32'hba816350),
	.w2(32'hbb38913a),
	.w3(32'h3ae84f7d),
	.w4(32'h3b8baeb0),
	.w5(32'hbaa07404),
	.w6(32'h3b1b5992),
	.w7(32'h3ba062bb),
	.w8(32'hba848435),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad66241),
	.w1(32'hbac100ed),
	.w2(32'h3ad07067),
	.w3(32'hbbc8d796),
	.w4(32'hbbf5e7f8),
	.w5(32'h39276a3f),
	.w6(32'hbba2e10b),
	.w7(32'h3a781d2a),
	.w8(32'h3bb454e2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc914b),
	.w1(32'h3b05490a),
	.w2(32'hbc387471),
	.w3(32'h3c672ee7),
	.w4(32'h3ae27a49),
	.w5(32'h3b02fa16),
	.w6(32'h3b952424),
	.w7(32'hbc17c7e1),
	.w8(32'hbbdce23f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e7b4d),
	.w1(32'hbb0f8bfa),
	.w2(32'hbb3b1299),
	.w3(32'hbb13054b),
	.w4(32'hbbb0d502),
	.w5(32'hbb42ed33),
	.w6(32'hbb8d428c),
	.w7(32'hbb57b08a),
	.w8(32'hbb9aa8a0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2351bc),
	.w1(32'h3b0b2cff),
	.w2(32'h3c002aa4),
	.w3(32'h39f6dd12),
	.w4(32'h3bae31b7),
	.w5(32'h3b31ea0d),
	.w6(32'h3b4a8aab),
	.w7(32'h3c01df80),
	.w8(32'h3bb125ce),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fd24a),
	.w1(32'hbb3271c2),
	.w2(32'h3a183f92),
	.w3(32'hbbe01977),
	.w4(32'hbb981a94),
	.w5(32'hbafbc9ab),
	.w6(32'hbb9aa4e9),
	.w7(32'hbb06a58c),
	.w8(32'hb99f7a4e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98971a),
	.w1(32'hba9feb21),
	.w2(32'h3c1d7ba0),
	.w3(32'hbb8ae970),
	.w4(32'hbc9e4aa7),
	.w5(32'hbb93ef05),
	.w6(32'hbb2588b0),
	.w7(32'h3bbcad1a),
	.w8(32'h3befcd16),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9a447),
	.w1(32'hbacb087d),
	.w2(32'hbb587cda),
	.w3(32'hb9cd8d9a),
	.w4(32'hbbc64587),
	.w5(32'hba35e497),
	.w6(32'hbc2dc273),
	.w7(32'hbbe10fec),
	.w8(32'hbbb4d8cd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6ac6a),
	.w1(32'h3c0809b0),
	.w2(32'h3b9c8010),
	.w3(32'h3bdc59a9),
	.w4(32'h3b4936b2),
	.w5(32'hbb08e081),
	.w6(32'h3c87a02b),
	.w7(32'h3c41a3ff),
	.w8(32'h3bf74181),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0195e),
	.w1(32'hbaf636d6),
	.w2(32'h3b9fcdd3),
	.w3(32'hba95a710),
	.w4(32'h3b967ab7),
	.w5(32'hba872bf2),
	.w6(32'hba117802),
	.w7(32'h3b7d0171),
	.w8(32'hbb791847),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac975e2),
	.w1(32'h3b380f65),
	.w2(32'h3b87fc44),
	.w3(32'hb91fd356),
	.w4(32'hbb0338c9),
	.w5(32'h3ac5dce6),
	.w6(32'hbc3f14a6),
	.w7(32'h3c3bb227),
	.w8(32'h3c067fe5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a62627),
	.w1(32'hbaf81bbc),
	.w2(32'hbb11eb51),
	.w3(32'h39fc2bd2),
	.w4(32'hbb8eba95),
	.w5(32'hbb3d6057),
	.w6(32'hbae80b59),
	.w7(32'hbb5a9121),
	.w8(32'hb95c46bf),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb924d3cc),
	.w1(32'h3afe274a),
	.w2(32'hba4de5d8),
	.w3(32'hba0a9ff2),
	.w4(32'h3a51c905),
	.w5(32'h3babf8a3),
	.w6(32'h381d166c),
	.w7(32'hbb2ea88f),
	.w8(32'h3b0cd4ab),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b05ba),
	.w1(32'hba81e6bd),
	.w2(32'hb937cf4b),
	.w3(32'h3a3ce907),
	.w4(32'hbad6de93),
	.w5(32'hbbaae1e7),
	.w6(32'h3acc4b2e),
	.w7(32'h3bd22843),
	.w8(32'hbad8fea5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb441233),
	.w1(32'hbb2a54da),
	.w2(32'hbb5a8c43),
	.w3(32'hbbe50b18),
	.w4(32'hbc19b732),
	.w5(32'hbbaed647),
	.w6(32'h3c015f70),
	.w7(32'h3bfe93d7),
	.w8(32'h3c446036),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c9512),
	.w1(32'hbad3118d),
	.w2(32'h3b9deffe),
	.w3(32'hbb487393),
	.w4(32'hbc3551fb),
	.w5(32'hbbd10b35),
	.w6(32'hbae168c5),
	.w7(32'hba961e8c),
	.w8(32'hb9ec0d9c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1dae2),
	.w1(32'hb9958a1f),
	.w2(32'h3c05c428),
	.w3(32'h3abbbf23),
	.w4(32'h3bad92b8),
	.w5(32'hbc36a7d3),
	.w6(32'hbb13f994),
	.w7(32'h3c2394c4),
	.w8(32'hbb98939f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb854efa),
	.w1(32'hbb5a1634),
	.w2(32'h3b813500),
	.w3(32'hbb147fee),
	.w4(32'hba641aaa),
	.w5(32'hbb314211),
	.w6(32'hbba91862),
	.w7(32'h3b895fc2),
	.w8(32'hbb90a3c9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b43a7),
	.w1(32'hbc82ee1f),
	.w2(32'hbc958cad),
	.w3(32'hbc230755),
	.w4(32'hbc3ccabb),
	.w5(32'hbc63c734),
	.w6(32'hbc452e04),
	.w7(32'hbc74845e),
	.w8(32'hbc881fe0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc881846),
	.w1(32'hb9e001bf),
	.w2(32'h3a84ec53),
	.w3(32'h39acc905),
	.w4(32'hbc029e84),
	.w5(32'hbae1c4cc),
	.w6(32'hba73e1fe),
	.w7(32'hbba071d1),
	.w8(32'h3ba1f1ed),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c183ddb),
	.w1(32'hba668830),
	.w2(32'hbab7db3e),
	.w3(32'hbb56fb87),
	.w4(32'hbba2d12d),
	.w5(32'hba2331d2),
	.w6(32'hbb94b652),
	.w7(32'hbb1a5ac3),
	.w8(32'h3a15ae01),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5292f),
	.w1(32'h3a2b67aa),
	.w2(32'hb83019b4),
	.w3(32'hba398e2b),
	.w4(32'h3a1cbf3b),
	.w5(32'h3af4ea7f),
	.w6(32'h3abeda7b),
	.w7(32'h3a09075d),
	.w8(32'h3b1077a7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48d7c9),
	.w1(32'hbad51fa7),
	.w2(32'h3acf5397),
	.w3(32'hba82ff58),
	.w4(32'hbb552099),
	.w5(32'hbba24d29),
	.w6(32'h3bdceaa2),
	.w7(32'h3b950256),
	.w8(32'h3af1ac05),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f7425),
	.w1(32'hbc1634a0),
	.w2(32'hbb819591),
	.w3(32'hbc36f94f),
	.w4(32'hbc6172d3),
	.w5(32'hbc4d0e5e),
	.w6(32'hbc557ee2),
	.w7(32'hbb3f56c1),
	.w8(32'h3b108b4e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68ebb3),
	.w1(32'h3ba4a9ed),
	.w2(32'hbba6c6df),
	.w3(32'h3c02a66e),
	.w4(32'hbc467c95),
	.w5(32'hbb8c99e3),
	.w6(32'hb9b3b290),
	.w7(32'hbc347a37),
	.w8(32'hb86070c6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb253bab),
	.w1(32'hba03e040),
	.w2(32'hb9a7c2d1),
	.w3(32'hbb1277a4),
	.w4(32'hbb38773f),
	.w5(32'h3a659c33),
	.w6(32'hbaea5511),
	.w7(32'hbae0e4bd),
	.w8(32'h3aa35287),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb9ea8),
	.w1(32'h3bb67a52),
	.w2(32'h3be3f162),
	.w3(32'hbbdcf88d),
	.w4(32'hbbcdc348),
	.w5(32'hba6849b4),
	.w6(32'h3ac843c9),
	.w7(32'h3b1ed6c0),
	.w8(32'h3c072be2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c821967),
	.w1(32'h3b94fd69),
	.w2(32'h3a886e82),
	.w3(32'hbb186ed8),
	.w4(32'hbb7c00b0),
	.w5(32'h3a86d1a8),
	.w6(32'hbad97e25),
	.w7(32'h395ba00e),
	.w8(32'h3b5f0155),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e5b48),
	.w1(32'h399b387d),
	.w2(32'h3a10dcc6),
	.w3(32'h3aaf835b),
	.w4(32'h3ab521bb),
	.w5(32'h3b31e91c),
	.w6(32'hba09b30b),
	.w7(32'hbac992e0),
	.w8(32'h3a1b49c8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b709f6e),
	.w1(32'hbad03f6d),
	.w2(32'h39dc6e21),
	.w3(32'h3b3bcbf3),
	.w4(32'hba1e0fdb),
	.w5(32'hbbb8dad7),
	.w6(32'h3b576e54),
	.w7(32'h3c227df4),
	.w8(32'hbb555e7d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd0b13),
	.w1(32'h3abbcb13),
	.w2(32'h3c267d6b),
	.w3(32'h3a6fe807),
	.w4(32'hbadb77b6),
	.w5(32'h39a972cf),
	.w6(32'hbaccaac1),
	.w7(32'h3becc6b4),
	.w8(32'h3b9ddebf),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c283c78),
	.w1(32'hba621891),
	.w2(32'hbb8789e0),
	.w3(32'h3ba24d20),
	.w4(32'hbc0c169b),
	.w5(32'hbadf7e0f),
	.w6(32'h3a80f712),
	.w7(32'hbbcc8a0c),
	.w8(32'h3a1775ec),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf700c3),
	.w1(32'hb9ac783f),
	.w2(32'hbbd94200),
	.w3(32'h3b9460cd),
	.w4(32'hba2c042a),
	.w5(32'h3b8d4485),
	.w6(32'h3a6e5f33),
	.w7(32'hbbf53fe7),
	.w8(32'hbaeb3fd3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc206c8),
	.w1(32'hbbfcbc30),
	.w2(32'h390896d7),
	.w3(32'hbb99f342),
	.w4(32'hbc133670),
	.w5(32'hbaf975a8),
	.w6(32'hbbed9118),
	.w7(32'hba114672),
	.w8(32'h3b04fddb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86acb2),
	.w1(32'h3ac3e079),
	.w2(32'h3bd544da),
	.w3(32'hbb6422c7),
	.w4(32'hbb0a69d9),
	.w5(32'h3b149971),
	.w6(32'hba6869bf),
	.w7(32'h3c0eaee8),
	.w8(32'h3b8dd1f0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1fc49),
	.w1(32'hbbbf645d),
	.w2(32'h3b28475f),
	.w3(32'hbc2547e5),
	.w4(32'hbb1663e5),
	.w5(32'hbb4b65cf),
	.w6(32'hbc130370),
	.w7(32'h3962d232),
	.w8(32'h394c7767),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7a2b2),
	.w1(32'hbca7f9c8),
	.w2(32'hbce1f2dc),
	.w3(32'hbc50177e),
	.w4(32'hbc9dcf35),
	.w5(32'hbc7aa8d7),
	.w6(32'hbc9e09fb),
	.w7(32'hbce258ce),
	.w8(32'hbca40631),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ced93),
	.w1(32'hbc96a6d6),
	.w2(32'hbc95f717),
	.w3(32'hbc485eeb),
	.w4(32'hbc9a4498),
	.w5(32'hbc884741),
	.w6(32'hbc8dcf7a),
	.w7(32'hbc9d7820),
	.w8(32'hbc629052),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d7069),
	.w1(32'h3acff8e8),
	.w2(32'h3b393a19),
	.w3(32'hbb25cf4a),
	.w4(32'hbb61e95b),
	.w5(32'h3ab6a820),
	.w6(32'hbac27004),
	.w7(32'h3bb18f0d),
	.w8(32'h3b67815a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6c256),
	.w1(32'hbbb215d3),
	.w2(32'h3ac2ab11),
	.w3(32'h3ae9e3d0),
	.w4(32'h3af1de83),
	.w5(32'hba0a6bb7),
	.w6(32'hbb382ea4),
	.w7(32'h3a95f232),
	.w8(32'hba477941),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68aa70),
	.w1(32'hbc5d452d),
	.w2(32'hbca504a8),
	.w3(32'hbc6e7b94),
	.w4(32'hbc97d1b8),
	.w5(32'hbc148f8b),
	.w6(32'hbca53b30),
	.w7(32'hbcd4dd39),
	.w8(32'hbc6f0359),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11c80d),
	.w1(32'hba318074),
	.w2(32'h3bd57b38),
	.w3(32'h3b272f7e),
	.w4(32'hb93ff4e8),
	.w5(32'h3ba17f88),
	.w6(32'h3b208936),
	.w7(32'h3c12d05a),
	.w8(32'h3ba376d5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12f0df),
	.w1(32'h388f4933),
	.w2(32'h3b8eb76e),
	.w3(32'hbb036973),
	.w4(32'h3a196dc4),
	.w5(32'hbab2047b),
	.w6(32'h3acadca1),
	.w7(32'h3b9fb121),
	.w8(32'h3ab379b8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad089cf),
	.w1(32'h3c01dbe7),
	.w2(32'h3c93fcdd),
	.w3(32'hbb22e405),
	.w4(32'h3bc86add),
	.w5(32'h3c516e40),
	.w6(32'h3c156ca2),
	.w7(32'h3c6f8c89),
	.w8(32'h3c5a9abd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22ee18),
	.w1(32'h3b9780aa),
	.w2(32'h3c251d86),
	.w3(32'h3b9a8296),
	.w4(32'h3b76c5ca),
	.w5(32'hbaab4e1b),
	.w6(32'h3c2a58f8),
	.w7(32'h3c4718e0),
	.w8(32'h3bc80e57),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b818439),
	.w1(32'hbb280ed4),
	.w2(32'hbb33f93b),
	.w3(32'h3b8f2418),
	.w4(32'h3bc2abc3),
	.w5(32'h3b0f59f2),
	.w6(32'h3b2f95dc),
	.w7(32'h3bd27c14),
	.w8(32'h397d3818),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab41b14),
	.w1(32'h3a974dd3),
	.w2(32'hbb618b89),
	.w3(32'h3c82f3b1),
	.w4(32'h3c6a819b),
	.w5(32'h3c7abefe),
	.w6(32'h3c9f8bb7),
	.w7(32'h3c9f8d13),
	.w8(32'h3c5662af),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d346c),
	.w1(32'h3d10f341),
	.w2(32'h3d28dc5b),
	.w3(32'h3d0ff38e),
	.w4(32'h3d1ea962),
	.w5(32'h3c01b2d2),
	.w6(32'h3d522ac7),
	.w7(32'h3d7534c2),
	.w8(32'h3cd28a89),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule