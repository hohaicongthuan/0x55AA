module layer_8_featuremap_232(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf2a22),
	.w1(32'hbb24d939),
	.w2(32'hbc0d3906),
	.w3(32'h3c03740e),
	.w4(32'h3b500c95),
	.w5(32'h39ae9178),
	.w6(32'h3b2dd9a5),
	.w7(32'hbaa011e3),
	.w8(32'h3b814b93),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9688a4),
	.w1(32'hbd9f8f69),
	.w2(32'h3c21a1da),
	.w3(32'hbadc109d),
	.w4(32'hbd6e7ccb),
	.w5(32'hbc14da65),
	.w6(32'hbd35687f),
	.w7(32'hbaf8fa07),
	.w8(32'h3cf034a3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dbb03ca),
	.w1(32'hbaddd6d0),
	.w2(32'h3b8248d2),
	.w3(32'h3d1fc3b0),
	.w4(32'hbb78760f),
	.w5(32'h3ba66f61),
	.w6(32'hbba5c62b),
	.w7(32'h3a9c73a1),
	.w8(32'h3b9a89e1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27eaab),
	.w1(32'h3b98f4b3),
	.w2(32'h3bd9079f),
	.w3(32'h3bf89fef),
	.w4(32'hbb59cdd4),
	.w5(32'h3bd60d4f),
	.w6(32'hba8bdc81),
	.w7(32'h3a0d57fe),
	.w8(32'h3ace168e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cf5ba),
	.w1(32'hbdec1063),
	.w2(32'h3c73e7df),
	.w3(32'h3b94d705),
	.w4(32'hbdb31d1f),
	.w5(32'hbbabaa60),
	.w6(32'hbd9703b4),
	.w7(32'hbc30ecd4),
	.w8(32'h3d3a3a39),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e06a912),
	.w1(32'h3a868228),
	.w2(32'hbc0d0214),
	.w3(32'h3d8652c3),
	.w4(32'hbb33b183),
	.w5(32'hbca46efc),
	.w6(32'h3b3a8156),
	.w7(32'hbc25a72c),
	.w8(32'hbbd3d550),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6eb21c),
	.w1(32'h3d0625fd),
	.w2(32'hbbf802ff),
	.w3(32'hbbcdd378),
	.w4(32'h3cdf1934),
	.w5(32'hb9b39634),
	.w6(32'h3c8e6e29),
	.w7(32'hbb53af6c),
	.w8(32'hbc7b81dc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd555192),
	.w1(32'h3a9add89),
	.w2(32'h3c36ff51),
	.w3(32'hbce8a668),
	.w4(32'h3b07f7fb),
	.w5(32'h3af13fb7),
	.w6(32'hbb20980f),
	.w7(32'hb8a18f58),
	.w8(32'hbbde14ed),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b448d55),
	.w1(32'hbdc0e2f5),
	.w2(32'h3cc54a7c),
	.w3(32'h3aa1f4e6),
	.w4(32'hbd8f74e1),
	.w5(32'h3ba9a1db),
	.w6(32'hbd5e2727),
	.w7(32'h3b036259),
	.w8(32'h3d4ed3cf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e00186f),
	.w1(32'hbb583dd0),
	.w2(32'hba87c162),
	.w3(32'h3d8497df),
	.w4(32'hbb052eda),
	.w5(32'h3bd834ba),
	.w6(32'hbb40fa60),
	.w7(32'hbb65b358),
	.w8(32'hbb212915),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24702e),
	.w1(32'h3c55d3d4),
	.w2(32'h3c6ad8c6),
	.w3(32'h3bd9afb1),
	.w4(32'h3c564b92),
	.w5(32'h3c8e9eda),
	.w6(32'h3b8827b2),
	.w7(32'hbb458797),
	.w8(32'hbbc9d2ea),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba886c82),
	.w1(32'hbb796db6),
	.w2(32'hbc09285e),
	.w3(32'h3b3523b0),
	.w4(32'h3a3eb2b9),
	.w5(32'hbbbcba44),
	.w6(32'hbb591df5),
	.w7(32'hbbdd0094),
	.w8(32'hbc180367),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97195e),
	.w1(32'h3a0b4d0c),
	.w2(32'hb9cb3189),
	.w3(32'hbc9490a8),
	.w4(32'h3bb32f1c),
	.w5(32'hbb6c007f),
	.w6(32'hbb3519ff),
	.w7(32'hbb0a2e9c),
	.w8(32'hbc1c670e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb50a2),
	.w1(32'hbc104cf9),
	.w2(32'hbb564478),
	.w3(32'hbb5831b5),
	.w4(32'hbabe8e49),
	.w5(32'h3b0a05c5),
	.w6(32'hbb2fd587),
	.w7(32'hbb5a959d),
	.w8(32'h39d740e9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1247d),
	.w1(32'h3d8ade16),
	.w2(32'hbcb508f6),
	.w3(32'h3b2710ef),
	.w4(32'h3d40105d),
	.w5(32'hbb8cfacb),
	.w6(32'h3d211ce9),
	.w7(32'hbb839c88),
	.w8(32'hbd2cfdac),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbddb0fe0),
	.w1(32'hbada54e9),
	.w2(32'hbaf7d3d3),
	.w3(32'hbd4f2479),
	.w4(32'hbb9096de),
	.w5(32'h3b99a66a),
	.w6(32'h3ad59281),
	.w7(32'h3a89b25a),
	.w8(32'h3ba08a63),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b37b6),
	.w1(32'h3b4f3f18),
	.w2(32'h39e4b86a),
	.w3(32'h3afa8616),
	.w4(32'h3c1d8a24),
	.w5(32'hba94ae1b),
	.w6(32'h3bb0be87),
	.w7(32'hbb9f7246),
	.w8(32'hbaa45616),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57f678),
	.w1(32'hbc1476f7),
	.w2(32'hbba093b1),
	.w3(32'hbb3d3723),
	.w4(32'hbbb602ef),
	.w5(32'hbbdb9c57),
	.w6(32'hbc4659d5),
	.w7(32'h3ad6b878),
	.w8(32'h3b5a265b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ac74f),
	.w1(32'hbaa2bfd4),
	.w2(32'hbb21dd96),
	.w3(32'h3b5a83c1),
	.w4(32'h3b4d63b8),
	.w5(32'hbb95455f),
	.w6(32'hbbb9884f),
	.w7(32'hbb92a7c7),
	.w8(32'hbc073f78),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc708c89),
	.w1(32'h3db3ca56),
	.w2(32'hbbef8a9a),
	.w3(32'hbbbca783),
	.w4(32'h3d82643b),
	.w5(32'h3bdc1e7d),
	.w6(32'h3d570e47),
	.w7(32'h3badd055),
	.w8(32'hbd20c726),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbddb71ed),
	.w1(32'h3c080adb),
	.w2(32'h3ab443e7),
	.w3(32'hbd60e641),
	.w4(32'h3bf164b7),
	.w5(32'h3b91bf64),
	.w6(32'h3ba7b789),
	.w7(32'hbb7cd164),
	.w8(32'h3b57a770),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d966a),
	.w1(32'hbc50f4f6),
	.w2(32'h3a40959f),
	.w3(32'hb9ccac13),
	.w4(32'hbb573a11),
	.w5(32'hbac6b76c),
	.w6(32'hbafa2c6f),
	.w7(32'hbc20bd64),
	.w8(32'h3a8c55b7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ee2ee),
	.w1(32'h3c5e0782),
	.w2(32'h3c8496d8),
	.w3(32'h397aa596),
	.w4(32'h3bc778e4),
	.w5(32'h3c34b08f),
	.w6(32'h3c022c08),
	.w7(32'h3c92ac24),
	.w8(32'h3c51b922),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be373fc),
	.w1(32'hbc2fe5b4),
	.w2(32'hbb9960f5),
	.w3(32'h3b9972df),
	.w4(32'hbbe1bc38),
	.w5(32'hbbac2d29),
	.w6(32'hbbce6780),
	.w7(32'hba0b84e0),
	.w8(32'h3aaa1c40),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a286b70),
	.w1(32'h3bb0455a),
	.w2(32'h3bf3d824),
	.w3(32'hbaeebfa0),
	.w4(32'h3bb2be96),
	.w5(32'h3a6cf9e4),
	.w6(32'hba5f74f5),
	.w7(32'h3ba4b1e2),
	.w8(32'hbb2e41df),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ffda9),
	.w1(32'hbb35cf97),
	.w2(32'hbc0836f5),
	.w3(32'hbbc2119d),
	.w4(32'hb8cbd257),
	.w5(32'h3b906066),
	.w6(32'h39e836bf),
	.w7(32'hbaeae675),
	.w8(32'hbadc3425),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1c314),
	.w1(32'hbbb8ec47),
	.w2(32'hbbca37b7),
	.w3(32'hbab2c38f),
	.w4(32'hbbc02425),
	.w5(32'hbc0697f7),
	.w6(32'hbba32760),
	.w7(32'hbb9a11f6),
	.w8(32'h3846e48e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50d185),
	.w1(32'hbc467dfb),
	.w2(32'hbb86347c),
	.w3(32'hba72329b),
	.w4(32'hbbf1d7f9),
	.w5(32'hbbab697d),
	.w6(32'hbc56e878),
	.w7(32'hbbc12f50),
	.w8(32'h3b60d52a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35a442),
	.w1(32'h3c000b48),
	.w2(32'hbadb2bac),
	.w3(32'hbbdc5bd9),
	.w4(32'h3c2bac14),
	.w5(32'hbb197c0f),
	.w6(32'h3bc594d5),
	.w7(32'h3b87057d),
	.w8(32'h3ba4e954),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace2a90),
	.w1(32'hbc067943),
	.w2(32'h3b255d7f),
	.w3(32'hbbc64ccd),
	.w4(32'hbc674455),
	.w5(32'hbbcc77e4),
	.w6(32'hbbe57c88),
	.w7(32'hbb9114c7),
	.w8(32'h3bfc15f6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c106492),
	.w1(32'h3b0dba3f),
	.w2(32'hbb47abb3),
	.w3(32'hbba3ce74),
	.w4(32'h3ba2fbf3),
	.w5(32'h3b39a278),
	.w6(32'hbad99358),
	.w7(32'h3a49ceb7),
	.w8(32'hbb7d97b6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4d156),
	.w1(32'h3b418f85),
	.w2(32'hba4e07ef),
	.w3(32'hbbc00dc0),
	.w4(32'hb9bce184),
	.w5(32'h3acc3d35),
	.w6(32'hbb71fd36),
	.w7(32'hbb63c6a8),
	.w8(32'h3be85aaa),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3faee8),
	.w1(32'h3c191ad4),
	.w2(32'h3c89dd1e),
	.w3(32'h3a0350f0),
	.w4(32'h3bfc0c72),
	.w5(32'h3c223b65),
	.w6(32'h3b40864c),
	.w7(32'h3c10f637),
	.w8(32'hbb8ebf54),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70c5ba),
	.w1(32'hba0f4ffd),
	.w2(32'h3bc09334),
	.w3(32'hbb00bc9c),
	.w4(32'h3a339dc4),
	.w5(32'h3abc17ce),
	.w6(32'h3c01f7d3),
	.w7(32'h3bb4a2d7),
	.w8(32'h3b1d97c0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69fcef),
	.w1(32'hbb498cf8),
	.w2(32'h3b9ed696),
	.w3(32'hbb1a340f),
	.w4(32'h3b7873ad),
	.w5(32'hb93de239),
	.w6(32'h3b5aeac0),
	.w7(32'h3bdcd4c9),
	.w8(32'h3b802983),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97a2c4),
	.w1(32'hbb63d623),
	.w2(32'hbb9d84ed),
	.w3(32'h3bd7a94b),
	.w4(32'hbacba041),
	.w5(32'h3b6b6954),
	.w6(32'hb9e0f038),
	.w7(32'hbb93012b),
	.w8(32'hbb9089a9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada5622),
	.w1(32'hbc26b82c),
	.w2(32'hbc6a2dd0),
	.w3(32'h3b8ca34c),
	.w4(32'hbbb5b4bc),
	.w5(32'hbc69463c),
	.w6(32'hbbfa5192),
	.w7(32'hbc01c0e9),
	.w8(32'h3b3fa8a1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8931a3),
	.w1(32'hbc28de8d),
	.w2(32'h3a9b1443),
	.w3(32'hbc117423),
	.w4(32'hbc44a20d),
	.w5(32'hbba31d91),
	.w6(32'hbae38ea4),
	.w7(32'h3b8dc66c),
	.w8(32'h3bd11b04),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c458311),
	.w1(32'hbbc9c0be),
	.w2(32'hbb354c16),
	.w3(32'h3bc3b3ed),
	.w4(32'hbb7a8c05),
	.w5(32'hbb3d6f60),
	.w6(32'hbb7c40fc),
	.w7(32'h3b336f36),
	.w8(32'h3b7295bd),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c044427),
	.w1(32'h3a98a307),
	.w2(32'hba3ff8e2),
	.w3(32'hb907b670),
	.w4(32'h3ac40eda),
	.w5(32'hb9e1067b),
	.w6(32'h3b33ba98),
	.w7(32'h3a8f1019),
	.w8(32'h3bd06c4a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5973d4),
	.w1(32'h3c4ba4ae),
	.w2(32'h3b01f4bc),
	.w3(32'h3b813cd7),
	.w4(32'h3ca32ebd),
	.w5(32'h3bf4190a),
	.w6(32'h3c69e26c),
	.w7(32'h3b44b782),
	.w8(32'h3b34699f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9169e),
	.w1(32'h3b47e3bd),
	.w2(32'hbbd36d27),
	.w3(32'h3bd340e6),
	.w4(32'h3ad7db82),
	.w5(32'hba22f94f),
	.w6(32'hba800174),
	.w7(32'hbbaf8db3),
	.w8(32'hbbc2e117),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdecb75),
	.w1(32'h3a08917f),
	.w2(32'hbc09d16e),
	.w3(32'hbae6eb68),
	.w4(32'h3b10c81c),
	.w5(32'hbbc68e2b),
	.w6(32'hbb18db6e),
	.w7(32'h3a91dddd),
	.w8(32'h3c461058),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b185986),
	.w1(32'hbc1e6231),
	.w2(32'hbbc747fd),
	.w3(32'h3afe8f08),
	.w4(32'hba89393d),
	.w5(32'hbbf22ac0),
	.w6(32'hbbe7ce8c),
	.w7(32'hbbf0aff4),
	.w8(32'hba7af983),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99cba4),
	.w1(32'h3b5b8f9a),
	.w2(32'h3bcb7290),
	.w3(32'hbb8de3e2),
	.w4(32'hbaa426d8),
	.w5(32'h3bafa27c),
	.w6(32'h3c01d81a),
	.w7(32'h39f72e17),
	.w8(32'hbb6c7bbe),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9634a8),
	.w1(32'h3d65e865),
	.w2(32'hbc210893),
	.w3(32'hb9c94848),
	.w4(32'h3d3bf97a),
	.w5(32'h3b873702),
	.w6(32'h3d02c9f9),
	.w7(32'hb9ea40b6),
	.w8(32'hbd2f37ae),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdb899ca),
	.w1(32'hbc0b38e3),
	.w2(32'hbb9eef37),
	.w3(32'hbd558373),
	.w4(32'hbbd7f029),
	.w5(32'hbbf9fcf6),
	.w6(32'hbc1814af),
	.w7(32'hbba91da2),
	.w8(32'hbbae7d63),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d27604),
	.w1(32'hbaca9e58),
	.w2(32'h3a434300),
	.w3(32'hbb71e7b9),
	.w4(32'hbbc327a5),
	.w5(32'h3a80b188),
	.w6(32'hba061c98),
	.w7(32'h3a9e9260),
	.w8(32'h3ba624dc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b260af4),
	.w1(32'hbbb8a5da),
	.w2(32'hbaba16e0),
	.w3(32'h3aca706a),
	.w4(32'hbb958279),
	.w5(32'hba32e625),
	.w6(32'hbb09b086),
	.w7(32'h3bd33751),
	.w8(32'h3b434119),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa17132),
	.w1(32'hbc08a64b),
	.w2(32'hbc463198),
	.w3(32'h3c171ada),
	.w4(32'hbbe304a4),
	.w5(32'hbc26bcd5),
	.w6(32'hbbbbe3c8),
	.w7(32'hbc694c08),
	.w8(32'hbb0035f6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc05a4),
	.w1(32'h3a2f734f),
	.w2(32'hbbd3e027),
	.w3(32'hbb9a9c5a),
	.w4(32'hbaaac05a),
	.w5(32'hbb6fdabd),
	.w6(32'h3abd448a),
	.w7(32'h3a2ec202),
	.w8(32'h3a7cf151),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfebbb1),
	.w1(32'h3c17a726),
	.w2(32'h3c4bdf96),
	.w3(32'h3b1c947a),
	.w4(32'h3c2922b5),
	.w5(32'h3c3c12e1),
	.w6(32'h3bbb8b6b),
	.w7(32'h3b9fb639),
	.w8(32'h3aa3a3e5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5090e),
	.w1(32'hbd2ef287),
	.w2(32'h3c29e9d6),
	.w3(32'h3bd955ef),
	.w4(32'hbcf1cd0d),
	.w5(32'hbb14b0c2),
	.w6(32'hbcb846c3),
	.w7(32'h3ae8d4fe),
	.w8(32'h3c92a164),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6b1685),
	.w1(32'h3bee81fd),
	.w2(32'h3c09bd24),
	.w3(32'h3cc62727),
	.w4(32'h3c023ad5),
	.w5(32'h3c498b4a),
	.w6(32'h3bdd2ab1),
	.w7(32'h3c01fbdd),
	.w8(32'h3ad8e0ab),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf82c20),
	.w1(32'h3b0b5cc0),
	.w2(32'h3c8a3bea),
	.w3(32'h3afa2393),
	.w4(32'h3b3b1b6c),
	.w5(32'h3cb67d14),
	.w6(32'h3bd160e5),
	.w7(32'h3c49b619),
	.w8(32'h3b980975),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c0f93),
	.w1(32'hbc089de5),
	.w2(32'hbc14918e),
	.w3(32'h3bf8754c),
	.w4(32'hbb8bd4ec),
	.w5(32'hbbc1c4f1),
	.w6(32'hbb3d0154),
	.w7(32'hbbb5e6e3),
	.w8(32'h3be6b430),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387bf82a),
	.w1(32'hbb7d41e7),
	.w2(32'hbb8c2df8),
	.w3(32'hb99e028b),
	.w4(32'hbb97fa35),
	.w5(32'h3b37d8dd),
	.w6(32'h3b87c919),
	.w7(32'h3ba17175),
	.w8(32'hbadf067f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb975636),
	.w1(32'hbc12a22a),
	.w2(32'hbcbf9840),
	.w3(32'h3b341e45),
	.w4(32'hbbbbcfcc),
	.w5(32'hbc937f6e),
	.w6(32'hbbaf55a4),
	.w7(32'hbc5b8ae1),
	.w8(32'h3b39db3f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e86c0),
	.w1(32'h3c41c964),
	.w2(32'h3b80cb45),
	.w3(32'hbb7799c6),
	.w4(32'h3c46bdce),
	.w5(32'h3b62a569),
	.w6(32'h3c1200cf),
	.w7(32'h3c0c6359),
	.w8(32'h3aa5eef0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bf5e6),
	.w1(32'hbb7ae9eb),
	.w2(32'h3b1148ad),
	.w3(32'hbc274646),
	.w4(32'hbb4666fb),
	.w5(32'h3aac40c8),
	.w6(32'hbc0b905d),
	.w7(32'hba24fe85),
	.w8(32'h3b05d385),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0daea1),
	.w1(32'hbc019279),
	.w2(32'hbb919457),
	.w3(32'hbaf59dff),
	.w4(32'hbc284f22),
	.w5(32'h3a0b052b),
	.w6(32'hbbb6f929),
	.w7(32'hbb9fc328),
	.w8(32'hbc2c20ac),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5d992),
	.w1(32'h38d60469),
	.w2(32'h3bca6441),
	.w3(32'hbb88f76a),
	.w4(32'h3c84f77b),
	.w5(32'h3b5b8b2c),
	.w6(32'hbc2955af),
	.w7(32'h3bbea208),
	.w8(32'h3c458163),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea9b2f),
	.w1(32'h3c1ac45d),
	.w2(32'hbb355ed2),
	.w3(32'hbc1effb4),
	.w4(32'h3bcd6cbd),
	.w5(32'hbac929bf),
	.w6(32'h3b976b9f),
	.w7(32'h3b416ab6),
	.w8(32'h3c58b82f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda60a2),
	.w1(32'hbb97c1b8),
	.w2(32'hbbd260db),
	.w3(32'hbb60b2a6),
	.w4(32'h3946e91a),
	.w5(32'hbb4fa21f),
	.w6(32'h3b6a5495),
	.w7(32'hba97a873),
	.w8(32'hbbf0de6e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4df6ae),
	.w1(32'h3d276b6d),
	.w2(32'hbac07a75),
	.w3(32'hbc2f016c),
	.w4(32'h3cfc6833),
	.w5(32'h3b03bfb2),
	.w6(32'h3ce42c01),
	.w7(32'h3bd493e9),
	.w8(32'hbc60ecdb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd13f4e8),
	.w1(32'h3b70b01f),
	.w2(32'hbb047c84),
	.w3(32'hbc97ad69),
	.w4(32'h3abf2aeb),
	.w5(32'hb9b6e39f),
	.w6(32'h3bb44279),
	.w7(32'h3ba0f13c),
	.w8(32'h3b32f054),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0fe0f),
	.w1(32'hbc1fa2ac),
	.w2(32'hbb2be3c9),
	.w3(32'h3be56720),
	.w4(32'hbabe7fe0),
	.w5(32'hbb833f97),
	.w6(32'hbb728e5b),
	.w7(32'hbbc90736),
	.w8(32'hbb9899e4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0c9d5),
	.w1(32'hbaf8bb19),
	.w2(32'hbc419131),
	.w3(32'h3a5e6cee),
	.w4(32'hbb3d185f),
	.w5(32'hbc256085),
	.w6(32'hbba9d662),
	.w7(32'hbc479685),
	.w8(32'hbc14b518),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53e710),
	.w1(32'hbc472c32),
	.w2(32'hbb0f893a),
	.w3(32'hbbdc35de),
	.w4(32'hbbf19e10),
	.w5(32'hbbefd157),
	.w6(32'hbc28b5c0),
	.w7(32'hb8e38e63),
	.w8(32'hbb26595a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf1737),
	.w1(32'hbb8f6c37),
	.w2(32'h3b4635b5),
	.w3(32'hbad0e1ff),
	.w4(32'hbaa3c320),
	.w5(32'h3b26fbba),
	.w6(32'hbb35b02a),
	.w7(32'h3bab5344),
	.w8(32'h3bdf6f88),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6104ef),
	.w1(32'h3ce0aa9e),
	.w2(32'h3d2fdd55),
	.w3(32'h3a3dfde3),
	.w4(32'h3c5790a9),
	.w5(32'h3d05e47a),
	.w6(32'h3cbe1519),
	.w7(32'h3d04aae0),
	.w8(32'h3c06b27d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26c1ee),
	.w1(32'hbb5b5072),
	.w2(32'h3bb690a1),
	.w3(32'h3c5e9ef1),
	.w4(32'hbb2af49a),
	.w5(32'h3b5e9a7c),
	.w6(32'hb9b079e9),
	.w7(32'h3c136945),
	.w8(32'h3c07ee3f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3ebfa),
	.w1(32'hbb45eda9),
	.w2(32'h3b8b1c25),
	.w3(32'h3bd8f6af),
	.w4(32'hbaea5d83),
	.w5(32'h3ab80c29),
	.w6(32'h3b673167),
	.w7(32'h3b69792f),
	.w8(32'h3bc29034),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55d009),
	.w1(32'hbb8ff5b1),
	.w2(32'h3b837f67),
	.w3(32'h3bfbed20),
	.w4(32'hbbc5ded0),
	.w5(32'h3b8d94dd),
	.w6(32'hbb119a78),
	.w7(32'h3a803560),
	.w8(32'h3bdae648),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d7975),
	.w1(32'h3c78bbcb),
	.w2(32'h3cb5f0f1),
	.w3(32'h3af2fda3),
	.w4(32'h3c8e38d1),
	.w5(32'h3c8bf025),
	.w6(32'h3b97496c),
	.w7(32'h3c755911),
	.w8(32'h3c0da1e4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ea172),
	.w1(32'hbc2a0e6b),
	.w2(32'h3ac769c4),
	.w3(32'h3bf5f4ef),
	.w4(32'hbc5ec13e),
	.w5(32'hbb56a47b),
	.w6(32'hbc5de63a),
	.w7(32'hbba7fe46),
	.w8(32'hba34cc8c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9444ce),
	.w1(32'h3b37f2b2),
	.w2(32'hbb2f4102),
	.w3(32'h3a454dfe),
	.w4(32'h3b40ab31),
	.w5(32'h3a99ab60),
	.w6(32'h3a2a56f2),
	.w7(32'hbb5f5fec),
	.w8(32'h3bf30ba8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a03e0),
	.w1(32'hbc4b016b),
	.w2(32'hbcabc028),
	.w3(32'h3c5d07e2),
	.w4(32'hbc4bae11),
	.w5(32'hbc7be705),
	.w6(32'hbc54c5bb),
	.w7(32'hbc7347a6),
	.w8(32'h3ac543e0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39477253),
	.w1(32'h3c415bb8),
	.w2(32'h3c28cfd1),
	.w3(32'h3b896a55),
	.w4(32'h3b6d26a8),
	.w5(32'h3c3789a8),
	.w6(32'h3b82361d),
	.w7(32'h3bd3d3fd),
	.w8(32'h3a70b465),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b437288),
	.w1(32'hb9f82a4a),
	.w2(32'h3c15ca63),
	.w3(32'h3bc42a1a),
	.w4(32'hbbbf8a75),
	.w5(32'h38e4b24b),
	.w6(32'hbb1499f6),
	.w7(32'h3ba2ad42),
	.w8(32'h3afac0f6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7330b3),
	.w1(32'hbbad8da7),
	.w2(32'hbb45b9b3),
	.w3(32'h3c18a7d3),
	.w4(32'hba813ca4),
	.w5(32'h3b751786),
	.w6(32'h3b2f68a6),
	.w7(32'h3ba7ec88),
	.w8(32'hbb0cb8c4),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25b689),
	.w1(32'hbb999042),
	.w2(32'hbb53a5d2),
	.w3(32'h3ba575f2),
	.w4(32'hbbee0ed8),
	.w5(32'hbba90861),
	.w6(32'hbb83c5e5),
	.w7(32'h3a897224),
	.w8(32'h3b2a59c7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01f9b5),
	.w1(32'hb907b5eb),
	.w2(32'h3ba0e170),
	.w3(32'h3a17114f),
	.w4(32'h3b5db9ad),
	.w5(32'h3b7d48c5),
	.w6(32'h3b9eef32),
	.w7(32'h3aaa6356),
	.w8(32'hbb49b127),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedef0a),
	.w1(32'h3c0968f9),
	.w2(32'h3c9f844c),
	.w3(32'hbaf0c4f5),
	.w4(32'h3c354ac4),
	.w5(32'h3bafd7c2),
	.w6(32'h3ba418d4),
	.w7(32'h3b73fdaf),
	.w8(32'h3bd870da),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94c3a9),
	.w1(32'h3b00b99e),
	.w2(32'h3b5831db),
	.w3(32'h3a4293f8),
	.w4(32'hbac2a263),
	.w5(32'h3b975374),
	.w6(32'hbb3e0cbe),
	.w7(32'hbb3fd8a5),
	.w8(32'h3b42fccb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c7f67),
	.w1(32'hbc2218a6),
	.w2(32'hbb8bb1b3),
	.w3(32'h3c26f149),
	.w4(32'hbc1178d8),
	.w5(32'hbbf0b478),
	.w6(32'hbbaf85f8),
	.w7(32'hbbb7db52),
	.w8(32'hbb998641),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17994a),
	.w1(32'h3b90f670),
	.w2(32'h3aa944f0),
	.w3(32'h3a056998),
	.w4(32'hbae9ab85),
	.w5(32'h3b2c4e52),
	.w6(32'h3bc39b9e),
	.w7(32'hbb3bbe2e),
	.w8(32'hbc070970),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8797df),
	.w1(32'h3b8191f9),
	.w2(32'hb8a777c8),
	.w3(32'h3ab1e645),
	.w4(32'h3b9ed645),
	.w5(32'hbabb6c36),
	.w6(32'h3bbb3ac0),
	.w7(32'h3b61c256),
	.w8(32'hbb1796ff),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeb014),
	.w1(32'hbbe334c4),
	.w2(32'hbb708e5b),
	.w3(32'hbbe4a8ff),
	.w4(32'hbb86385c),
	.w5(32'hb9e81b6d),
	.w6(32'hbbe82134),
	.w7(32'hbbda0c60),
	.w8(32'hbbf1cda5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae780f8),
	.w1(32'hbb88f8c3),
	.w2(32'h3b70ab3a),
	.w3(32'hbb15a616),
	.w4(32'h3a2e6c74),
	.w5(32'h3bf58460),
	.w6(32'h3a7b7d1f),
	.w7(32'h3c2edd6f),
	.w8(32'h3c0ff53b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ecda2),
	.w1(32'hbb52a666),
	.w2(32'h3b588f74),
	.w3(32'h3bde73b3),
	.w4(32'h3a162d0c),
	.w5(32'hba3c5a9c),
	.w6(32'hbb20eef0),
	.w7(32'hbb314b2f),
	.w8(32'hbabf6798),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba9cba),
	.w1(32'h3bb87584),
	.w2(32'h3b87a3bf),
	.w3(32'h3bbe763c),
	.w4(32'h38497dea),
	.w5(32'h3b31ad17),
	.w6(32'h3bc390eb),
	.w7(32'h3b7c6a59),
	.w8(32'h3b695d40),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a348c),
	.w1(32'hbca193fe),
	.w2(32'h3a0d3592),
	.w3(32'h3bf2f34c),
	.w4(32'hbc472daa),
	.w5(32'hba6182f1),
	.w6(32'hbbefed75),
	.w7(32'hbb1806ab),
	.w8(32'h3ba6820e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82ef25),
	.w1(32'hbd043298),
	.w2(32'h3a07154e),
	.w3(32'h3be4c576),
	.w4(32'hbc9d8e20),
	.w5(32'hbbd506ef),
	.w6(32'hbc74e00d),
	.w7(32'hbb69cc25),
	.w8(32'h3c09311e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d02f760),
	.w1(32'hbb9ce20f),
	.w2(32'hbb7f99dc),
	.w3(32'h3c07904f),
	.w4(32'hbc1ca236),
	.w5(32'hbba1cf44),
	.w6(32'h3a867588),
	.w7(32'h3b09fb05),
	.w8(32'hbaa10ef0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d59ab),
	.w1(32'hbc7444df),
	.w2(32'hbc70aa81),
	.w3(32'hbb48da7c),
	.w4(32'hbbee7ecd),
	.w5(32'hbbfb102a),
	.w6(32'hbc13cceb),
	.w7(32'hbc112444),
	.w8(32'h3b9176b2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a580a50),
	.w1(32'hbb1f105e),
	.w2(32'h3c557c97),
	.w3(32'h3b9748b3),
	.w4(32'hbaa6ee8c),
	.w5(32'h3c6a2ec6),
	.w6(32'h3ab38c06),
	.w7(32'h3c299a77),
	.w8(32'h3c167d4d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dab22),
	.w1(32'hbb857554),
	.w2(32'h3c2e56e9),
	.w3(32'h3b5dae3f),
	.w4(32'hbbdbd1f9),
	.w5(32'h3b6a15f6),
	.w6(32'hbb6e09ac),
	.w7(32'hb9aa0b4d),
	.w8(32'h3af6f3c3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb2864),
	.w1(32'hbc11d9d7),
	.w2(32'hbc1c9700),
	.w3(32'h3c0691ec),
	.w4(32'hbc345397),
	.w5(32'hbbdd0985),
	.w6(32'hbc5fe4e2),
	.w7(32'hbbf42131),
	.w8(32'hb9abdddb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdd519),
	.w1(32'h3adda76c),
	.w2(32'h3bc8557b),
	.w3(32'h39c3cfc9),
	.w4(32'hba796ccd),
	.w5(32'h3bb74134),
	.w6(32'h3bbd569c),
	.w7(32'h3a616898),
	.w8(32'h3a1c54f0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f9e92),
	.w1(32'h3b99db4c),
	.w2(32'h3b19cb1c),
	.w3(32'hbb7d2d70),
	.w4(32'h3ba84c85),
	.w5(32'h3a9a4bf4),
	.w6(32'hbbad4494),
	.w7(32'h3aaee29c),
	.w8(32'hbbb3e748),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba893fd8),
	.w1(32'h3c72a1d1),
	.w2(32'h3acd6fd4),
	.w3(32'hbbbcc5d6),
	.w4(32'h3c2f9f4d),
	.w5(32'h3ab599b3),
	.w6(32'h3c3932cd),
	.w7(32'hbb769425),
	.w8(32'hbba69ad3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18ade2),
	.w1(32'hbb6aac44),
	.w2(32'hbb440b69),
	.w3(32'hbbad242f),
	.w4(32'hbb2875b4),
	.w5(32'hb9eaa99d),
	.w6(32'h3a9815f6),
	.w7(32'h3a93a27d),
	.w8(32'h39bd01e9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50ab48),
	.w1(32'hbbc3d833),
	.w2(32'hbb8888d9),
	.w3(32'hbbb5eba7),
	.w4(32'hbbb2ec39),
	.w5(32'hbaf9d95c),
	.w6(32'h3b1a178e),
	.w7(32'h3b893630),
	.w8(32'hba0a8517),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94799a),
	.w1(32'h3adf0ad1),
	.w2(32'h3c22bc2a),
	.w3(32'h3bb5ed4e),
	.w4(32'hbac5eeb2),
	.w5(32'h3be011cc),
	.w6(32'h3b40c7a0),
	.w7(32'h3b6ad606),
	.w8(32'hbae2a63e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9017b9),
	.w1(32'h3d835358),
	.w2(32'hbbfe3dea),
	.w3(32'h3b4876e5),
	.w4(32'h3d453410),
	.w5(32'h3c0b6cb1),
	.w6(32'h3d191e84),
	.w7(32'h3bf34a2d),
	.w8(32'hbd02c6fb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdb1825d),
	.w1(32'hbc35b435),
	.w2(32'hbb8114c1),
	.w3(32'hbd21b3fa),
	.w4(32'hbc3f2ff7),
	.w5(32'hbbb7538c),
	.w6(32'hbc337533),
	.w7(32'hbc6bccf8),
	.w8(32'hbc59cc27),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc14599),
	.w1(32'hbbd88ed5),
	.w2(32'hbc46e1d1),
	.w3(32'hbb7abf4b),
	.w4(32'hbb326de6),
	.w5(32'hbc46cd2b),
	.w6(32'hbbf27949),
	.w7(32'h3b2761d7),
	.w8(32'h3bf774f2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc8b96),
	.w1(32'hbbffcad3),
	.w2(32'hbc202f76),
	.w3(32'hbbc25e5d),
	.w4(32'hbb956ae9),
	.w5(32'hbbc552e2),
	.w6(32'hbb0091f1),
	.w7(32'hbbeaaf4e),
	.w8(32'hbb339780),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf882b4),
	.w1(32'hbd2622b9),
	.w2(32'h3c294181),
	.w3(32'hbb52f854),
	.w4(32'hbcf994e7),
	.w5(32'hbb4fc19b),
	.w6(32'hbcc41ec3),
	.w7(32'h3b86e45d),
	.w8(32'h3cc33903),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d688708),
	.w1(32'hb98742c9),
	.w2(32'h3b08399b),
	.w3(32'h3cc03d38),
	.w4(32'hbab6429f),
	.w5(32'hb9b7a5d8),
	.w6(32'h3b91086c),
	.w7(32'hbb2266e5),
	.w8(32'h39fb8ec1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d8910),
	.w1(32'h3d0e69aa),
	.w2(32'h3b447983),
	.w3(32'h3b130c80),
	.w4(32'h3ce18421),
	.w5(32'h3c053de1),
	.w6(32'h3cb28bbf),
	.w7(32'h3af0930c),
	.w8(32'hbc5c5544),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7abbe),
	.w1(32'hbc439a1f),
	.w2(32'hbbe7b139),
	.w3(32'hbc50e820),
	.w4(32'hbc3a1343),
	.w5(32'hbbcfd030),
	.w6(32'hbc8ac257),
	.w7(32'hbbb76eba),
	.w8(32'hbc19fa98),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8ecf3),
	.w1(32'h3b0a2270),
	.w2(32'hbb19f880),
	.w3(32'hbbe3b2ed),
	.w4(32'h3b801e81),
	.w5(32'h3b89e4f2),
	.w6(32'hbba963fa),
	.w7(32'h3aaf17d8),
	.w8(32'h3bed528b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cf3d3),
	.w1(32'h3bc6c88c),
	.w2(32'h3c28805c),
	.w3(32'h3abb1d82),
	.w4(32'h3c0f69e5),
	.w5(32'h3c729d25),
	.w6(32'h3bad4faa),
	.w7(32'h3b9c4673),
	.w8(32'h3b0667f9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8ed68),
	.w1(32'hbcafffe6),
	.w2(32'h3aea826d),
	.w3(32'h3bff2b0e),
	.w4(32'hbc931384),
	.w5(32'hbbdf67d1),
	.w6(32'hbc512ad5),
	.w7(32'h3b168c60),
	.w8(32'h3c2c6f57),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdd9d2f),
	.w1(32'h3b39d91a),
	.w2(32'h3c02cd1f),
	.w3(32'h3c0d2344),
	.w4(32'hbc3b12b7),
	.w5(32'hba7d7d1b),
	.w6(32'hba458770),
	.w7(32'hbb375a63),
	.w8(32'h395e7b62),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c090e8f),
	.w1(32'hbc002111),
	.w2(32'hba8fde2d),
	.w3(32'hbacf7e23),
	.w4(32'hbbee202b),
	.w5(32'hbb93d7a3),
	.w6(32'hbc1092eb),
	.w7(32'hbb44d367),
	.w8(32'hba4974dd),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98908c),
	.w1(32'hbc0fc81e),
	.w2(32'hbc21b122),
	.w3(32'hbb3fac38),
	.w4(32'h3a1a1730),
	.w5(32'h3a7f6968),
	.w6(32'hbbf8467f),
	.w7(32'hbbbc4da6),
	.w8(32'h3b6a7b52),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbef58),
	.w1(32'h3bed2bb0),
	.w2(32'h3c4d6c6f),
	.w3(32'h3a80fc61),
	.w4(32'h3be39629),
	.w5(32'h3c0984bc),
	.w6(32'h3a02a409),
	.w7(32'h3b4e6cdd),
	.w8(32'h3b7c2eb7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f6112),
	.w1(32'hbc123aa8),
	.w2(32'h3995cf9f),
	.w3(32'h3bd255b5),
	.w4(32'hbbc52ca3),
	.w5(32'hbb7a2d44),
	.w6(32'hbbbcf2a6),
	.w7(32'hbb10715d),
	.w8(32'h386c7abf),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12c0c8),
	.w1(32'h3c281220),
	.w2(32'h3c858112),
	.w3(32'h3ae1a399),
	.w4(32'h3c280235),
	.w5(32'h3c382bae),
	.w6(32'h3c5426c2),
	.w7(32'h3c3c4253),
	.w8(32'h3bf91756),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa0069),
	.w1(32'hbd4096ee),
	.w2(32'h3a0a5ca2),
	.w3(32'h3c69c8dd),
	.w4(32'hbcf04ee5),
	.w5(32'hbc3bc43a),
	.w6(32'hbcc1fe02),
	.w7(32'hbc24481a),
	.w8(32'h3b657724),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d298a10),
	.w1(32'hbbbb41aa),
	.w2(32'hbb502ad7),
	.w3(32'h3c1ac05e),
	.w4(32'hbc117459),
	.w5(32'hbbbf5667),
	.w6(32'hbbf584d8),
	.w7(32'hbbdedeac),
	.w8(32'hbc0e3ce5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18fa98),
	.w1(32'hbbacb889),
	.w2(32'h3a4ad6e2),
	.w3(32'hbbff5d78),
	.w4(32'hbb991cd2),
	.w5(32'hbb0c642f),
	.w6(32'hbc037dda),
	.w7(32'hbb89ea4c),
	.w8(32'hba141b0a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f98e9c),
	.w1(32'hbbdad07a),
	.w2(32'h3a8e34e1),
	.w3(32'h3bb8e7e1),
	.w4(32'hbb6003b5),
	.w5(32'h3bafcb8f),
	.w6(32'h39b04292),
	.w7(32'hbb4eb6c1),
	.w8(32'h3a6d62cc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397f40da),
	.w1(32'hba8a4020),
	.w2(32'h3b62d0f8),
	.w3(32'hb7251e84),
	.w4(32'h3b07b10b),
	.w5(32'h3b6997fc),
	.w6(32'h3b1571be),
	.w7(32'h3b85bd3f),
	.w8(32'h3b14a73a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b9906),
	.w1(32'hba102efa),
	.w2(32'hbae10eb4),
	.w3(32'h3a1b939f),
	.w4(32'h3a365b4b),
	.w5(32'h3bd7c1e5),
	.w6(32'hbb436564),
	.w7(32'hbbee8dcd),
	.w8(32'hbafe060f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule