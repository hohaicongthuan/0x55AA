module layer_10_featuremap_170(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8052fa),
	.w1(32'hb99b75b0),
	.w2(32'hba01e3ec),
	.w3(32'hbabe98a9),
	.w4(32'h3aba8080),
	.w5(32'h3a903fa7),
	.w6(32'hb89e61e7),
	.w7(32'hb67c4d02),
	.w8(32'hb9837472),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31c137),
	.w1(32'hb9086b2c),
	.w2(32'h3a2c00e9),
	.w3(32'h39f92fc0),
	.w4(32'hb9847818),
	.w5(32'h3a037448),
	.w6(32'hba205690),
	.w7(32'hb82418cf),
	.w8(32'h3954495f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35a641),
	.w1(32'hbad6ef4c),
	.w2(32'hbad02beb),
	.w3(32'h3a11eab5),
	.w4(32'hbb034a02),
	.w5(32'hbae5ee0f),
	.w6(32'hbad657ae),
	.w7(32'hba82591a),
	.w8(32'hba4f1788),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0fdc1),
	.w1(32'h3a971563),
	.w2(32'h3acb5fef),
	.w3(32'hbad285d8),
	.w4(32'hba9781fd),
	.w5(32'hbacccd32),
	.w6(32'h3a983722),
	.w7(32'h3aafb34e),
	.w8(32'h389b27c4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b72726),
	.w1(32'h39e074d3),
	.w2(32'hb7ab89f1),
	.w3(32'hbac61e3d),
	.w4(32'h3a0fc359),
	.w5(32'h3a525474),
	.w6(32'h3a0870bc),
	.w7(32'hb7c252ef),
	.w8(32'h3ae4320d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf4ec6),
	.w1(32'hba64c944),
	.w2(32'hba6d2c71),
	.w3(32'h39cf3301),
	.w4(32'hbab9cb8f),
	.w5(32'hbad7b462),
	.w6(32'hba2d6e24),
	.w7(32'hba9d6285),
	.w8(32'hbaae5db4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba0bef),
	.w1(32'h39c6148e),
	.w2(32'h3a83e1ff),
	.w3(32'hbade2b27),
	.w4(32'h39a6d97c),
	.w5(32'h3a787ee6),
	.w6(32'hb9ba4e71),
	.w7(32'hb8626332),
	.w8(32'h3a540bac),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf6564),
	.w1(32'h39de31a7),
	.w2(32'hb890f2e4),
	.w3(32'h3aad7b5a),
	.w4(32'hb981fdad),
	.w5(32'hba901882),
	.w6(32'h3a3c2d40),
	.w7(32'h38dc9283),
	.w8(32'hb9ba6bd7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6201d2),
	.w1(32'hb72764a5),
	.w2(32'hba2261e9),
	.w3(32'hbac3f828),
	.w4(32'hb91d2485),
	.w5(32'hba930e71),
	.w6(32'h38cba2a4),
	.w7(32'hb9cb094d),
	.w8(32'hba301b72),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c5236),
	.w1(32'hba717231),
	.w2(32'h39542d9f),
	.w3(32'hba72559c),
	.w4(32'hba1d3f63),
	.w5(32'h399fca26),
	.w6(32'hbb1283f8),
	.w7(32'hbaad90a1),
	.w8(32'hba03b62a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59f7a4),
	.w1(32'hba881cc7),
	.w2(32'hbafc154a),
	.w3(32'h3a6cb86f),
	.w4(32'hbab50877),
	.w5(32'hbb0944d7),
	.w6(32'h39af0d2f),
	.w7(32'h3a801401),
	.w8(32'h3a554415),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09c82f),
	.w1(32'hbaeb9c8c),
	.w2(32'hbada3519),
	.w3(32'hbb0a1e98),
	.w4(32'hba9c0c28),
	.w5(32'hbaeb50a6),
	.w6(32'hb9cf2cb8),
	.w7(32'h391223d1),
	.w8(32'hb8df219c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb068c33),
	.w1(32'hb97046ad),
	.w2(32'hba41c1cd),
	.w3(32'hbaa5e239),
	.w4(32'hb8c5e1f5),
	.w5(32'hba4a471f),
	.w6(32'h39a60b33),
	.w7(32'hb9e94ab8),
	.w8(32'hba0476b3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba486042),
	.w1(32'h3a8ef098),
	.w2(32'h3a1921a6),
	.w3(32'hba46a565),
	.w4(32'hb831622e),
	.w5(32'hba9051cc),
	.w6(32'h3ac62ffa),
	.w7(32'h3a51f6c2),
	.w8(32'hba813d02),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa82f1),
	.w1(32'hbb22e1ab),
	.w2(32'hbb067da3),
	.w3(32'hbb2949da),
	.w4(32'hba4a363e),
	.w5(32'hbade0fff),
	.w6(32'hb9a45ec0),
	.w7(32'h3a272300),
	.w8(32'h3ac1fb5a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02475e),
	.w1(32'h39c646d0),
	.w2(32'hb90c04d0),
	.w3(32'hbab7360a),
	.w4(32'hb824dcc7),
	.w5(32'hba1ceeca),
	.w6(32'h3a000c0e),
	.w7(32'h383d94e7),
	.w8(32'hb9e879d6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47fe6c),
	.w1(32'hba9130cb),
	.w2(32'hba3271a5),
	.w3(32'hba3462ae),
	.w4(32'h38b5c1da),
	.w5(32'h3a2258bc),
	.w6(32'hbaf10c8c),
	.w7(32'hbad1ca8a),
	.w8(32'h3a610f88),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cd1e3),
	.w1(32'hba1ed984),
	.w2(32'h38e8f181),
	.w3(32'h3b03feb3),
	.w4(32'hb9dc48f1),
	.w5(32'h399d59ae),
	.w6(32'hbacfb6e0),
	.w7(32'hba83a7f8),
	.w8(32'h3910dc4c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50f8a7),
	.w1(32'hba6a2ee1),
	.w2(32'hba495da3),
	.w3(32'h3a28c651),
	.w4(32'hba662fdb),
	.w5(32'hba3bd907),
	.w6(32'hba9621ba),
	.w7(32'hba609d72),
	.w8(32'hb8b3683d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97133ba),
	.w1(32'hba286a1d),
	.w2(32'hbab88db1),
	.w3(32'hb995e9c8),
	.w4(32'hba0cd98d),
	.w5(32'hbac4eabf),
	.w6(32'hba087dce),
	.w7(32'hba8f82df),
	.w8(32'hba8a1e03),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fdb21),
	.w1(32'h3b01e111),
	.w2(32'h3ad3b3c6),
	.w3(32'hba87d8cf),
	.w4(32'h3a793a13),
	.w5(32'h39d3f049),
	.w6(32'h3b528cb6),
	.w7(32'h3b06fdbd),
	.w8(32'h3a916f99),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5aed7),
	.w1(32'hba8a1182),
	.w2(32'hbabd12af),
	.w3(32'h397aa0dd),
	.w4(32'hb9e0caaa),
	.w5(32'hba650bb5),
	.w6(32'hbac34ce4),
	.w7(32'hba6e18c1),
	.w8(32'hbab7dae8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade86c2),
	.w1(32'h3bba06d0),
	.w2(32'h3bb625c5),
	.w3(32'hbb0819ec),
	.w4(32'h3aae1acc),
	.w5(32'h3b0e225b),
	.w6(32'h3b818851),
	.w7(32'h3b94c9c7),
	.w8(32'h3b9c0a83),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2a00c),
	.w1(32'h39c42d64),
	.w2(32'hb9299a9b),
	.w3(32'h3b476d2b),
	.w4(32'hb8e6486d),
	.w5(32'hba74e7b4),
	.w6(32'h3a6c08d1),
	.w7(32'h39cf99b2),
	.w8(32'hb9afbe66),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c9f55),
	.w1(32'hb95cf4fe),
	.w2(32'hb9690968),
	.w3(32'hbaa24a5d),
	.w4(32'hb99e5a6b),
	.w5(32'hba2d69c5),
	.w6(32'h39c6d489),
	.w7(32'h3a0536a9),
	.w8(32'h3a4a2b88),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3fdae),
	.w1(32'h393a9435),
	.w2(32'h39dd8752),
	.w3(32'hb9d220f7),
	.w4(32'h3add76d8),
	.w5(32'h3aaff2d9),
	.w6(32'hbb0e16bf),
	.w7(32'hbaf0c6bb),
	.w8(32'h38dafbea),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a950caf),
	.w1(32'hb9dc4b78),
	.w2(32'hba85aaa2),
	.w3(32'h3b1655cc),
	.w4(32'hb9d5b403),
	.w5(32'hbaa08cc3),
	.w6(32'hb91d222e),
	.w7(32'hba2ea0c6),
	.w8(32'hba05a2cd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49ca0b),
	.w1(32'hbaf41d83),
	.w2(32'hbafab2fa),
	.w3(32'hba16d422),
	.w4(32'hbaddedef),
	.w5(32'hbb0feae9),
	.w6(32'hbaa94b7c),
	.w7(32'hba999592),
	.w8(32'hba86535b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9e808),
	.w1(32'h3baf9089),
	.w2(32'h3b3f14e3),
	.w3(32'hbad916cf),
	.w4(32'h3b61e160),
	.w5(32'h3a9bde3b),
	.w6(32'h3bb57896),
	.w7(32'h3b622d26),
	.w8(32'h3b95a612),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7faeb9),
	.w1(32'h3b06a8aa),
	.w2(32'h3b08ea66),
	.w3(32'h3b506e19),
	.w4(32'h3b4a4150),
	.w5(32'h3b86266f),
	.w6(32'h3a52ef9e),
	.w7(32'h398407c5),
	.w8(32'hb78c1742),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b132f63),
	.w1(32'h3a3b3c70),
	.w2(32'h39df2ceb),
	.w3(32'h3b4b30d1),
	.w4(32'h39a22f39),
	.w5(32'h363f57b1),
	.w6(32'h3aaf7c51),
	.w7(32'h3a53cfc8),
	.w8(32'h39ce973d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e65012),
	.w1(32'h3a1d70b5),
	.w2(32'h380b0cde),
	.w3(32'h369b4db8),
	.w4(32'h394bd576),
	.w5(32'hb9e9327d),
	.w6(32'h3a9bdab4),
	.w7(32'h3977b6fd),
	.w8(32'h395e6ee3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d75e3),
	.w1(32'hbaea62cc),
	.w2(32'hbb141515),
	.w3(32'hb9927542),
	.w4(32'hbac91261),
	.w5(32'hbade480a),
	.w6(32'hbab93372),
	.w7(32'hbb013147),
	.w8(32'hba9dc7d8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4697a),
	.w1(32'h39f98796),
	.w2(32'hbb0c8c7f),
	.w3(32'hba81fc20),
	.w4(32'hb84914db),
	.w5(32'hbb1487a1),
	.w6(32'h3ac498c3),
	.w7(32'hbab5edf6),
	.w8(32'h39eae254),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39652c8b),
	.w1(32'hbadfb835),
	.w2(32'hbab0cf56),
	.w3(32'h3a02b55a),
	.w4(32'hbac1b62d),
	.w5(32'hba96d256),
	.w6(32'hbb0abba4),
	.w7(32'hbae90a52),
	.w8(32'hba2063fe),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99bdb87),
	.w1(32'hb91f0084),
	.w2(32'hb8b31343),
	.w3(32'h392c5a45),
	.w4(32'hb9ff6ec5),
	.w5(32'hba5bed7c),
	.w6(32'h398324fc),
	.w7(32'h38e17022),
	.w8(32'h398a78de),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff446e),
	.w1(32'hbaa52ea5),
	.w2(32'hb9e73cc9),
	.w3(32'hba591496),
	.w4(32'hba705c5f),
	.w5(32'hb912e6ba),
	.w6(32'hbaaaf7a8),
	.w7(32'hba84f33d),
	.w8(32'h392dd601),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39955e11),
	.w1(32'hb9b4e0d3),
	.w2(32'h398f7db4),
	.w3(32'h39c0bcdd),
	.w4(32'hb84675f7),
	.w5(32'h3a534bba),
	.w6(32'hba4b710c),
	.w7(32'hb9c07bd3),
	.w8(32'h380ce4b0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32ca21),
	.w1(32'h39d7b0d9),
	.w2(32'hb988d50d),
	.w3(32'h3a7a07ac),
	.w4(32'hb82c4666),
	.w5(32'hba65a719),
	.w6(32'h3a716e9e),
	.w7(32'h393c3c18),
	.w8(32'hb9d0c804),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba350680),
	.w1(32'hb97cc135),
	.w2(32'h393193f0),
	.w3(32'hba84b203),
	.w4(32'hb9e5ff64),
	.w5(32'hb9b9e9a5),
	.w6(32'hb9d7d9bc),
	.w7(32'hb9834691),
	.w8(32'h394e7ccc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c86298),
	.w1(32'h3b4af1cd),
	.w2(32'h3b8ed5c8),
	.w3(32'hb8e59bb5),
	.w4(32'h3b3d5c90),
	.w5(32'h3ba85707),
	.w6(32'h3aee7407),
	.w7(32'h3ae384a9),
	.w8(32'h381eebea),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b713748),
	.w1(32'hba939869),
	.w2(32'hbaa4ff42),
	.w3(32'h3b794c69),
	.w4(32'hbada95b4),
	.w5(32'hbadfecaf),
	.w6(32'hba7ab770),
	.w7(32'hb9ee5fa9),
	.w8(32'hb9de4dd4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba999bb5),
	.w1(32'h3a1aa352),
	.w2(32'hb8fd1975),
	.w3(32'hbaba0f45),
	.w4(32'h39438fd2),
	.w5(32'hba2f2a23),
	.w6(32'h3a4ee0e2),
	.w7(32'hb906b7f5),
	.w8(32'h38fac000),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cfb3ad),
	.w1(32'hba1d91f5),
	.w2(32'h3ab2a3e5),
	.w3(32'hb99481dd),
	.w4(32'hba0f7190),
	.w5(32'h3a99ef5c),
	.w6(32'hbb48aaf3),
	.w7(32'hbacf1423),
	.w8(32'hbaa19ce3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa702d),
	.w1(32'hb9f13853),
	.w2(32'hb9bd2bdf),
	.w3(32'h39fc4c4a),
	.w4(32'hb8aba25e),
	.w5(32'hb7601553),
	.w6(32'hba5c37e0),
	.w7(32'hba4e22c4),
	.w8(32'hba37cc9a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8d1b4),
	.w1(32'hbacfdf68),
	.w2(32'hbabccb41),
	.w3(32'hba407df9),
	.w4(32'hba9b1ef4),
	.w5(32'hba4cad3c),
	.w6(32'hbaed87a5),
	.w7(32'hbad2a11a),
	.w8(32'hba4deec9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba246c69),
	.w1(32'hb9a27c93),
	.w2(32'h397c1dac),
	.w3(32'hb9f78641),
	.w4(32'h3a824985),
	.w5(32'h39de55b8),
	.w6(32'h3ae37d2b),
	.w7(32'h3b1ce37b),
	.w8(32'h3b306401),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea35c8),
	.w1(32'h3b198c71),
	.w2(32'h3a95489b),
	.w3(32'h3a4acdfc),
	.w4(32'h3a9bda08),
	.w5(32'h38575077),
	.w6(32'h3b83c6a6),
	.w7(32'h3b51dd4f),
	.w8(32'h3baa361f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b710990),
	.w1(32'hba14a74c),
	.w2(32'hba9c2cfe),
	.w3(32'h3b68a1c6),
	.w4(32'hba2d30d8),
	.w5(32'hbabdbafb),
	.w6(32'hb956ff6e),
	.w7(32'hba7294d6),
	.w8(32'hb9e2b255),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba787122),
	.w1(32'h3a515587),
	.w2(32'h39fb70ce),
	.w3(32'hba3ebd01),
	.w4(32'h394b26da),
	.w5(32'hb9de69ee),
	.w6(32'h3a9c4fcb),
	.w7(32'h3a400708),
	.w8(32'hb94f1ace),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02f0af),
	.w1(32'hba23fd7f),
	.w2(32'hb999177f),
	.w3(32'hba9d8ee9),
	.w4(32'hba503256),
	.w5(32'hba2fef86),
	.w6(32'hbacf5729),
	.w7(32'hba99d3f8),
	.w8(32'hba3f8cda),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1344a),
	.w1(32'hb9ed811c),
	.w2(32'hbadeeea2),
	.w3(32'hba4f66b9),
	.w4(32'hba429d75),
	.w5(32'hbab1a628),
	.w6(32'h3a6c05cf),
	.w7(32'hb987a4df),
	.w8(32'hba8025c1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00522e),
	.w1(32'h3981f18c),
	.w2(32'h3a1b1817),
	.w3(32'hba0f84ca),
	.w4(32'hb901dcfd),
	.w5(32'h399b3db4),
	.w6(32'hb9d0ffc9),
	.w7(32'hba13ed57),
	.w8(32'hba6ab6de),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c7e0b),
	.w1(32'hb9a86530),
	.w2(32'h3729314b),
	.w3(32'hb8c3016f),
	.w4(32'hb91d7625),
	.w5(32'h3a34b636),
	.w6(32'hb8f90f37),
	.w7(32'hba0b08c3),
	.w8(32'h3a26b840),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97768b),
	.w1(32'hba2da7ad),
	.w2(32'h39963dd6),
	.w3(32'h39cc8f68),
	.w4(32'h390d195b),
	.w5(32'h3aa46c9f),
	.w6(32'hbabcf319),
	.w7(32'hba17f47d),
	.w8(32'h393c466b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53d0d9),
	.w1(32'h3b1caca4),
	.w2(32'h3b1b686c),
	.w3(32'h3ab85f51),
	.w4(32'h3b2ca7d5),
	.w5(32'h3b4989ac),
	.w6(32'h3a88bbe6),
	.w7(32'h3a8d739d),
	.w8(32'hba378acb),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00a7b3),
	.w1(32'hba1a9290),
	.w2(32'hb92c5651),
	.w3(32'h3b0b2e59),
	.w4(32'hb9f6ca18),
	.w5(32'h398e6770),
	.w6(32'hb9a94a39),
	.w7(32'hb9e92bf9),
	.w8(32'hb9b72cf7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c9281),
	.w1(32'hbaf37678),
	.w2(32'hbb1c5c01),
	.w3(32'h3a0bfb5c),
	.w4(32'hbaeaa324),
	.w5(32'hbaca8cb8),
	.w6(32'hbaf004b6),
	.w7(32'hbb0ef077),
	.w8(32'h392cf888),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3295a0),
	.w1(32'h39a3e127),
	.w2(32'h3a0f4ec9),
	.w3(32'hba66a2f8),
	.w4(32'hb7e65203),
	.w5(32'hb75bfca1),
	.w6(32'hb99d7b2a),
	.w7(32'hb908ef61),
	.w8(32'h3908468f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a68092),
	.w1(32'h39a3479e),
	.w2(32'hb970a2d8),
	.w3(32'hb88088a9),
	.w4(32'hb96e24e9),
	.w5(32'hba8357ee),
	.w6(32'h3a579f9c),
	.w7(32'h39878989),
	.w8(32'hb9ab947d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58ba91),
	.w1(32'hbabf251d),
	.w2(32'hba9ccf4d),
	.w3(32'hba999a25),
	.w4(32'hbadf7c78),
	.w5(32'hbacdad6e),
	.w6(32'hbaf8b695),
	.w7(32'hbad84209),
	.w8(32'hbaa285e2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba911a5b),
	.w1(32'h399a4c5c),
	.w2(32'h38f16af7),
	.w3(32'hbaacaf82),
	.w4(32'h39cf6bb5),
	.w5(32'h38550e27),
	.w6(32'h3a3da5c9),
	.w7(32'h3a29e5bd),
	.w8(32'h3645c81b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ff12e),
	.w1(32'hbaff84c0),
	.w2(32'hbb46324e),
	.w3(32'hba64b1e4),
	.w4(32'hbaaa68b6),
	.w5(32'hbb06c56e),
	.w6(32'hbae03c98),
	.w7(32'hbb300ff5),
	.w8(32'hbb273bf5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11ab25),
	.w1(32'hba3bcf30),
	.w2(32'h3a1c9e83),
	.w3(32'hbac6d273),
	.w4(32'hba39587a),
	.w5(32'h39fcdc69),
	.w6(32'hbb108278),
	.w7(32'hbaa97550),
	.w8(32'hba62bd38),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31be88),
	.w1(32'hba3aeb8b),
	.w2(32'hb9cfd14d),
	.w3(32'h39462a3c),
	.w4(32'hba389e30),
	.w5(32'hba37c25d),
	.w6(32'hba3e7b6b),
	.w7(32'hba389cf1),
	.w8(32'h386edf3b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a86360),
	.w1(32'hbaa27a6e),
	.w2(32'hbaeac40d),
	.w3(32'hb8d471a5),
	.w4(32'hbad73144),
	.w5(32'hbac4a156),
	.w6(32'hba79e8eb),
	.w7(32'hbabd4f84),
	.w8(32'hba0ce56c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9093b1),
	.w1(32'hb9a9ed66),
	.w2(32'h3a5d16e5),
	.w3(32'hbab6da87),
	.w4(32'h3a1e51cd),
	.w5(32'h3b3ec757),
	.w6(32'hbac5bec8),
	.w7(32'hba2f0872),
	.w8(32'hb8a272a5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b217a27),
	.w1(32'h3bec5e8a),
	.w2(32'h3c02531d),
	.w3(32'h3b7fec71),
	.w4(32'h3b69f955),
	.w5(32'h3bb2175d),
	.w6(32'h3bd76090),
	.w7(32'h3bd0921e),
	.w8(32'h3ba5d9a9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdff661),
	.w1(32'h39dbdc08),
	.w2(32'h3947796b),
	.w3(32'h3bbd5986),
	.w4(32'h39198fa1),
	.w5(32'h38a2532b),
	.w6(32'h3a40ce38),
	.w7(32'h39c97ec0),
	.w8(32'hb9bb37d9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba202615),
	.w1(32'hba41e324),
	.w2(32'hba91bbd6),
	.w3(32'hba163b34),
	.w4(32'hba610dc9),
	.w5(32'hbabfc78e),
	.w6(32'hbab1074d),
	.w7(32'hbab3edf5),
	.w8(32'hba34e135),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba011fb6),
	.w1(32'hba3befbc),
	.w2(32'hb969b7a7),
	.w3(32'hbab677a5),
	.w4(32'hba3c5528),
	.w5(32'hb90de45f),
	.w6(32'hba9aaf98),
	.w7(32'hba5692e6),
	.w8(32'hb9506243),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934361f),
	.w1(32'hb924ea27),
	.w2(32'hba17803e),
	.w3(32'h39254030),
	.w4(32'hba13d953),
	.w5(32'hba6c4211),
	.w6(32'h39b0042e),
	.w7(32'hb95c1b75),
	.w8(32'hba31dbb7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76db63),
	.w1(32'h39b10f12),
	.w2(32'hb918fd68),
	.w3(32'hbaa2fddc),
	.w4(32'hb96f1201),
	.w5(32'hba5f8ecc),
	.w6(32'h3a54a1f8),
	.w7(32'h3980ffdf),
	.w8(32'hb9885911),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba321f66),
	.w1(32'h39fcc833),
	.w2(32'h396a6093),
	.w3(32'hba7f1898),
	.w4(32'hb793255b),
	.w5(32'hba2741c3),
	.w6(32'h3aa1e266),
	.w7(32'h3a078946),
	.w8(32'h3a254d39),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c0fae1),
	.w1(32'hb95b1f84),
	.w2(32'hb91028fb),
	.w3(32'hb9b9df80),
	.w4(32'hba487518),
	.w5(32'hba1c00b1),
	.w6(32'hb992f705),
	.w7(32'hb8bcf68f),
	.w8(32'h38c8667c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0944b6),
	.w1(32'hbb3e6511),
	.w2(32'hbb21d941),
	.w3(32'hba2714d5),
	.w4(32'hba83b407),
	.w5(32'hba9d29b7),
	.w6(32'hbb090aa1),
	.w7(32'hbab4705b),
	.w8(32'hbaedea3e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51b1c8),
	.w1(32'h3a115b2d),
	.w2(32'h394f1e97),
	.w3(32'hba26f031),
	.w4(32'hb9bc34d8),
	.w5(32'hba8189b8),
	.w6(32'h3a33a417),
	.w7(32'h394fbbac),
	.w8(32'hba1b41b9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41fcc3),
	.w1(32'hba94c947),
	.w2(32'hbabed050),
	.w3(32'hbae848d9),
	.w4(32'hbaa2c5f4),
	.w5(32'hbab470a4),
	.w6(32'hbaade29f),
	.w7(32'hbac66aaa),
	.w8(32'hba3a8b52),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ba941),
	.w1(32'hba7c3733),
	.w2(32'h3a85374d),
	.w3(32'hba4a5fe9),
	.w4(32'h3992f933),
	.w5(32'h3ab04e87),
	.w6(32'hbb33d983),
	.w7(32'hba3a94a0),
	.w8(32'h3ad013b5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16b59f),
	.w1(32'h3ae2561c),
	.w2(32'h3a908fdf),
	.w3(32'h3b4aafdd),
	.w4(32'h3a95a17e),
	.w5(32'h39963b15),
	.w6(32'h3b17f2a4),
	.w7(32'h3aac3433),
	.w8(32'h3a283d71),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381bf5f3),
	.w1(32'h3ba18c17),
	.w2(32'h3ba1f47b),
	.w3(32'h39108164),
	.w4(32'h3b1af85e),
	.w5(32'h3b3966be),
	.w6(32'h3bdce941),
	.w7(32'h3bb71acb),
	.w8(32'h3b9b555c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6f8a3),
	.w1(32'h391ef4fe),
	.w2(32'h39e42f9f),
	.w3(32'h3b916041),
	.w4(32'hb962d2d4),
	.w5(32'h38d307b9),
	.w6(32'hb926be35),
	.w7(32'hb553ff95),
	.w8(32'h390e7e1e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fbbf9d),
	.w1(32'h3a2094ee),
	.w2(32'h3a4c4aa1),
	.w3(32'h39a41ddd),
	.w4(32'h3953f7cc),
	.w5(32'h395829ff),
	.w6(32'h39cc0d6b),
	.w7(32'h3a68d41d),
	.w8(32'h3a4b0dbd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d71821),
	.w1(32'h39c56d49),
	.w2(32'h39d67a9b),
	.w3(32'hb7318016),
	.w4(32'h3997b7c4),
	.w5(32'h39a9cead),
	.w6(32'hb9e7c01b),
	.w7(32'hb9e4bdb4),
	.w8(32'hb8cb2418),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad6703),
	.w1(32'h3aa08bb9),
	.w2(32'hb9a521b7),
	.w3(32'h39b3d5de),
	.w4(32'hb9b0469d),
	.w5(32'hbacdb61d),
	.w6(32'h3bb27942),
	.w7(32'h3b872508),
	.w8(32'h3bb57ea4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a8f65),
	.w1(32'hb92016c7),
	.w2(32'h39b33880),
	.w3(32'h3b3ea0cc),
	.w4(32'h39882567),
	.w5(32'h3a98ef5f),
	.w6(32'hba05554d),
	.w7(32'hb98264ab),
	.w8(32'hb8bfc542),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55a038),
	.w1(32'hba69ac29),
	.w2(32'hbacb360e),
	.w3(32'h3a9e0a15),
	.w4(32'hba51d5a6),
	.w5(32'hbad0fc3c),
	.w6(32'hb97c5ebc),
	.w7(32'hba2b52f1),
	.w8(32'hba9112e4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0a901),
	.w1(32'h3a8b7dc8),
	.w2(32'h3a739ccb),
	.w3(32'hbaa9d5ee),
	.w4(32'h3a443dd4),
	.w5(32'h39f30345),
	.w6(32'h3af0bcf7),
	.w7(32'h3aa9a040),
	.w8(32'h3a56efe2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be2483),
	.w1(32'hb9dfc347),
	.w2(32'hb8a41324),
	.w3(32'h39953722),
	.w4(32'h389bbc25),
	.w5(32'h3a476a91),
	.w6(32'hba80a665),
	.w7(32'hba345579),
	.w8(32'hb9ed6074),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375ee8ae),
	.w1(32'h3ac9b627),
	.w2(32'h3a9ea1ee),
	.w3(32'h3a21505b),
	.w4(32'h3a6a422f),
	.w5(32'h39d37112),
	.w6(32'h3b16b1be),
	.w7(32'h3abb8975),
	.w8(32'h3a752106),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398cc221),
	.w1(32'h3aae81c9),
	.w2(32'h3a5891ef),
	.w3(32'h39b27c5c),
	.w4(32'h39be87ed),
	.w5(32'hb95b0807),
	.w6(32'h3b1dd4d6),
	.w7(32'h3ad88005),
	.w8(32'h3aa39a40),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d70b3),
	.w1(32'hb9988d7d),
	.w2(32'h39e56b54),
	.w3(32'hb9a464c6),
	.w4(32'h3928e4ac),
	.w5(32'h3a94e12e),
	.w6(32'hbab066ef),
	.w7(32'hba52b1ea),
	.w8(32'hb98222b5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7fc040),
	.w1(32'hba299f5b),
	.w2(32'hb96daf89),
	.w3(32'h3a97344c),
	.w4(32'hba03dc55),
	.w5(32'h39071f2a),
	.w6(32'hba60ca97),
	.w7(32'hba2b3d50),
	.w8(32'hb9f73a17),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b99fd6),
	.w1(32'h3ba6ac0a),
	.w2(32'h3b99a56a),
	.w3(32'h38f49dbe),
	.w4(32'h3b43a36c),
	.w5(32'h3b49cc3a),
	.w6(32'h3bcc2c84),
	.w7(32'h3b9db544),
	.w8(32'h3b860939),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ca8c2),
	.w1(32'hba981a00),
	.w2(32'hbabd2a9c),
	.w3(32'h3b4dff42),
	.w4(32'hbad1a5a6),
	.w5(32'hbad22f04),
	.w6(32'hbaf661ec),
	.w7(32'hbac9263d),
	.w8(32'hbac52cc3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbd7ee),
	.w1(32'hba5cedc8),
	.w2(32'hba36593a),
	.w3(32'hbab89f8e),
	.w4(32'hb9a8cf14),
	.w5(32'h3875825a),
	.w6(32'hb9914a22),
	.w7(32'hb9ce3e4a),
	.w8(32'hba2a16a0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8862db8),
	.w1(32'h3b7ea8b0),
	.w2(32'h3b9a574f),
	.w3(32'hb8b57316),
	.w4(32'h3abcdcde),
	.w5(32'h3b3d0409),
	.w6(32'h3a81c3c3),
	.w7(32'h3b18948c),
	.w8(32'h3b15de34),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a52de),
	.w1(32'hb7dbf7ae),
	.w2(32'hba121071),
	.w3(32'h3b4b00cb),
	.w4(32'h3916ac39),
	.w5(32'hb9e67d7e),
	.w6(32'hb874570d),
	.w7(32'hb9ac8e0a),
	.w8(32'hbac7ff3e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2c690),
	.w1(32'hba8fbb6a),
	.w2(32'hb9af9351),
	.w3(32'hba88ec20),
	.w4(32'hba99f5d8),
	.w5(32'hba44ce2f),
	.w6(32'hbac2442c),
	.w7(32'hba72f7cd),
	.w8(32'hba07e657),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c23dd),
	.w1(32'h3ac172d5),
	.w2(32'h3aff9e8f),
	.w3(32'hb9bc482a),
	.w4(32'h3a80b3ef),
	.w5(32'h3aaa173a),
	.w6(32'h3a73cafd),
	.w7(32'h3a883b41),
	.w8(32'h3a8ac425),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8458b8),
	.w1(32'hbb36058a),
	.w2(32'hbac985a3),
	.w3(32'h3a9b44cd),
	.w4(32'hbb059aba),
	.w5(32'hb8019687),
	.w6(32'hbb5781e2),
	.w7(32'hbb1cd1cf),
	.w8(32'hba8e9979),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e492bf),
	.w1(32'hba491d2a),
	.w2(32'hbaf9903a),
	.w3(32'hba881732),
	.w4(32'hba936691),
	.w5(32'hb9c8ac18),
	.w6(32'hba245e00),
	.w7(32'hbafa2711),
	.w8(32'hba9fafc1),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1384a5),
	.w1(32'h3a40ee79),
	.w2(32'h399daf30),
	.w3(32'hb8a37aa4),
	.w4(32'hba0c1e0a),
	.w5(32'hbabd7cb0),
	.w6(32'h3a85e027),
	.w7(32'h398e1558),
	.w8(32'hba681743),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa04b2d),
	.w1(32'hb99a1f3f),
	.w2(32'hba17aa35),
	.w3(32'hbb30b960),
	.w4(32'hb9fa912b),
	.w5(32'hba73cd47),
	.w6(32'h3896cbeb),
	.w7(32'hb9b67db3),
	.w8(32'hba46e779),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f3565),
	.w1(32'h399743a7),
	.w2(32'h37b4b237),
	.w3(32'hbab500f1),
	.w4(32'hb9c441c6),
	.w5(32'hba5ae3f5),
	.w6(32'h39f87e3b),
	.w7(32'h388eac11),
	.w8(32'hba0ffc73),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba281583),
	.w1(32'hb9b02bb5),
	.w2(32'hba8984a0),
	.w3(32'hbab9926b),
	.w4(32'hb9a57fcc),
	.w5(32'hbab7d698),
	.w6(32'hb9b8106a),
	.w7(32'hba446999),
	.w8(32'hba0203c5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba350cf3),
	.w1(32'hbab4f623),
	.w2(32'hbadcaf85),
	.w3(32'hba1b1546),
	.w4(32'hbae00abb),
	.w5(32'hbad65111),
	.w6(32'hbaca2dc4),
	.w7(32'hbab4756d),
	.w8(32'hba70dab3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3962a),
	.w1(32'h3af90e8c),
	.w2(32'h3ad0824b),
	.w3(32'hbac09f7b),
	.w4(32'h3a12b243),
	.w5(32'h39306c33),
	.w6(32'h3b4042d5),
	.w7(32'h3b15c38d),
	.w8(32'h3ac82f54),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bca94),
	.w1(32'h3a07050b),
	.w2(32'h3915a561),
	.w3(32'h378bb657),
	.w4(32'hb94a284f),
	.w5(32'hba465088),
	.w6(32'h3a107f4d),
	.w7(32'h394aa349),
	.w8(32'hb9fe7a18),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31ceb1),
	.w1(32'hba492e28),
	.w2(32'hb9aae780),
	.w3(32'hbac20c97),
	.w4(32'hba4bab32),
	.w5(32'hba230077),
	.w6(32'hbab7d65e),
	.w7(32'hbaa52297),
	.w8(32'hbabc4c61),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72975d),
	.w1(32'h39a59ec1),
	.w2(32'hb887fd82),
	.w3(32'hba682c98),
	.w4(32'hba1dc8a9),
	.w5(32'hba923f9f),
	.w6(32'h3a74e235),
	.w7(32'h39f06282),
	.w8(32'hb86d82ea),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51b2ba),
	.w1(32'hba8c9c0c),
	.w2(32'hbb0befae),
	.w3(32'hba63321f),
	.w4(32'hb98a3f8a),
	.w5(32'hba8b3771),
	.w6(32'hb9050ebf),
	.w7(32'hba9230bc),
	.w8(32'hbae84c10),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f3c24),
	.w1(32'h39d127e4),
	.w2(32'h390aebfb),
	.w3(32'hbad0b3f3),
	.w4(32'hb895a216),
	.w5(32'hba123644),
	.w6(32'h3a718209),
	.w7(32'h39e8432c),
	.w8(32'h38d60f4b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fccceb),
	.w1(32'hba9a1682),
	.w2(32'hbaecf7d6),
	.w3(32'hba1cc310),
	.w4(32'hba9004f7),
	.w5(32'hbabfe15a),
	.w6(32'hba985e8f),
	.w7(32'hba6d974d),
	.w8(32'hba2e61ff),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd3b52),
	.w1(32'hba19f32d),
	.w2(32'hbaa745d4),
	.w3(32'hba99d115),
	.w4(32'hba01a423),
	.w5(32'hba88a301),
	.w6(32'h387e6970),
	.w7(32'hba7080eb),
	.w8(32'hba3519b9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2a727),
	.w1(32'h3a2f9a26),
	.w2(32'h39769a8d),
	.w3(32'hba9dce7e),
	.w4(32'hb9bfd392),
	.w5(32'hba92b093),
	.w6(32'h3a531ab1),
	.w7(32'h399bbc17),
	.w8(32'hba28721e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ef8b9),
	.w1(32'hb8775e21),
	.w2(32'hba0c422c),
	.w3(32'hbb0474c5),
	.w4(32'hba034d42),
	.w5(32'hba89a262),
	.w6(32'h39be2ae6),
	.w7(32'hb8e6176c),
	.w8(32'hba0bf02a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba889c39),
	.w1(32'hb6b4d7fa),
	.w2(32'hba0d7c4f),
	.w3(32'hbaaaf8ff),
	.w4(32'hba107b0c),
	.w5(32'hba9d4504),
	.w6(32'h39eaeb9d),
	.w7(32'hb8a20898),
	.w8(32'hba0bef30),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba964f72),
	.w1(32'hbaee3b7a),
	.w2(32'hbac4abdf),
	.w3(32'hbabed4fd),
	.w4(32'hba611fed),
	.w5(32'hba26075e),
	.w6(32'hba7d9371),
	.w7(32'hb9d459a5),
	.w8(32'hba878fcc),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb107397),
	.w1(32'hbb019508),
	.w2(32'hbaf8b7bd),
	.w3(32'hbab4889a),
	.w4(32'hbb004be7),
	.w5(32'hbac47013),
	.w6(32'hbb149e13),
	.w7(32'hbaf6e200),
	.w8(32'hb895695b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994ed04),
	.w1(32'hba8c0916),
	.w2(32'hbae5ff15),
	.w3(32'hb9954547),
	.w4(32'hbac42a4d),
	.w5(32'hbb0f1261),
	.w6(32'hba1bf26c),
	.w7(32'hba90f546),
	.w8(32'hba87992d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9c8c6),
	.w1(32'hba203676),
	.w2(32'hbaade73b),
	.w3(32'hbaee70b8),
	.w4(32'hba02a362),
	.w5(32'hba94d29f),
	.w6(32'hba221a4a),
	.w7(32'hba870f45),
	.w8(32'hbacd95b0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9cfee),
	.w1(32'h3a02f7cf),
	.w2(32'hb785f9ee),
	.w3(32'hbaa83eea),
	.w4(32'hb8a1857c),
	.w5(32'hba56597e),
	.w6(32'h3a801195),
	.w7(32'h39e7affc),
	.w8(32'hb96f0377),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fc326),
	.w1(32'hbadb296b),
	.w2(32'hbaa9354d),
	.w3(32'hbaa335ad),
	.w4(32'hba20089c),
	.w5(32'h3a30c4c2),
	.w6(32'hba981828),
	.w7(32'hba7308c0),
	.w8(32'hbac49b12),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c7a84),
	.w1(32'h3895a811),
	.w2(32'h3964cc05),
	.w3(32'h3a244ae2),
	.w4(32'hb9ef767f),
	.w5(32'h38a19433),
	.w6(32'hb964b46a),
	.w7(32'hba85bc61),
	.w8(32'hba82a23c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8519553),
	.w1(32'h3ad3aa06),
	.w2(32'h3a88d8af),
	.w3(32'hb912e6b4),
	.w4(32'h3a7610c2),
	.w5(32'hb81a110a),
	.w6(32'h3b31aec2),
	.w7(32'h3ae1a6b8),
	.w8(32'h3a8d0633),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d53e6),
	.w1(32'hb9ffddf3),
	.w2(32'hb990c827),
	.w3(32'hb7fb01a6),
	.w4(32'hb9f5694d),
	.w5(32'hb90ba24f),
	.w6(32'hb9def646),
	.w7(32'hb8d44f14),
	.w8(32'hb9166030),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b74a72),
	.w1(32'hba46c41f),
	.w2(32'hba2d150d),
	.w3(32'hb908a0d6),
	.w4(32'hba3dd199),
	.w5(32'hba4026f6),
	.w6(32'hba3c0f08),
	.w7(32'hba4d616a),
	.w8(32'hba40fb6d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ae910),
	.w1(32'hb9c1ef2d),
	.w2(32'hb9e2bb3a),
	.w3(32'hba24ded1),
	.w4(32'h396d8dd9),
	.w5(32'hb912fb1e),
	.w6(32'hb9600cf2),
	.w7(32'h39cbd9f5),
	.w8(32'h39de0d2f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b61e1a),
	.w1(32'h3919356d),
	.w2(32'h39b2ace3),
	.w3(32'hba72c6de),
	.w4(32'hb71e637a),
	.w5(32'h390022af),
	.w6(32'h3950429c),
	.w7(32'h399c7192),
	.w8(32'h393c619e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe8453),
	.w1(32'hb775469c),
	.w2(32'h392694de),
	.w3(32'h38fe18e1),
	.w4(32'hb91e2bc4),
	.w5(32'hb8a64b88),
	.w6(32'hb7740fa1),
	.w7(32'hb95bb99a),
	.w8(32'hb9b620cc),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9936eee),
	.w1(32'hba5603fa),
	.w2(32'hba1dc30a),
	.w3(32'hb97a843e),
	.w4(32'h39b431ee),
	.w5(32'hb90952c9),
	.w6(32'h39951bb0),
	.w7(32'hb9d96d13),
	.w8(32'hb9b584eb),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9193f10),
	.w1(32'h39a03564),
	.w2(32'hb8db8dd4),
	.w3(32'hb9819ca1),
	.w4(32'h3a09821e),
	.w5(32'hba2177c0),
	.w6(32'h393c7682),
	.w7(32'hb93acb77),
	.w8(32'h39f01428),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c47d2),
	.w1(32'hb913b5c8),
	.w2(32'hb8201e43),
	.w3(32'hb8015143),
	.w4(32'hb8615d72),
	.w5(32'hb942b800),
	.w6(32'hb95d2fda),
	.w7(32'hb926fdb8),
	.w8(32'hb9701a4e),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cae74c),
	.w1(32'hb8079f0e),
	.w2(32'h395f4763),
	.w3(32'hb97287cf),
	.w4(32'hb9968c58),
	.w5(32'hb8c26be8),
	.w6(32'h37b7bced),
	.w7(32'h3943730c),
	.w8(32'h39917003),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b09b6),
	.w1(32'hb9e4c820),
	.w2(32'hb9c1ed5a),
	.w3(32'h392bbe40),
	.w4(32'hb977a5fb),
	.w5(32'hb96e7773),
	.w6(32'hb9de0195),
	.w7(32'hb99aa9b1),
	.w8(32'hb9b69582),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edcdc2),
	.w1(32'hba32324b),
	.w2(32'hb9da8836),
	.w3(32'hb95e5638),
	.w4(32'hba355fa5),
	.w5(32'hba094914),
	.w6(32'hba125ce0),
	.w7(32'hb9fa2e18),
	.w8(32'hb9929a8b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a1a98),
	.w1(32'h391d828a),
	.w2(32'h399b6e5e),
	.w3(32'hb9c6177e),
	.w4(32'h37eb8362),
	.w5(32'h398641af),
	.w6(32'h39358aa3),
	.w7(32'h39c29804),
	.w8(32'h3a70887d),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a204a6b),
	.w1(32'hb9cdf62a),
	.w2(32'hb935f226),
	.w3(32'h3a0674f3),
	.w4(32'h39649237),
	.w5(32'h3a29cdca),
	.w6(32'hba4ba980),
	.w7(32'hba273eaf),
	.w8(32'hba54dd80),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4ec79),
	.w1(32'hba052b3b),
	.w2(32'hb9273d4c),
	.w3(32'h399e375e),
	.w4(32'hba1a6931),
	.w5(32'hba336795),
	.w6(32'hba4438cd),
	.w7(32'hba4699a3),
	.w8(32'hba2b3e54),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b4329d),
	.w1(32'hba262617),
	.w2(32'hba10ab97),
	.w3(32'hba14f135),
	.w4(32'hba0cdc7e),
	.w5(32'hb9b3bf43),
	.w6(32'hba30f9cf),
	.w7(32'hb9fd9902),
	.w8(32'hb9e071a0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0f422),
	.w1(32'hba1da77b),
	.w2(32'hb81f6bc8),
	.w3(32'hb99e1a09),
	.w4(32'hb960caf9),
	.w5(32'h38961752),
	.w6(32'hb97a310b),
	.w7(32'h37f3c80d),
	.w8(32'h3888cbed),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a62d8a),
	.w1(32'hba97819a),
	.w2(32'hb9df76c0),
	.w3(32'h39ae6051),
	.w4(32'h394a55bc),
	.w5(32'hbab96c0a),
	.w6(32'hbab2a407),
	.w7(32'hba96a6d8),
	.w8(32'hba23af29),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2da573),
	.w1(32'hba2e0eea),
	.w2(32'hba0d86f1),
	.w3(32'hba6e9021),
	.w4(32'hba3c2e47),
	.w5(32'hba065eaf),
	.w6(32'hba242035),
	.w7(32'hba12d37c),
	.w8(32'hb9f0550b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba319012),
	.w1(32'h3a77cdeb),
	.w2(32'h3a8e6898),
	.w3(32'hb9ad6462),
	.w4(32'h3a1846dc),
	.w5(32'h3a017584),
	.w6(32'h39a482ad),
	.w7(32'h39033c15),
	.w8(32'h3716b89f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12abe5),
	.w1(32'hb7077023),
	.w2(32'h3995edf1),
	.w3(32'h39c6a96b),
	.w4(32'hb9441921),
	.w5(32'h371d4c8e),
	.w6(32'hb96538c7),
	.w7(32'hb9104cc1),
	.w8(32'hb94fefdf),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968feb7),
	.w1(32'hb9733e09),
	.w2(32'h38e86f6e),
	.w3(32'hb8e55250),
	.w4(32'hba061495),
	.w5(32'hb9abf6e1),
	.w6(32'hb950320c),
	.w7(32'hb89b9abf),
	.w8(32'hb92ce083),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987706d),
	.w1(32'hb99df6fd),
	.w2(32'hb91bcce6),
	.w3(32'hb9925202),
	.w4(32'hb9c4576a),
	.w5(32'hb8f82591),
	.w6(32'hb9a5a132),
	.w7(32'hb9880cdb),
	.w8(32'hb91d6daa),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9beba),
	.w1(32'hb91c944e),
	.w2(32'h39124d95),
	.w3(32'hb93cb9cb),
	.w4(32'h3937bcc7),
	.w5(32'h3a0dc33e),
	.w6(32'h38d692ef),
	.w7(32'h398d3633),
	.w8(32'h39e1998b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974549f),
	.w1(32'hbaa65671),
	.w2(32'hb9a78fb0),
	.w3(32'h39e13efa),
	.w4(32'hba25d14d),
	.w5(32'hb9dda147),
	.w6(32'h3895064b),
	.w7(32'h39805886),
	.w8(32'hba7c129f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb935b5ec),
	.w1(32'h397b6f15),
	.w2(32'h3a3ee0c8),
	.w3(32'hba5772b5),
	.w4(32'hb906c3d9),
	.w5(32'h39a5c023),
	.w6(32'h3981bd43),
	.w7(32'h39e4f9df),
	.w8(32'hb98b2a73),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1320f),
	.w1(32'hba146314),
	.w2(32'hb99c7ed4),
	.w3(32'hba192c97),
	.w4(32'hb9f632a6),
	.w5(32'hb9a0315f),
	.w6(32'hba0fdd6e),
	.w7(32'hb9d2ba6c),
	.w8(32'hb9b99a20),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d148c5),
	.w1(32'h39113b5c),
	.w2(32'hb834408d),
	.w3(32'hb9308c47),
	.w4(32'h397f39c8),
	.w5(32'h39a5cc0d),
	.w6(32'h39f22502),
	.w7(32'h398f845e),
	.w8(32'h39334568),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9678348),
	.w1(32'hba222c24),
	.w2(32'hb9bee69a),
	.w3(32'h39b6cf30),
	.w4(32'hb9a7d1ac),
	.w5(32'hb9bc546d),
	.w6(32'hba81376c),
	.w7(32'hba42850e),
	.w8(32'hba8ae6a9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5db24d),
	.w1(32'hba469052),
	.w2(32'hb9e2c77b),
	.w3(32'hba5ca362),
	.w4(32'hb9db6740),
	.w5(32'hb9a7a159),
	.w6(32'hba03d5fe),
	.w7(32'hb96660ea),
	.w8(32'hb992477d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ced9c),
	.w1(32'hba83fd5a),
	.w2(32'hba8b1420),
	.w3(32'hb9b74aa5),
	.w4(32'hba3f9ce2),
	.w5(32'hba76681e),
	.w6(32'hba4e1379),
	.w7(32'hba3171b1),
	.w8(32'hba40ec0d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1bbb6),
	.w1(32'hb9b8469d),
	.w2(32'h3a5727b3),
	.w3(32'hba68b3f6),
	.w4(32'hba12842a),
	.w5(32'h3a19e3d3),
	.w6(32'h38674a92),
	.w7(32'h3a4ac172),
	.w8(32'h3943a453),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c629bb),
	.w1(32'h3aac126f),
	.w2(32'h3ac3ab5e),
	.w3(32'hb74d5f4d),
	.w4(32'h3a56cbfc),
	.w5(32'h3a7f1c9d),
	.w6(32'h3a33ffb3),
	.w7(32'h3a2db36d),
	.w8(32'h3a1201b7),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf288c),
	.w1(32'hb8618157),
	.w2(32'h3830e526),
	.w3(32'h3a886729),
	.w4(32'h39516982),
	.w5(32'h39a9e06b),
	.w6(32'h38288e32),
	.w7(32'h38a6ed41),
	.w8(32'h39587532),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a5f30c),
	.w1(32'hba00746e),
	.w2(32'hb9728043),
	.w3(32'h3943a82b),
	.w4(32'hb9ef2491),
	.w5(32'hb97b3788),
	.w6(32'hb9e6fd07),
	.w7(32'hb9b368a3),
	.w8(32'hb9c27eba),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e96ba0),
	.w1(32'hba36cedb),
	.w2(32'h37d335ae),
	.w3(32'hb9c083bb),
	.w4(32'hba192534),
	.w5(32'hb9979307),
	.w6(32'hb9f950b2),
	.w7(32'hb9454f95),
	.w8(32'h3937c1b9),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39009cb3),
	.w1(32'hba216017),
	.w2(32'hb9924ee3),
	.w3(32'h397629be),
	.w4(32'hba5048a4),
	.w5(32'hb8cabfc3),
	.w6(32'hba8e3f1f),
	.w7(32'hba28e86a),
	.w8(32'hba70ad91),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62e931),
	.w1(32'hb92249e8),
	.w2(32'h386f1b3e),
	.w3(32'hba87d04f),
	.w4(32'hb98b5448),
	.w5(32'hb7b0fcb0),
	.w6(32'hb8573194),
	.w7(32'h396a0f88),
	.w8(32'h39ed5990),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81b9282),
	.w1(32'hb98c2b53),
	.w2(32'hb8883a3e),
	.w3(32'h38972f08),
	.w4(32'hb73aa5ec),
	.w5(32'h38c9f371),
	.w6(32'hb9952d5b),
	.w7(32'hb994f277),
	.w8(32'hb9cf7cc6),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9859937),
	.w1(32'h39c25838),
	.w2(32'h3a595a3a),
	.w3(32'h37584980),
	.w4(32'h39ccef63),
	.w5(32'h39d91866),
	.w6(32'h3938eb30),
	.w7(32'h39ed5862),
	.w8(32'h3a0b08a3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a421863),
	.w1(32'h39044e03),
	.w2(32'h39f2a47a),
	.w3(32'h3a28d657),
	.w4(32'hb8052a1e),
	.w5(32'h392511d3),
	.w6(32'h38a2891a),
	.w7(32'h398d8094),
	.w8(32'h389cf5de),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ab3082),
	.w1(32'hba3e86cd),
	.w2(32'hba0bf151),
	.w3(32'h3820abd6),
	.w4(32'hba1d3385),
	.w5(32'hba0d7904),
	.w6(32'hba1d79d8),
	.w7(32'hba0c29b5),
	.w8(32'hba17c9f3),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba490083),
	.w1(32'hb8ef1d0d),
	.w2(32'h39125023),
	.w3(32'hba1b6c88),
	.w4(32'hb99a734c),
	.w5(32'hb959d238),
	.w6(32'hb8080895),
	.w7(32'h392d7256),
	.w8(32'h38eb760c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37364b75),
	.w1(32'h3a6783b7),
	.w2(32'h3a828f59),
	.w3(32'h37bcb960),
	.w4(32'h3a3ae074),
	.w5(32'h3a3cb9f3),
	.w6(32'h3a2f595a),
	.w7(32'h3a4aee76),
	.w8(32'h3a384d24),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91a800),
	.w1(32'h3978c21a),
	.w2(32'h39ca3b93),
	.w3(32'h3a640c85),
	.w4(32'h39921fb9),
	.w5(32'h39e816e7),
	.w6(32'h36ee8f73),
	.w7(32'h374ba7f3),
	.w8(32'hb98fb22b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398cb472),
	.w1(32'hba338582),
	.w2(32'hb9d4b347),
	.w3(32'h398b1c1d),
	.w4(32'hba354370),
	.w5(32'hb9f20d40),
	.w6(32'hba4887e6),
	.w7(32'hba0b401a),
	.w8(32'hba2befee),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ff381),
	.w1(32'h3a1e5eff),
	.w2(32'h3a1113ea),
	.w3(32'hba0a599b),
	.w4(32'h3a3dc5bb),
	.w5(32'h3a2dadda),
	.w6(32'h3a527a6f),
	.w7(32'h3a40d804),
	.w8(32'h3aa2ee8f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e5281),
	.w1(32'hb9bc3640),
	.w2(32'h39427ccd),
	.w3(32'h3a9d31d1),
	.w4(32'hb8abd03a),
	.w5(32'h39a80d80),
	.w6(32'h399e7d74),
	.w7(32'h39d121c0),
	.w8(32'h395f8da6),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373b4999),
	.w1(32'hba5757e8),
	.w2(32'hba9b25f2),
	.w3(32'h3a482953),
	.w4(32'hba685522),
	.w5(32'hba6b95fe),
	.w6(32'hb9b7edf9),
	.w7(32'hba061f62),
	.w8(32'hba3934f3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba880aff),
	.w1(32'hba2c2c68),
	.w2(32'h39e6bcf0),
	.w3(32'hb9db657c),
	.w4(32'h3856b312),
	.w5(32'hba22ab2d),
	.w6(32'h397b3962),
	.w7(32'hb883243b),
	.w8(32'h38042061),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bf703),
	.w1(32'h39aba4fc),
	.w2(32'h3a707afe),
	.w3(32'hba3f779c),
	.w4(32'h37a77645),
	.w5(32'h3a43ecc5),
	.w6(32'h396c2941),
	.w7(32'h39aa248c),
	.w8(32'h392f7022),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3957ac64),
	.w1(32'hba0066ab),
	.w2(32'hb8c39574),
	.w3(32'h389b57d0),
	.w4(32'hba1d1da6),
	.w5(32'hb95a7c96),
	.w6(32'hba12268d),
	.w7(32'hb99ce524),
	.w8(32'hb97c4a05),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8600a),
	.w1(32'hb9d5bda0),
	.w2(32'hb999f699),
	.w3(32'hb9dda9b0),
	.w4(32'hb943c392),
	.w5(32'hb8f2b02b),
	.w6(32'hb9b0eedf),
	.w7(32'hb9609510),
	.w8(32'hb98692e0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9927eef),
	.w1(32'h396d0904),
	.w2(32'hb8986c95),
	.w3(32'h37871421),
	.w4(32'h39a7d59d),
	.w5(32'h39252aa2),
	.w6(32'hb71aef15),
	.w7(32'h3694227b),
	.w8(32'h39ae5f95),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378375c0),
	.w1(32'h39b39d2b),
	.w2(32'hb955e9e7),
	.w3(32'h38932ae3),
	.w4(32'hb9f03cdc),
	.w5(32'hb95aac67),
	.w6(32'h39d3e548),
	.w7(32'h39f9d74a),
	.w8(32'hba0e2f2b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5823e),
	.w1(32'h3984f79b),
	.w2(32'h39022908),
	.w3(32'hb9874821),
	.w4(32'h39b1e198),
	.w5(32'h392fe3f9),
	.w6(32'h39a5040f),
	.w7(32'h399f0c14),
	.w8(32'h39d740f6),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e5477c),
	.w1(32'h39777f9d),
	.w2(32'h3a107764),
	.w3(32'h39d23a1f),
	.w4(32'h39803309),
	.w5(32'h392b8561),
	.w6(32'h3997db32),
	.w7(32'h39f7e856),
	.w8(32'h3a090669),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a542d2a),
	.w1(32'hb962909a),
	.w2(32'h39a96efc),
	.w3(32'h3a0231e4),
	.w4(32'hb92deb66),
	.w5(32'h382fd551),
	.w6(32'h3892a038),
	.w7(32'h39402c7f),
	.w8(32'hb77949e7),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38059dd9),
	.w1(32'h3a830ff4),
	.w2(32'h3a8a578d),
	.w3(32'hb929a730),
	.w4(32'h3a5aab6e),
	.w5(32'h3a74e4b7),
	.w6(32'h3aa7fdcb),
	.w7(32'h3a723dd4),
	.w8(32'h3a1e8639),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28b730),
	.w1(32'hb9b5b475),
	.w2(32'hb9ce6a16),
	.w3(32'h3a2d99f7),
	.w4(32'hb917aa10),
	.w5(32'hb98843d5),
	.w6(32'hb914b6a9),
	.w7(32'hb9b9429e),
	.w8(32'hba367aa1),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba817380),
	.w1(32'h392a2612),
	.w2(32'hba7d9104),
	.w3(32'hba028cc6),
	.w4(32'hb95ace03),
	.w5(32'hbaa29f5f),
	.w6(32'hb9c384a5),
	.w7(32'hba3435e9),
	.w8(32'hba2c0fdc),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15a76b),
	.w1(32'hb85750e7),
	.w2(32'h399ba70b),
	.w3(32'hba63a074),
	.w4(32'hb9695b9c),
	.w5(32'h38bd67ab),
	.w6(32'h392ac654),
	.w7(32'h398ebda0),
	.w8(32'h389f8c17),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9125483),
	.w1(32'hba5a44a1),
	.w2(32'hba08b26f),
	.w3(32'h3715a784),
	.w4(32'hba2d1c13),
	.w5(32'hba0d5fbf),
	.w6(32'hba3b71fb),
	.w7(32'hba02a863),
	.w8(32'hb9fc84bc),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3239dc),
	.w1(32'hb951d3e0),
	.w2(32'h3939b451),
	.w3(32'hb9f3dbfb),
	.w4(32'hb9bc283e),
	.w5(32'hb9b70758),
	.w6(32'hb915f38e),
	.w7(32'h38f0181d),
	.w8(32'hb98a7b1d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cabb97),
	.w1(32'hb9f0a7ac),
	.w2(32'h38905d5c),
	.w3(32'hb9d59dd0),
	.w4(32'hb894abe0),
	.w5(32'h38f07943),
	.w6(32'hb9234dff),
	.w7(32'h394e0a62),
	.w8(32'h394ad753),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3845f7f9),
	.w1(32'hba95e0bd),
	.w2(32'hb9a11a9f),
	.w3(32'h390bb79f),
	.w4(32'hbac8b0ef),
	.w5(32'hba95028d),
	.w6(32'hba55a1d0),
	.w7(32'hb8fb63a7),
	.w8(32'hba37fd58),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba779494),
	.w1(32'h39815daa),
	.w2(32'h397a31a3),
	.w3(32'hba447cfe),
	.w4(32'h398ca25e),
	.w5(32'h3971920b),
	.w6(32'h39c95570),
	.w7(32'h39b8c810),
	.w8(32'h3a464710),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b45d0),
	.w1(32'hb9990be9),
	.w2(32'h38d35e9a),
	.w3(32'h3a3275be),
	.w4(32'hb9dc8c91),
	.w5(32'hb9a8408b),
	.w6(32'hb958d1a1),
	.w7(32'hb9074f1f),
	.w8(32'hb95df728),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946b99a),
	.w1(32'hba0c5c54),
	.w2(32'hbaa173f3),
	.w3(32'hb9822cc7),
	.w4(32'hba3c59fa),
	.w5(32'hba82135d),
	.w6(32'hba115a3a),
	.w7(32'hba31ae30),
	.w8(32'hba90b46a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba850e8e),
	.w1(32'h3a39a94c),
	.w2(32'h3a42453b),
	.w3(32'hba49bd88),
	.w4(32'h3a042f14),
	.w5(32'h396c61dc),
	.w6(32'h39a3c620),
	.w7(32'h396ae915),
	.w8(32'h38f4abfa),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6aa3d6),
	.w1(32'h39657c4a),
	.w2(32'h39f6a5a1),
	.w3(32'h39bad2bf),
	.w4(32'h38331a28),
	.w5(32'h39cc8e65),
	.w6(32'h39a3f93d),
	.w7(32'h3a038a9d),
	.w8(32'h3915a78e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce5567),
	.w1(32'hba4f2b13),
	.w2(32'hba2fab82),
	.w3(32'hb7c735c7),
	.w4(32'hba0bc879),
	.w5(32'hba1d692d),
	.w6(32'hba344cc3),
	.w7(32'hba3a9b3d),
	.w8(32'hba3d08ee),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41df4b),
	.w1(32'h39a92026),
	.w2(32'hba14ff73),
	.w3(32'hb9f26bec),
	.w4(32'h39a9be3f),
	.w5(32'hb848b7cb),
	.w6(32'hb7bd6898),
	.w7(32'hb9106d04),
	.w8(32'h38a3d56b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977423e),
	.w1(32'h38a2720b),
	.w2(32'h39de6883),
	.w3(32'h39032a6e),
	.w4(32'hb9166874),
	.w5(32'h3908aaca),
	.w6(32'hb563a1e7),
	.w7(32'h382b9019),
	.w8(32'hb85d2f55),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368f172d),
	.w1(32'hba1e3c4b),
	.w2(32'hba079bc9),
	.w3(32'h3872eae0),
	.w4(32'hb9f199a6),
	.w5(32'hba0da82c),
	.w6(32'hba0fb118),
	.w7(32'hba26c34d),
	.w8(32'hba30c6c5),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c05b2),
	.w1(32'hba2cb16c),
	.w2(32'hb9f23c72),
	.w3(32'hb9fdc43e),
	.w4(32'hba1b66a9),
	.w5(32'hba0d78b6),
	.w6(32'hba10a19e),
	.w7(32'hba028445),
	.w8(32'hba09ea31),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25adae),
	.w1(32'hb9c935f4),
	.w2(32'hb8b82e30),
	.w3(32'hba055dea),
	.w4(32'hb90f6027),
	.w5(32'h38a9d813),
	.w6(32'hb9b762e6),
	.w7(32'hb99571e8),
	.w8(32'hb9c418e0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d82763),
	.w1(32'h395b614f),
	.w2(32'h39a9b08a),
	.w3(32'hb8d76d84),
	.w4(32'h375f05d2),
	.w5(32'h3994ac6a),
	.w6(32'h392f34ae),
	.w7(32'h39bfa53a),
	.w8(32'hb899c233),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb909cf3f),
	.w1(32'hba43e10e),
	.w2(32'hba1204f3),
	.w3(32'h3986b8ed),
	.w4(32'hba4dda37),
	.w5(32'hb9f45d47),
	.w6(32'hba6d4de9),
	.w7(32'hbac73255),
	.w8(32'hbb10ee95),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a49b15),
	.w1(32'hb9e7cbdd),
	.w2(32'hb9b900d2),
	.w3(32'hba64967b),
	.w4(32'hb7d2b629),
	.w5(32'hb74bf5aa),
	.w6(32'hb966992b),
	.w7(32'hb8c036b8),
	.w8(32'h3681acfc),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9009d86),
	.w1(32'hb9dc77fa),
	.w2(32'h374a708e),
	.w3(32'h396e9305),
	.w4(32'hba05cf34),
	.w5(32'hb9a7c7a6),
	.w6(32'hb9687414),
	.w7(32'hb8f4135f),
	.w8(32'hb994168a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d99a59),
	.w1(32'hb9717025),
	.w2(32'h39b0a12c),
	.w3(32'hb9652cb5),
	.w4(32'hb9bddf98),
	.w5(32'h390e7dc8),
	.w6(32'hb6c0603b),
	.w7(32'h39a1c8be),
	.w8(32'h37613bbe),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984bcf7),
	.w1(32'hb986fab9),
	.w2(32'hb814f208),
	.w3(32'hb9f7fd77),
	.w4(32'h37f69239),
	.w5(32'h395d8c06),
	.w6(32'hb88fb62c),
	.w7(32'h38d22924),
	.w8(32'h395c4815),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67ad78f),
	.w1(32'h3a01f261),
	.w2(32'h39f171e2),
	.w3(32'h392b6f0e),
	.w4(32'h396fb7e1),
	.w5(32'h39c49bbe),
	.w6(32'h3a2e9e93),
	.w7(32'h3a33c7de),
	.w8(32'h399607da),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908f5ca),
	.w1(32'h39e236d6),
	.w2(32'h381a186c),
	.w3(32'h390fde0f),
	.w4(32'h39978cad),
	.w5(32'h3912cd46),
	.w6(32'h3a396271),
	.w7(32'h3a009868),
	.w8(32'h39a834df),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9338718),
	.w1(32'h39aec84d),
	.w2(32'h39943812),
	.w3(32'h34d91522),
	.w4(32'h390094d4),
	.w5(32'h39a16651),
	.w6(32'h39d31d81),
	.w7(32'h38bf30e5),
	.w8(32'h3816ca1f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8077f0c),
	.w1(32'h38b79e9a),
	.w2(32'h39866aab),
	.w3(32'h39a7fae2),
	.w4(32'hb89046ea),
	.w5(32'h392dec4f),
	.w6(32'h393dc4ca),
	.w7(32'h39bd5e63),
	.w8(32'h381ac493),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb814fce8),
	.w1(32'h394ce7f2),
	.w2(32'h39fe1f55),
	.w3(32'h37db0044),
	.w4(32'hb8982c12),
	.w5(32'h3a140929),
	.w6(32'hb95c6a7b),
	.w7(32'h399736b7),
	.w8(32'hb73cc1b7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39510e20),
	.w1(32'h3a1cfb3a),
	.w2(32'h39eea1bb),
	.w3(32'h38805380),
	.w4(32'h3a3371bc),
	.w5(32'h3a037050),
	.w6(32'h3a23f482),
	.w7(32'h39ed5a3f),
	.w8(32'hb7330bec),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396cc55d),
	.w1(32'hb99f399b),
	.w2(32'h38002976),
	.w3(32'h39a7b364),
	.w4(32'hb9d20e72),
	.w5(32'hb92decdc),
	.w6(32'hb9d72481),
	.w7(32'hb9d62e86),
	.w8(32'hba25f9f1),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef771c),
	.w1(32'hb8e93c92),
	.w2(32'hb829dfc7),
	.w3(32'hba0e4fac),
	.w4(32'h38d3b35a),
	.w5(32'h39636051),
	.w6(32'hb80895e0),
	.w7(32'h36b8de52),
	.w8(32'h38b0541c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ba619e),
	.w1(32'h3910fbb0),
	.w2(32'h3a0f4ae2),
	.w3(32'h391b5949),
	.w4(32'h38bd4981),
	.w5(32'h39886c0b),
	.w6(32'h39d845c9),
	.w7(32'h3a18b0ca),
	.w8(32'h39abf36b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a74ad),
	.w1(32'hba03a4c9),
	.w2(32'hb9727381),
	.w3(32'h387df963),
	.w4(32'hb95bacdc),
	.w5(32'h379581e0),
	.w6(32'hb9892d27),
	.w7(32'hb8fd8b8f),
	.w8(32'hb88a1fe7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d046a),
	.w1(32'hb99507ab),
	.w2(32'hb95878aa),
	.w3(32'hb8e792d7),
	.w4(32'hb911395f),
	.w5(32'h38a88941),
	.w6(32'hb9aae85f),
	.w7(32'hb98d5aa0),
	.w8(32'hb8c12884),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9835697),
	.w1(32'h39ef1ad4),
	.w2(32'h3a35714f),
	.w3(32'hb8be3560),
	.w4(32'h39b69bba),
	.w5(32'h3a110e56),
	.w6(32'h39d814e4),
	.w7(32'h39fcc505),
	.w8(32'h3a00fb36),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a05f4),
	.w1(32'h3a054d57),
	.w2(32'h3a1d89cb),
	.w3(32'h3a15ee25),
	.w4(32'h39eba53e),
	.w5(32'h3a1e6cf1),
	.w6(32'h3a33544d),
	.w7(32'h3a5af658),
	.w8(32'h3a512323),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44fac6),
	.w1(32'h3a19bfe6),
	.w2(32'h3a38c7c3),
	.w3(32'h3a5468b4),
	.w4(32'h39c781bd),
	.w5(32'h3a2c6c9e),
	.w6(32'h3a814f22),
	.w7(32'h3a9346f7),
	.w8(32'h3a05d2c6),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b724b),
	.w1(32'hb7c05ff0),
	.w2(32'h38ff4601),
	.w3(32'h390954ad),
	.w4(32'hb94edb4c),
	.w5(32'hb9270bdd),
	.w6(32'hb895a134),
	.w7(32'hb88d80e2),
	.w8(32'hb9401828),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c04f7),
	.w1(32'hb6de3d9a),
	.w2(32'hb783c084),
	.w3(32'hb94dd5ff),
	.w4(32'hb947fbea),
	.w5(32'hb970d0ce),
	.w6(32'h379c09d9),
	.w7(32'hb8e8e2f5),
	.w8(32'hb68b7572),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915414e),
	.w1(32'h38d5f50e),
	.w2(32'h3a4d1d8b),
	.w3(32'hb9d140b9),
	.w4(32'hb9c1d7fd),
	.w5(32'h39f7a1ac),
	.w6(32'hb9498953),
	.w7(32'h3a43b52e),
	.w8(32'hb97da06e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca0baf),
	.w1(32'hb9e09d1e),
	.w2(32'hba39447b),
	.w3(32'hba1302ec),
	.w4(32'hb9fa63c7),
	.w5(32'hba089600),
	.w6(32'hb9e98112),
	.w7(32'hb96fd3b8),
	.w8(32'hb96e79a5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15bfee),
	.w1(32'h384948d6),
	.w2(32'h385af997),
	.w3(32'hb9a18ffc),
	.w4(32'hb95fb7a5),
	.w5(32'hb92b113b),
	.w6(32'h39484b78),
	.w7(32'h394d7629),
	.w8(32'h38d316e4),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd3700),
	.w1(32'h3a29e091),
	.w2(32'h39ceca36),
	.w3(32'hb9c6d3c7),
	.w4(32'h3a4037e4),
	.w5(32'h3a4a8f11),
	.w6(32'h3a54776f),
	.w7(32'h3a62f2cb),
	.w8(32'h3a5eafad),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fba3f9),
	.w1(32'h39fd0af9),
	.w2(32'hba729bff),
	.w3(32'h3a3e2ef4),
	.w4(32'hb8fc13e0),
	.w5(32'hbad083e7),
	.w6(32'hb911f687),
	.w7(32'hb90c38ac),
	.w8(32'hbaa3067e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35eb5a),
	.w1(32'h39a1eea1),
	.w2(32'hba88d6da),
	.w3(32'hba8b8b67),
	.w4(32'h3706113a),
	.w5(32'hba1f3046),
	.w6(32'h3995894d),
	.w7(32'hba562420),
	.w8(32'hbab9a4b6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c5b86),
	.w1(32'hba2f11e1),
	.w2(32'hb9d70b97),
	.w3(32'hb8eea0c6),
	.w4(32'hb909d7b3),
	.w5(32'h38b048ab),
	.w6(32'hb9dd5e0f),
	.w7(32'hb97ea9fb),
	.w8(32'h38a238b4),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ce2d9),
	.w1(32'hba0419af),
	.w2(32'hb9cfc068),
	.w3(32'h39af6646),
	.w4(32'hb98d05d9),
	.w5(32'hb9ec12f1),
	.w6(32'hb9caced4),
	.w7(32'hb9e7b11e),
	.w8(32'hba10b7c0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0552bd),
	.w1(32'hb9a6fb79),
	.w2(32'hb9488d78),
	.w3(32'hb9e2272c),
	.w4(32'hb86ba03a),
	.w5(32'h3681ba84),
	.w6(32'hb92f47a8),
	.w7(32'hb88c5b1e),
	.w8(32'h3865c430),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f0a04d),
	.w1(32'hba10006e),
	.w2(32'hb97ad542),
	.w3(32'h3919e5d7),
	.w4(32'hba090f5f),
	.w5(32'hb98c9f4a),
	.w6(32'hba06e948),
	.w7(32'hb9b8ae3b),
	.w8(32'hb954ff8b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f40952),
	.w1(32'hb956d9ca),
	.w2(32'hb667be26),
	.w3(32'hb97b10b1),
	.w4(32'hb9c32623),
	.w5(32'hb9aafebd),
	.w6(32'h38bba1d0),
	.w7(32'hb7ee3c18),
	.w8(32'hb9d3736f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04ee0f),
	.w1(32'h38d322a5),
	.w2(32'h3987081e),
	.w3(32'hb9d2c402),
	.w4(32'h39bac103),
	.w5(32'h3a24652c),
	.w6(32'h395c94ce),
	.w7(32'h398f0230),
	.w8(32'h39bc174c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921aa95),
	.w1(32'hb995e9b2),
	.w2(32'hb948bc1c),
	.w3(32'h39cf1270),
	.w4(32'hb6ef7250),
	.w5(32'h383f6f19),
	.w6(32'hb900abd2),
	.w7(32'hb85dd60c),
	.w8(32'h384e359c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d05d7d),
	.w1(32'hb9e8ad41),
	.w2(32'hb9021084),
	.w3(32'h39488be5),
	.w4(32'hb9c14266),
	.w5(32'hb9bd9bce),
	.w6(32'hb98f6237),
	.w7(32'hb9a6a7cc),
	.w8(32'hba2a0b39),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43f903),
	.w1(32'hba84da0f),
	.w2(32'hba71b69f),
	.w3(32'hba172c26),
	.w4(32'hba897f4e),
	.w5(32'hba4fbafb),
	.w6(32'hba5cb76b),
	.w7(32'hba40fd39),
	.w8(32'hba506800),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97667d),
	.w1(32'hbaa6c49a),
	.w2(32'hb9ed5811),
	.w3(32'hba3cddaa),
	.w4(32'hbae00d72),
	.w5(32'hba924806),
	.w6(32'hb9e95172),
	.w7(32'h394156bc),
	.w8(32'hb9c7504d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba130e21),
	.w1(32'hba5dddf7),
	.w2(32'hba4a9d4a),
	.w3(32'hba062a69),
	.w4(32'hba4498cf),
	.w5(32'hba45131e),
	.w6(32'hba4d73d6),
	.w7(32'hba4e34fe),
	.w8(32'hba4bece3),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba890a86),
	.w1(32'h39c4ef3d),
	.w2(32'h39c67127),
	.w3(32'hba302f25),
	.w4(32'h393bdb5d),
	.w5(32'h3904aae3),
	.w6(32'hb8f3d03b),
	.w7(32'hb910bd50),
	.w8(32'hb9df9964),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a517b),
	.w1(32'hba8cbb5d),
	.w2(32'hba149ce9),
	.w3(32'hb95a71c7),
	.w4(32'hba2e75f7),
	.w5(32'hb974cb8f),
	.w6(32'hba49ca5b),
	.w7(32'hba259dbe),
	.w8(32'hb99abcbd),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9774fc4),
	.w1(32'hb9e99190),
	.w2(32'hb9912ad4),
	.w3(32'h38f86e1f),
	.w4(32'hb84c9236),
	.w5(32'h38378177),
	.w6(32'hb969424e),
	.w7(32'hb8b41973),
	.w8(32'h38b28a6e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e87e1),
	.w1(32'hb9292cd2),
	.w2(32'hb8975b79),
	.w3(32'h398be1c0),
	.w4(32'hb8832afb),
	.w5(32'hb87aaee0),
	.w6(32'hb935447e),
	.w7(32'hb8d7fa55),
	.w8(32'hb9192208),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9714209),
	.w1(32'hb97243a8),
	.w2(32'hb93ec804),
	.w3(32'hb87c4c94),
	.w4(32'hb8a498f2),
	.w5(32'hb8c7ec4b),
	.w6(32'hb9627ffb),
	.w7(32'hb9062bc6),
	.w8(32'hb8820881),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9888d2b),
	.w1(32'hbaaabe22),
	.w2(32'hba37bd46),
	.w3(32'hb5b16216),
	.w4(32'hba4e6e9e),
	.w5(32'hba375052),
	.w6(32'hba317e8e),
	.w7(32'hb9955f8a),
	.w8(32'hb9ac21da),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc8cc5),
	.w1(32'hba32020f),
	.w2(32'hb9d17c42),
	.w3(32'hb98c0b84),
	.w4(32'hba864ac8),
	.w5(32'hba339e55),
	.w6(32'hba6ae204),
	.w7(32'hba0a6dd8),
	.w8(32'hba563b8c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55be9b),
	.w1(32'hb99dcd06),
	.w2(32'hb9821db2),
	.w3(32'hba258026),
	.w4(32'hb7527867),
	.w5(32'hb9850322),
	.w6(32'hb8072a8c),
	.w7(32'hb807c901),
	.w8(32'h3796df15),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba072882),
	.w1(32'hb63dc5b6),
	.w2(32'hb9151854),
	.w3(32'hb8e9f021),
	.w4(32'hb94b6820),
	.w5(32'hb9313fb0),
	.w6(32'hb85788e8),
	.w7(32'hb6fac2d6),
	.w8(32'h396b8b19),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2db02),
	.w1(32'hba18bc49),
	.w2(32'hb9bedfda),
	.w3(32'hb8b3c977),
	.w4(32'hb9ffb503),
	.w5(32'hb9be2938),
	.w6(32'hba0a4a66),
	.w7(32'hb9d03940),
	.w8(32'hb9bb99b3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f260b9),
	.w1(32'hba4e814e),
	.w2(32'hba3d8aa5),
	.w3(32'hb9962ab0),
	.w4(32'hba6dccbc),
	.w5(32'hba9c1d39),
	.w6(32'h39435456),
	.w7(32'h38f730ba),
	.w8(32'hb9ca97ad),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1c229),
	.w1(32'hb8f75259),
	.w2(32'hb6d2e77b),
	.w3(32'hba5e9fad),
	.w4(32'hb887bd56),
	.w5(32'hb95f9104),
	.w6(32'hb9022828),
	.w7(32'hb90948e1),
	.w8(32'h392f2580),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe3281),
	.w1(32'hb927d3d9),
	.w2(32'h37d7dd6f),
	.w3(32'hb93795d9),
	.w4(32'h391bed50),
	.w5(32'h39b3d24f),
	.w6(32'h36d1b4fa),
	.w7(32'h38c64e4e),
	.w8(32'h39543d76),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8952fa4),
	.w1(32'hb94d5313),
	.w2(32'hba2cc283),
	.w3(32'h397353c7),
	.w4(32'h39392810),
	.w5(32'h398c84be),
	.w6(32'hb996c51f),
	.w7(32'hbaacd838),
	.w8(32'hba081e20),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396592cd),
	.w1(32'hbab3661a),
	.w2(32'hbae883a7),
	.w3(32'h39acb398),
	.w4(32'hba08d8a9),
	.w5(32'hbaa9b9b9),
	.w6(32'hba8a4c6c),
	.w7(32'hbac9488f),
	.w8(32'hba6f818d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule