module layer_8_featuremap_44(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf91bba),
	.w1(32'hbb35bf6d),
	.w2(32'hbaaa43f3),
	.w3(32'hbb2afdce),
	.w4(32'hbb68b8bb),
	.w5(32'hbac43671),
	.w6(32'hbb21a752),
	.w7(32'hbacecf9e),
	.w8(32'h38e24e0f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdbc1d),
	.w1(32'hba9c6926),
	.w2(32'hba730c51),
	.w3(32'hbad45019),
	.w4(32'hba60e216),
	.w5(32'hb97a8ccc),
	.w6(32'h368e5aee),
	.w7(32'h39706d67),
	.w8(32'h3a4c5530),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb807f1a),
	.w1(32'hb9cc994e),
	.w2(32'h3a8d0418),
	.w3(32'hbb964b99),
	.w4(32'hbab8fa3d),
	.w5(32'h3a048928),
	.w6(32'hbbc8be40),
	.w7(32'hbb82ca2d),
	.w8(32'hbad7e33d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb522def),
	.w1(32'hbae3576d),
	.w2(32'hbb0548e9),
	.w3(32'hbb586161),
	.w4(32'hbb26ad24),
	.w5(32'hbaac1bf5),
	.w6(32'hbb299479),
	.w7(32'hbaacc0ff),
	.w8(32'hbaecd7c0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cf48a),
	.w1(32'hbbb1d644),
	.w2(32'hbb1cd685),
	.w3(32'hbb640b97),
	.w4(32'hbb73bb95),
	.w5(32'hbae8c301),
	.w6(32'hbaf02cbd),
	.w7(32'hbac0f144),
	.w8(32'h3944c010),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2824c8),
	.w1(32'h3ba0433f),
	.w2(32'h3abe6b41),
	.w3(32'h3a7f980a),
	.w4(32'h3b40907a),
	.w5(32'h387120b7),
	.w6(32'hba9d131a),
	.w7(32'h3ab33154),
	.w8(32'hba900977),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9ad40),
	.w1(32'hb9a4cd86),
	.w2(32'hb9a49c2c),
	.w3(32'hb9008b5b),
	.w4(32'hb9680279),
	.w5(32'h38571bf3),
	.w6(32'h390f0ec7),
	.w7(32'h37c54ce3),
	.w8(32'h38664607),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5de23),
	.w1(32'hbb7d895a),
	.w2(32'hb8be5f2e),
	.w3(32'hbbcd542c),
	.w4(32'hbb99119e),
	.w5(32'hba5868af),
	.w6(32'hbb673313),
	.w7(32'hba52cd01),
	.w8(32'h3b25aaf8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd30229),
	.w1(32'hbb91d5a6),
	.w2(32'hba5dc2cd),
	.w3(32'hbbcd2f53),
	.w4(32'hbbbf9e0d),
	.w5(32'hb9fde88e),
	.w6(32'hbb6e0fd0),
	.w7(32'hba963c9b),
	.w8(32'h3b0de730),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc3f3d),
	.w1(32'hbab44c68),
	.w2(32'h3a946acc),
	.w3(32'hbb7126a2),
	.w4(32'hbb07d02a),
	.w5(32'h3a313188),
	.w6(32'hbb11a7a6),
	.w7(32'hb9aaf810),
	.w8(32'h3b07c18c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba27de9),
	.w1(32'hbbec9406),
	.w2(32'hbb8c5ead),
	.w3(32'hbb923446),
	.w4(32'hbbbfa71a),
	.w5(32'hbb7d0092),
	.w6(32'hbb819653),
	.w7(32'hbb4310a8),
	.w8(32'hbb0eb503),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb118fcd),
	.w1(32'hbaf29103),
	.w2(32'hbacceea2),
	.w3(32'hbb7180a7),
	.w4(32'hbb077ba3),
	.w5(32'hbae3ce63),
	.w6(32'hbb62d97a),
	.w7(32'hbb09f9b2),
	.w8(32'hbae72bea),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade8a2e),
	.w1(32'h3aafee7e),
	.w2(32'h3afbbc37),
	.w3(32'hbb89777f),
	.w4(32'hba91075c),
	.w5(32'h3a74358c),
	.w6(32'hba6e0dc8),
	.w7(32'h3aafd849),
	.w8(32'h3b2c8b6a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8faefed),
	.w1(32'h3587970f),
	.w2(32'h388c4983),
	.w3(32'h38392b0f),
	.w4(32'h3989cab4),
	.w5(32'hb66db263),
	.w6(32'h38814ec8),
	.w7(32'hb897d110),
	.w8(32'hb8582f34),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e79c5e),
	.w1(32'hb90bc79f),
	.w2(32'hb912e449),
	.w3(32'hb911d3e2),
	.w4(32'hb8f80e59),
	.w5(32'hb90e28c5),
	.w6(32'hb8fa3472),
	.w7(32'hb9035e83),
	.w8(32'hb91d99b9),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a7938),
	.w1(32'hba3e4058),
	.w2(32'hb98075be),
	.w3(32'hbacd18e3),
	.w4(32'hbab19653),
	.w5(32'hb9df012b),
	.w6(32'hbaaf8edd),
	.w7(32'hbab8f759),
	.w8(32'hba9c3ef0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39245136),
	.w1(32'hba344469),
	.w2(32'h3a2034eb),
	.w3(32'hbaaed67a),
	.w4(32'hba2398ed),
	.w5(32'h38a8fa2e),
	.w6(32'hbadbaaef),
	.w7(32'hba93f6e0),
	.w8(32'hb92a68a4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb59ae1),
	.w1(32'hbb15f6ba),
	.w2(32'hba3142e7),
	.w3(32'hbc0e9238),
	.w4(32'hbbd0bf4c),
	.w5(32'hbb3bf481),
	.w6(32'hbbea2a72),
	.w7(32'hbba30068),
	.w8(32'hbb4116f5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95bdd4),
	.w1(32'hbc77990f),
	.w2(32'hbade8503),
	.w3(32'hbc5af8af),
	.w4(32'hbc45a5fe),
	.w5(32'hba9f8ee4),
	.w6(32'hbc6241b1),
	.w7(32'hbc17b849),
	.w8(32'h3ac540ed),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14d567),
	.w1(32'hbbefc18a),
	.w2(32'hbbac6a92),
	.w3(32'hbc3741be),
	.w4(32'hbc038f08),
	.w5(32'hbb97afa9),
	.w6(32'hbbd414a9),
	.w7(32'hbbb27ee1),
	.w8(32'hbaf0a0ce),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26ce5f),
	.w1(32'h3a1aaba2),
	.w2(32'hbb0d388b),
	.w3(32'hba59e461),
	.w4(32'hb9cb721a),
	.w5(32'hbb4737df),
	.w6(32'hb9992e05),
	.w7(32'hb9514feb),
	.w8(32'h3838a853),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41685a),
	.w1(32'h3b8f7e1d),
	.w2(32'hb83e75e9),
	.w3(32'hbb0be0a2),
	.w4(32'h3b9812c5),
	.w5(32'h3b4c5f21),
	.w6(32'h3b763f38),
	.w7(32'h3bc88699),
	.w8(32'h3b4feed2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2aca9e),
	.w1(32'hbc78731f),
	.w2(32'hbae7a913),
	.w3(32'hbc2b3e22),
	.w4(32'hbc63b7fd),
	.w5(32'h3a684327),
	.w6(32'hbbcaaabb),
	.w7(32'hbbbc7595),
	.w8(32'h3bc2d23d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fbb175),
	.w1(32'h383bda2c),
	.w2(32'hb926c511),
	.w3(32'hbac689ba),
	.w4(32'hbb0466c9),
	.w5(32'hbabff931),
	.w6(32'hbac1d5d4),
	.w7(32'hbb3d0411),
	.w8(32'hbb2e98a3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0158fa),
	.w1(32'h3a2b9bc2),
	.w2(32'hb898d222),
	.w3(32'h394293e8),
	.w4(32'hbaa7cff8),
	.w5(32'hb9fb156b),
	.w6(32'h3ab4e80f),
	.w7(32'h3b0dff2d),
	.w8(32'h3b210b12),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dd9cf),
	.w1(32'hbbf2912b),
	.w2(32'hbb88532f),
	.w3(32'hbb50f568),
	.w4(32'hbb9d89bf),
	.w5(32'hbb202180),
	.w6(32'hbafc39e0),
	.w7(32'hbb70a0f0),
	.w8(32'hbab77bd8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4e3d1),
	.w1(32'h3a97f9d3),
	.w2(32'h3a9e557f),
	.w3(32'h3ad481f4),
	.w4(32'h3aa6c8a2),
	.w5(32'h3a9a3677),
	.w6(32'h3aa78b9a),
	.w7(32'h3a87e142),
	.w8(32'h3a8504fa),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcea30f0),
	.w1(32'hbcce44c1),
	.w2(32'hbbd7d776),
	.w3(32'hbcd071a1),
	.w4(32'hbc814ff7),
	.w5(32'h39a60c1f),
	.w6(32'hbc1be452),
	.w7(32'hbbb46941),
	.w8(32'h3c77b844),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f5c8d),
	.w1(32'hbb71c103),
	.w2(32'hbadada68),
	.w3(32'hbb895225),
	.w4(32'hbb7ec946),
	.w5(32'hbad2e5fd),
	.w6(32'hbabd9d10),
	.w7(32'hb9eb3b66),
	.w8(32'h3a96b2c2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb037fe7),
	.w1(32'hba1372bd),
	.w2(32'hb98b9362),
	.w3(32'hbacbd864),
	.w4(32'hba2f5928),
	.w5(32'hb9c1deba),
	.w6(32'hbac00473),
	.w7(32'hba541d55),
	.w8(32'hba7ab7dd),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39e22b),
	.w1(32'h3b844a42),
	.w2(32'h3a9d7891),
	.w3(32'h3b7ba049),
	.w4(32'h3b9c14fb),
	.w5(32'h3aeb221f),
	.w6(32'h3b7af917),
	.w7(32'h3b8d71f2),
	.w8(32'h3b2fc9bc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97b5b0),
	.w1(32'hba84de8d),
	.w2(32'hbb01bc5b),
	.w3(32'hbaa5dafc),
	.w4(32'hba4e3c41),
	.w5(32'hba8d9e8d),
	.w6(32'h3aa3693c),
	.w7(32'h3af0148f),
	.w8(32'h3adbf1c1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9706e82),
	.w1(32'hb9bb532e),
	.w2(32'hb98d04d8),
	.w3(32'hb907a836),
	.w4(32'hb9581cc8),
	.w5(32'hb964b0d7),
	.w6(32'hb8f37b3d),
	.w7(32'hb938a814),
	.w8(32'hb9368dd8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dd80b0),
	.w1(32'hb89432cf),
	.w2(32'hb89e9858),
	.w3(32'h3802cef6),
	.w4(32'hb83faa4f),
	.w5(32'hb8132d9f),
	.w6(32'h38b07c5b),
	.w7(32'h33585c20),
	.w8(32'h378bf198),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc1d96),
	.w1(32'h3b739513),
	.w2(32'h3b27f850),
	.w3(32'hba8bed10),
	.w4(32'h3a584319),
	.w5(32'hba472b66),
	.w6(32'hba128404),
	.w7(32'h393d741d),
	.w8(32'hbabb7c02),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16a321),
	.w1(32'hbbb374e2),
	.w2(32'hbb07aaab),
	.w3(32'hbae2cd8b),
	.w4(32'hbb48fefc),
	.w5(32'hbb21bbee),
	.w6(32'hbaec7766),
	.w7(32'hbb1fff39),
	.w8(32'hba9db995),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af1f26),
	.w1(32'hb9131c55),
	.w2(32'h39da0de7),
	.w3(32'hb9db922e),
	.w4(32'hb93b0a06),
	.w5(32'h399382c8),
	.w6(32'hba1530ee),
	.w7(32'hba031931),
	.w8(32'hb919fd60),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb851367),
	.w1(32'hbae0ebc7),
	.w2(32'hbaae2f2c),
	.w3(32'hbafeafe7),
	.w4(32'hb9b2b338),
	.w5(32'h39d34de9),
	.w6(32'h3a22c5ec),
	.w7(32'h3b1b1435),
	.w8(32'h3b177ef8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39993cba),
	.w1(32'hb8536681),
	.w2(32'hb869c29b),
	.w3(32'h38b4f5dd),
	.w4(32'hb80818e6),
	.w5(32'hb88f9630),
	.w6(32'hb9674691),
	.w7(32'hb9a7639d),
	.w8(32'hba07c56a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ebe24),
	.w1(32'h3a31251d),
	.w2(32'h3a38c82e),
	.w3(32'h3a7a55f7),
	.w4(32'h3a5cefda),
	.w5(32'h3a874619),
	.w6(32'h3ab62df5),
	.w7(32'h3aad689f),
	.w8(32'h3ac22a03),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4d769),
	.w1(32'hbaa3a1bf),
	.w2(32'hbb0a06bd),
	.w3(32'hbc57136b),
	.w4(32'hbbf9589e),
	.w5(32'hbc0ae99b),
	.w6(32'hbc309b44),
	.w7(32'hbbac5a5d),
	.w8(32'hbbf547fb),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebcfff),
	.w1(32'hba9b7604),
	.w2(32'h3b44256a),
	.w3(32'hbb4a216a),
	.w4(32'hbb199f6c),
	.w5(32'h3a855b4d),
	.w6(32'hbb1a4480),
	.w7(32'h3942c385),
	.w8(32'hbb2b138d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa5d72),
	.w1(32'hb9e19145),
	.w2(32'h3a749e61),
	.w3(32'hbbab2c33),
	.w4(32'h3a66a6b5),
	.w5(32'h3a291d58),
	.w6(32'h3b80810e),
	.w7(32'hb9114b21),
	.w8(32'h395a9337),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d79c0),
	.w1(32'hbb201558),
	.w2(32'hbaf78922),
	.w3(32'hbb84730b),
	.w4(32'hbb49b2c1),
	.w5(32'hbb4c55fc),
	.w6(32'hbb7036be),
	.w7(32'hbb086068),
	.w8(32'hbb2d11dd),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b41f7),
	.w1(32'hbc0c8e93),
	.w2(32'hbb062a2e),
	.w3(32'hbc103be4),
	.w4(32'hbbf77b08),
	.w5(32'hbb396fae),
	.w6(32'hbbef88b5),
	.w7(32'hbb3c9baa),
	.w8(32'h3b5c33ed),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b041b0c),
	.w1(32'h3b5f0701),
	.w2(32'h3bd05f4c),
	.w3(32'h3b06ed2a),
	.w4(32'h3b75f436),
	.w5(32'h3bb90fec),
	.w6(32'hb81c7c1d),
	.w7(32'h3b81c82f),
	.w8(32'hba287eb2),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb023139),
	.w1(32'h3ae2ff84),
	.w2(32'hbb070e17),
	.w3(32'hbb33743a),
	.w4(32'h3b9f79d5),
	.w5(32'hba22bcd8),
	.w6(32'hbaef80e9),
	.w7(32'hbaa1dfe6),
	.w8(32'h3a6a2710),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd96da6),
	.w1(32'hbbff99e0),
	.w2(32'hb7ca298f),
	.w3(32'hbbb0728a),
	.w4(32'hbb45ede6),
	.w5(32'h3b3f49db),
	.w6(32'hbbb678c6),
	.w7(32'hbb7d03ae),
	.w8(32'hba8f0bfd),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49065a),
	.w1(32'hb91af4b5),
	.w2(32'h3b1d8a32),
	.w3(32'hbb7bccd2),
	.w4(32'hbad00b0b),
	.w5(32'h39e57f75),
	.w6(32'hbb30d9cf),
	.w7(32'hb8ea1418),
	.w8(32'hba99983f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d4ed8),
	.w1(32'hbb9f3781),
	.w2(32'hba900694),
	.w3(32'hbbacb048),
	.w4(32'hbb9c62f2),
	.w5(32'hbae7deeb),
	.w6(32'hbb99fd38),
	.w7(32'hbb30b6db),
	.w8(32'hba9eea9f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b3d50),
	.w1(32'h3bf8cef5),
	.w2(32'h3b95bc78),
	.w3(32'h3a895983),
	.w4(32'h3c038567),
	.w5(32'h3bc23b44),
	.w6(32'h3bad9727),
	.w7(32'h3c3ef93e),
	.w8(32'h3c1b8a35),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82d88a),
	.w1(32'hbc777b35),
	.w2(32'hbc062ef0),
	.w3(32'hbca19faa),
	.w4(32'hbc9df441),
	.w5(32'hbc35f123),
	.w6(32'hbc76d09f),
	.w7(32'hbc457dd1),
	.w8(32'hbbbe7a60),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00ec65),
	.w1(32'hbbbae059),
	.w2(32'hbb274c46),
	.w3(32'hbb815a14),
	.w4(32'hbbad6b2d),
	.w5(32'h3a262798),
	.w6(32'hbb25c8c7),
	.w7(32'hbb8eb4cd),
	.w8(32'hb771b566),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba696ea),
	.w1(32'hbbacf00f),
	.w2(32'hbb525ed6),
	.w3(32'hbbfcd2e8),
	.w4(32'hbbfc9321),
	.w5(32'hbbb53b77),
	.w6(32'hbc10cd53),
	.w7(32'hbbb285ec),
	.w8(32'h3b11a387),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51042e),
	.w1(32'hbae06c88),
	.w2(32'hbb8875d2),
	.w3(32'h3ae7b819),
	.w4(32'h3b1dc3ee),
	.w5(32'hba15a33b),
	.w6(32'h394c8831),
	.w7(32'hbb90c0ea),
	.w8(32'hb9ae45dd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42b9f8),
	.w1(32'hbaf192e3),
	.w2(32'hbb190a35),
	.w3(32'hbb9f5538),
	.w4(32'hbbbf9760),
	.w5(32'hba31dc83),
	.w6(32'hbba0fd16),
	.w7(32'hba80139e),
	.w8(32'h39d32753),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b729a1),
	.w1(32'h3b665bd7),
	.w2(32'hba4dc5ed),
	.w3(32'hbb29e80d),
	.w4(32'hb9c13de1),
	.w5(32'hbacd42fc),
	.w6(32'h3a85a646),
	.w7(32'hba5d4aec),
	.w8(32'h3ad39727),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5d8c6),
	.w1(32'h3ad4778b),
	.w2(32'h3b501a77),
	.w3(32'hbb9b6e6b),
	.w4(32'hbb708c34),
	.w5(32'h398cfc0c),
	.w6(32'h39f48b8e),
	.w7(32'h391f9908),
	.w8(32'hba0e8eed),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b13f9),
	.w1(32'hbb5b2593),
	.w2(32'hb92924c6),
	.w3(32'hbba8978b),
	.w4(32'hbb4673c3),
	.w5(32'hba62536e),
	.w6(32'hbabf95ed),
	.w7(32'h3a0b9b9c),
	.w8(32'h3a975342),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba193753),
	.w1(32'hbb3881c2),
	.w2(32'h38b28e91),
	.w3(32'hba4e3b76),
	.w4(32'hbb13e7dd),
	.w5(32'hbaa88a59),
	.w6(32'hbb3979ed),
	.w7(32'hba81618d),
	.w8(32'hbbac02e2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2f4d2),
	.w1(32'h39ffebbc),
	.w2(32'hbb9ec640),
	.w3(32'hbb33e07d),
	.w4(32'hba9b1936),
	.w5(32'hbb68dda9),
	.w6(32'hbaa81066),
	.w7(32'hbbf0aaaa),
	.w8(32'h3a8060ea),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f9f52),
	.w1(32'h3b098719),
	.w2(32'h3b4b78b8),
	.w3(32'h3b30731b),
	.w4(32'h3b489941),
	.w5(32'h3b7f329a),
	.w6(32'hb99778b1),
	.w7(32'h3b059676),
	.w8(32'hbb418cb5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3e7bd),
	.w1(32'hbafd4659),
	.w2(32'hba9583dd),
	.w3(32'hbc1d514c),
	.w4(32'hbbc0dce5),
	.w5(32'hbb59b6cf),
	.w6(32'hbc0144d9),
	.w7(32'hbb269786),
	.w8(32'h3b1ea4b2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d36d2),
	.w1(32'h395e924b),
	.w2(32'hb7c5d4bc),
	.w3(32'hba8fb320),
	.w4(32'hba6758f1),
	.w5(32'hbb7f13f9),
	.w6(32'hba0cd054),
	.w7(32'hbb8c0c46),
	.w8(32'hbb73e5d0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7564cb),
	.w1(32'h3a283c37),
	.w2(32'h3a4be0e7),
	.w3(32'h3a1a0101),
	.w4(32'hb97a0b23),
	.w5(32'hb89ca171),
	.w6(32'h3aae59cd),
	.w7(32'h3881a07c),
	.w8(32'h3a825005),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba852dcf),
	.w1(32'hba64d7f8),
	.w2(32'h3ac42dff),
	.w3(32'hbaf4d269),
	.w4(32'hba9dd841),
	.w5(32'h3a18d246),
	.w6(32'hbb0a9b24),
	.w7(32'hba0c42fb),
	.w8(32'h3a259134),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87bdaf),
	.w1(32'hbb5bad55),
	.w2(32'hbaaa0529),
	.w3(32'hbb8e01fe),
	.w4(32'hbb4bfc68),
	.w5(32'hbab313b8),
	.w6(32'hbb9ee975),
	.w7(32'hbb2ac7b6),
	.w8(32'h39b00f60),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6481cb),
	.w1(32'h3b785a06),
	.w2(32'h3b4f2249),
	.w3(32'hba27ea18),
	.w4(32'h3b894788),
	.w5(32'h3b84b8b1),
	.w6(32'hbb0716e4),
	.w7(32'h39e52ef4),
	.w8(32'h3aecd5c4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b673d),
	.w1(32'hbacd028f),
	.w2(32'hb9254362),
	.w3(32'hbb058be9),
	.w4(32'hbb0a1eaf),
	.w5(32'hb9dddcb5),
	.w6(32'hbb30385a),
	.w7(32'hbaaaa4ea),
	.w8(32'hbb3daae8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc064226),
	.w1(32'hbc504503),
	.w2(32'hbbdb7608),
	.w3(32'hbc2526b2),
	.w4(32'hbc28745f),
	.w5(32'hbbeecd05),
	.w6(32'hbc10fe09),
	.w7(32'hbbfd4ba6),
	.w8(32'hbb926775),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a099dc2),
	.w1(32'h38903cf4),
	.w2(32'h39c3826e),
	.w3(32'hb92e5816),
	.w4(32'hb9cc8c5f),
	.w5(32'hb892e039),
	.w6(32'hb9e41cd1),
	.w7(32'h3a073782),
	.w8(32'h38d364d0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba8e5b),
	.w1(32'hbbc55ca8),
	.w2(32'hbb208ee4),
	.w3(32'hbbf18dab),
	.w4(32'hbbe1f101),
	.w5(32'hbb30e3d1),
	.w6(32'hbbbec651),
	.w7(32'hbb9d8e86),
	.w8(32'hbb217b6a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba681e9e),
	.w1(32'hbaa4a20c),
	.w2(32'h399083ef),
	.w3(32'hbad450ac),
	.w4(32'hbb06aefb),
	.w5(32'hba403d8f),
	.w6(32'hbb5f64a6),
	.w7(32'hba8931b5),
	.w8(32'h3ae87899),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b390d),
	.w1(32'hbb6fa3d3),
	.w2(32'hbb9c1a1f),
	.w3(32'hbbaedd73),
	.w4(32'hbb647582),
	.w5(32'h38ab22a6),
	.w6(32'hbb5e45f1),
	.w7(32'hba79dca5),
	.w8(32'h3a40632b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a330df3),
	.w1(32'hb9ff5149),
	.w2(32'h389f79ae),
	.w3(32'hb97aa145),
	.w4(32'hbaa16b88),
	.w5(32'hba4f8261),
	.w6(32'hba737c87),
	.w7(32'hb97fba00),
	.w8(32'hba260a0f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0df66d),
	.w1(32'hbb4039db),
	.w2(32'hba5eee1a),
	.w3(32'hbb07dbaa),
	.w4(32'hbb0c91ef),
	.w5(32'h38f7b1b8),
	.w6(32'hb951e368),
	.w7(32'h3a7f26cc),
	.w8(32'h3a849ff1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397313c2),
	.w1(32'hb89dd14e),
	.w2(32'h39f8362b),
	.w3(32'hba04d192),
	.w4(32'hba22a1ee),
	.w5(32'hb9403a17),
	.w6(32'hba989d81),
	.w7(32'hb900ce30),
	.w8(32'hbb798929),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24a01f),
	.w1(32'hbbffe814),
	.w2(32'hbb5913a9),
	.w3(32'hbc2e3df6),
	.w4(32'hbbea837a),
	.w5(32'hbb3b6918),
	.w6(32'hbb9ecba4),
	.w7(32'hbb23d8bd),
	.w8(32'hbb600148),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7a677),
	.w1(32'hba929a35),
	.w2(32'h3a842599),
	.w3(32'hbba70afa),
	.w4(32'hbaf88420),
	.w5(32'h3adf3890),
	.w6(32'hbadfad71),
	.w7(32'hba0278e4),
	.w8(32'h3a8926a0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5887a2),
	.w1(32'hba7cab4c),
	.w2(32'hbafa5243),
	.w3(32'hbac1bd2c),
	.w4(32'h390a7056),
	.w5(32'hba82dffc),
	.w6(32'h39802813),
	.w7(32'hba0d87e5),
	.w8(32'h3b4693e8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabab000),
	.w1(32'h3b3655d1),
	.w2(32'hba5cb776),
	.w3(32'hb9ca8e63),
	.w4(32'h3a584748),
	.w5(32'hbaa8af8a),
	.w6(32'h3b7905d0),
	.w7(32'h3b106821),
	.w8(32'h39c30ba7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb122cd3),
	.w1(32'hbb3db27e),
	.w2(32'hba97ed07),
	.w3(32'hbb98ab69),
	.w4(32'hbba953d3),
	.w5(32'hbb7e3ff6),
	.w6(32'hbb9d8902),
	.w7(32'hbb497176),
	.w8(32'hbb1b09e5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0be79),
	.w1(32'hbbe50fc3),
	.w2(32'hbb03a62b),
	.w3(32'hbbf535b4),
	.w4(32'hbbe55d75),
	.w5(32'hbb458dc1),
	.w6(32'hbbc9a310),
	.w7(32'hbb1993d3),
	.w8(32'hbb76e425),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc308a22),
	.w1(32'h3a9a0312),
	.w2(32'hbb98fbd5),
	.w3(32'hbc83aa0b),
	.w4(32'hbb6c9e28),
	.w5(32'hbc2d22b4),
	.w6(32'hbc7e2728),
	.w7(32'hbb940e53),
	.w8(32'hbc071513),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b0b79),
	.w1(32'hbc36ff58),
	.w2(32'h37faab43),
	.w3(32'hbc8320ad),
	.w4(32'hbc5eb207),
	.w5(32'hbadfed5e),
	.w6(32'hbc7ab136),
	.w7(32'hbbfef05f),
	.w8(32'h3a4b8d00),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d4288),
	.w1(32'hbbfeb856),
	.w2(32'hbbe5c486),
	.w3(32'hbbc52869),
	.w4(32'hbc47bbd3),
	.w5(32'hbc1c4667),
	.w6(32'hbbe8e8e1),
	.w7(32'hbbe54978),
	.w8(32'hbbeeda5b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c0aae),
	.w1(32'h3a321a0f),
	.w2(32'h3b136aa2),
	.w3(32'hb9f5b66f),
	.w4(32'h3941ad45),
	.w5(32'h3aa4c6c3),
	.w6(32'h3a340c3d),
	.w7(32'h3ac61784),
	.w8(32'hba86a95a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fef08a),
	.w1(32'hba731f28),
	.w2(32'hb90441f5),
	.w3(32'h38f6f4f7),
	.w4(32'h399ebe24),
	.w5(32'h3a538416),
	.w6(32'hbaa6a29d),
	.w7(32'hba619e27),
	.w8(32'h3a20a517),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c91ce),
	.w1(32'hbac4a088),
	.w2(32'h3ab231b7),
	.w3(32'h3a968018),
	.w4(32'h38af8d2e),
	.w5(32'h3ab79b1c),
	.w6(32'hb510caa1),
	.w7(32'h3a8fd2f0),
	.w8(32'hbb18b485),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ea1b3),
	.w1(32'hba007adc),
	.w2(32'h3a948067),
	.w3(32'h3a5a4b70),
	.w4(32'hbab74f57),
	.w5(32'hb957457e),
	.w6(32'h3b27e38d),
	.w7(32'h3aba28dc),
	.w8(32'hba8e33a7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14c9bd),
	.w1(32'h391912a6),
	.w2(32'h3a66a775),
	.w3(32'hbb7dad21),
	.w4(32'hbb2ace93),
	.w5(32'hbaab7fbb),
	.w6(32'hbaf98e09),
	.w7(32'h39caf5fc),
	.w8(32'hbb325cba),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba931e73),
	.w1(32'hbb4d7736),
	.w2(32'hbae1dc58),
	.w3(32'hbb158bb1),
	.w4(32'hbb752e8e),
	.w5(32'hbb76a26a),
	.w6(32'hbb49b59b),
	.w7(32'hba8bd569),
	.w8(32'hbacadcb0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d4752),
	.w1(32'h3b90bb6d),
	.w2(32'h3ad3b2bf),
	.w3(32'hbb63476a),
	.w4(32'h3b4569c5),
	.w5(32'hb9c22580),
	.w6(32'h3b7acc3c),
	.w7(32'hb9b9197e),
	.w8(32'h3b04a348),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6b7de),
	.w1(32'hbb954c7d),
	.w2(32'hba3e4b01),
	.w3(32'hbc12697b),
	.w4(32'hbbf90da5),
	.w5(32'hbb5f31b7),
	.w6(32'hbc033b44),
	.w7(32'hbbc1f1f8),
	.w8(32'hbb9eb008),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb92cbd),
	.w1(32'hba9616eb),
	.w2(32'hbb6de634),
	.w3(32'hba9079eb),
	.w4(32'h399f035b),
	.w5(32'hb8e8d3ed),
	.w6(32'hbaa629ab),
	.w7(32'hbb0a6a2d),
	.w8(32'hbb633949),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e58fed),
	.w1(32'h3a612f07),
	.w2(32'h3bb5aee4),
	.w3(32'h3aa7ec97),
	.w4(32'hba87ceee),
	.w5(32'h3adce1b4),
	.w6(32'hba312878),
	.w7(32'h3b8a6c9d),
	.w8(32'h3bc853c8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09add7),
	.w1(32'hbb60d7c9),
	.w2(32'hba84488c),
	.w3(32'hbc4e91bc),
	.w4(32'hbc1c1dc6),
	.w5(32'hbaa67aaf),
	.w6(32'hbb8616db),
	.w7(32'hbb81900c),
	.w8(32'hba87ff0c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc536c4),
	.w1(32'hbb5b5948),
	.w2(32'hbb82dbb5),
	.w3(32'hbb454396),
	.w4(32'hba649ff8),
	.w5(32'hbb7fc101),
	.w6(32'hbbe70f89),
	.w7(32'hbb923bfd),
	.w8(32'hbb47edbd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb714f59),
	.w1(32'hba2af11d),
	.w2(32'h3936062e),
	.w3(32'hbb8155f5),
	.w4(32'hb9baa07b),
	.w5(32'h3a9c42b5),
	.w6(32'h399221df),
	.w7(32'h3ab06aad),
	.w8(32'hba7f52d3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380c81e3),
	.w1(32'hbaad3722),
	.w2(32'hba618af5),
	.w3(32'hba034d6c),
	.w4(32'hba118f5b),
	.w5(32'hb9559e07),
	.w6(32'hbaa394fb),
	.w7(32'hba66737a),
	.w8(32'h3a8d5411),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05cfb7),
	.w1(32'hb91df261),
	.w2(32'hba5784f7),
	.w3(32'h3b1d63d4),
	.w4(32'h3a66afff),
	.w5(32'hbab798ab),
	.w6(32'h3ab1525a),
	.w7(32'hb9caf621),
	.w8(32'hba6025b2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20c634),
	.w1(32'hbb548503),
	.w2(32'hbb471939),
	.w3(32'hbae437ef),
	.w4(32'hbb30fd5d),
	.w5(32'hbb13f61c),
	.w6(32'h394c144c),
	.w7(32'h3a83dc2a),
	.w8(32'hba6bd097),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb73220),
	.w1(32'h399357e2),
	.w2(32'h38c04347),
	.w3(32'hbbe1a907),
	.w4(32'hba5d17d6),
	.w5(32'h3b422b8f),
	.w6(32'hba9b2df4),
	.w7(32'h3b010363),
	.w8(32'h3b27225e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a997d),
	.w1(32'hbab8a98a),
	.w2(32'h3b20df9e),
	.w3(32'hbbbe2a1e),
	.w4(32'hbb4d3afa),
	.w5(32'hba452d81),
	.w6(32'hbb8a5926),
	.w7(32'hba9564ed),
	.w8(32'hb9a43fb6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6eb67b3),
	.w1(32'h3aa3f146),
	.w2(32'h3a26c353),
	.w3(32'hba2fcc3d),
	.w4(32'h39a420d8),
	.w5(32'hb9850267),
	.w6(32'hb9a30326),
	.w7(32'h3a1ca16b),
	.w8(32'hbab86fb9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84a235),
	.w1(32'hbba64988),
	.w2(32'h3b603e77),
	.w3(32'hbc163127),
	.w4(32'hbc051381),
	.w5(32'hbac96a6a),
	.w6(32'hbc4d5e62),
	.w7(32'hbc0022fb),
	.w8(32'hbb0f23e6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba707fe0),
	.w1(32'hbbaf22a4),
	.w2(32'hbb3b3df0),
	.w3(32'h3a029586),
	.w4(32'hbb8550da),
	.w5(32'hbaa737d4),
	.w6(32'hbafe5c2b),
	.w7(32'hbab9072e),
	.w8(32'hba601519),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ea6d7),
	.w1(32'hbaac9032),
	.w2(32'h3a844d7a),
	.w3(32'hbb83c34d),
	.w4(32'hbb28bdf1),
	.w5(32'hba7c7884),
	.w6(32'hbb737467),
	.w7(32'hbacce3ee),
	.w8(32'hbaf1a6e4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad84531),
	.w1(32'h3a9cd0fe),
	.w2(32'hbac0a507),
	.w3(32'h3adc9205),
	.w4(32'h3abfddd9),
	.w5(32'hbab661f1),
	.w6(32'h3a744a2b),
	.w7(32'h3a12b098),
	.w8(32'hba5c8739),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a503a),
	.w1(32'hbbe56033),
	.w2(32'hbb0cc7c3),
	.w3(32'hbbdf5406),
	.w4(32'hbbb51882),
	.w5(32'hb9a1dd07),
	.w6(32'hbb70494a),
	.w7(32'hbb362a19),
	.w8(32'h3a593282),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb299423),
	.w1(32'h3a3b749b),
	.w2(32'h3b5b2de5),
	.w3(32'hbac6d38e),
	.w4(32'h3a547568),
	.w5(32'h3b032bff),
	.w6(32'hbaba0304),
	.w7(32'h3b35fd60),
	.w8(32'h3ae7301b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb961b51),
	.w1(32'h3a5c7ebc),
	.w2(32'h39bdbdc0),
	.w3(32'hbb97c448),
	.w4(32'h39e57d4b),
	.w5(32'h399029a9),
	.w6(32'hbb4f384b),
	.w7(32'h39ea6d01),
	.w8(32'h3b1aade6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedc53e),
	.w1(32'h3b50350e),
	.w2(32'h3b18a778),
	.w3(32'h3b1bf279),
	.w4(32'h3a7bf8a7),
	.w5(32'h3a415c43),
	.w6(32'h39dde79f),
	.w7(32'h3abc8e85),
	.w8(32'hbb262338),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8da0b),
	.w1(32'hba8c6688),
	.w2(32'hba9a5248),
	.w3(32'hb9cd519c),
	.w4(32'hba9a7b56),
	.w5(32'hbab53a8e),
	.w6(32'hba242911),
	.w7(32'hbabbbbaf),
	.w8(32'hba677261),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ef7d8),
	.w1(32'hbab64182),
	.w2(32'hba9c2ec4),
	.w3(32'hbaae73c7),
	.w4(32'hbb011186),
	.w5(32'hbaab43e5),
	.w6(32'hba86a1c4),
	.w7(32'hbaeb5d16),
	.w8(32'hbaf48db4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba077175),
	.w1(32'hb80b39f3),
	.w2(32'hb9987e52),
	.w3(32'hba104b7a),
	.w4(32'hb97bb0c3),
	.w5(32'hb96b53ed),
	.w6(32'h3a07a6fe),
	.w7(32'h3a704518),
	.w8(32'h3a53e6bf),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04021b),
	.w1(32'h3aa0ce17),
	.w2(32'h3a89b052),
	.w3(32'hba508573),
	.w4(32'h3a3c4d0e),
	.w5(32'h39f2c1ad),
	.w6(32'hb68d008c),
	.w7(32'h3a730b67),
	.w8(32'h3a33c08c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63bb92),
	.w1(32'hbb06724f),
	.w2(32'hb9e9185a),
	.w3(32'hbb8a4c5f),
	.w4(32'hbacce78d),
	.w5(32'hbaaf2c9d),
	.w6(32'hbb7e0c25),
	.w7(32'hba792609),
	.w8(32'h3890adab),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21c302),
	.w1(32'h39413bce),
	.w2(32'h3a835dff),
	.w3(32'hb8cf737f),
	.w4(32'hba08046b),
	.w5(32'h3a0715cf),
	.w6(32'hba0af956),
	.w7(32'h3a4d0078),
	.w8(32'h393f10ea),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f46363),
	.w1(32'hb822605c),
	.w2(32'hb9e51b29),
	.w3(32'hb95a5358),
	.w4(32'hb909ec5d),
	.w5(32'hb92f39db),
	.w6(32'hb8afb83e),
	.w7(32'hb9af9fbd),
	.w8(32'h3a88413a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b206ff9),
	.w1(32'h3aeb0059),
	.w2(32'h3b2f42b2),
	.w3(32'hbb5a6a73),
	.w4(32'hbb81afe2),
	.w5(32'hba676f5f),
	.w6(32'hba3ac865),
	.w7(32'h391b2bd9),
	.w8(32'h3ad47c47),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb784909),
	.w1(32'hbb91a273),
	.w2(32'hbb1c0714),
	.w3(32'hbaf5091b),
	.w4(32'hbb8b95dc),
	.w5(32'hbab1869b),
	.w6(32'hbae0377b),
	.w7(32'hbb28c2d0),
	.w8(32'hbadee0a9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba757f2d),
	.w1(32'hbace564d),
	.w2(32'hbacf6bf8),
	.w3(32'hba8cbe1a),
	.w4(32'hbac9c02e),
	.w5(32'hbabbf309),
	.w6(32'hba510e50),
	.w7(32'hba355e08),
	.w8(32'hb96b5d0d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9343b7),
	.w1(32'h3abaf40d),
	.w2(32'hb9e850ee),
	.w3(32'h3ad30be4),
	.w4(32'h3aef4e4f),
	.w5(32'hb93c46ee),
	.w6(32'h3a9355e7),
	.w7(32'h3b098efa),
	.w8(32'hba645ccd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85eec1),
	.w1(32'hbac52276),
	.w2(32'hba70ca10),
	.w3(32'hbb3e72ba),
	.w4(32'hba82e459),
	.w5(32'h3a7d3c0e),
	.w6(32'hbabb73d8),
	.w7(32'hba2dc77f),
	.w8(32'h3abd4b60),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2e565),
	.w1(32'h3aa16517),
	.w2(32'h3a04a742),
	.w3(32'hba33fdb2),
	.w4(32'hb8dbbfcb),
	.w5(32'h39c3acb5),
	.w6(32'h3ac834c1),
	.w7(32'h39d6f775),
	.w8(32'h3a6cbcfb),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31d0c1),
	.w1(32'hbaaf2ca6),
	.w2(32'hba9035ea),
	.w3(32'hbaceeff6),
	.w4(32'hba8ff0a1),
	.w5(32'hb939fa46),
	.w6(32'h38f81ba1),
	.w7(32'h3933d1d7),
	.w8(32'h3b0aa7fd),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5cb7d),
	.w1(32'hb70fd6bd),
	.w2(32'h3a8be5e8),
	.w3(32'h3932f90f),
	.w4(32'h3aa70005),
	.w5(32'h3a7844da),
	.w6(32'h3a076363),
	.w7(32'h3a5a8707),
	.w8(32'h3b0ef852),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule