module layer_8_featuremap_254(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d95e27),
	.w1(32'hb9e79fb6),
	.w2(32'hb8c06bfb),
	.w3(32'h3a35f696),
	.w4(32'hba0ad495),
	.w5(32'h39d15885),
	.w6(32'h39d70d2f),
	.w7(32'hb7afb662),
	.w8(32'hba095ad5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e7e49),
	.w1(32'h3938791c),
	.w2(32'h3874f66a),
	.w3(32'h39b74cbd),
	.w4(32'h38b7edf0),
	.w5(32'hb8b2794b),
	.w6(32'hb80554e7),
	.w7(32'h37bd4e8a),
	.w8(32'hb7a32159),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb839d3ec),
	.w1(32'h37c8cdff),
	.w2(32'hb7b8ad00),
	.w3(32'hb91c9f56),
	.w4(32'hb97d512d),
	.w5(32'hb9a3724c),
	.w6(32'hb9a8784d),
	.w7(32'hb9318501),
	.w8(32'hb98164c5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968f904),
	.w1(32'hb8848ecd),
	.w2(32'hb951dd7a),
	.w3(32'hba0b6212),
	.w4(32'hba13b606),
	.w5(32'hba0e0e87),
	.w6(32'h3936f9c9),
	.w7(32'hb9afc25a),
	.w8(32'hba0f536d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b71a6f),
	.w1(32'hb787735d),
	.w2(32'h38934125),
	.w3(32'h3a09a9ae),
	.w4(32'hb797e2c3),
	.w5(32'h3936a36f),
	.w6(32'hb86d6d94),
	.w7(32'hb7cf2a74),
	.w8(32'h36d68437),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e1afb),
	.w1(32'h3a21fca2),
	.w2(32'hb8d4c8bf),
	.w3(32'h3a336f93),
	.w4(32'hb8a49fee),
	.w5(32'hba7cb281),
	.w6(32'hb9bb344d),
	.w7(32'h38886649),
	.w8(32'h3731f988),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f44de),
	.w1(32'hb90ea3d5),
	.w2(32'h37ab76d5),
	.w3(32'hb9d23b17),
	.w4(32'h379bcea5),
	.w5(32'h394fce71),
	.w6(32'h35831e81),
	.w7(32'hb855cb95),
	.w8(32'hb7c05edc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb924196f),
	.w1(32'h3a5f9788),
	.w2(32'h3a99ca08),
	.w3(32'hb8b56ca4),
	.w4(32'h397df2a0),
	.w5(32'h3a17dbff),
	.w6(32'hb92e8ac5),
	.w7(32'hb7741d6a),
	.w8(32'hb88ff97e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396183ae),
	.w1(32'hb9a48a9e),
	.w2(32'h3963a9f1),
	.w3(32'h3894e2c3),
	.w4(32'h36a56346),
	.w5(32'h39c2da64),
	.w6(32'hb9a5af63),
	.w7(32'hb8d7f137),
	.w8(32'hb9371e91),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16b90e),
	.w1(32'h394bc930),
	.w2(32'h376b5de0),
	.w3(32'hb9297a33),
	.w4(32'hb91862dd),
	.w5(32'h3a3f352c),
	.w6(32'h3a3179a8),
	.w7(32'hb8f1a526),
	.w8(32'hb9b76af4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68064c),
	.w1(32'hba0bc038),
	.w2(32'hba1ac858),
	.w3(32'h3958740f),
	.w4(32'hb94e606d),
	.w5(32'hba1c7ad4),
	.w6(32'h3a31997e),
	.w7(32'h3a1756c2),
	.w8(32'h3a2d049d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b03463),
	.w1(32'h39400c0c),
	.w2(32'h3a0a7a59),
	.w3(32'h39172caf),
	.w4(32'hb9a857ee),
	.w5(32'hb85110ac),
	.w6(32'hb90c1c9c),
	.w7(32'hb97ee6ab),
	.w8(32'hb9dabb32),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900bc3f),
	.w1(32'h39905a79),
	.w2(32'hb94676b3),
	.w3(32'hb987df1c),
	.w4(32'hb907d276),
	.w5(32'h39855dc1),
	.w6(32'h39d5e3f2),
	.w7(32'hb8b9d9a8),
	.w8(32'hb95de992),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab25b8),
	.w1(32'h394d625d),
	.w2(32'h39489572),
	.w3(32'h398c676d),
	.w4(32'hb98daf36),
	.w5(32'hb7a5bbfe),
	.w6(32'h390505b7),
	.w7(32'hb7b3ec56),
	.w8(32'h3910b777),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999dc14),
	.w1(32'hb9b18f5c),
	.w2(32'h37d813bc),
	.w3(32'h37c9bdf2),
	.w4(32'hb90006df),
	.w5(32'h3926bb02),
	.w6(32'hb98c1c67),
	.w7(32'hb931e3e9),
	.w8(32'hb96e39e1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92915f0),
	.w1(32'hb87b74d5),
	.w2(32'h386c5702),
	.w3(32'hb8a1b568),
	.w4(32'hb8006064),
	.w5(32'h395ffdcb),
	.w6(32'h38a48371),
	.w7(32'h3856f802),
	.w8(32'h3923144b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9969d23),
	.w1(32'hb9e2e6b5),
	.w2(32'hb99d69a7),
	.w3(32'hb94d3ab7),
	.w4(32'hb8d5e28e),
	.w5(32'h3a0c4755),
	.w6(32'h37cabac6),
	.w7(32'hb99efee4),
	.w8(32'h390948e8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d089d4),
	.w1(32'hb99b72fc),
	.w2(32'h382b9cba),
	.w3(32'h371b8c12),
	.w4(32'hba16d6c4),
	.w5(32'hb9ff50d2),
	.w6(32'hb9a0b34e),
	.w7(32'hb9e661d1),
	.w8(32'hba93c23a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f54a9),
	.w1(32'hb90fa5b9),
	.w2(32'h3ac04655),
	.w3(32'h3b1cee9f),
	.w4(32'h3acda949),
	.w5(32'h3ae3ff9a),
	.w6(32'h3af3a8c3),
	.w7(32'h3a29597d),
	.w8(32'h39b9c2b2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394114fe),
	.w1(32'h3a131c39),
	.w2(32'h39f5d045),
	.w3(32'hba2174bc),
	.w4(32'h39d9fb3d),
	.w5(32'h39898b20),
	.w6(32'h378c4603),
	.w7(32'h38002f7b),
	.w8(32'hb997fcd9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb881e8dd),
	.w1(32'hba9ecf94),
	.w2(32'hba156e27),
	.w3(32'hb94ec6ac),
	.w4(32'hba5ecb74),
	.w5(32'h38c27471),
	.w6(32'hba0803ef),
	.w7(32'hba5af1ee),
	.w8(32'hb9836c39),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7457cac),
	.w1(32'h3a0a590c),
	.w2(32'hb9329056),
	.w3(32'h3a2efabc),
	.w4(32'h3778f9be),
	.w5(32'h398271a7),
	.w6(32'h3a6c091f),
	.w7(32'h3a3b22d3),
	.w8(32'hb81070a2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff7d90),
	.w1(32'hb9d9ecdd),
	.w2(32'hba9b09f6),
	.w3(32'hba338fcd),
	.w4(32'hbad2d6b0),
	.w5(32'hbadf6843),
	.w6(32'h3b0c3166),
	.w7(32'h3a970f23),
	.w8(32'hb99b6a25),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883c7f7),
	.w1(32'h3971b3f7),
	.w2(32'h3a1074d9),
	.w3(32'h3998e237),
	.w4(32'h39548250),
	.w5(32'hb878df46),
	.w6(32'h37d11307),
	.w7(32'h39226876),
	.w8(32'h383dd8a0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bf598f),
	.w1(32'h39a6890b),
	.w2(32'h398a68b4),
	.w3(32'h39a2ebca),
	.w4(32'hb85c3af7),
	.w5(32'hb99b77f5),
	.w6(32'h373c1191),
	.w7(32'h36fd59e9),
	.w8(32'hb8846828),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3889170c),
	.w1(32'hb99e747b),
	.w2(32'h39bb18b8),
	.w3(32'hb9ec9309),
	.w4(32'hba4e2e13),
	.w5(32'hb9e4cee4),
	.w6(32'hba184dd1),
	.w7(32'h38a6758e),
	.w8(32'hb945f327),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e23c1a),
	.w1(32'h398c1aa9),
	.w2(32'h39fc9e4b),
	.w3(32'hb9b08abd),
	.w4(32'h39c6c6e9),
	.w5(32'h39479dd8),
	.w6(32'hba238f8e),
	.w7(32'hb9f5ee0b),
	.w8(32'hb960a472),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915c53e),
	.w1(32'hb9f311fc),
	.w2(32'h3a07838f),
	.w3(32'hbaec3836),
	.w4(32'hbaeb6d71),
	.w5(32'h39ccf8fe),
	.w6(32'hb8d16f74),
	.w7(32'h3af8a41b),
	.w8(32'h3ac24909),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb917bec4),
	.w1(32'hb90816e1),
	.w2(32'hb999170c),
	.w3(32'h3849412f),
	.w4(32'hb9db7b19),
	.w5(32'hb9bf38d8),
	.w6(32'h397a65f0),
	.w7(32'hb8e2d0fd),
	.w8(32'hb91a9414),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e190b4),
	.w1(32'h390d9030),
	.w2(32'h395b02ec),
	.w3(32'h3a144855),
	.w4(32'hb8d56e7b),
	.w5(32'hb711ae65),
	.w6(32'h38a65dd3),
	.w7(32'h38f47ad3),
	.w8(32'h39262687),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944acef),
	.w1(32'h362fb627),
	.w2(32'hb9ba53e4),
	.w3(32'h37b9c623),
	.w4(32'hb988c7fb),
	.w5(32'hb80cabe6),
	.w6(32'h3a1446fc),
	.w7(32'h38b61ce4),
	.w8(32'h39711c99),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d97eaf),
	.w1(32'hb9e6ab1d),
	.w2(32'hba6501e9),
	.w3(32'h3957e0a4),
	.w4(32'h3933e2d0),
	.w5(32'hb8f3a1a0),
	.w6(32'hb9ff2070),
	.w7(32'hb9194581),
	.w8(32'hb81b8df5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcbbb6),
	.w1(32'hb9b344db),
	.w2(32'h396f41f8),
	.w3(32'hb98ecc80),
	.w4(32'h38ac1c53),
	.w5(32'h39ba138c),
	.w6(32'h38f541cf),
	.w7(32'h39800140),
	.w8(32'h393a733a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382642e0),
	.w1(32'hb9520fff),
	.w2(32'hb9a2ffb5),
	.w3(32'h39a2b059),
	.w4(32'hb979dba1),
	.w5(32'hb9bca728),
	.w6(32'hb96cde0c),
	.w7(32'hb9969d38),
	.w8(32'hb857abf8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14499e),
	.w1(32'h39dccd1b),
	.w2(32'h39982fe4),
	.w3(32'h3a0982b3),
	.w4(32'h39cf0d8f),
	.w5(32'h39e0eff8),
	.w6(32'h3995a6ad),
	.w7(32'h391f47b8),
	.w8(32'hb89a64cc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397f8237),
	.w1(32'hb78cca5f),
	.w2(32'h3a1ae5f6),
	.w3(32'h3a0e43b1),
	.w4(32'h36a968af),
	.w5(32'h39fd2628),
	.w6(32'h37612352),
	.w7(32'h3979c64a),
	.w8(32'h391599c5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384a015c),
	.w1(32'hb6b74553),
	.w2(32'h390097ce),
	.w3(32'hb867b439),
	.w4(32'hb7c67315),
	.w5(32'h388c2f54),
	.w6(32'hb9015fd6),
	.w7(32'hb8b9b88d),
	.w8(32'h3792cc1c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab8e6d),
	.w1(32'hb9abc131),
	.w2(32'h38fbf2a0),
	.w3(32'h39a50a31),
	.w4(32'hb8975274),
	.w5(32'h3979c173),
	.w6(32'hb963f0c4),
	.w7(32'hb8c5153a),
	.w8(32'hb96fd141),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b4dd4),
	.w1(32'hb85e80c9),
	.w2(32'h396b0890),
	.w3(32'hb830564a),
	.w4(32'h377a1f31),
	.w5(32'h393f5382),
	.w6(32'hb7f3a5d2),
	.w7(32'h397d4b9e),
	.w8(32'hb9513baa),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e4e0a6),
	.w1(32'h39351d2e),
	.w2(32'h398aaf8b),
	.w3(32'h391c86af),
	.w4(32'h3999042e),
	.w5(32'h3859be68),
	.w6(32'h39a40f78),
	.w7(32'h399e3d98),
	.w8(32'h396bd1d6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d1db8),
	.w1(32'hba445af3),
	.w2(32'hba31bfdf),
	.w3(32'hba995244),
	.w4(32'hbac2ac00),
	.w5(32'hbacd67fc),
	.w6(32'hb9e54c2c),
	.w7(32'hba2b0849),
	.w8(32'hba8a1605),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb965fc0e),
	.w1(32'h3a01207b),
	.w2(32'h39e8290c),
	.w3(32'hb99140f7),
	.w4(32'h3a1ef4ad),
	.w5(32'h3a2cb53c),
	.w6(32'h39fa1183),
	.w7(32'h38c8663d),
	.w8(32'h3988130e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0d7f3),
	.w1(32'hb9078c5a),
	.w2(32'hb882da76),
	.w3(32'hb9b32591),
	.w4(32'hb973b91a),
	.w5(32'hb9438c7e),
	.w6(32'hb8add0d2),
	.w7(32'hb922f79f),
	.w8(32'hb8a15bd4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d3b26),
	.w1(32'hba0eafcf),
	.w2(32'hb9b111c9),
	.w3(32'hb9a7b926),
	.w4(32'hb9fc0ffb),
	.w5(32'hb992fe0f),
	.w6(32'hba0ab9c8),
	.w7(32'hb8014417),
	.w8(32'hb94a19b8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6aa678),
	.w1(32'hb9db366b),
	.w2(32'hb7fbcc1a),
	.w3(32'hba3b63ff),
	.w4(32'hba4c7e7e),
	.w5(32'hb96fda62),
	.w6(32'hb7ed99fb),
	.w7(32'h3a2cbca5),
	.w8(32'h3a1792ec),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97885ae),
	.w1(32'hb92cc5d0),
	.w2(32'h3a18f51f),
	.w3(32'hb9cdbe64),
	.w4(32'h39056862),
	.w5(32'h3a72c473),
	.w6(32'hb886192a),
	.w7(32'hb881641a),
	.w8(32'h39bd5226),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75f4932),
	.w1(32'h38881041),
	.w2(32'hb71cac80),
	.w3(32'h37afa2c8),
	.w4(32'hb80f56ca),
	.w5(32'h374d88e9),
	.w6(32'h3906a9a2),
	.w7(32'h389ccc40),
	.w8(32'hb81d4a37),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd048c),
	.w1(32'hb89ef28a),
	.w2(32'h3a954249),
	.w3(32'h3a46e9f6),
	.w4(32'h3a6e26f7),
	.w5(32'h3a9a7d8f),
	.w6(32'h39a3912c),
	.w7(32'h3ab8716e),
	.w8(32'h3ab052a1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912fd35),
	.w1(32'h396c209c),
	.w2(32'hb98cde33),
	.w3(32'hb9476c1d),
	.w4(32'hba25e742),
	.w5(32'hba0317ae),
	.w6(32'h39e43918),
	.w7(32'h39135985),
	.w8(32'h38ddf0a4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2c10a),
	.w1(32'h39088555),
	.w2(32'hb99295a8),
	.w3(32'hba3942b1),
	.w4(32'hb9f4b6c5),
	.w5(32'hba8a9708),
	.w6(32'h38adc2ff),
	.w7(32'hb9880100),
	.w8(32'hba3f1633),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6795d),
	.w1(32'hb9cf6b0e),
	.w2(32'hba0cf0c4),
	.w3(32'hb83a4bab),
	.w4(32'hb944d931),
	.w5(32'hb94ada1f),
	.w6(32'hba4b0749),
	.w7(32'hba8f95e5),
	.w8(32'hba5b9d98),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46a97d),
	.w1(32'h3886e8a7),
	.w2(32'hba509dc6),
	.w3(32'hbae936c7),
	.w4(32'hbab73711),
	.w5(32'hba9cb040),
	.w6(32'hba257320),
	.w7(32'h38828f78),
	.w8(32'hb9913b09),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11d33e),
	.w1(32'hb90b2e62),
	.w2(32'hb91036ae),
	.w3(32'hb9f48826),
	.w4(32'hb9c6347f),
	.w5(32'hb9548456),
	.w6(32'h37c6ebf6),
	.w7(32'h390c4dc0),
	.w8(32'hb7c23a48),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c24cff),
	.w1(32'h398e9be6),
	.w2(32'h391d8645),
	.w3(32'hba57beff),
	.w4(32'hb96a51ed),
	.w5(32'hb8b39049),
	.w6(32'h38c3603a),
	.w7(32'hb9829a94),
	.w8(32'hba19ddaa),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87a26f4),
	.w1(32'hba15d0a7),
	.w2(32'h39ea2f2f),
	.w3(32'h394b19cd),
	.w4(32'hba0096e0),
	.w5(32'h39cd5409),
	.w6(32'hb9b6ef64),
	.w7(32'h39e66718),
	.w8(32'hb8b32255),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a96ce),
	.w1(32'h39fef777),
	.w2(32'h3adf33f9),
	.w3(32'h3ab38ebf),
	.w4(32'h3a7d9be5),
	.w5(32'h3ae00037),
	.w6(32'hba7e2ac4),
	.w7(32'h39b27674),
	.w8(32'hb7878f80),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e539a),
	.w1(32'hba6df622),
	.w2(32'h3948cdf6),
	.w3(32'hb98762ae),
	.w4(32'hb997f251),
	.w5(32'h3a1c5b6d),
	.w6(32'hb86db49b),
	.w7(32'h385025d4),
	.w8(32'hb905ab73),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ccfd9f),
	.w1(32'hb861ef7e),
	.w2(32'hb68c54e0),
	.w3(32'hb93487c4),
	.w4(32'hba091742),
	.w5(32'hb84dff33),
	.w6(32'hb96dd1bf),
	.w7(32'hb8e274d0),
	.w8(32'hb4c655a0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8271dad),
	.w1(32'h39500b18),
	.w2(32'h38c895cb),
	.w3(32'hb88da5c2),
	.w4(32'hb9423ca6),
	.w5(32'h38716041),
	.w6(32'h3a1078ff),
	.w7(32'h3a25e4d8),
	.w8(32'h3a4e5363),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39267c31),
	.w1(32'hb7f5ec0f),
	.w2(32'h38854612),
	.w3(32'hba4f3d1c),
	.w4(32'hb9d98278),
	.w5(32'hbaba10b7),
	.w6(32'h38f389b4),
	.w7(32'h39c83297),
	.w8(32'hb9e5d7f7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0d9cf),
	.w1(32'h38d4b5c5),
	.w2(32'h39a2f0ce),
	.w3(32'hb997184e),
	.w4(32'h3938abf8),
	.w5(32'hb8bfef8f),
	.w6(32'hb9df2a42),
	.w7(32'h38e478ee),
	.w8(32'hb9ab6892),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39387fb7),
	.w1(32'h39414f04),
	.w2(32'h3a20a19e),
	.w3(32'hb9f7445f),
	.w4(32'h398b1820),
	.w5(32'h38cc1c9d),
	.w6(32'hb9986d47),
	.w7(32'h394310ca),
	.w8(32'h39054773),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ca0b0),
	.w1(32'hb8c78e0d),
	.w2(32'h399b2572),
	.w3(32'h39c761b6),
	.w4(32'h391d6cd6),
	.w5(32'h39831372),
	.w6(32'hb9183519),
	.w7(32'hb9d61811),
	.w8(32'hb9ded24f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb688cd73),
	.w1(32'h38784989),
	.w2(32'hb91b63d6),
	.w3(32'hb8388e7f),
	.w4(32'hb89ad299),
	.w5(32'hb9463b08),
	.w6(32'h37fe587e),
	.w7(32'hb827d456),
	.w8(32'h3732f34a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb693760c),
	.w1(32'h395783f1),
	.w2(32'hb8b7ae75),
	.w3(32'hb80d8498),
	.w4(32'h379eca48),
	.w5(32'hb92a0eab),
	.w6(32'h390675c6),
	.w7(32'hb815f639),
	.w8(32'hb6a99ca2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cb9e8a),
	.w1(32'h3762b6af),
	.w2(32'h36f15274),
	.w3(32'h37cdcaac),
	.w4(32'hb813ea6e),
	.w5(32'h3994a8ca),
	.w6(32'h391aab8d),
	.w7(32'h3957d2e2),
	.w8(32'h38a82bfe),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941747c),
	.w1(32'h37d205c8),
	.w2(32'hb9c39854),
	.w3(32'hb892ce85),
	.w4(32'hb5a2e798),
	.w5(32'hba2b73d0),
	.w6(32'h37d93516),
	.w7(32'hb9878ec8),
	.w8(32'h39896abd),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3d43e),
	.w1(32'h39dea681),
	.w2(32'h3a56f70f),
	.w3(32'h39c44141),
	.w4(32'h3a3bd321),
	.w5(32'h3a3aab2c),
	.w6(32'hba1aecd3),
	.w7(32'hb9b68215),
	.w8(32'hb9ba19de),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82f5343),
	.w1(32'h371fe6e5),
	.w2(32'h394d72b8),
	.w3(32'hb8f50f43),
	.w4(32'h387dbe60),
	.w5(32'h3729d9aa),
	.w6(32'h38f2447c),
	.w7(32'h37b6b3e6),
	.w8(32'hb8edc0d2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f2e67),
	.w1(32'hbaa66b7f),
	.w2(32'hbac2ee6e),
	.w3(32'hba57bc7b),
	.w4(32'hbae88166),
	.w5(32'hba880ba3),
	.w6(32'h39f08a27),
	.w7(32'h3b1017d0),
	.w8(32'h3a0ee128),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01177e),
	.w1(32'h393d4f06),
	.w2(32'h39dd01db),
	.w3(32'hb958f4b4),
	.w4(32'h39fc9a24),
	.w5(32'h3a22ba12),
	.w6(32'hb8162f95),
	.w7(32'h38bb7307),
	.w8(32'hba155f52),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e3fc4),
	.w1(32'hb886199e),
	.w2(32'hb8e1cc7c),
	.w3(32'hba0eb5ba),
	.w4(32'hb8b57777),
	.w5(32'hb91a6f44),
	.w6(32'h3a5d262b),
	.w7(32'h3a1d0bb3),
	.w8(32'h3a3eafbe),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39672268),
	.w1(32'h391df01e),
	.w2(32'h3923b974),
	.w3(32'h38b308ff),
	.w4(32'hba019c5a),
	.w5(32'hba37dcb9),
	.w6(32'hb9a4a4f7),
	.w7(32'hb7bbbae7),
	.w8(32'hb8aab1ee),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2375c9),
	.w1(32'h3953de1e),
	.w2(32'h39f47196),
	.w3(32'hb9fb4043),
	.w4(32'h39b3cc4a),
	.w5(32'h39abda08),
	.w6(32'hb93ec01a),
	.w7(32'hb8e043f2),
	.w8(32'hb9fbd903),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e17e8),
	.w1(32'h39f3c114),
	.w2(32'h399bd6db),
	.w3(32'h392352bd),
	.w4(32'h396d3e87),
	.w5(32'hb7f367cc),
	.w6(32'h389b361e),
	.w7(32'h391e32eb),
	.w8(32'hb9632178),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aced53),
	.w1(32'hb93c5991),
	.w2(32'hb9e82593),
	.w3(32'hba22a7e0),
	.w4(32'hb8ecb106),
	.w5(32'hb9a6854d),
	.w6(32'hb9382e43),
	.w7(32'hb8571bd0),
	.w8(32'hb953e1c1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b7db6),
	.w1(32'hb9253ffc),
	.w2(32'hb8f60e4b),
	.w3(32'h386f8128),
	.w4(32'hb900916f),
	.w5(32'h37660f23),
	.w6(32'hb74fb008),
	.w7(32'hb7d1cca0),
	.w8(32'hb898ae65),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26f424),
	.w1(32'hba8e5891),
	.w2(32'hba05b751),
	.w3(32'h39dc3ebd),
	.w4(32'h37b17f4e),
	.w5(32'h39e7bd7f),
	.w6(32'h3a159da7),
	.w7(32'h3a0d1435),
	.w8(32'h3998d29b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a430cb5),
	.w1(32'h3a296bea),
	.w2(32'h3a96a263),
	.w3(32'h39760b5f),
	.w4(32'h3a053cae),
	.w5(32'h3ac378c1),
	.w6(32'hb9627044),
	.w7(32'h391fc4b2),
	.w8(32'h39d13e3f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba208f5b),
	.w1(32'hb9b69378),
	.w2(32'hb90dd83e),
	.w3(32'hb949b92a),
	.w4(32'h3872a50a),
	.w5(32'hb9d96eb9),
	.w6(32'hb9486315),
	.w7(32'hb980dd71),
	.w8(32'h39288ed5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39856678),
	.w1(32'h39023a37),
	.w2(32'h39f14a44),
	.w3(32'hb90524de),
	.w4(32'hb981d734),
	.w5(32'hb950ac02),
	.w6(32'h3953175e),
	.w7(32'h391f3d9a),
	.w8(32'h3a001e03),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999cec4),
	.w1(32'hb8456f3e),
	.w2(32'hb994b439),
	.w3(32'hba715e8e),
	.w4(32'hba85ef00),
	.w5(32'hba5049fc),
	.w6(32'hb7cf2caf),
	.w7(32'h3a1278e8),
	.w8(32'h3a4a0746),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f0d664),
	.w1(32'h389c5e1e),
	.w2(32'h381f0135),
	.w3(32'h3902fb84),
	.w4(32'h3a4213d1),
	.w5(32'h39b0ea52),
	.w6(32'h39af286b),
	.w7(32'h398e95fb),
	.w8(32'h3942f9fa),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb876e7d8),
	.w1(32'hb8189740),
	.w2(32'hb840fb52),
	.w3(32'hba8cc618),
	.w4(32'hbafc9549),
	.w5(32'hba8e43b2),
	.w6(32'hba7f9c09),
	.w7(32'hbae22175),
	.w8(32'hbb449df5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7e2f8),
	.w1(32'h3938da19),
	.w2(32'h3a0a66ef),
	.w3(32'hb98d98a0),
	.w4(32'hb98de895),
	.w5(32'h3a1c21f8),
	.w6(32'h38aa2cde),
	.w7(32'h3a4de757),
	.w8(32'h380f21d7),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b5957),
	.w1(32'h3a05bb32),
	.w2(32'hb8a53b73),
	.w3(32'hba0bb407),
	.w4(32'hbab65743),
	.w5(32'hbade4bc8),
	.w6(32'h3a0268eb),
	.w7(32'h3961474b),
	.w8(32'hb996c698),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8827721),
	.w1(32'hb78bd66e),
	.w2(32'hb9149027),
	.w3(32'h3962237d),
	.w4(32'h37513821),
	.w5(32'h390a3bcc),
	.w6(32'h3935cd74),
	.w7(32'hb91787dc),
	.w8(32'hb915071b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec211f),
	.w1(32'h39c5d22c),
	.w2(32'h39948a83),
	.w3(32'h38999683),
	.w4(32'h391e8d27),
	.w5(32'hb9928e14),
	.w6(32'hb98816ea),
	.w7(32'hb88b086f),
	.w8(32'hb847b6ef),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a000603),
	.w1(32'hb8e3041a),
	.w2(32'hb964aa0f),
	.w3(32'h381f7ca7),
	.w4(32'hb996e1cb),
	.w5(32'hb8a5753f),
	.w6(32'h397f8c3f),
	.w7(32'h353034f2),
	.w8(32'h3757d35a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb907abe3),
	.w1(32'h398b31c0),
	.w2(32'h38aae7fb),
	.w3(32'h38048aab),
	.w4(32'h38f71dbe),
	.w5(32'h3722d169),
	.w6(32'h392300eb),
	.w7(32'hb9401fda),
	.w8(32'h3894c634),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39142e5c),
	.w1(32'h39a72596),
	.w2(32'h39ba3924),
	.w3(32'hb9b51752),
	.w4(32'hba286036),
	.w5(32'hb9c662a9),
	.w6(32'hb976c80c),
	.w7(32'hb998a913),
	.w8(32'hb9bc21fa),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397ed3ac),
	.w1(32'hb8fbe53e),
	.w2(32'h392ef7a4),
	.w3(32'hb973165c),
	.w4(32'hb8aed752),
	.w5(32'h399c10e8),
	.w6(32'hb76908b7),
	.w7(32'hb8fb9c2c),
	.w8(32'hb861de8a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90578b1),
	.w1(32'h390bc4c2),
	.w2(32'hb925fb10),
	.w3(32'hba365cb9),
	.w4(32'hba2371c4),
	.w5(32'hba539233),
	.w6(32'h38227e65),
	.w7(32'hb8b5fd20),
	.w8(32'h37d2f3e0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b84a5),
	.w1(32'h395e414c),
	.w2(32'h391fa250),
	.w3(32'hb8f55fd8),
	.w4(32'h378340c2),
	.w5(32'h38e2b799),
	.w6(32'hb73a34b9),
	.w7(32'h3817691e),
	.w8(32'h375341e3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39faa25b),
	.w1(32'h39bce8e3),
	.w2(32'h39b42d34),
	.w3(32'h39ac383b),
	.w4(32'h3a29652a),
	.w5(32'h3a87b932),
	.w6(32'h39a18c23),
	.w7(32'hb94fb8e8),
	.w8(32'h39053d91),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90fee96),
	.w1(32'hb9573739),
	.w2(32'h3a19e601),
	.w3(32'hb88e9c58),
	.w4(32'h390815a6),
	.w5(32'h3a891d36),
	.w6(32'h38859564),
	.w7(32'h3929fc19),
	.w8(32'h3a12786e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38575271),
	.w1(32'hb87537fb),
	.w2(32'h38bf806d),
	.w3(32'h39981361),
	.w4(32'h3a38832d),
	.w5(32'h39d9eece),
	.w6(32'h399b58ac),
	.w7(32'hb9901a2b),
	.w8(32'h39bdd9b4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81abc87),
	.w1(32'hb7863007),
	.w2(32'h391026af),
	.w3(32'hb89a6af4),
	.w4(32'h3995501c),
	.w5(32'h399cf8ef),
	.w6(32'hb86d359c),
	.w7(32'h3897137c),
	.w8(32'hba22b370),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26fcb7),
	.w1(32'h390a62ad),
	.w2(32'hb9bbead6),
	.w3(32'hba2d2b53),
	.w4(32'h39391369),
	.w5(32'hb8d74da9),
	.w6(32'h38baa152),
	.w7(32'hb9833bf0),
	.w8(32'hb92e23db),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a0f10d),
	.w1(32'h39b64e36),
	.w2(32'hb80bcd3f),
	.w3(32'hb691420b),
	.w4(32'hb9851154),
	.w5(32'hba106e51),
	.w6(32'h39d61c98),
	.w7(32'h39203168),
	.w8(32'h39368f01),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfef7e),
	.w1(32'h39a60555),
	.w2(32'hb98fc0cf),
	.w3(32'h39d3812b),
	.w4(32'h3a01df3b),
	.w5(32'hb882479e),
	.w6(32'h37f61d4e),
	.w7(32'hb96946ae),
	.w8(32'h397e427e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f7b1bb),
	.w1(32'h37bf2adf),
	.w2(32'h398223ec),
	.w3(32'h3902c06d),
	.w4(32'h392666e6),
	.w5(32'h395a4d6e),
	.w6(32'h39a922da),
	.w7(32'h38df9207),
	.w8(32'h389311f0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ebef60),
	.w1(32'h39ac9b00),
	.w2(32'h3a12ca29),
	.w3(32'h37700cc8),
	.w4(32'h39b4a86b),
	.w5(32'h3879404a),
	.w6(32'hb8422094),
	.w7(32'h39a8f31f),
	.w8(32'h39620fd6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391983c5),
	.w1(32'hb98cb29a),
	.w2(32'hb8492365),
	.w3(32'hb9c095dd),
	.w4(32'hb8941c56),
	.w5(32'hb923ec97),
	.w6(32'hba1b527f),
	.w7(32'hb921207e),
	.w8(32'h38c0b2ff),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb658a29b),
	.w1(32'h39fb6aea),
	.w2(32'hba513391),
	.w3(32'hb8d3c8b4),
	.w4(32'h3a1a9f31),
	.w5(32'hba2683bb),
	.w6(32'h39ba8f30),
	.w7(32'hb9d46100),
	.w8(32'h38d5c0a8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99233a5),
	.w1(32'hb861af09),
	.w2(32'hb9241a55),
	.w3(32'hb9b827f1),
	.w4(32'hba2dae31),
	.w5(32'hba17a9c1),
	.w6(32'hb99a4040),
	.w7(32'h3a24cabb),
	.w8(32'h395cb7ac),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01683a),
	.w1(32'hba165001),
	.w2(32'hba5d64f7),
	.w3(32'hb9ae7f1b),
	.w4(32'hba3fed8d),
	.w5(32'hb9d4518a),
	.w6(32'hb8b270c8),
	.w7(32'hb9f40e91),
	.w8(32'hb98b90ce),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930f19c),
	.w1(32'h39afea3f),
	.w2(32'h39caedf5),
	.w3(32'h39ae64d0),
	.w4(32'hb907473c),
	.w5(32'hb9396c82),
	.w6(32'hb89f9f21),
	.w7(32'h37f4c314),
	.w8(32'h38aa1d8d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b7899),
	.w1(32'h38e2647f),
	.w2(32'h3926fb49),
	.w3(32'h39460ac2),
	.w4(32'h38f4ca0f),
	.w5(32'h38aa527f),
	.w6(32'h38d7351e),
	.w7(32'h38484f28),
	.w8(32'hb927e875),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07e445),
	.w1(32'h39861910),
	.w2(32'h3974bc02),
	.w3(32'h39d534d7),
	.w4(32'h393a3004),
	.w5(32'h3949db74),
	.w6(32'h39ca8063),
	.w7(32'h3913fc81),
	.w8(32'h399ce810),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cdad05),
	.w1(32'h38fb2072),
	.w2(32'h3931400d),
	.w3(32'h3850d0c6),
	.w4(32'h38a0e7cb),
	.w5(32'hb98daefa),
	.w6(32'hb99b314e),
	.w7(32'hba138f0a),
	.w8(32'hb96928d1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39947f74),
	.w1(32'h38686c30),
	.w2(32'hb91494c4),
	.w3(32'h39a63573),
	.w4(32'h397082c1),
	.w5(32'h38b442b4),
	.w6(32'h38c7385e),
	.w7(32'hb8941495),
	.w8(32'h3895f472),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c4e7a),
	.w1(32'hb8e785ac),
	.w2(32'hb94d735e),
	.w3(32'h39a37932),
	.w4(32'h38302b08),
	.w5(32'hb8fbfe20),
	.w6(32'h3924e95b),
	.w7(32'hb93ba508),
	.w8(32'hb9add105),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86f4754),
	.w1(32'hb9b605a3),
	.w2(32'hba01f64c),
	.w3(32'hb8f06695),
	.w4(32'hb946fbf4),
	.w5(32'hb7da5a3e),
	.w6(32'h39ee3e87),
	.w7(32'h3a30173e),
	.w8(32'h38719c89),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e5b42),
	.w1(32'h394303fa),
	.w2(32'hb8c77c2e),
	.w3(32'hb8ea8a90),
	.w4(32'hb9dc6db4),
	.w5(32'hb975e982),
	.w6(32'h39b7a030),
	.w7(32'hb7fc0212),
	.w8(32'hb8666e9c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f31c9),
	.w1(32'h3977d6e0),
	.w2(32'hb65f4dea),
	.w3(32'hb8e8c0d3),
	.w4(32'h38c21dcd),
	.w5(32'hb88daeaa),
	.w6(32'h3944a0a5),
	.w7(32'h388574df),
	.w8(32'h38a5e5f3),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c5118e),
	.w1(32'h38152da3),
	.w2(32'hb7f96206),
	.w3(32'hb9136110),
	.w4(32'h38ecdc4a),
	.w5(32'hb928a73b),
	.w6(32'hb92deb99),
	.w7(32'h38b4a381),
	.w8(32'h369cd254),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39093786),
	.w1(32'h3803e675),
	.w2(32'h399e1cea),
	.w3(32'hb9ad2e4b),
	.w4(32'hb860ace1),
	.w5(32'h39e3a76c),
	.w6(32'hb9e9dfdc),
	.w7(32'hb9c3ac9a),
	.w8(32'hb9a48426),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b2a45),
	.w1(32'h39110c7f),
	.w2(32'hb89f2435),
	.w3(32'hb80c24f5),
	.w4(32'h38b41353),
	.w5(32'h3918a9cb),
	.w6(32'h387c6e95),
	.w7(32'hb8ed41f7),
	.w8(32'h39e0e3c8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad4b4f),
	.w1(32'h3991fbf1),
	.w2(32'h39b542da),
	.w3(32'hb9a3f548),
	.w4(32'h3952b27b),
	.w5(32'h3958bdf4),
	.w6(32'hb7819244),
	.w7(32'hb69cc5c6),
	.w8(32'hb6d30a51),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01fa4b),
	.w1(32'h39851686),
	.w2(32'h3a24fba8),
	.w3(32'hba8579e0),
	.w4(32'hba2286b0),
	.w5(32'hba3c0699),
	.w6(32'hb9f9ed36),
	.w7(32'hb9fecae6),
	.w8(32'hba5a5714),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382f6868),
	.w1(32'h39945d41),
	.w2(32'hb99893f0),
	.w3(32'h38d3b639),
	.w4(32'h3994a5d6),
	.w5(32'hb924150a),
	.w6(32'h393b79d4),
	.w7(32'hb902f674),
	.w8(32'h38bb3ad9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9213b56),
	.w1(32'h3749843f),
	.w2(32'hb924f810),
	.w3(32'hb91c54e6),
	.w4(32'hb83c8bd7),
	.w5(32'hb95b8b77),
	.w6(32'h38568657),
	.w7(32'hb877e67b),
	.w8(32'hb7ae9673),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dc6145),
	.w1(32'h367fe5ca),
	.w2(32'hb802e908),
	.w3(32'hb8f149a0),
	.w4(32'hb8e1988f),
	.w5(32'h368d835a),
	.w6(32'h39641df2),
	.w7(32'hb968b38b),
	.w8(32'hb93003f5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d3d5e1),
	.w1(32'hba07ec57),
	.w2(32'hba26761f),
	.w3(32'hb83dc469),
	.w4(32'h393ff767),
	.w5(32'h380a279c),
	.w6(32'h396f230a),
	.w7(32'h398928a9),
	.w8(32'h39c02fc3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908f683),
	.w1(32'h39ad777f),
	.w2(32'h3a2434bb),
	.w3(32'hb8c82b0e),
	.w4(32'h39691f1f),
	.w5(32'h379b87b4),
	.w6(32'hb8349eaf),
	.w7(32'h3a363c21),
	.w8(32'h3a1498be),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f7849),
	.w1(32'hbb13a8db),
	.w2(32'hbb93cfe8),
	.w3(32'hb90d034f),
	.w4(32'h39b29639),
	.w5(32'h3af3ecd1),
	.w6(32'hbb9aa74c),
	.w7(32'hbb81ccee),
	.w8(32'hbab7f25d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba236c61),
	.w1(32'h3c884c9d),
	.w2(32'h3ce7451f),
	.w3(32'hb9791fe0),
	.w4(32'h3c061512),
	.w5(32'h3c22fc6a),
	.w6(32'h3bbf9779),
	.w7(32'h3cc2abbd),
	.w8(32'h3cabd2fe),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule