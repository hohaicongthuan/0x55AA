module layer_10_featuremap_293(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4352c3),
	.w1(32'hbaef6ed9),
	.w2(32'h3b6167be),
	.w3(32'hbabf8955),
	.w4(32'h3c1be440),
	.w5(32'hbb5972c4),
	.w6(32'h3ab719ef),
	.w7(32'h3bdff202),
	.w8(32'hbc0a1944),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacf302),
	.w1(32'hbb29e1de),
	.w2(32'h3c2da084),
	.w3(32'h3b2e254f),
	.w4(32'h3aaba833),
	.w5(32'h3bbd5582),
	.w6(32'hbab52fca),
	.w7(32'h3c45c8e1),
	.w8(32'h3c447792),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eeb1d),
	.w1(32'h3aaf603c),
	.w2(32'hbbf4a544),
	.w3(32'h3b6f9189),
	.w4(32'hbbe1a29b),
	.w5(32'h3b208031),
	.w6(32'h3b6d8f33),
	.w7(32'hbc2d33ec),
	.w8(32'hbb93c6a8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9e041),
	.w1(32'hba071fb1),
	.w2(32'hbb35a755),
	.w3(32'h3b88efd5),
	.w4(32'h3ab3bf8e),
	.w5(32'h3be8d03c),
	.w6(32'hba678538),
	.w7(32'h3b4ac664),
	.w8(32'h3c80acaa),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e1591),
	.w1(32'hbc99d723),
	.w2(32'h3c4da35a),
	.w3(32'hbcaa7a8d),
	.w4(32'h3c547826),
	.w5(32'hbc1c4586),
	.w6(32'hbc41428d),
	.w7(32'h3ca1ef51),
	.w8(32'hbcec90e7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca47828),
	.w1(32'hbb1a2792),
	.w2(32'h3c87660e),
	.w3(32'h3c269133),
	.w4(32'h3ccf9ceb),
	.w5(32'hbc226cc7),
	.w6(32'hbb550d2e),
	.w7(32'h3cc1f895),
	.w8(32'hbc97db05),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12f293),
	.w1(32'h3b17a432),
	.w2(32'h3cb4497c),
	.w3(32'h3b39d050),
	.w4(32'h3c841247),
	.w5(32'hbcb88fbb),
	.w6(32'hbb0277c3),
	.w7(32'h3cb29b83),
	.w8(32'hbd010e50),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c2a3c),
	.w1(32'h3a6dd31a),
	.w2(32'h3c78b7e7),
	.w3(32'hbc02ed20),
	.w4(32'hbaba0edc),
	.w5(32'hbd0bfb8d),
	.w6(32'hbbd27d5b),
	.w7(32'h3c8db3c9),
	.w8(32'hbd43e9a9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1a8a21),
	.w1(32'hbc1ceb81),
	.w2(32'h3cb3b69b),
	.w3(32'hbb4ef9ea),
	.w4(32'h3cc7a816),
	.w5(32'hbc15364e),
	.w6(32'hbbee9fc9),
	.w7(32'h3d073e4f),
	.w8(32'hbce167ff),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc805d4),
	.w1(32'hbc010c52),
	.w2(32'h3c4ad2b6),
	.w3(32'h3ba00a64),
	.w4(32'h3cadc17b),
	.w5(32'hbb3a0e12),
	.w6(32'hbc1b3754),
	.w7(32'h3c982746),
	.w8(32'hbc677f2c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085f95),
	.w1(32'h3b194997),
	.w2(32'h3c282dea),
	.w3(32'h3b6f922c),
	.w4(32'h3c13625f),
	.w5(32'h3a452a2e),
	.w6(32'hbb641208),
	.w7(32'h3c4c8759),
	.w8(32'h3c608106),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88c225),
	.w1(32'h3a09fc0a),
	.w2(32'h3bb51d34),
	.w3(32'hba51662f),
	.w4(32'hbc476ad7),
	.w5(32'h3a3ae0e0),
	.w6(32'hbb7a4b23),
	.w7(32'hbc0136ef),
	.w8(32'hb9994e82),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ecbbb),
	.w1(32'hbb0a43a2),
	.w2(32'hbc2089e3),
	.w3(32'hbc7eb2d6),
	.w4(32'hbc87b89a),
	.w5(32'hbc236dfd),
	.w6(32'hbbb47598),
	.w7(32'hbb5c6977),
	.w8(32'hba838cf9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad3047),
	.w1(32'hbc1ddc4a),
	.w2(32'h3b67ecba),
	.w3(32'hbc72f843),
	.w4(32'h3b509ae5),
	.w5(32'hbb7dbbb5),
	.w6(32'h38bb3a61),
	.w7(32'h3a875282),
	.w8(32'hbc5f48cd),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b8d0f),
	.w1(32'h3bfdb6b1),
	.w2(32'h3bae944a),
	.w3(32'hbb2b3049),
	.w4(32'h3b0852ed),
	.w5(32'hbb4f9f6f),
	.w6(32'h38c84bc6),
	.w7(32'h3c1a5180),
	.w8(32'hbc11d0d8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2836f4),
	.w1(32'hbbd4cf50),
	.w2(32'h3c1b13ba),
	.w3(32'h39f5a9c4),
	.w4(32'h3ca9ff2e),
	.w5(32'hbc5488f6),
	.w6(32'hbc066129),
	.w7(32'h3cc24c08),
	.w8(32'hbcae3838),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc648729),
	.w1(32'h3b988e2a),
	.w2(32'h3cd4bf75),
	.w3(32'h3b53a16e),
	.w4(32'h3cbf9376),
	.w5(32'h3c779f08),
	.w6(32'hba81a09d),
	.w7(32'h3cfd1b54),
	.w8(32'h3cb6fbcd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb736c),
	.w1(32'hbc0d7ba4),
	.w2(32'hbced8bb0),
	.w3(32'hbc2f302c),
	.w4(32'hbcef14f9),
	.w5(32'h3c6cb378),
	.w6(32'hbb377380),
	.w7(32'hbcdee220),
	.w8(32'h3ccdd3c8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99fe7f),
	.w1(32'hbb530775),
	.w2(32'hbcdd7d37),
	.w3(32'hb9e1cf3b),
	.w4(32'hbcc8b99e),
	.w5(32'hbbcf4981),
	.w6(32'h3ae2b76e),
	.w7(32'hbd189ac1),
	.w8(32'hbc1cb5bd),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe9167),
	.w1(32'hbbc2a0e9),
	.w2(32'hbc0bf9a2),
	.w3(32'h3990a296),
	.w4(32'h3b175531),
	.w5(32'hbc09536a),
	.w6(32'h3a98e1ea),
	.w7(32'hba75ba0e),
	.w8(32'hbbdd68f8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e10b6),
	.w1(32'hbbc4f4b7),
	.w2(32'hba8a21fc),
	.w3(32'hba908b8c),
	.w4(32'h3c1f3075),
	.w5(32'hbc80535b),
	.w6(32'hbaedf785),
	.w7(32'h3c3faf7d),
	.w8(32'hbc98e601),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8395d2),
	.w1(32'h3bd83bd0),
	.w2(32'h3c9db56c),
	.w3(32'h3c20fcaa),
	.w4(32'h3ca4a5e8),
	.w5(32'h3b2d1b9a),
	.w6(32'h3b62723c),
	.w7(32'h3cb9cb1f),
	.w8(32'h3b5026af),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb88f8),
	.w1(32'hbc2aad77),
	.w2(32'hbc5e14a7),
	.w3(32'hbbd9420d),
	.w4(32'hbc093fef),
	.w5(32'hbc4acd63),
	.w6(32'hbb8b4f5a),
	.w7(32'hbc2a1d71),
	.w8(32'hbcae6600),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc452aa8),
	.w1(32'hbc1faa62),
	.w2(32'h3bc45d2a),
	.w3(32'hbc06a62e),
	.w4(32'h3c50cfad),
	.w5(32'h3c563269),
	.w6(32'h3b3ee14c),
	.w7(32'h3c627df2),
	.w8(32'h3c54b28f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6edfd),
	.w1(32'h3bd3aebf),
	.w2(32'hbc05e28a),
	.w3(32'h3bdb8aaf),
	.w4(32'h3aff0293),
	.w5(32'hbb1b0f9c),
	.w6(32'h3a88f23a),
	.w7(32'hbc53a6b9),
	.w8(32'hbc5c3978),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca0518),
	.w1(32'h3b894b3c),
	.w2(32'h3c24a222),
	.w3(32'h3ad6e7e8),
	.w4(32'h3c3d351a),
	.w5(32'hba610db3),
	.w6(32'h3b0b9d3b),
	.w7(32'h3c684258),
	.w8(32'hbbd4e2e7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39977a),
	.w1(32'hbbb51722),
	.w2(32'h3c2a075b),
	.w3(32'hbb86528a),
	.w4(32'h3c41862e),
	.w5(32'hbc8b6936),
	.w6(32'hbbd11d0f),
	.w7(32'h3c730738),
	.w8(32'hbce7ce81),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd8f123),
	.w1(32'hbac1eb1b),
	.w2(32'h3c8a9950),
	.w3(32'h3bbdd5c0),
	.w4(32'h3d049b5f),
	.w5(32'hb9d9e312),
	.w6(32'h3b6cfd90),
	.w7(32'h3cd07680),
	.w8(32'h3b1d4aca),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd59825),
	.w1(32'hbae843d2),
	.w2(32'hbc42dc45),
	.w3(32'hba5ca8b0),
	.w4(32'h3b6d6f91),
	.w5(32'hbbd93caf),
	.w6(32'h3b8e0288),
	.w7(32'hbbbf0c79),
	.w8(32'hbbd8c4ad),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaacabd),
	.w1(32'h3913b220),
	.w2(32'h3c1468f4),
	.w3(32'hbaaffb0b),
	.w4(32'h3c58b6e4),
	.w5(32'h3c08a838),
	.w6(32'hbbecdec1),
	.w7(32'h3c4f788e),
	.w8(32'h3be907de),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc124595),
	.w1(32'hbc182394),
	.w2(32'hba52895b),
	.w3(32'hbc9a6699),
	.w4(32'hbcb7b0fb),
	.w5(32'hbc34feab),
	.w6(32'hbbdc1cd2),
	.w7(32'hbbb33f7a),
	.w8(32'h39a10a9b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fe700),
	.w1(32'hbb5d2a06),
	.w2(32'hbc519f84),
	.w3(32'hba1f5190),
	.w4(32'hba2c7e7e),
	.w5(32'h3c3f977d),
	.w6(32'hbb2a2d88),
	.w7(32'hbbcd8e99),
	.w8(32'h3c3e7939),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62c8bf),
	.w1(32'hbbb3f34c),
	.w2(32'hbb20931b),
	.w3(32'hbb4cf519),
	.w4(32'hbcc720fa),
	.w5(32'h3c19e620),
	.w6(32'h3ab37d86),
	.w7(32'hbc95cf17),
	.w8(32'h3cb89fae),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62d8ab),
	.w1(32'h3a58efb3),
	.w2(32'hbc6370e0),
	.w3(32'hbbdc5f62),
	.w4(32'hbc6d8508),
	.w5(32'hbb85953c),
	.w6(32'hbb2ffbbc),
	.w7(32'hbc657ee2),
	.w8(32'hbb4e2f8f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52599e),
	.w1(32'hba51fc24),
	.w2(32'hbbbae0b6),
	.w3(32'h3a952d5b),
	.w4(32'h3c3140ef),
	.w5(32'h3c5c81fe),
	.w6(32'h3b38f4b1),
	.w7(32'hbac3e8ee),
	.w8(32'h3c01f102),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca7351),
	.w1(32'hbb23ad2d),
	.w2(32'hbc4fbbd4),
	.w3(32'h3b435fb3),
	.w4(32'hbc7a0647),
	.w5(32'h3c2a36b1),
	.w6(32'h3b8c8774),
	.w7(32'hbc84102b),
	.w8(32'h3c886bff),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3dbd08),
	.w1(32'hbc7bc32f),
	.w2(32'hbc807c4b),
	.w3(32'hbc2262bb),
	.w4(32'hbc3ff862),
	.w5(32'h3adb0fd5),
	.w6(32'hbba1af14),
	.w7(32'hbc61cbc8),
	.w8(32'hbc84d870),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9137b6),
	.w1(32'h3c532199),
	.w2(32'h3bc7afd4),
	.w3(32'h3c795ed0),
	.w4(32'h3c9f59d9),
	.w5(32'h38d8f46a),
	.w6(32'h3b6fad2c),
	.w7(32'h3c5aa897),
	.w8(32'hbc67804d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aade215),
	.w1(32'h3c3653e9),
	.w2(32'h3be86fdc),
	.w3(32'h3c89fbc2),
	.w4(32'h3c84734c),
	.w5(32'hb9b2a7db),
	.w6(32'h3c88c7de),
	.w7(32'h3c92673a),
	.w8(32'h3ce96758),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e670c),
	.w1(32'hba593909),
	.w2(32'hbc959ff0),
	.w3(32'hbb15235e),
	.w4(32'hbb77fa47),
	.w5(32'h3ba5f7a6),
	.w6(32'hba404f25),
	.w7(32'hbcbd18ac),
	.w8(32'h3c22f080),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d0892),
	.w1(32'hb9c1d3c4),
	.w2(32'hb80d85a1),
	.w3(32'hba866388),
	.w4(32'hbb93f7f2),
	.w5(32'hbb815407),
	.w6(32'h3ba2ac7f),
	.w7(32'hbb8d48ea),
	.w8(32'hbc5f00c0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9addc0),
	.w1(32'hba6ffe22),
	.w2(32'h3c0181ef),
	.w3(32'h3c1a486f),
	.w4(32'h3c3bbf3b),
	.w5(32'h3c956539),
	.w6(32'hba3a0b11),
	.w7(32'h3c67eaa4),
	.w8(32'h3ceaa5cf),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f4644),
	.w1(32'h3a9a82e2),
	.w2(32'hbc9ed495),
	.w3(32'h3a6881eb),
	.w4(32'hbc3c9d0c),
	.w5(32'h3ad9789e),
	.w6(32'h3b88cbcf),
	.w7(32'hbcb7a0dd),
	.w8(32'hbc260fbf),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbfc04),
	.w1(32'h3ae33444),
	.w2(32'h3c10d08d),
	.w3(32'hbbacf6d8),
	.w4(32'h3c01c753),
	.w5(32'h3c94f0ef),
	.w6(32'hbbc91ced),
	.w7(32'h3c8e94d7),
	.w8(32'h3d14bdec),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9fb67c),
	.w1(32'hbbd53d0e),
	.w2(32'hbd180866),
	.w3(32'hbb935c2a),
	.w4(32'hbccb177c),
	.w5(32'h3b865db2),
	.w6(32'hbc323ca7),
	.w7(32'hbd3ed94a),
	.w8(32'h3c5023d4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b088ad4),
	.w1(32'hba388582),
	.w2(32'hbabc4f87),
	.w3(32'h3b6abb8e),
	.w4(32'h3ae9d17f),
	.w5(32'h3cc44247),
	.w6(32'hba5ba2b0),
	.w7(32'hbc038b7a),
	.w8(32'h3ce44049),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90aff6),
	.w1(32'hbbf72ebd),
	.w2(32'hbc8bc0a9),
	.w3(32'hbbef38be),
	.w4(32'hbc1ac3d7),
	.w5(32'hbd1f05c2),
	.w6(32'hbc8abd94),
	.w7(32'hbcd53e69),
	.w8(32'hbd5b988e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd555515),
	.w1(32'hbcad6478),
	.w2(32'h3cfbd8d8),
	.w3(32'hbbbf5081),
	.w4(32'h3cf8bd18),
	.w5(32'hbc6e7bcd),
	.w6(32'hbbaae0cd),
	.w7(32'h3d735bcb),
	.w8(32'hbc5a09b4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5389a8),
	.w1(32'h3bd0a62b),
	.w2(32'h3ae7b23d),
	.w3(32'hbba579d0),
	.w4(32'hbc141858),
	.w5(32'hbc86553b),
	.w6(32'h3be63db3),
	.w7(32'h3bc0e0b9),
	.w8(32'hbcc9debe),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb52951),
	.w1(32'hba6876b4),
	.w2(32'h3c9fd168),
	.w3(32'h3b672fe0),
	.w4(32'h3cc1b276),
	.w5(32'h3ba58caa),
	.w6(32'hbb5fd6c7),
	.w7(32'h3cd924d8),
	.w8(32'h3b85559d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc834603),
	.w1(32'hbcaefb4e),
	.w2(32'h3bcd2c1f),
	.w3(32'hbc140064),
	.w4(32'h3a41d730),
	.w5(32'h3c50404d),
	.w6(32'hbc5bac1e),
	.w7(32'h3a21ae81),
	.w8(32'h3ce57aaf),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8832e8),
	.w1(32'h3c02c81a),
	.w2(32'hbca3dbea),
	.w3(32'hbb095147),
	.w4(32'hbc10ea0c),
	.w5(32'h3c47c8d2),
	.w6(32'h3bebd336),
	.w7(32'hbcacc478),
	.w8(32'h3b3cdc46),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb284506),
	.w1(32'h399a30aa),
	.w2(32'hbafd851e),
	.w3(32'h3b5c3e1b),
	.w4(32'hbba43f33),
	.w5(32'hbb90ae57),
	.w6(32'h3a9dd544),
	.w7(32'hbbae1e11),
	.w8(32'h3c574c7a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c850b3),
	.w1(32'hbbeb91a8),
	.w2(32'hb96aca1f),
	.w3(32'hbc0025dc),
	.w4(32'hbc7c57fb),
	.w5(32'h3b9a1b90),
	.w6(32'hbc0a6382),
	.w7(32'hbb0cc07e),
	.w8(32'h3c1b2803),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1205c),
	.w1(32'hba744024),
	.w2(32'hbc476f91),
	.w3(32'h3b9100eb),
	.w4(32'h3b409917),
	.w5(32'hbb648c7d),
	.w6(32'h3b75548f),
	.w7(32'hbb8df017),
	.w8(32'h38805938),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb1e8f),
	.w1(32'hbb7e4cd6),
	.w2(32'hbb88b6fc),
	.w3(32'hbb6c48b8),
	.w4(32'h3bac5394),
	.w5(32'hbba484ee),
	.w6(32'h3a32bdb3),
	.w7(32'hb98bab3d),
	.w8(32'h39b3c241),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb056915),
	.w1(32'h3b0014ba),
	.w2(32'hba80743e),
	.w3(32'h37fc950a),
	.w4(32'hbb1521cc),
	.w5(32'hbb399643),
	.w6(32'h3c171a62),
	.w7(32'hbb118929),
	.w8(32'hbb335fb8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2136e0),
	.w1(32'hbc087051),
	.w2(32'h3b839bf9),
	.w3(32'hbc38325d),
	.w4(32'h39b2de34),
	.w5(32'hbca1b7f8),
	.w6(32'hbc790d7d),
	.w7(32'h3b5d26f8),
	.w8(32'hbcf64301),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc2f068),
	.w1(32'hbb4f998f),
	.w2(32'h3cbedd19),
	.w3(32'h39e19919),
	.w4(32'h3cd119f4),
	.w5(32'hb964ae3d),
	.w6(32'hbbc79c75),
	.w7(32'h3ce1d713),
	.w8(32'h3bcd5d16),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfa1b2),
	.w1(32'h3c26d428),
	.w2(32'h3ab4d599),
	.w3(32'h3c2a5725),
	.w4(32'h38dc2007),
	.w5(32'hbc051a9e),
	.w6(32'h3c4e713c),
	.w7(32'hbbdc4705),
	.w8(32'hbc21fc1d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26a796),
	.w1(32'h39e8cea4),
	.w2(32'h3ac2a0c9),
	.w3(32'h3acf4f89),
	.w4(32'h3bcf8a6e),
	.w5(32'hbb8949f2),
	.w6(32'h3b0a3204),
	.w7(32'h3c0d658f),
	.w8(32'hbc7e25c0),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae538b),
	.w1(32'hbb9f58cb),
	.w2(32'h3bfa1d47),
	.w3(32'hba01ce9d),
	.w4(32'h3c24c7c6),
	.w5(32'h3c0d6746),
	.w6(32'hbadb4fa4),
	.w7(32'h3c6631d7),
	.w8(32'h3bd3c242),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc24711),
	.w1(32'h3b49302e),
	.w2(32'hb9f1c730),
	.w3(32'h3c020285),
	.w4(32'h3c682805),
	.w5(32'hba227862),
	.w6(32'h3c0a20ee),
	.w7(32'h3b7d0b06),
	.w8(32'h3c0c47a4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09aef4),
	.w1(32'hbc07c89e),
	.w2(32'hbc04968e),
	.w3(32'hbc32e32c),
	.w4(32'hbb9c57f4),
	.w5(32'h3a557671),
	.w6(32'h3a9ed434),
	.w7(32'hbc1f42cc),
	.w8(32'h3bac88fb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f6aca),
	.w1(32'hbbb4e99c),
	.w2(32'hbac8e10a),
	.w3(32'hbbcad421),
	.w4(32'h3c1ddbab),
	.w5(32'h3c42935a),
	.w6(32'hb980ed1d),
	.w7(32'h3b8782a9),
	.w8(32'h3b931399),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a644d70),
	.w1(32'h3aab26ee),
	.w2(32'hbb2a2fcf),
	.w3(32'h3c116a30),
	.w4(32'h3bc8b405),
	.w5(32'hbc5deed5),
	.w6(32'h39a2000b),
	.w7(32'hbacfbf25),
	.w8(32'hbcb0ae30),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9fae92),
	.w1(32'h3c57a62c),
	.w2(32'h3c240a24),
	.w3(32'hbb7d0591),
	.w4(32'h3b383444),
	.w5(32'hbc8b175d),
	.w6(32'h3bd2cb96),
	.w7(32'h3c8277a2),
	.w8(32'hbd2306e1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c0fba),
	.w1(32'hbc689e6e),
	.w2(32'h3cb7ff98),
	.w3(32'hbba0295f),
	.w4(32'h3ca13bd2),
	.w5(32'hbbedd3bb),
	.w6(32'hbc620265),
	.w7(32'h3ce704a1),
	.w8(32'hbc19a8a5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e4b39),
	.w1(32'hbd03e3a9),
	.w2(32'h3a949c29),
	.w3(32'hbc81c154),
	.w4(32'h3bef8ce1),
	.w5(32'h3ba88a40),
	.w6(32'hbcb2c534),
	.w7(32'h3aecadd3),
	.w8(32'h3b5b77a8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c7f85),
	.w1(32'h3c80fa16),
	.w2(32'hbbe652bc),
	.w3(32'h3a9499a5),
	.w4(32'hbc19dbd4),
	.w5(32'h3c853e19),
	.w6(32'h3ac848a0),
	.w7(32'hbc3522a5),
	.w8(32'h3c517962),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb7896),
	.w1(32'h3b5f7177),
	.w2(32'hbc24b5ac),
	.w3(32'h3ae3ff13),
	.w4(32'hbc0188fa),
	.w5(32'hbbacb375),
	.w6(32'hb9cdafda),
	.w7(32'hbc58ec34),
	.w8(32'hbc19e1f5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25ecbb),
	.w1(32'h39df0aa2),
	.w2(32'h3ba874f5),
	.w3(32'hbb0f1f4e),
	.w4(32'h3b4f8a84),
	.w5(32'hbb5e69b5),
	.w6(32'hb983fb78),
	.w7(32'h3c9c0a9a),
	.w8(32'hbc55596a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5dfddc),
	.w1(32'h3b4d21ac),
	.w2(32'h3c2c4c9b),
	.w3(32'hbb1760f2),
	.w4(32'h3ae60392),
	.w5(32'h3ba637ca),
	.w6(32'h3c0ef0f8),
	.w7(32'h3c840975),
	.w8(32'h3cd94366),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c198704),
	.w1(32'h3a98b2a8),
	.w2(32'hbc8bd797),
	.w3(32'hbc3df8d1),
	.w4(32'hbcb6fed6),
	.w5(32'hbc8e8dba),
	.w6(32'h3babd590),
	.w7(32'hbc5fef90),
	.w8(32'hbcbb640b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c7841),
	.w1(32'h3c0cdd4d),
	.w2(32'h3c041d8a),
	.w3(32'h3ba139a4),
	.w4(32'h3c0c393e),
	.w5(32'h3c848270),
	.w6(32'h3c0da473),
	.w7(32'h3c9b78e3),
	.w8(32'h3d148bed),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae96ae),
	.w1(32'hbc24671a),
	.w2(32'hbd021b5a),
	.w3(32'hbc93f6e8),
	.w4(32'hbd1b7942),
	.w5(32'h3c2a2b41),
	.w6(32'h3aff6b53),
	.w7(32'hbd0a35e2),
	.w8(32'h3bb68a1d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd272e1),
	.w1(32'hbc7187ff),
	.w2(32'hbbefee3a),
	.w3(32'h3bc18d9a),
	.w4(32'hbbfeee6e),
	.w5(32'h3c80f97b),
	.w6(32'hbbd31a72),
	.w7(32'hbc38e8eb),
	.w8(32'h3cfcd0e1),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc28d91),
	.w1(32'hbbff39f9),
	.w2(32'hbcdc2cc6),
	.w3(32'hbc625c17),
	.w4(32'hbc8f6564),
	.w5(32'h3c319ac9),
	.w6(32'hbc7b2ea1),
	.w7(32'hbd07db59),
	.w8(32'h3ca378ec),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55ec1b),
	.w1(32'hba64abcc),
	.w2(32'hbca3c09b),
	.w3(32'hbbb369b0),
	.w4(32'hbc71c687),
	.w5(32'hbc96832d),
	.w6(32'h3b4d6daf),
	.w7(32'hbc9065cc),
	.w8(32'hbd1155d0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd85129),
	.w1(32'h396ce916),
	.w2(32'h3ccf1514),
	.w3(32'h3c0d28d3),
	.w4(32'h3cc1d897),
	.w5(32'hbbf76d49),
	.w6(32'h3b7008c3),
	.w7(32'h3d1638d8),
	.w8(32'h3bb34ecb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9f966),
	.w1(32'h3b63dc34),
	.w2(32'hbb3f1ee8),
	.w3(32'hbc06b252),
	.w4(32'hbc53ceed),
	.w5(32'h3c685e39),
	.w6(32'h3b103a96),
	.w7(32'hbc6c0576),
	.w8(32'h3cdc3fed),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cf02d),
	.w1(32'hbada55f1),
	.w2(32'hbccc9094),
	.w3(32'hbbce9719),
	.w4(32'hbd09de14),
	.w5(32'h3b2758fb),
	.w6(32'h3c2e6b62),
	.w7(32'hbcc82b51),
	.w8(32'hba603f12),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb904a15),
	.w1(32'hbc717d50),
	.w2(32'h3b899304),
	.w3(32'hbbd65285),
	.w4(32'hbb4330ab),
	.w5(32'h3af18cb9),
	.w6(32'hbbf3fa4f),
	.w7(32'hbbc6e77e),
	.w8(32'hbbdf2741),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a000dc4),
	.w1(32'hbbad827a),
	.w2(32'h3baa31a1),
	.w3(32'h3ba07f32),
	.w4(32'h3bbd8faa),
	.w5(32'h3ba2d7fe),
	.w6(32'h3b100c9e),
	.w7(32'h3c9480ca),
	.w8(32'h3b97d487),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb862623),
	.w1(32'hbbb596b1),
	.w2(32'hbb7f8360),
	.w3(32'h3b5a60ec),
	.w4(32'hba7d0fbc),
	.w5(32'hbb1dbba5),
	.w6(32'h3b25a5bb),
	.w7(32'hbbb25a54),
	.w8(32'hbbe5addb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c2dcf),
	.w1(32'hbb066b5b),
	.w2(32'h3b08a4c9),
	.w3(32'h3b8bcdd7),
	.w4(32'h3c2ff023),
	.w5(32'h3b17ea7f),
	.w6(32'h3b2a82d4),
	.w7(32'h3b263833),
	.w8(32'h3b9ca21f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8b271),
	.w1(32'hba9c04f6),
	.w2(32'hbbb381d2),
	.w3(32'hbc027562),
	.w4(32'h3b37e6a0),
	.w5(32'h3c4e1bce),
	.w6(32'hbc3e7038),
	.w7(32'h39f48fc4),
	.w8(32'h3a8900d2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ac808),
	.w1(32'hbb792e7a),
	.w2(32'hbb118285),
	.w3(32'h3c008d97),
	.w4(32'h3c239254),
	.w5(32'hbc814a34),
	.w6(32'h3b02f664),
	.w7(32'h3b17ff9e),
	.w8(32'hbcd296f5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95dbae),
	.w1(32'h3b09b6ae),
	.w2(32'h3ccd2520),
	.w3(32'h3b916bd3),
	.w4(32'h3cb1acb5),
	.w5(32'hbbca1afe),
	.w6(32'hbb150099),
	.w7(32'h3cf9a3cf),
	.w8(32'hbc80fe20),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48bfe6),
	.w1(32'hbc3eaa00),
	.w2(32'hbbbc966d),
	.w3(32'hbbf901b0),
	.w4(32'h3b363b8e),
	.w5(32'hbc2e4e6d),
	.w6(32'hbc10bd51),
	.w7(32'hbb7bd5db),
	.w8(32'hbc1e7a38),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac08801),
	.w1(32'hbba74759),
	.w2(32'h3b8c6ce7),
	.w3(32'hbbbbaba4),
	.w4(32'h3b8ce1d5),
	.w5(32'h3addc108),
	.w6(32'h3ae3de63),
	.w7(32'h3c144c7e),
	.w8(32'h3bb8931f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb636299),
	.w1(32'hbcc4e1a9),
	.w2(32'hbc60c44a),
	.w3(32'hbc20665c),
	.w4(32'h3b8ca7a6),
	.w5(32'hbbce8efc),
	.w6(32'hbc8281c0),
	.w7(32'hba2bc3af),
	.w8(32'hbb3a8d88),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be82fae),
	.w1(32'hbc440a03),
	.w2(32'hbbf42638),
	.w3(32'hbb95b4df),
	.w4(32'h3bc58282),
	.w5(32'h3a5b050f),
	.w6(32'hbbd26e80),
	.w7(32'h3b8a7cad),
	.w8(32'h3bcc5a11),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea729e),
	.w1(32'hbc40d6b1),
	.w2(32'hbcadcc85),
	.w3(32'hbcacb567),
	.w4(32'hbccda4ba),
	.w5(32'hba12d049),
	.w6(32'hbc671c50),
	.w7(32'hbcbbdcd0),
	.w8(32'hbc0d85cf),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda50ae),
	.w1(32'h3ba16c7e),
	.w2(32'h3aac6932),
	.w3(32'h3b9c8ade),
	.w4(32'h3c2234ac),
	.w5(32'h3b009ab0),
	.w6(32'hbaecc566),
	.w7(32'h3b8ce5cb),
	.w8(32'h3c8fa6e2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cafea5f),
	.w1(32'h3c37f896),
	.w2(32'hbc9c310b),
	.w3(32'h3bcbf6c1),
	.w4(32'h3bd55f37),
	.w5(32'h3c44fe2b),
	.w6(32'h3aa1233a),
	.w7(32'hbc854c75),
	.w8(32'h3d150825),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf736a),
	.w1(32'h3abf33be),
	.w2(32'hbcd06ca5),
	.w3(32'h36866f9e),
	.w4(32'hbc3458fc),
	.w5(32'h3ac81229),
	.w6(32'h3c21453b),
	.w7(32'hbd01bb54),
	.w8(32'hbc50dcff),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0750d),
	.w1(32'hbc6cfd39),
	.w2(32'h3bb7306b),
	.w3(32'hbc6f2489),
	.w4(32'hbb25b920),
	.w5(32'h3a5302bc),
	.w6(32'hbb280aec),
	.w7(32'hbb2e74d6),
	.w8(32'h39b96713),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e821d),
	.w1(32'hbab5a92f),
	.w2(32'h3a08f8f3),
	.w3(32'hb9bc2759),
	.w4(32'h3b2ad77c),
	.w5(32'h38fc506e),
	.w6(32'h3a223edb),
	.w7(32'hba902121),
	.w8(32'hbb45c8d3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7edddd),
	.w1(32'hbc4bcc32),
	.w2(32'hbbfe7993),
	.w3(32'hba4add1f),
	.w4(32'hbc1d0f01),
	.w5(32'hbbae6783),
	.w6(32'hbb5670e0),
	.w7(32'hbb90cb04),
	.w8(32'hbb3d0350),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe5ac6),
	.w1(32'h3a84b2fa),
	.w2(32'hbb8a9a3d),
	.w3(32'h3ae61737),
	.w4(32'h3b9d4987),
	.w5(32'hbb9f0750),
	.w6(32'hba784b03),
	.w7(32'h3c1839cd),
	.w8(32'h3bb03220),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8119a1),
	.w1(32'h3b63d1b3),
	.w2(32'h3add52da),
	.w3(32'h3b117b8d),
	.w4(32'h3baff756),
	.w5(32'h3b70dcca),
	.w6(32'hba974b88),
	.w7(32'h3b2d5c3c),
	.w8(32'h3b943ca3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb508593),
	.w1(32'hbbf702e2),
	.w2(32'hbbc29846),
	.w3(32'hba238e70),
	.w4(32'hbb7407b7),
	.w5(32'hbb84541e),
	.w6(32'h3af1ac63),
	.w7(32'h3a83dd55),
	.w8(32'hbb3c2bb1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1b312),
	.w1(32'h3ac28317),
	.w2(32'h386deb21),
	.w3(32'hba18cb03),
	.w4(32'h3b164fab),
	.w5(32'h3ab70b8c),
	.w6(32'h39951436),
	.w7(32'h3b0520c5),
	.w8(32'h3aafccbf),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce4f34),
	.w1(32'hbc92f189),
	.w2(32'hbc840f38),
	.w3(32'hbbfa84b8),
	.w4(32'hbc5d1606),
	.w5(32'hbc17b42d),
	.w6(32'hbbbd37c3),
	.w7(32'hbc1c3394),
	.w8(32'hbbcc3e8b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b702152),
	.w1(32'hb9f07ba1),
	.w2(32'h3a69d466),
	.w3(32'h3b984ad6),
	.w4(32'h3a90aec3),
	.w5(32'hb98bd8d4),
	.w6(32'h3b7b89fb),
	.w7(32'h3a72fd5d),
	.w8(32'h3ae02e8a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08993a),
	.w1(32'hb81238ba),
	.w2(32'hb9abd0af),
	.w3(32'h3a4e4faf),
	.w4(32'h395980ed),
	.w5(32'hba253da9),
	.w6(32'h39ca51d9),
	.w7(32'hb9730783),
	.w8(32'hba1d7e2c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba203796),
	.w1(32'h38796924),
	.w2(32'hb9ef7fad),
	.w3(32'hba413cab),
	.w4(32'h3a2880f3),
	.w5(32'hb804bd85),
	.w6(32'hba9dedd7),
	.w7(32'hb867e98e),
	.w8(32'hb9448fea),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8df03b),
	.w1(32'h3b224740),
	.w2(32'h3a8d3069),
	.w3(32'h39fa4e27),
	.w4(32'h3b31bc62),
	.w5(32'h3b2b1b80),
	.w6(32'h3b07b4c1),
	.w7(32'h3b0f688f),
	.w8(32'h3b1a3021),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84034a),
	.w1(32'h3ba04b42),
	.w2(32'h3a7b50d4),
	.w3(32'h3b8e5f0d),
	.w4(32'h3be753c0),
	.w5(32'h3b92485f),
	.w6(32'h3b63df39),
	.w7(32'h3b80babf),
	.w8(32'h3b531f27),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab94b4b),
	.w1(32'hb945f4a5),
	.w2(32'hbb60cdda),
	.w3(32'hbad8d2a8),
	.w4(32'h39d1d914),
	.w5(32'hba43d626),
	.w6(32'hbab960a3),
	.w7(32'hb99dde7d),
	.w8(32'h39b2d812),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a7758),
	.w1(32'hba3a768e),
	.w2(32'hb989af5a),
	.w3(32'hbb83c503),
	.w4(32'hbb59ba61),
	.w5(32'hba01a864),
	.w6(32'hbb5d40d0),
	.w7(32'hbb460eab),
	.w8(32'hba585406),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01f0e7),
	.w1(32'h3adc23b2),
	.w2(32'h3b6cbff7),
	.w3(32'h3ac6417d),
	.w4(32'h3b1dc9e4),
	.w5(32'h3b0cab48),
	.w6(32'h39e4156a),
	.w7(32'h3b3e09c1),
	.w8(32'h3b8a1207),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb512015),
	.w1(32'hba911974),
	.w2(32'hba707435),
	.w3(32'hbb959be1),
	.w4(32'hbae13726),
	.w5(32'hb9cc8466),
	.w6(32'hbb93868b),
	.w7(32'hbad69fb7),
	.w8(32'h3a97f2e8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b651d),
	.w1(32'hb8d07029),
	.w2(32'hb8114b2d),
	.w3(32'h39b63efc),
	.w4(32'h3a54355e),
	.w5(32'h3a44e695),
	.w6(32'h39ed2902),
	.w7(32'h39b69baa),
	.w8(32'h3a7cd93c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9828664),
	.w1(32'hb92aff25),
	.w2(32'hb9194963),
	.w3(32'hb99ac315),
	.w4(32'hb94d01e9),
	.w5(32'hb954f982),
	.w6(32'hb99aea3f),
	.w7(32'hb9994cb1),
	.w8(32'hb8f37485),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3853d349),
	.w1(32'h38f15b1f),
	.w2(32'hb8cf8edb),
	.w3(32'hb8d6b783),
	.w4(32'hb6b7405f),
	.w5(32'h389a054b),
	.w6(32'hb852a0a2),
	.w7(32'h39129c10),
	.w8(32'h39460e91),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374bea2e),
	.w1(32'hb7644705),
	.w2(32'h38181475),
	.w3(32'hb771b764),
	.w4(32'hb7677366),
	.w5(32'h3398e57c),
	.w6(32'h37e2fc08),
	.w7(32'h380116d6),
	.w8(32'h37db0779),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b335996),
	.w1(32'h3b1c1bf5),
	.w2(32'h3b6a8517),
	.w3(32'h3b31526e),
	.w4(32'h3b3a62c3),
	.w5(32'h3b2cd2dd),
	.w6(32'h3a864af7),
	.w7(32'h3a89c6dc),
	.w8(32'h3ac7f804),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e9c5c),
	.w1(32'h3b6ba0f5),
	.w2(32'h3b56d9f6),
	.w3(32'h3af9d5ff),
	.w4(32'h3b64b961),
	.w5(32'h3b7308fb),
	.w6(32'h39a06cd2),
	.w7(32'h3b19eca8),
	.w8(32'h3ba0088b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba238348),
	.w1(32'hba5a8b3e),
	.w2(32'hba9ee577),
	.w3(32'h394bbfd2),
	.w4(32'h3a41fce7),
	.w5(32'hba58308b),
	.w6(32'h3a9681e5),
	.w7(32'h3a95f692),
	.w8(32'h39888884),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec81f1),
	.w1(32'hbb2e498c),
	.w2(32'hba33427a),
	.w3(32'hb9985dee),
	.w4(32'hba19085e),
	.w5(32'h3a643e48),
	.w6(32'hb816d509),
	.w7(32'h3a26a0f5),
	.w8(32'h3a05ac06),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b173773),
	.w1(32'h3ba9c1f6),
	.w2(32'h3b142eff),
	.w3(32'h3b1b8e58),
	.w4(32'h3b395f3a),
	.w5(32'h3828afb9),
	.w6(32'h39ad8587),
	.w7(32'h3a0b120f),
	.w8(32'hba397bf3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962453a),
	.w1(32'h3921f714),
	.w2(32'h3852f578),
	.w3(32'h39228c93),
	.w4(32'h35cb97da),
	.w5(32'hb9892a88),
	.w6(32'h38a83b86),
	.w7(32'h37941723),
	.w8(32'hb88f21c4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373b88b8),
	.w1(32'hb8b524c2),
	.w2(32'hb99a7c55),
	.w3(32'h39daf565),
	.w4(32'h38a2a9f5),
	.w5(32'hb9efafb0),
	.w6(32'h39ecc020),
	.w7(32'h39322250),
	.w8(32'hb9fd446b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c0eff3),
	.w1(32'h38482965),
	.w2(32'h388c95fb),
	.w3(32'h3845fc91),
	.w4(32'h3889eb67),
	.w5(32'h38c0f3c4),
	.w6(32'h38051614),
	.w7(32'h38b8b66b),
	.w8(32'h389217b3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e268f),
	.w1(32'h3a5f0137),
	.w2(32'h3a0aa087),
	.w3(32'h3ab7d1ed),
	.w4(32'h3aac7ba8),
	.w5(32'h3a084dfb),
	.w6(32'h3aa187c2),
	.w7(32'h3a9994d4),
	.w8(32'h3a00cd28),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36b0ee),
	.w1(32'hbacac63e),
	.w2(32'h3b254496),
	.w3(32'h3b6ef180),
	.w4(32'h3a48b8c2),
	.w5(32'hb9e01369),
	.w6(32'hbad38dac),
	.w7(32'h3a6a822f),
	.w8(32'h3b08ec18),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35ebfb),
	.w1(32'hbae7916f),
	.w2(32'hb957268a),
	.w3(32'hbb445a26),
	.w4(32'hba09cb98),
	.w5(32'h3b158fc9),
	.w6(32'hbab87389),
	.w7(32'h3aa177d3),
	.w8(32'h3b8de0f1),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c53ea5),
	.w1(32'hba836b99),
	.w2(32'hba6fc4c9),
	.w3(32'hba237910),
	.w4(32'hba8ede89),
	.w5(32'hba39d9dd),
	.w6(32'hb9832983),
	.w7(32'hb933d36d),
	.w8(32'hba0e4609),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b97cd),
	.w1(32'hbab5e4ed),
	.w2(32'h38b26c7e),
	.w3(32'hb9be29de),
	.w4(32'hb99f281c),
	.w5(32'hb8c13a18),
	.w6(32'hba81d303),
	.w7(32'hb9274dcf),
	.w8(32'hba61fb12),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84dc8da),
	.w1(32'h39a7a412),
	.w2(32'h39c67e8b),
	.w3(32'h399202fb),
	.w4(32'h39db46fe),
	.w5(32'h39d19ecd),
	.w6(32'h3997a2d3),
	.w7(32'h390ff2a7),
	.w8(32'h3a226c58),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba018da7),
	.w1(32'h38127d0b),
	.w2(32'h399d4852),
	.w3(32'hba74338c),
	.w4(32'h38b81afd),
	.w5(32'h3a952f54),
	.w6(32'hb9988809),
	.w7(32'h39c19e93),
	.w8(32'h3a857318),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d78e1),
	.w1(32'h3aeb855c),
	.w2(32'h3ac2fe08),
	.w3(32'hbb4f09e4),
	.w4(32'h39af4129),
	.w5(32'h3b265a2d),
	.w6(32'hbb27b905),
	.w7(32'hb9aa28b8),
	.w8(32'h3a4804ef),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c8b25),
	.w1(32'hbbdf1c47),
	.w2(32'hbb9154a3),
	.w3(32'hbb7dcc9f),
	.w4(32'hbbb3bc03),
	.w5(32'hbb20951c),
	.w6(32'hbb2056cf),
	.w7(32'hbb13a8e0),
	.w8(32'hbb398d20),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a307b63),
	.w1(32'h3a86d26a),
	.w2(32'hb9a3e525),
	.w3(32'hb9b490af),
	.w4(32'h39970074),
	.w5(32'h39d1943c),
	.w6(32'hba18101e),
	.w7(32'hba70a6b3),
	.w8(32'h3aa7f524),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03dd82),
	.w1(32'h38b855f7),
	.w2(32'hb98a75ea),
	.w3(32'hba7e17dc),
	.w4(32'h39aec611),
	.w5(32'hb79fa644),
	.w6(32'hbb31caf4),
	.w7(32'hbabe1594),
	.w8(32'hb96ab43c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb56ef5),
	.w1(32'hbbbdfca5),
	.w2(32'hbb82ba7f),
	.w3(32'hbb56e019),
	.w4(32'hbb9c8f7e),
	.w5(32'hbb10751b),
	.w6(32'h37cddf3e),
	.w7(32'h3aa4f6fb),
	.w8(32'hbb27fe19),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a273134),
	.w1(32'h3a4884d9),
	.w2(32'hb9dbe8e6),
	.w3(32'h3ae40fe5),
	.w4(32'h3ac52904),
	.w5(32'hba390a19),
	.w6(32'hb9c279be),
	.w7(32'h3ab07e93),
	.w8(32'h3acf450f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35ee49),
	.w1(32'hba83b7a3),
	.w2(32'h39991b6b),
	.w3(32'hbb081d6d),
	.w4(32'hba37e968),
	.w5(32'h3adc849b),
	.w6(32'hba5d95ac),
	.w7(32'h3961ea4f),
	.w8(32'h3ae88ab1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d0525),
	.w1(32'hb8b7665f),
	.w2(32'hb96f2c9f),
	.w3(32'hb9920314),
	.w4(32'h3979ccd8),
	.w5(32'h39bd100e),
	.w6(32'hb9a0336b),
	.w7(32'h38cce355),
	.w8(32'h39df6b7c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba327ee),
	.w1(32'h3b47514f),
	.w2(32'hb9700723),
	.w3(32'h3bae1093),
	.w4(32'h3b44df95),
	.w5(32'hbaff8c43),
	.w6(32'h3b334a3f),
	.w7(32'h3b1ecfbe),
	.w8(32'hba1ce747),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb092742),
	.w1(32'hba90af07),
	.w2(32'hba3f9cf1),
	.w3(32'hbb301fc4),
	.w4(32'hb9ec1edc),
	.w5(32'h3a005c83),
	.w6(32'hbb3ce565),
	.w7(32'hba93e0c6),
	.w8(32'h3a5ac2c5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79ce0ae),
	.w1(32'hb89a391d),
	.w2(32'hb7d53acd),
	.w3(32'hb614ecb2),
	.w4(32'hb7412467),
	.w5(32'hb7c36d0a),
	.w6(32'h383a1b11),
	.w7(32'h38b6d639),
	.w8(32'h388b5601),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c9dd14),
	.w1(32'hb816cea5),
	.w2(32'h37d0ae1b),
	.w3(32'h37e258f9),
	.w4(32'hb6201fef),
	.w5(32'hb7e1c0e1),
	.w6(32'h38172d85),
	.w7(32'h3538a394),
	.w8(32'h3808b6fe),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39367ff2),
	.w1(32'h39e69c03),
	.w2(32'h3a2b27b5),
	.w3(32'h3a3d9623),
	.w4(32'h39bf2620),
	.w5(32'h3996c2f9),
	.w6(32'h3a19994f),
	.w7(32'h3a07646d),
	.w8(32'h3a81c19b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4fe95),
	.w1(32'h3aba8aa3),
	.w2(32'hbaeff781),
	.w3(32'h3a22ae30),
	.w4(32'hb8c7bc71),
	.w5(32'hba23c570),
	.w6(32'hbb4dc7b9),
	.w7(32'hbb0c824b),
	.w8(32'h39dfe688),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f81ff),
	.w1(32'hb9b5c4b0),
	.w2(32'h3a9ca47d),
	.w3(32'hba9227d8),
	.w4(32'hb8792ce1),
	.w5(32'h3b1ccb21),
	.w6(32'h3a23dea6),
	.w7(32'h38caf0a6),
	.w8(32'h3b0a2232),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb878b8d7),
	.w1(32'hb800b72f),
	.w2(32'h356010cc),
	.w3(32'hb8327af5),
	.w4(32'hb8181abc),
	.w5(32'hb7107768),
	.w6(32'hb79eb8f9),
	.w7(32'hb810fe9e),
	.w8(32'hb7a7fd45),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9392ad),
	.w1(32'hba8cb642),
	.w2(32'hba07f86f),
	.w3(32'hbb15c4f7),
	.w4(32'hb8bde2ef),
	.w5(32'h3b159632),
	.w6(32'hba4001a3),
	.w7(32'hba84ab84),
	.w8(32'h3b1e8704),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58619e),
	.w1(32'h3a6fd61b),
	.w2(32'h37f7489d),
	.w3(32'h3b61edba),
	.w4(32'h3b2355a6),
	.w5(32'h3a71d55a),
	.w6(32'hb91ad6df),
	.w7(32'hbb02556d),
	.w8(32'h3a85694e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a7f7),
	.w1(32'hbba98297),
	.w2(32'hbbb1a0d3),
	.w3(32'h3acaf995),
	.w4(32'hbadcb92a),
	.w5(32'hbb2e8e0e),
	.w6(32'h39c9988a),
	.w7(32'hb580f45e),
	.w8(32'hbb36d904),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5f9af),
	.w1(32'h3b68ead3),
	.w2(32'h3a6b7882),
	.w3(32'h3b148b17),
	.w4(32'h3b7733d9),
	.w5(32'h3b1cbac1),
	.w6(32'h39bb6673),
	.w7(32'h397543c6),
	.w8(32'h3a00e324),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c77d48),
	.w1(32'h3a25fd83),
	.w2(32'h395bdc14),
	.w3(32'hba74175a),
	.w4(32'hb9f6b91d),
	.w5(32'hba55cb5b),
	.w6(32'hba3ddad6),
	.w7(32'hb9c3ad14),
	.w8(32'hbae239e7),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a613d83),
	.w1(32'h3a3dbf30),
	.w2(32'hb9c88115),
	.w3(32'h3b0173c4),
	.w4(32'h3ae621a3),
	.w5(32'h3aa59f2d),
	.w6(32'h3b0b1d47),
	.w7(32'h3b1f166f),
	.w8(32'h3a6a0b82),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959c5c9),
	.w1(32'h3a6539a6),
	.w2(32'hb99bc511),
	.w3(32'h390791e2),
	.w4(32'h3afc5706),
	.w5(32'h3a097559),
	.w6(32'hba718782),
	.w7(32'h3abb4d4c),
	.w8(32'h3a9d8d12),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7dea6),
	.w1(32'h39935b3f),
	.w2(32'h3adb7de6),
	.w3(32'hb9cf95a9),
	.w4(32'hb9c98dca),
	.w5(32'hba23e9cb),
	.w6(32'hbb7cc13c),
	.w7(32'hbb8338a6),
	.w8(32'hb92ba69d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44eb0c),
	.w1(32'h3b6a0a7a),
	.w2(32'h3b2056ba),
	.w3(32'h3b339c53),
	.w4(32'h3b49b89f),
	.w5(32'h3b03d35a),
	.w6(32'h3aca64ed),
	.w7(32'h3a9546b2),
	.w8(32'h3a4b312f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a3c05),
	.w1(32'hbad90967),
	.w2(32'hba48699c),
	.w3(32'hba6eb3e3),
	.w4(32'hbac0c0f9),
	.w5(32'hba0557de),
	.w6(32'hb926e7eb),
	.w7(32'hb93989de),
	.w8(32'hb9faee04),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392e80d0),
	.w1(32'h392fa12b),
	.w2(32'h38684574),
	.w3(32'h396913e0),
	.w4(32'h39f7b6fb),
	.w5(32'h3980cd82),
	.w6(32'h39a82449),
	.w7(32'h39676221),
	.w8(32'h38e6c672),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe0fa7),
	.w1(32'hbb20f536),
	.w2(32'h3a12626e),
	.w3(32'hbb1cf810),
	.w4(32'hba1965a3),
	.w5(32'h3b1ac5c2),
	.w6(32'hbb12f162),
	.w7(32'hb9039687),
	.w8(32'h3afb988d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d12e25),
	.w1(32'h372f04e6),
	.w2(32'h3908cbe6),
	.w3(32'h3a46b2d7),
	.w4(32'h39fee6fd),
	.w5(32'h384a69eb),
	.w6(32'h39fce605),
	.w7(32'h39831ad7),
	.w8(32'h38ef199c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8014ee7),
	.w1(32'h3abc8857),
	.w2(32'h3abeee31),
	.w3(32'hba2079ba),
	.w4(32'h3aee43f3),
	.w5(32'h3ad0de14),
	.w6(32'hbacb546d),
	.w7(32'h390a74e0),
	.w8(32'h3b04fc78),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394298e8),
	.w1(32'hb8df115d),
	.w2(32'hb9d069dc),
	.w3(32'h39d7446c),
	.w4(32'h394720e1),
	.w5(32'hba30f056),
	.w6(32'h38c901fb),
	.w7(32'h397c1d8e),
	.w8(32'hb9c4022e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c027b13),
	.w1(32'h3b1d213f),
	.w2(32'h3b361ef3),
	.w3(32'h3c00cb77),
	.w4(32'h3aee69ef),
	.w5(32'h3abc4674),
	.w6(32'h3bc883d4),
	.w7(32'hb93d9d73),
	.w8(32'hb9ffbdaf),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e9a4dd),
	.w1(32'hb8106743),
	.w2(32'h38176be8),
	.w3(32'h36c6eb26),
	.w4(32'hb942693f),
	.w5(32'h381fecbb),
	.w6(32'h36f5bb7e),
	.w7(32'h39435c30),
	.w8(32'h3908efbd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bfe291),
	.w1(32'hba2a3440),
	.w2(32'hba303316),
	.w3(32'h39929748),
	.w4(32'hba1161cd),
	.w5(32'hba573e81),
	.w6(32'hb94ca697),
	.w7(32'hba13b9bb),
	.w8(32'hba6ca940),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa64eb7),
	.w1(32'hb9c3882e),
	.w2(32'hba9323c1),
	.w3(32'hbb0b5dd4),
	.w4(32'hb9e5454a),
	.w5(32'h3ab94547),
	.w6(32'hbaa467dc),
	.w7(32'hba17ff81),
	.w8(32'h3b2f2053),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b97a46),
	.w1(32'hbb2645d4),
	.w2(32'hbabaf5b9),
	.w3(32'hbab6a9eb),
	.w4(32'hb90ac3b7),
	.w5(32'h38df3240),
	.w6(32'hbc16168d),
	.w7(32'hba95acbd),
	.w8(32'h3b3fdb16),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae53e6e),
	.w1(32'h3ac377e8),
	.w2(32'h3a47b20f),
	.w3(32'h3b31060b),
	.w4(32'h3ab067d4),
	.w5(32'hb98b7a7e),
	.w6(32'h3b37d088),
	.w7(32'h3b153547),
	.w8(32'h37e7e014),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72a6fb),
	.w1(32'hbb5e19d9),
	.w2(32'hbbccd77d),
	.w3(32'hb9db94c2),
	.w4(32'hbb79a186),
	.w5(32'hbbafe795),
	.w6(32'h3a6ccf26),
	.w7(32'hbb1d6554),
	.w8(32'hbb5ab0a6),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9269f),
	.w1(32'h3a5296d8),
	.w2(32'hb9cadcc0),
	.w3(32'hb87cfdff),
	.w4(32'h39e358d2),
	.w5(32'hb98a50fe),
	.w6(32'hb8afe833),
	.w7(32'hb9163b99),
	.w8(32'hb9cf864d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4f1e5),
	.w1(32'h3aa6e551),
	.w2(32'h3a87bddf),
	.w3(32'h3af1bda9),
	.w4(32'h3b437a6d),
	.w5(32'h3b272ac1),
	.w6(32'h3b1eca46),
	.w7(32'h3b3fa071),
	.w8(32'h3b326be5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb072171),
	.w1(32'hbb0ab253),
	.w2(32'hbb222674),
	.w3(32'hbaae9dfe),
	.w4(32'hba414fb8),
	.w5(32'hba9928d0),
	.w6(32'hbaa11f8e),
	.w7(32'hba176fea),
	.w8(32'hba85397d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42ba3b),
	.w1(32'hbae16e9a),
	.w2(32'hbadde322),
	.w3(32'hbb8b9c2f),
	.w4(32'hba9baa24),
	.w5(32'h39d3dc4a),
	.w6(32'hbb774715),
	.w7(32'hbb133fa8),
	.w8(32'hb9cfc7cc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c7c4d),
	.w1(32'h3a66c1b5),
	.w2(32'h3a26fb50),
	.w3(32'h3a39660e),
	.w4(32'h3ab42635),
	.w5(32'h3adea92e),
	.w6(32'h3a15dca2),
	.w7(32'h3ae2b8e4),
	.w8(32'h3b10578e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1163eb),
	.w1(32'hba84c5c5),
	.w2(32'h39a525a6),
	.w3(32'hbb4c3341),
	.w4(32'hb9b854e1),
	.w5(32'h3a97dc28),
	.w6(32'hbb1ed890),
	.w7(32'hba041b52),
	.w8(32'h3acb27bf),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f7a923),
	.w1(32'h3747bae4),
	.w2(32'h386ebd86),
	.w3(32'h384a7b36),
	.w4(32'hb6364f51),
	.w5(32'h37ca9cea),
	.w6(32'h38a2f612),
	.w7(32'h37c26770),
	.w8(32'h37f63841),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e0b7c),
	.w1(32'hb91480d5),
	.w2(32'h3a10e018),
	.w3(32'h39e4a7a8),
	.w4(32'h3a20b621),
	.w5(32'h3a5316ff),
	.w6(32'h3a37bbc7),
	.w7(32'h3a416abd),
	.w8(32'h39c7a348),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82409ca),
	.w1(32'h38d850d5),
	.w2(32'h385260e4),
	.w3(32'h38a729cc),
	.w4(32'h39213c9e),
	.w5(32'hb9a0aa51),
	.w6(32'hb94094ca),
	.w7(32'hb874f6eb),
	.w8(32'hb9ae4b82),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd1d15),
	.w1(32'h39c9b773),
	.w2(32'hb9e73cc3),
	.w3(32'hb9eeb631),
	.w4(32'h3a602d71),
	.w5(32'h398575ae),
	.w6(32'hba3589c6),
	.w7(32'hb990e0bd),
	.w8(32'h398515fb),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35db9e2b),
	.w1(32'hb7dd3e6b),
	.w2(32'h38130272),
	.w3(32'hb7b94f4a),
	.w4(32'h37b1bd0b),
	.w5(32'hb0e219de),
	.w6(32'hb7951b17),
	.w7(32'h37e181a9),
	.w8(32'h362a5caa),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1417a),
	.w1(32'hb9ab3ca9),
	.w2(32'hb9832dcc),
	.w3(32'hb8d31a93),
	.w4(32'h388a01a1),
	.w5(32'h38c3393b),
	.w6(32'hb88cbfd8),
	.w7(32'h38e00805),
	.w8(32'hb87d72ed),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ec0a7),
	.w1(32'hb98a6df8),
	.w2(32'h39288703),
	.w3(32'h3a7b0b3d),
	.w4(32'h3ae29aca),
	.w5(32'h3a0d97fd),
	.w6(32'hba837a79),
	.w7(32'h388d8e0e),
	.w8(32'h38e8405b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4eb76),
	.w1(32'hbab2647a),
	.w2(32'hba52872a),
	.w3(32'h3b7a5aba),
	.w4(32'h3b47b435),
	.w5(32'h3b06c848),
	.w6(32'h3b4412bc),
	.w7(32'hb9d0e78f),
	.w8(32'hba7da064),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d6119),
	.w1(32'hbabd7a7f),
	.w2(32'h39aa1af8),
	.w3(32'hba741857),
	.w4(32'hb9b3dd2c),
	.w5(32'h3a1d1b70),
	.w6(32'hb984a9c7),
	.w7(32'h39a1c29c),
	.w8(32'h3a14110f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bb595),
	.w1(32'hbb18cc3a),
	.w2(32'hbb03a2c5),
	.w3(32'hba809686),
	.w4(32'hba94601a),
	.w5(32'hbb29a31d),
	.w6(32'h39ce922b),
	.w7(32'hba14459e),
	.w8(32'hbb103f98),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc10cd8),
	.w1(32'hbbd06689),
	.w2(32'hbb1c9a9a),
	.w3(32'hbb38d72d),
	.w4(32'hba17de6b),
	.w5(32'h3a54b4aa),
	.w6(32'hba107bbe),
	.w7(32'hb85ba91e),
	.w8(32'h3a3c16ac),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb853ebd),
	.w1(32'h3b6efe33),
	.w2(32'hb9ce3814),
	.w3(32'hbac2d2a7),
	.w4(32'h3bb79fc0),
	.w5(32'h3b59dce7),
	.w6(32'hba3095b1),
	.w7(32'h3b065ea8),
	.w8(32'h3b15454b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad9e04),
	.w1(32'h381c2237),
	.w2(32'h3951c77f),
	.w3(32'h3a8c049a),
	.w4(32'h39eb250d),
	.w5(32'h39b9e3cb),
	.w6(32'h3a9ec478),
	.w7(32'h3a417f04),
	.w8(32'h390f1354),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896bb55),
	.w1(32'hb8929e82),
	.w2(32'hb83a2fc5),
	.w3(32'hb80f2d99),
	.w4(32'hb88407ee),
	.w5(32'hb8e87760),
	.w6(32'hb8ba31b2),
	.w7(32'hb8928e99),
	.w8(32'hb8da7dd1),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ccf95),
	.w1(32'hb7dc45a3),
	.w2(32'hb9b65ba6),
	.w3(32'hb923fb83),
	.w4(32'h39a4bb0f),
	.w5(32'hb978dbdc),
	.w6(32'h393eae58),
	.w7(32'h39aa6e08),
	.w8(32'hb99b2210),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a0dedf),
	.w1(32'h383a52b2),
	.w2(32'h38541dc2),
	.w3(32'h385bfdc2),
	.w4(32'hb560bcd2),
	.w5(32'hb6c6c357),
	.w6(32'h3866a4c9),
	.w7(32'h379f501a),
	.w8(32'h38028cc6),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68f16a),
	.w1(32'h38be1feb),
	.w2(32'h3a0acfec),
	.w3(32'h39dd8a08),
	.w4(32'hba1e86f4),
	.w5(32'h3a1f7df8),
	.w6(32'h39efdac5),
	.w7(32'h39e44bb2),
	.w8(32'h39c27bda),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39672f),
	.w1(32'hbb7b850e),
	.w2(32'hbb27250b),
	.w3(32'hba934e97),
	.w4(32'hbb3b4b5b),
	.w5(32'hbb174a14),
	.w6(32'hbb1dfc02),
	.w7(32'hbb1023ec),
	.w8(32'hbb0e3add),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9371fe),
	.w1(32'h3b4b5509),
	.w2(32'h3b318808),
	.w3(32'h3aedb2ea),
	.w4(32'h3b414cc2),
	.w5(32'h3b937bc1),
	.w6(32'h3aa8abab),
	.w7(32'h3b4b0ef1),
	.w8(32'h3bafdafa),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e48002),
	.w1(32'hba7d8027),
	.w2(32'hb9a06f77),
	.w3(32'hb97c14dd),
	.w4(32'h37139998),
	.w5(32'hb9a2786a),
	.w6(32'hb9d8d173),
	.w7(32'h3783a507),
	.w8(32'h39f93d11),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980a860),
	.w1(32'hb994cd5a),
	.w2(32'hbb6529e3),
	.w3(32'h3ab743b2),
	.w4(32'h3996b069),
	.w5(32'hbb1a60e8),
	.w6(32'h3b7996ce),
	.w7(32'h3aa8334c),
	.w8(32'hbaa2271e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa8c06),
	.w1(32'hba60b8ad),
	.w2(32'hb9712c7e),
	.w3(32'h3a999945),
	.w4(32'h39cd3dc5),
	.w5(32'h3a19f1cd),
	.w6(32'h3a810c10),
	.w7(32'h3a83cc18),
	.w8(32'h3aadc9a2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382507e9),
	.w1(32'h388e97d9),
	.w2(32'h39020d20),
	.w3(32'h358098fe),
	.w4(32'h3868025b),
	.w5(32'h38f69929),
	.w6(32'h37639074),
	.w7(32'h387033f9),
	.w8(32'h390911ce),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d04d6),
	.w1(32'hbb0d4fdd),
	.w2(32'hbab4cbce),
	.w3(32'hba6c8308),
	.w4(32'hba14a2fc),
	.w5(32'hb9b0b291),
	.w6(32'hba2d0162),
	.w7(32'h39ae198a),
	.w8(32'h39e54c76),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38378ed7),
	.w1(32'hb787e034),
	.w2(32'h392c09d3),
	.w3(32'h3734b16b),
	.w4(32'hb7945cc7),
	.w5(32'h39035643),
	.w6(32'h38c5a293),
	.w7(32'h385acbbd),
	.w8(32'h394da71b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefe479),
	.w1(32'hbade32c2),
	.w2(32'hba92bcb8),
	.w3(32'hbadb7ba4),
	.w4(32'hb8febfaa),
	.w5(32'hb8d5675c),
	.w6(32'h3a09e648),
	.w7(32'h38d64f07),
	.w8(32'hb8bce83e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba8bf8),
	.w1(32'h3aad1577),
	.w2(32'h3ab42295),
	.w3(32'h3a572330),
	.w4(32'h3b05216f),
	.w5(32'h3b4c4548),
	.w6(32'hba2be127),
	.w7(32'hba89ca46),
	.w8(32'h39d7111a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c6e23),
	.w1(32'h3a4df3f8),
	.w2(32'hbab867fc),
	.w3(32'h3aa27321),
	.w4(32'h3aaf74ca),
	.w5(32'hb97a6dd1),
	.w6(32'h3ab05e43),
	.w7(32'h39ee0188),
	.w8(32'hb8ad6031),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a630d1),
	.w1(32'h39ed9370),
	.w2(32'hba0b64dd),
	.w3(32'h3aaab782),
	.w4(32'h39b68371),
	.w5(32'hba891786),
	.w6(32'h3ab97870),
	.w7(32'h3a323856),
	.w8(32'hba87cb05),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aade8e9),
	.w1(32'h3b26f54d),
	.w2(32'h3982d8a5),
	.w3(32'h3a8ade6c),
	.w4(32'h3a9fdbb7),
	.w5(32'h3abf493f),
	.w6(32'h3aad387b),
	.w7(32'h3a9375cc),
	.w8(32'h3ad76e51),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d0074b),
	.w1(32'hba20997f),
	.w2(32'hba043460),
	.w3(32'hbac25228),
	.w4(32'hb9f37639),
	.w5(32'h3aea2074),
	.w6(32'hbaee0dd9),
	.w7(32'hba39d144),
	.w8(32'h3b21b434),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa924da),
	.w1(32'h376c1c35),
	.w2(32'h3adf86f5),
	.w3(32'hba7ed95c),
	.w4(32'hb944cb7f),
	.w5(32'h3b227307),
	.w6(32'hbaa74d72),
	.w7(32'hb924723e),
	.w8(32'h3b1a255d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38662861),
	.w1(32'h38445e4f),
	.w2(32'h38b99c9b),
	.w3(32'h3892fa31),
	.w4(32'h38a5607d),
	.w5(32'h390061fc),
	.w6(32'h390b3f91),
	.w7(32'h38fa0b87),
	.w8(32'h38f6593a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c3aa66),
	.w1(32'hb7d2a5a1),
	.w2(32'hb7d6eba0),
	.w3(32'hb92df8f3),
	.w4(32'hb9587e79),
	.w5(32'hb8d7852b),
	.w6(32'h38f2a884),
	.w7(32'hb8a20ae1),
	.w8(32'hb89e014f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03390a),
	.w1(32'h3a8955b6),
	.w2(32'h3a7eec6b),
	.w3(32'h3bab5a0a),
	.w4(32'h3b060dcd),
	.w5(32'h3b07face),
	.w6(32'h398e0327),
	.w7(32'h3a838ce4),
	.w8(32'h3ad7dc2f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a8655),
	.w1(32'hbbd53642),
	.w2(32'hbb96e166),
	.w3(32'hbaf80557),
	.w4(32'h3abd3811),
	.w5(32'h3ae3b7a9),
	.w6(32'hbc04a3f1),
	.w7(32'hbb807490),
	.w8(32'hba2ea138),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3386e9),
	.w1(32'h3aaf62e1),
	.w2(32'h3b2b1faf),
	.w3(32'h3a933715),
	.w4(32'h3b33ac50),
	.w5(32'h3b5205b2),
	.w6(32'hba281830),
	.w7(32'h3a806e32),
	.w8(32'h3b3d323b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e99f2),
	.w1(32'hb988aeeb),
	.w2(32'h3aebc5db),
	.w3(32'h3a32bf94),
	.w4(32'h3ad5bbf8),
	.w5(32'h3b552ce4),
	.w6(32'h3b2c589d),
	.w7(32'h39602e2b),
	.w8(32'hba183e7b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d8e94a),
	.w1(32'h397965b2),
	.w2(32'h38bc9c50),
	.w3(32'hb92683f6),
	.w4(32'hb8c6ea15),
	.w5(32'hb940db02),
	.w6(32'hb9b903e4),
	.w7(32'hb92fa966),
	.w8(32'hb8f7b303),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba362be1),
	.w1(32'hba2a945d),
	.w2(32'h393076d2),
	.w3(32'hba6fcf50),
	.w4(32'hba4aa9b0),
	.w5(32'h3a04c83c),
	.w6(32'hba7ed848),
	.w7(32'hb95ab7c7),
	.w8(32'h3a2c52c4),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5cb9d),
	.w1(32'hbac78329),
	.w2(32'hb9b38075),
	.w3(32'h3b8979e8),
	.w4(32'hbaf5fb8d),
	.w5(32'hbae11c59),
	.w6(32'h3a913390),
	.w7(32'h3a84932a),
	.w8(32'hba38591f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde3dde),
	.w1(32'hbc13af3b),
	.w2(32'hbb4b50fb),
	.w3(32'hbbba31ac),
	.w4(32'hbbc2fb49),
	.w5(32'hbab5d7dd),
	.w6(32'hbb1138d8),
	.w7(32'hbb456058),
	.w8(32'hbb1b40e9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01a241),
	.w1(32'hbb5de483),
	.w2(32'hbb3ac7a1),
	.w3(32'h39f5467f),
	.w4(32'hbb82602c),
	.w5(32'hbb186e0a),
	.w6(32'hb9bdcb47),
	.w7(32'h39bc5b9b),
	.w8(32'hb87873b2),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e56c7),
	.w1(32'h3b0fc39e),
	.w2(32'h3a76b44d),
	.w3(32'h3a987be4),
	.w4(32'h3addea2f),
	.w5(32'h3a1fb31a),
	.w6(32'h39884f00),
	.w7(32'h38f71dc7),
	.w8(32'h389543c8),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fd6da),
	.w1(32'h3b236296),
	.w2(32'h3a407ab3),
	.w3(32'hbaabecad),
	.w4(32'h3b177da1),
	.w5(32'h3afba460),
	.w6(32'hbb06ffd3),
	.w7(32'hba64a8fd),
	.w8(32'h3a9c26a7),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3809d9b7),
	.w1(32'h381f5d3b),
	.w2(32'h388654a6),
	.w3(32'h37f9ba94),
	.w4(32'h37f86279),
	.w5(32'h3835b392),
	.w6(32'h3833b939),
	.w7(32'h380df30b),
	.w8(32'h3815e372),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381ecd71),
	.w1(32'h381f30d0),
	.w2(32'h38859c8f),
	.w3(32'h37fc9710),
	.w4(32'h37826025),
	.w5(32'h38135a2e),
	.w6(32'h376d0c83),
	.w7(32'h37364dca),
	.w8(32'h384ca2e7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e42167),
	.w1(32'h3a4cc064),
	.w2(32'h3a5abe68),
	.w3(32'hb8f69a9f),
	.w4(32'h38026e2f),
	.w5(32'hb9c18c43),
	.w6(32'hb8e44a78),
	.w7(32'hb9486118),
	.w8(32'hb9731396),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e9c3a4),
	.w1(32'hb7322d62),
	.w2(32'h37117935),
	.w3(32'hb8075f3c),
	.w4(32'hb80f3186),
	.w5(32'h3b1a5299),
	.w6(32'h37944275),
	.w7(32'hb78edf9e),
	.w8(32'hb905425d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cad967),
	.w1(32'hbadfeb72),
	.w2(32'hba045f1a),
	.w3(32'h3b2efb59),
	.w4(32'h3b5c2465),
	.w5(32'hbbbbf393),
	.w6(32'h3ac3a43f),
	.w7(32'h3a87254f),
	.w8(32'hbb0cd412),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80cc93),
	.w1(32'hbbd7787c),
	.w2(32'hbbd2e8f6),
	.w3(32'hbc600add),
	.w4(32'hbb8b1af2),
	.w5(32'h3aa583f2),
	.w6(32'hbc0aceb7),
	.w7(32'hbc547f83),
	.w8(32'hbb4db479),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae0e66),
	.w1(32'hbbaa7874),
	.w2(32'hbb3d4d5c),
	.w3(32'h3aaa5d4a),
	.w4(32'h3b759095),
	.w5(32'h3c1e355f),
	.w6(32'hbb2b1f6c),
	.w7(32'hbb59ff5f),
	.w8(32'h39591a1a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fcd55),
	.w1(32'hbbd56086),
	.w2(32'hbb2169b2),
	.w3(32'h3c35d995),
	.w4(32'hbb170d8b),
	.w5(32'hb986bbf8),
	.w6(32'hbb8d3e47),
	.w7(32'h3a80c218),
	.w8(32'hba54ff79),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ecefe),
	.w1(32'hbbed9637),
	.w2(32'hbaf09a86),
	.w3(32'hbad60a9b),
	.w4(32'hbb454d5c),
	.w5(32'hbb999297),
	.w6(32'h3a470e4a),
	.w7(32'h3abf24a6),
	.w8(32'hbb06305b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca5ef),
	.w1(32'hbb25f280),
	.w2(32'hbb3e9b8d),
	.w3(32'hbb259b30),
	.w4(32'hbb362c7c),
	.w5(32'hbaabf79d),
	.w6(32'h3a2f3813),
	.w7(32'hbb0279e7),
	.w8(32'h395785ee),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1109d),
	.w1(32'h3ad8b910),
	.w2(32'h3b5d206c),
	.w3(32'h3b1af5c5),
	.w4(32'h3b58fbad),
	.w5(32'hbbfd0f60),
	.w6(32'hbbbb7333),
	.w7(32'hb9a419ec),
	.w8(32'hbadb1db7),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb770034),
	.w1(32'h3c1af3fa),
	.w2(32'h3a95ad53),
	.w3(32'hbc2f9baa),
	.w4(32'hbc243bda),
	.w5(32'hbb41da42),
	.w6(32'h3a92ba09),
	.w7(32'hbba18e13),
	.w8(32'hbc21d6af),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb825a02),
	.w1(32'hbabf5f95),
	.w2(32'h3a8ed697),
	.w3(32'hbb16411c),
	.w4(32'hbae100e7),
	.w5(32'hbb10308f),
	.w6(32'hbb3734ce),
	.w7(32'hbb087276),
	.w8(32'h389708f1),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60646bb),
	.w1(32'h3afe686c),
	.w2(32'hbb36b07f),
	.w3(32'hbaf7a8f0),
	.w4(32'h3b8e43ff),
	.w5(32'h3bb1cbbc),
	.w6(32'h3b0dcd5c),
	.w7(32'hbad505dd),
	.w8(32'h3a7374ac),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb200288),
	.w1(32'hbb733df9),
	.w2(32'hbae44c0c),
	.w3(32'h3b5a5ea4),
	.w4(32'h3ba9e435),
	.w5(32'h3b206bf2),
	.w6(32'h39c53827),
	.w7(32'h395ad34d),
	.w8(32'h3adfefc5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf449b3),
	.w1(32'hbae54c03),
	.w2(32'hbb8e232e),
	.w3(32'h3afcfb21),
	.w4(32'h3b0c2f72),
	.w5(32'h3b2f9cca),
	.w6(32'h38ed67d5),
	.w7(32'hbb2dab75),
	.w8(32'hbad66082),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58f9c2),
	.w1(32'hba948436),
	.w2(32'h3ab6d063),
	.w3(32'hbb5cf25a),
	.w4(32'hbbf883d8),
	.w5(32'h3a9c751b),
	.w6(32'h3b475c91),
	.w7(32'hbb6712b5),
	.w8(32'hb86151a3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0129b6),
	.w1(32'hbba99a34),
	.w2(32'hbbcb3259),
	.w3(32'hbb8f7799),
	.w4(32'h3ad75343),
	.w5(32'h3bd285ff),
	.w6(32'hbb8040ec),
	.w7(32'hbb85b764),
	.w8(32'h3bbb4f6e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc058ae0),
	.w1(32'hbbbe1402),
	.w2(32'hbb51cae0),
	.w3(32'hbb9589ae),
	.w4(32'hbb3edaab),
	.w5(32'h3aabce38),
	.w6(32'h3a51025f),
	.w7(32'h3b53bcf5),
	.w8(32'hb86c2a58),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8f135),
	.w1(32'h39f00bc9),
	.w2(32'h3b7acff4),
	.w3(32'hbbb9e3f1),
	.w4(32'hbae90c5d),
	.w5(32'hbb44f78a),
	.w6(32'hba9da61e),
	.w7(32'hba31c2bc),
	.w8(32'hbba1b31c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39572f05),
	.w1(32'h3aa1a3bc),
	.w2(32'hbba9b973),
	.w3(32'h3b9f034f),
	.w4(32'h3c338b73),
	.w5(32'h3bb2ee40),
	.w6(32'hbb2f30d3),
	.w7(32'hba9b71f2),
	.w8(32'h3bb93f5a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34485d),
	.w1(32'hbba8e49a),
	.w2(32'hbbc09626),
	.w3(32'h3b855ff1),
	.w4(32'hbaaeca28),
	.w5(32'h3a6a449a),
	.w6(32'hbab3a80b),
	.w7(32'hbb79d64c),
	.w8(32'h3b237370),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22eeac),
	.w1(32'hba536fc4),
	.w2(32'h3a3253bd),
	.w3(32'h3950b3ec),
	.w4(32'hbb1a3f15),
	.w5(32'hbb877832),
	.w6(32'hb9e52366),
	.w7(32'hbaceec33),
	.w8(32'hbba90d0a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9f8f1),
	.w1(32'hbbf4daea),
	.w2(32'hbb30518b),
	.w3(32'h3aa0705d),
	.w4(32'hbb23ca09),
	.w5(32'h3a319829),
	.w6(32'hbb9cdd63),
	.w7(32'h3be5627a),
	.w8(32'h3aa31218),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb882d06),
	.w1(32'hbb3229e6),
	.w2(32'hbb40922c),
	.w3(32'hbb58dd6c),
	.w4(32'hba265367),
	.w5(32'h3bca2b89),
	.w6(32'h38a510fb),
	.w7(32'hbaa3e99d),
	.w8(32'hbb4b3657),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32a7c3),
	.w1(32'h39604149),
	.w2(32'h3aa7c038),
	.w3(32'h3b7acc95),
	.w4(32'h3c341c64),
	.w5(32'h3b1ae45e),
	.w6(32'hbac61318),
	.w7(32'h3b89bd47),
	.w8(32'h3ab17596),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2abd19),
	.w1(32'hbb31a1b0),
	.w2(32'hbb838e9e),
	.w3(32'h3be791c0),
	.w4(32'h3b37ade9),
	.w5(32'hbb17f2e2),
	.w6(32'h3b85e867),
	.w7(32'hb996972a),
	.w8(32'h3b7a1024),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80f5c5),
	.w1(32'h3981466c),
	.w2(32'hbc023a01),
	.w3(32'h3b6223c1),
	.w4(32'h3b8a8d58),
	.w5(32'hba7ae55a),
	.w6(32'h3b26fdff),
	.w7(32'hb94addbe),
	.w8(32'hbb2f9d23),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba15da7),
	.w1(32'h3b56369c),
	.w2(32'hbb4293ec),
	.w3(32'hba1fda0c),
	.w4(32'hbbc2ca23),
	.w5(32'hbafef16c),
	.w6(32'hbc0ea80f),
	.w7(32'hbb1524c0),
	.w8(32'h3a27ccb8),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badc6a3),
	.w1(32'h3b13840c),
	.w2(32'h3a959b59),
	.w3(32'h3b813db0),
	.w4(32'h3ac7156d),
	.w5(32'h3add9b08),
	.w6(32'h3b208f17),
	.w7(32'h3b6da1da),
	.w8(32'h3ac25233),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02c2f5),
	.w1(32'h3bcf8c23),
	.w2(32'h3ad6330b),
	.w3(32'hbb46a85d),
	.w4(32'hbb47d4a8),
	.w5(32'h3bf7fc88),
	.w6(32'hbbec3cb7),
	.w7(32'hba2e1c08),
	.w8(32'hbab6f6d7),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37de36),
	.w1(32'hbbcf5d61),
	.w2(32'hbc09d787),
	.w3(32'hbb1d2a3c),
	.w4(32'hbabc02bf),
	.w5(32'hbb2ca704),
	.w6(32'hbba1db7c),
	.w7(32'hbb9c08ce),
	.w8(32'hbb51414b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87b9c1),
	.w1(32'hbbbfa039),
	.w2(32'hbb0150db),
	.w3(32'h3b5fa4c3),
	.w4(32'h3af0d790),
	.w5(32'hba321e27),
	.w6(32'hbb401888),
	.w7(32'hbb75ec46),
	.w8(32'hbb2eaabd),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9933e25),
	.w1(32'hbbb0c7cf),
	.w2(32'hbb154d4a),
	.w3(32'hb90f6c5f),
	.w4(32'h3b8c7a54),
	.w5(32'h3b15a28f),
	.w6(32'hbbc552a7),
	.w7(32'hba877cbe),
	.w8(32'h3acae6a0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule