module layer_10_featuremap_500(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3679ed),
	.w1(32'hba30f704),
	.w2(32'h3acf090d),
	.w3(32'hbb867463),
	.w4(32'hbb8f1fe1),
	.w5(32'h3af5584c),
	.w6(32'hbbcf664d),
	.w7(32'h3a80d124),
	.w8(32'h3b28503d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a85a9),
	.w1(32'hbb2800d6),
	.w2(32'hbb75e750),
	.w3(32'hbb005db6),
	.w4(32'h3b3aae99),
	.w5(32'h3b70fd0e),
	.w6(32'h3b866bc3),
	.w7(32'hbb4b7d41),
	.w8(32'hbb3df981),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f0952),
	.w1(32'hbb2386e6),
	.w2(32'hbbac323d),
	.w3(32'hb810ab1f),
	.w4(32'h3bba3f0c),
	.w5(32'h3ba89f4f),
	.w6(32'hbb43b734),
	.w7(32'h3c06db4b),
	.w8(32'h3be993f8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30968e),
	.w1(32'hbb87cb0e),
	.w2(32'h3b62876c),
	.w3(32'hbb6899fc),
	.w4(32'hbb942c95),
	.w5(32'hbbb5e947),
	.w6(32'h3b974376),
	.w7(32'hbb519e20),
	.w8(32'h3a81a5ba),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40c65e),
	.w1(32'hbae48eef),
	.w2(32'h39f2a4c5),
	.w3(32'hbb466299),
	.w4(32'h3b24c989),
	.w5(32'hbb774ef3),
	.w6(32'h3b8af64a),
	.w7(32'h3b958ab1),
	.w8(32'hb98dcbb5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1474a),
	.w1(32'h3b91656e),
	.w2(32'hbbc7172d),
	.w3(32'hbb8305d5),
	.w4(32'h3c906d87),
	.w5(32'h3b16ec1f),
	.w6(32'h39b45e79),
	.w7(32'h3c944596),
	.w8(32'h3c8de8b8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4f696),
	.w1(32'hbb88a181),
	.w2(32'h3ab95337),
	.w3(32'h3bb2ed17),
	.w4(32'hbb94d328),
	.w5(32'hbb039e72),
	.w6(32'hba959264),
	.w7(32'hba00366a),
	.w8(32'h3bc29120),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69ad4d),
	.w1(32'hb9311e34),
	.w2(32'h3a89fdb9),
	.w3(32'hbc04a70b),
	.w4(32'h3c479953),
	.w5(32'hbb37a170),
	.w6(32'h3aad4ac3),
	.w7(32'h3a2333ff),
	.w8(32'h3adb0db4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4468e8),
	.w1(32'hbaf7614b),
	.w2(32'h3bdcdc0b),
	.w3(32'hbb699958),
	.w4(32'hb9b36f84),
	.w5(32'h3b8d24ad),
	.w6(32'h3b56a78c),
	.w7(32'h3b22fbee),
	.w8(32'h3be62956),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b877b8d),
	.w1(32'hbad03ce0),
	.w2(32'hbb901891),
	.w3(32'hbb266e5e),
	.w4(32'hba774162),
	.w5(32'hbb644913),
	.w6(32'h3b144256),
	.w7(32'h3bd5dc25),
	.w8(32'hb8ef7301),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefee18),
	.w1(32'hba0eed6a),
	.w2(32'hbb2544ae),
	.w3(32'hbaa08481),
	.w4(32'hbc0507c4),
	.w5(32'h3b8e5fb8),
	.w6(32'h3bb66640),
	.w7(32'hb9529560),
	.w8(32'h3a521278),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e9c3e),
	.w1(32'hbc32eac8),
	.w2(32'h3aa580e6),
	.w3(32'hbc0c90bf),
	.w4(32'hbb709aa7),
	.w5(32'h3a5fde73),
	.w6(32'hbb94b23f),
	.w7(32'hbad4a271),
	.w8(32'hba7a6cce),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe26615),
	.w1(32'h3b4bf911),
	.w2(32'hbb8265a8),
	.w3(32'hbbba0929),
	.w4(32'h3bbca41f),
	.w5(32'h3b19adb9),
	.w6(32'hbc07a13b),
	.w7(32'h3babc0de),
	.w8(32'h3b031c6c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f9129),
	.w1(32'h3aa12526),
	.w2(32'h3b38d5a7),
	.w3(32'h3b1085b0),
	.w4(32'h3bcb1f99),
	.w5(32'h3c36af1a),
	.w6(32'hbbd92ae1),
	.w7(32'hba89e975),
	.w8(32'h3b832878),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b463113),
	.w1(32'hbbaf97f5),
	.w2(32'hbc121322),
	.w3(32'h3bae92c2),
	.w4(32'hbad6e701),
	.w5(32'hbbf7b7ac),
	.w6(32'h3b5d3d08),
	.w7(32'h3a6c75a9),
	.w8(32'hbb4951fb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d0eda),
	.w1(32'hbad0456c),
	.w2(32'hb9ffeb33),
	.w3(32'hbba069c4),
	.w4(32'hbbc5217c),
	.w5(32'hbba6137a),
	.w6(32'hbb884fd2),
	.w7(32'hbb611c3c),
	.w8(32'hbbde6bff),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f0132),
	.w1(32'hbbaf629c),
	.w2(32'hbb1e9945),
	.w3(32'hbb13b686),
	.w4(32'hbc12cbcf),
	.w5(32'hbb31290d),
	.w6(32'hbbc8b343),
	.w7(32'hbc300cf9),
	.w8(32'hbc077b47),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ee878),
	.w1(32'h3ae0decd),
	.w2(32'h3b5cd40b),
	.w3(32'hbb156b38),
	.w4(32'h3ba35417),
	.w5(32'h3c7c36d4),
	.w6(32'hbbc6b8a2),
	.w7(32'hba70e769),
	.w8(32'h3bdba10c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbac4d9),
	.w1(32'hb8658f5a),
	.w2(32'hbb3bba4a),
	.w3(32'h3ad44e5d),
	.w4(32'h3a82a7e3),
	.w5(32'h3b3bb72a),
	.w6(32'h3c2de720),
	.w7(32'h3b9fc11a),
	.w8(32'h3b42a51d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb052f14),
	.w1(32'hbbf37e90),
	.w2(32'hbba358ed),
	.w3(32'h3b0b249b),
	.w4(32'hbc02738f),
	.w5(32'h3bd7cdf4),
	.w6(32'hba08224f),
	.w7(32'hbc60f429),
	.w8(32'hbb644266),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fe118),
	.w1(32'h3ae7e22a),
	.w2(32'hbc335fbd),
	.w3(32'hbba2e17d),
	.w4(32'h3c88fa1f),
	.w5(32'hbc172be6),
	.w6(32'hbc29cf01),
	.w7(32'h3b827d83),
	.w8(32'hbbc70ed3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e7088),
	.w1(32'h3a47d848),
	.w2(32'hbc14314d),
	.w3(32'hbbf792b3),
	.w4(32'h3c0e832a),
	.w5(32'hbbdeb1fc),
	.w6(32'hbc28fe29),
	.w7(32'h3ba44b55),
	.w8(32'h3bbb6ee4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b5647),
	.w1(32'h3b9ba839),
	.w2(32'h3c8d8131),
	.w3(32'hbbf94c64),
	.w4(32'h3b9f0290),
	.w5(32'hbc1608da),
	.w6(32'hbb6be50a),
	.w7(32'h3b58bbd2),
	.w8(32'h3ca7d5bd),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba810aa7),
	.w1(32'hbbc916bf),
	.w2(32'hbbd4a5e4),
	.w3(32'h3c073d30),
	.w4(32'h3b5e22b8),
	.w5(32'hbba48768),
	.w6(32'h3c123607),
	.w7(32'hba7b9bba),
	.w8(32'hba01527c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb25e29),
	.w1(32'h3aa708b7),
	.w2(32'h3ba0172c),
	.w3(32'hba9bd063),
	.w4(32'h3c08c635),
	.w5(32'h3c84265e),
	.w6(32'h3bbd2fcc),
	.w7(32'h3c473f29),
	.w8(32'h3c7c163b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd52d0),
	.w1(32'h3bcbbee5),
	.w2(32'hbbc03411),
	.w3(32'h3c6010c6),
	.w4(32'h3c8e096c),
	.w5(32'hbb67da46),
	.w6(32'h3c138aeb),
	.w7(32'h3c4d2c3f),
	.w8(32'h3c2bfeab),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc031b70),
	.w1(32'hbbcc0ad6),
	.w2(32'hbaba3fd6),
	.w3(32'h3c0c1e75),
	.w4(32'hba926984),
	.w5(32'hbb9389cb),
	.w6(32'h3c3ca4aa),
	.w7(32'hbbe627a1),
	.w8(32'hbbc93cc3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bb29b),
	.w1(32'hbacf6ee2),
	.w2(32'h3be28a09),
	.w3(32'hbb53a982),
	.w4(32'hba689c1c),
	.w5(32'hba1e7175),
	.w6(32'hbb0cc05b),
	.w7(32'h3bd4a2a8),
	.w8(32'h3bc89dfb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ec608),
	.w1(32'hbb5192a8),
	.w2(32'hbbc42a99),
	.w3(32'h38caf3d1),
	.w4(32'hbba591a7),
	.w5(32'hbc421e11),
	.w6(32'h3b37005b),
	.w7(32'hbc5cef23),
	.w8(32'hbc50b9d7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0286f9),
	.w1(32'hbc052339),
	.w2(32'hbc2c1fa9),
	.w3(32'hbc930d71),
	.w4(32'hba594fa3),
	.w5(32'hbcb0f2b4),
	.w6(32'hba80d847),
	.w7(32'h3c2c37a5),
	.w8(32'hbc013327),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5f95f),
	.w1(32'hbbd1a012),
	.w2(32'hbbe713a2),
	.w3(32'hbbac6aac),
	.w4(32'hbc0a2912),
	.w5(32'hbb5aa2e8),
	.w6(32'hbc2b04f8),
	.w7(32'hbc124e8c),
	.w8(32'hbc179f97),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc344bb5),
	.w1(32'hba2b05d3),
	.w2(32'h3ab40953),
	.w3(32'hbc398fa3),
	.w4(32'h3b6d0965),
	.w5(32'hb9c4a744),
	.w6(32'hbc002510),
	.w7(32'h3bb3f52c),
	.w8(32'hbba4f424),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2121b4),
	.w1(32'h3adb3a33),
	.w2(32'h3a911349),
	.w3(32'h39c91545),
	.w4(32'hbb0f302d),
	.w5(32'h3bc4737a),
	.w6(32'hbacf00d5),
	.w7(32'h3b31ce0b),
	.w8(32'hb9da7f38),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc738e2),
	.w1(32'hba81cbd5),
	.w2(32'h3b10131c),
	.w3(32'hbba58ffa),
	.w4(32'hbae24bed),
	.w5(32'hbbc7ccda),
	.w6(32'h3b27310a),
	.w7(32'h3bf23fd1),
	.w8(32'h3ac79558),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adba369),
	.w1(32'hbb9757f4),
	.w2(32'hbbe9cabe),
	.w3(32'hba96f871),
	.w4(32'h3b97d2ef),
	.w5(32'hbc485f54),
	.w6(32'h3bf857af),
	.w7(32'h3bb75a70),
	.w8(32'h3ab1e64a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7b176),
	.w1(32'hbaf96e2b),
	.w2(32'h3bcda43c),
	.w3(32'hbbc9723a),
	.w4(32'hbab837bb),
	.w5(32'h3b064fc0),
	.w6(32'hbb5b4b6b),
	.w7(32'hbbf15aff),
	.w8(32'hbaefa3c9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4cf39),
	.w1(32'hbc3d196b),
	.w2(32'h3ba99097),
	.w3(32'hba46b06c),
	.w4(32'hbc6ef882),
	.w5(32'h3c40c78c),
	.w6(32'h3ac258a3),
	.w7(32'hbb3ff85c),
	.w8(32'h3b931792),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94149b),
	.w1(32'hbb27b23e),
	.w2(32'hbb5b69c8),
	.w3(32'h3aac6f8d),
	.w4(32'hbafc7d34),
	.w5(32'h3ae0a426),
	.w6(32'h3b592e41),
	.w7(32'h3b9b2261),
	.w8(32'h3be5db48),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb414052),
	.w1(32'hb9a8889a),
	.w2(32'hbaa9450b),
	.w3(32'hbb0e5b28),
	.w4(32'h36d63f67),
	.w5(32'h3baf9abf),
	.w6(32'h3b8dd2fe),
	.w7(32'hbb2f7aae),
	.w8(32'h3b98e6b8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e544b),
	.w1(32'h3b02dd5d),
	.w2(32'h3c20b8a2),
	.w3(32'hbac743aa),
	.w4(32'hbbc82eee),
	.w5(32'h3a9760e4),
	.w6(32'h3b7f56ca),
	.w7(32'hbb486c16),
	.w8(32'h3b8eca6d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23c833),
	.w1(32'h398d9331),
	.w2(32'h3c2e222e),
	.w3(32'h3bb26dca),
	.w4(32'h39fbd468),
	.w5(32'h3bb0f84c),
	.w6(32'h3c169af3),
	.w7(32'hba204255),
	.w8(32'h3b23c6b5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e7e19),
	.w1(32'hbb1e9fd8),
	.w2(32'hbb7e19ca),
	.w3(32'h3b5b4a99),
	.w4(32'h3bc61245),
	.w5(32'h3bca1909),
	.w6(32'hbb242c8c),
	.w7(32'h3b9213e1),
	.w8(32'h3a472d05),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb939e16),
	.w1(32'h39b21b26),
	.w2(32'h3b004e50),
	.w3(32'h3ad530c4),
	.w4(32'hba9ac506),
	.w5(32'hba8f2dce),
	.w6(32'hbb54bd17),
	.w7(32'h3a57a083),
	.w8(32'hba84959a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4499f),
	.w1(32'hbbd9ae47),
	.w2(32'hbc1401df),
	.w3(32'h3b8a4476),
	.w4(32'hbab5dbd4),
	.w5(32'hbb0d9257),
	.w6(32'h3bf4df34),
	.w7(32'h3b5007be),
	.w8(32'h3bb74a93),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c310c),
	.w1(32'hbbdcb7e2),
	.w2(32'hbbf3299a),
	.w3(32'hbbc00085),
	.w4(32'hbc270c0e),
	.w5(32'hbb77f72f),
	.w6(32'hbabe3bc3),
	.w7(32'h3a4932db),
	.w8(32'h3891b988),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae79de1),
	.w1(32'hbbc0a14c),
	.w2(32'h3b75539b),
	.w3(32'hbbf17645),
	.w4(32'hbc2ed5db),
	.w5(32'hbbc45d0c),
	.w6(32'hbb70f11e),
	.w7(32'hbc010d8f),
	.w8(32'hbc420b66),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8e106),
	.w1(32'h3bddfc69),
	.w2(32'hbb1420a2),
	.w3(32'hbbb756fe),
	.w4(32'h3bb26f2c),
	.w5(32'h3bd29f12),
	.w6(32'hbbf5b35f),
	.w7(32'h3c20bf87),
	.w8(32'h3c035252),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ae036),
	.w1(32'h3a893c7e),
	.w2(32'h3c00a33e),
	.w3(32'h3baee2df),
	.w4(32'h3b186384),
	.w5(32'h3bbabed6),
	.w6(32'h3c129dd5),
	.w7(32'hbb5e6f55),
	.w8(32'h3b77a193),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ad2d7),
	.w1(32'h3bf179cf),
	.w2(32'h3a7300d5),
	.w3(32'hbba0c426),
	.w4(32'h3ba3d231),
	.w5(32'hbb22fd0a),
	.w6(32'hbb106a4a),
	.w7(32'hbbdc0154),
	.w8(32'hbb992850),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c230caf),
	.w1(32'h3ae4b82c),
	.w2(32'h3ad7f112),
	.w3(32'h3a9c4b82),
	.w4(32'h3b1520ff),
	.w5(32'hbbdd4fc4),
	.w6(32'h3a3b8b8e),
	.w7(32'h3ad68a95),
	.w8(32'hbbe0d09d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbcc0f),
	.w1(32'hba4844f8),
	.w2(32'hbb1283ac),
	.w3(32'h3c77e971),
	.w4(32'h3c066c4e),
	.w5(32'hbc347604),
	.w6(32'hba776eb1),
	.w7(32'h3bad6355),
	.w8(32'h3a76fc02),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06cb63),
	.w1(32'hbb5d5944),
	.w2(32'hbc0b3e2b),
	.w3(32'hbae601f9),
	.w4(32'hbaa25f56),
	.w5(32'hba188c7e),
	.w6(32'h3a30e894),
	.w7(32'hbb145ee8),
	.w8(32'hbb61705d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96eb34),
	.w1(32'h3ae32c56),
	.w2(32'hbb3c2132),
	.w3(32'hbbb0ea02),
	.w4(32'h3ab87603),
	.w5(32'hbb9587fd),
	.w6(32'hb99bb34b),
	.w7(32'h3b4e91cf),
	.w8(32'h3b8fb1b4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba8f42),
	.w1(32'h3ba859c3),
	.w2(32'h3b2f7fe4),
	.w3(32'h3c04874d),
	.w4(32'h3c5bd719),
	.w5(32'hbab035f3),
	.w6(32'h3bf76e32),
	.w7(32'h3bad07fb),
	.w8(32'h3b8dccc0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89c09a),
	.w1(32'hbbb1c02f),
	.w2(32'h3bc974c2),
	.w3(32'h3b5361fd),
	.w4(32'hbb8f6031),
	.w5(32'h3b821625),
	.w6(32'h3b255de9),
	.w7(32'hbc354b9a),
	.w8(32'hbbcd9ed1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb858c2e),
	.w1(32'h3a9a022b),
	.w2(32'hbb72e817),
	.w3(32'h3b63b2dc),
	.w4(32'h3bb22877),
	.w5(32'h3b81c108),
	.w6(32'h3b717a06),
	.w7(32'hbb28cf0c),
	.w8(32'h3b62eb6c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f73b9),
	.w1(32'h3b9c4c37),
	.w2(32'h3c1b0c41),
	.w3(32'hbbaecacb),
	.w4(32'h3c1be91e),
	.w5(32'h3beca5cc),
	.w6(32'hbb0694d5),
	.w7(32'h3c585364),
	.w8(32'h3b9e4dac),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51e167),
	.w1(32'hbb55c251),
	.w2(32'hbb1f5f63),
	.w3(32'h3a99b28a),
	.w4(32'hbb341f4e),
	.w5(32'hbbfc0268),
	.w6(32'h394a54dc),
	.w7(32'h3b9e5c1a),
	.w8(32'hbb9ea663),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a05eb),
	.w1(32'hbbe04a6d),
	.w2(32'hbbd54510),
	.w3(32'hbbba6cc2),
	.w4(32'hbbc0f72c),
	.w5(32'h39c5987a),
	.w6(32'hbb0d038c),
	.w7(32'hbb821d17),
	.w8(32'hbb6e6b03),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b768826),
	.w1(32'h3c8d1014),
	.w2(32'h3cf1b50e),
	.w3(32'hbb32482a),
	.w4(32'h3be92943),
	.w5(32'h3cbe7796),
	.w6(32'h3c0e868d),
	.w7(32'h3c5593a6),
	.w8(32'h3c585fd9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19d0d5),
	.w1(32'h3b88387f),
	.w2(32'h3c0e9693),
	.w3(32'h3c9fac41),
	.w4(32'h3c453a78),
	.w5(32'h3c6c2436),
	.w6(32'h3c45035d),
	.w7(32'h3bba3444),
	.w8(32'h3892037a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb903cd3a),
	.w1(32'h3a333a70),
	.w2(32'h3b68cd6c),
	.w3(32'h3c5c71cd),
	.w4(32'hbb7d4953),
	.w5(32'hbb7bfee5),
	.w6(32'h3bfc20ab),
	.w7(32'hba044d2b),
	.w8(32'hbb0cc032),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0a9b7),
	.w1(32'h3b50d750),
	.w2(32'hb8b9a30a),
	.w3(32'hbbdd14b3),
	.w4(32'h3b1da33b),
	.w5(32'hba9c9445),
	.w6(32'hbbd7320f),
	.w7(32'hbb5be78a),
	.w8(32'hbbbfec42),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf43167),
	.w1(32'h3a9b9134),
	.w2(32'h3b44b5db),
	.w3(32'h3a0673a4),
	.w4(32'h38a6d3a6),
	.w5(32'h3ad14061),
	.w6(32'h3b6eb4e9),
	.w7(32'h3944f9d8),
	.w8(32'h3b80dbfd),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79f7ba),
	.w1(32'h3b68533b),
	.w2(32'h3a22988b),
	.w3(32'hba6060c7),
	.w4(32'h3ba0012f),
	.w5(32'h3b8b2e6e),
	.w6(32'h3b83d43c),
	.w7(32'h3bb7b1ed),
	.w8(32'h3bec8d73),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf62df5),
	.w1(32'h3ae850d8),
	.w2(32'hbb53ac35),
	.w3(32'h3be0566e),
	.w4(32'hba4a2560),
	.w5(32'hba0d9e88),
	.w6(32'h3c11dd3c),
	.w7(32'hbbc5b9de),
	.w8(32'hbb76328b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb0529),
	.w1(32'hbad5158c),
	.w2(32'hbb564880),
	.w3(32'hbbcaff98),
	.w4(32'h3a8ba0a6),
	.w5(32'hbc11c211),
	.w6(32'hbb348f25),
	.w7(32'h3be70f58),
	.w8(32'h3c3c6439),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf5189),
	.w1(32'h3c2e2735),
	.w2(32'h3bfc026d),
	.w3(32'h3a892a95),
	.w4(32'h3b8ec2ee),
	.w5(32'hbac0f221),
	.w6(32'hb9c3c1be),
	.w7(32'hbc246577),
	.w8(32'hbb60806c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c811f70),
	.w1(32'h3a1e9761),
	.w2(32'hbb936fea),
	.w3(32'h3be9dba9),
	.w4(32'hbbffd66b),
	.w5(32'hbc16ed4a),
	.w6(32'h3ad7639e),
	.w7(32'hbc35a636),
	.w8(32'hbbcda5a3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73db5d),
	.w1(32'hb8be8bfc),
	.w2(32'h3b22a6a9),
	.w3(32'hbc589af3),
	.w4(32'hbb3ae06b),
	.w5(32'hbb86178d),
	.w6(32'hbbe824ed),
	.w7(32'h3c0c7d41),
	.w8(32'h3b8c92f3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8ba8b),
	.w1(32'h3a8b9a24),
	.w2(32'h3ac84ecf),
	.w3(32'h3b4b1dda),
	.w4(32'hbb09fbe4),
	.w5(32'hbba553b2),
	.w6(32'h3b9ba793),
	.w7(32'hbc1b8bd8),
	.w8(32'hbc36f4cb),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2e753),
	.w1(32'h3a8c6a33),
	.w2(32'hbb537183),
	.w3(32'hbc1de070),
	.w4(32'h3b5a0e5e),
	.w5(32'hbac868d6),
	.w6(32'hbbffe99d),
	.w7(32'hbbbaada2),
	.w8(32'hbc79baf2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bc371),
	.w1(32'hbbac698e),
	.w2(32'hbb0fa1b1),
	.w3(32'hbb8042a9),
	.w4(32'hbc07da3e),
	.w5(32'hbbbce592),
	.w6(32'hbc3f9de0),
	.w7(32'hbb1e46d8),
	.w8(32'hbad7302e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86835a),
	.w1(32'hbc865bb0),
	.w2(32'hbc1b41b9),
	.w3(32'h3b66aef5),
	.w4(32'hbaf906c4),
	.w5(32'h3ba8e254),
	.w6(32'h3ac5a2b2),
	.w7(32'h3b2ff1aa),
	.w8(32'h3c4c3d01),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77a081),
	.w1(32'hba9e367b),
	.w2(32'hbbf91ba2),
	.w3(32'h3b16b043),
	.w4(32'hb8db60a4),
	.w5(32'h3ae8512b),
	.w6(32'h3b9ede42),
	.w7(32'hbb318f34),
	.w8(32'hbbbd50a2),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6c26d),
	.w1(32'hba0c38c8),
	.w2(32'h3a48b523),
	.w3(32'h3b5cd0bb),
	.w4(32'h3bccdd2f),
	.w5(32'h3ad77146),
	.w6(32'hbb9349bb),
	.w7(32'h3c03fc49),
	.w8(32'h3bbb335b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93932d),
	.w1(32'h3bf1b186),
	.w2(32'h3c17de03),
	.w3(32'h3b92cc67),
	.w4(32'h3ab6a953),
	.w5(32'h3bb4614e),
	.w6(32'h3b747f22),
	.w7(32'h3c143057),
	.w8(32'h3c11a949),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad5d17),
	.w1(32'hbc708dcf),
	.w2(32'hbc927083),
	.w3(32'hbb95c375),
	.w4(32'h3c34fcd2),
	.w5(32'hbb1afa64),
	.w6(32'h3b44bcbe),
	.w7(32'h3c4a151b),
	.w8(32'h3bf6d7af),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd00a06),
	.w1(32'h3a8acf9f),
	.w2(32'hbbe6328f),
	.w3(32'h3bca19ee),
	.w4(32'h3c586d1a),
	.w5(32'h3b499430),
	.w6(32'h3c6e96c6),
	.w7(32'h3bf6f80f),
	.w8(32'hbaab4293),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0610e8),
	.w1(32'hbbc38b58),
	.w2(32'hbb88cd4c),
	.w3(32'hb9a72b9b),
	.w4(32'hba5bbdd7),
	.w5(32'hbb282a95),
	.w6(32'hbb182b41),
	.w7(32'h3b4b3b19),
	.w8(32'h3a76c848),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb005c7e),
	.w1(32'hbaf73c8f),
	.w2(32'hbbe3b527),
	.w3(32'hbb055b56),
	.w4(32'h3b97cc8f),
	.w5(32'h3c19a37d),
	.w6(32'hbab659e2),
	.w7(32'h3b5ce73c),
	.w8(32'hbb0cf2fd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad21013),
	.w1(32'h3a27fea7),
	.w2(32'h3b5da4c5),
	.w3(32'h3bf6c6cb),
	.w4(32'hbae8cb43),
	.w5(32'hbb0646da),
	.w6(32'h3b0fcfb6),
	.w7(32'hbac567dd),
	.w8(32'h3abf5de0),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa00c9),
	.w1(32'h3bd6c03c),
	.w2(32'h3c015a67),
	.w3(32'hba6cf8a1),
	.w4(32'h3c05980d),
	.w5(32'h3bffadbf),
	.w6(32'h3b82b986),
	.w7(32'hbc368e38),
	.w8(32'hbcbeabd8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd11c83),
	.w1(32'h3a38d00f),
	.w2(32'h3a0a28da),
	.w3(32'h39f5d1a2),
	.w4(32'h3a0e51de),
	.w5(32'h3aee7b98),
	.w6(32'hbc9790fd),
	.w7(32'hbb5aecec),
	.w8(32'h3a6b2c7d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7f620),
	.w1(32'hbb760915),
	.w2(32'hbbf5521c),
	.w3(32'hbae635e5),
	.w4(32'hbba5e733),
	.w5(32'hbc11a9e7),
	.w6(32'h3b9bdda3),
	.w7(32'hbb98a969),
	.w8(32'hbc1f51a5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5707e4),
	.w1(32'hbbfc08b3),
	.w2(32'hb9c12a1f),
	.w3(32'hbbe9a3dc),
	.w4(32'hbb592ff0),
	.w5(32'h3a81cb7e),
	.w6(32'hbc70ddd0),
	.w7(32'h3bf206e0),
	.w8(32'h3c12b1d7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dba52),
	.w1(32'hbc5f8bf2),
	.w2(32'hbbf91c3e),
	.w3(32'h3a891a32),
	.w4(32'hbbcb376d),
	.w5(32'hbc371c1f),
	.w6(32'h3b3f8ff1),
	.w7(32'h3bb67736),
	.w8(32'h3b2dbe46),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81c1e7),
	.w1(32'hbade08c1),
	.w2(32'hbb226805),
	.w3(32'hbae07114),
	.w4(32'h3c361004),
	.w5(32'h3b5b1fc7),
	.w6(32'h3b49f710),
	.w7(32'h3c786028),
	.w8(32'h3c583995),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe64841),
	.w1(32'h3be3b097),
	.w2(32'h3b5dd415),
	.w3(32'hba8ba30a),
	.w4(32'hbb18db1f),
	.w5(32'h3b7d3913),
	.w6(32'h3c399783),
	.w7(32'hba62acc6),
	.w8(32'hbaea7c79),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc79ec4),
	.w1(32'hbb812751),
	.w2(32'h3b693ac6),
	.w3(32'h3c040cc4),
	.w4(32'h3bdfc856),
	.w5(32'h3bcc00b8),
	.w6(32'h39db8bb4),
	.w7(32'h3bed7867),
	.w8(32'h3c5ec80e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ba1ce),
	.w1(32'hbb8ef138),
	.w2(32'h3b35b342),
	.w3(32'hbc154dd8),
	.w4(32'hbc417e67),
	.w5(32'hbbfbe882),
	.w6(32'hbb91651a),
	.w7(32'hbc09e399),
	.w8(32'hbaacc0ac),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85859a),
	.w1(32'h3ada5802),
	.w2(32'h3c028554),
	.w3(32'hbb9a7e89),
	.w4(32'hbbd0bae2),
	.w5(32'hbb6c2d70),
	.w6(32'hbb756bae),
	.w7(32'hbb67d84e),
	.w8(32'h3a2811fd),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6f193),
	.w1(32'h3cac89ad),
	.w2(32'h3ca48a3c),
	.w3(32'h3ba9803d),
	.w4(32'h3c3c8a9f),
	.w5(32'h3c6bc643),
	.w6(32'h3ad0920a),
	.w7(32'hbcddef0e),
	.w8(32'hbd023940),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba08b8),
	.w1(32'h3b19354d),
	.w2(32'hbb8eea0c),
	.w3(32'h3c233a6d),
	.w4(32'h3c087dc3),
	.w5(32'h3bb98c55),
	.w6(32'hbcd55551),
	.w7(32'h3bbe76f1),
	.w8(32'hbb045135),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5794af),
	.w1(32'h39f92905),
	.w2(32'hbaa49b70),
	.w3(32'h3b8442b5),
	.w4(32'hbae72703),
	.w5(32'h3a47b7d4),
	.w6(32'h3ac71dfc),
	.w7(32'h3b2cdaad),
	.w8(32'h3bad1ae7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ec9b6),
	.w1(32'hba2cf629),
	.w2(32'h3af753f7),
	.w3(32'h3c00f30b),
	.w4(32'hbaeeb341),
	.w5(32'h3b9c8af8),
	.w6(32'h3ba8c921),
	.w7(32'h3b3bde55),
	.w8(32'h3c387b33),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d6307),
	.w1(32'hba142b7c),
	.w2(32'hbbc225bf),
	.w3(32'h3c5a541b),
	.w4(32'hbbf04e6b),
	.w5(32'hbc182e48),
	.w6(32'hbb5c7c1f),
	.w7(32'hbaa925d7),
	.w8(32'h3bbe1735),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7278b4),
	.w1(32'h3b90e59e),
	.w2(32'hbaf0a684),
	.w3(32'hbbe1a73b),
	.w4(32'h3bca5817),
	.w5(32'hbb8df4e3),
	.w6(32'hba26facb),
	.w7(32'h3b2a960a),
	.w8(32'hbba63b09),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb937172),
	.w1(32'hbb65f08e),
	.w2(32'h3b1e89a1),
	.w3(32'hbbfad010),
	.w4(32'hbc76c5aa),
	.w5(32'hbcb9bebb),
	.w6(32'hbbf8e42f),
	.w7(32'hb9e246a5),
	.w8(32'h3bb6bcce),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5156d8),
	.w1(32'h3a135267),
	.w2(32'h3c03bbac),
	.w3(32'hbc338a1f),
	.w4(32'hbb3f2c64),
	.w5(32'h3c333b8f),
	.w6(32'h3bfea6d1),
	.w7(32'h397363f7),
	.w8(32'h3c4ce2e3),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fbd7e),
	.w1(32'hbcae1045),
	.w2(32'hbc862901),
	.w3(32'hbb4bd99f),
	.w4(32'hbc99638b),
	.w5(32'hbc7ab371),
	.w6(32'h3c0cb70e),
	.w7(32'hbc05daf3),
	.w8(32'h3b6150a3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99c43d),
	.w1(32'hbba9256f),
	.w2(32'hbc162e79),
	.w3(32'hbc5d6191),
	.w4(32'hbb537bcb),
	.w5(32'h3a8ec6e0),
	.w6(32'h3ac2e637),
	.w7(32'hbbbbb822),
	.w8(32'hbc40a029),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44b299),
	.w1(32'h3c896835),
	.w2(32'h3c2cfc4f),
	.w3(32'h3b289014),
	.w4(32'h3b45768c),
	.w5(32'hbb5daa92),
	.w6(32'hbc4ce489),
	.w7(32'h3c14741a),
	.w8(32'h3bbd26e6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f3511),
	.w1(32'hbc10c315),
	.w2(32'hbbae8b4f),
	.w3(32'hbb8ceae9),
	.w4(32'hbb5da4ad),
	.w5(32'hbc04e1f8),
	.w6(32'h3af26a11),
	.w7(32'hbbee913f),
	.w8(32'hbbcbeeef),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b509c68),
	.w1(32'h3c69c766),
	.w2(32'h3caac148),
	.w3(32'h3acf5d5a),
	.w4(32'h3b9026fd),
	.w5(32'h3c5ecb07),
	.w6(32'hbb2f7673),
	.w7(32'hbba6eb37),
	.w8(32'hbb5df0cd),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cedc2),
	.w1(32'hbc9e4454),
	.w2(32'hbc569019),
	.w3(32'h3c127cd8),
	.w4(32'hbc764b06),
	.w5(32'hbbc9fc11),
	.w6(32'hba21d7f5),
	.w7(32'h3b2291eb),
	.w8(32'h3c3748c8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd48d9),
	.w1(32'h3c93dd1c),
	.w2(32'h3c452dd6),
	.w3(32'hbb537e71),
	.w4(32'h3caa72f3),
	.w5(32'h3b9a5bfa),
	.w6(32'h3b9fd50e),
	.w7(32'h3bcf353d),
	.w8(32'hbb5d42bc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c295868),
	.w1(32'h3a226dc8),
	.w2(32'h3b9e01ab),
	.w3(32'hba517e2a),
	.w4(32'hbb646f73),
	.w5(32'h3a679349),
	.w6(32'h3a89e4e8),
	.w7(32'h3b119331),
	.w8(32'h3baa5403),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9816f38),
	.w1(32'h3b4942f3),
	.w2(32'h3b4a43dd),
	.w3(32'h3b318a0f),
	.w4(32'hbc094698),
	.w5(32'hbb840d38),
	.w6(32'h3788dfa1),
	.w7(32'hbc064c57),
	.w8(32'hbc57a9a4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27bfa4),
	.w1(32'h3b8d9011),
	.w2(32'hbba6e17f),
	.w3(32'hbaf5f08f),
	.w4(32'h3b9530af),
	.w5(32'h3befc95b),
	.w6(32'hbbdabbb8),
	.w7(32'h3b4d8e59),
	.w8(32'h395a5d01),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2686c),
	.w1(32'h3b639466),
	.w2(32'h3c18cd31),
	.w3(32'h3c41de86),
	.w4(32'h3b2e99ed),
	.w5(32'hb8df4273),
	.w6(32'hbb671c82),
	.w7(32'h39b00428),
	.w8(32'h3b8feb36),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a6c3b),
	.w1(32'h3a702b42),
	.w2(32'h3c0f1bb7),
	.w3(32'hbb294840),
	.w4(32'hbc008379),
	.w5(32'hb8c51805),
	.w6(32'h388252da),
	.w7(32'hba2b1fe0),
	.w8(32'h3b9cca65),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b680a79),
	.w1(32'hbc69ab8a),
	.w2(32'hbc4288d6),
	.w3(32'hbb9040f7),
	.w4(32'hbc3eac38),
	.w5(32'h3aa88f78),
	.w6(32'hbb124e91),
	.w7(32'h3a9d6505),
	.w8(32'h3c29c05a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02318b),
	.w1(32'hbb1dd918),
	.w2(32'hbbaf67cd),
	.w3(32'h3ba0103e),
	.w4(32'h3b8baba5),
	.w5(32'hbb06fed8),
	.w6(32'h3c55a302),
	.w7(32'hbc0eb6e8),
	.w8(32'hbc91059c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54e157),
	.w1(32'hbb26473e),
	.w2(32'hbbc7c0c6),
	.w3(32'hbc6d8ad5),
	.w4(32'h3b9cbfcd),
	.w5(32'hbbad5b05),
	.w6(32'hbc7f41bc),
	.w7(32'h398b013f),
	.w8(32'hbb1b8cb0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe441c3),
	.w1(32'hbc551302),
	.w2(32'hbc28edf9),
	.w3(32'hbb3471be),
	.w4(32'hbc160d25),
	.w5(32'hbbaaeb71),
	.w6(32'hbb5b63d7),
	.w7(32'hbb914785),
	.w8(32'hbab35d2e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf813fe),
	.w1(32'h3ba42039),
	.w2(32'h3bc13d94),
	.w3(32'hbb6743f5),
	.w4(32'h3b0f5c45),
	.w5(32'h3b07a016),
	.w6(32'hbb839c2c),
	.w7(32'h3b1659aa),
	.w8(32'hbb103d3d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa0c6a),
	.w1(32'h3ca93a05),
	.w2(32'h3cc8a2cf),
	.w3(32'h3b97a2d4),
	.w4(32'h3c19da34),
	.w5(32'h3c075402),
	.w6(32'hbbe4e8e1),
	.w7(32'hbc72a92b),
	.w8(32'hbcb080dd),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1a140),
	.w1(32'hbcb35d2c),
	.w2(32'hbc969dd8),
	.w3(32'h3abc3774),
	.w4(32'hbb0e6460),
	.w5(32'h3aa775b0),
	.w6(32'hbc95f8f5),
	.w7(32'h3a892aca),
	.w8(32'h3b9fea34),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca25ed4),
	.w1(32'hbc2683a5),
	.w2(32'hbc2c99b1),
	.w3(32'hba4278d6),
	.w4(32'hbc240193),
	.w5(32'hbc7db08c),
	.w6(32'h3b724ab6),
	.w7(32'hbc10e7c3),
	.w8(32'hbc379d8c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb75b1),
	.w1(32'h3a1f2847),
	.w2(32'hbb2d78d3),
	.w3(32'hbbc8bec4),
	.w4(32'h3b86f0ae),
	.w5(32'h3b411840),
	.w6(32'hbc33db73),
	.w7(32'hba965ab9),
	.w8(32'hbb28ddc3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d4a5c),
	.w1(32'h3a1b871b),
	.w2(32'h3b12baf1),
	.w3(32'hb9cf2e02),
	.w4(32'h3ad7257f),
	.w5(32'h3befb4bb),
	.w6(32'hbafe2780),
	.w7(32'hba3b51f0),
	.w8(32'h3bc9c959),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb642b69),
	.w1(32'h3a936732),
	.w2(32'hbad1ea7f),
	.w3(32'hbade9174),
	.w4(32'hba91e163),
	.w5(32'hbb3e8e31),
	.w6(32'h3bbe0532),
	.w7(32'h3b3a2ba8),
	.w8(32'h3af2b70b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2767),
	.w1(32'hbb742c93),
	.w2(32'h397d1897),
	.w3(32'hbb5e411d),
	.w4(32'h3a90defd),
	.w5(32'h3c370750),
	.w6(32'h3ac4a75a),
	.w7(32'hbba5808d),
	.w8(32'h397be325),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16e774),
	.w1(32'h3c593bb6),
	.w2(32'h3c51e5c0),
	.w3(32'h3c88b005),
	.w4(32'h3ba06151),
	.w5(32'h3c02e4ee),
	.w6(32'h3a4a05f0),
	.w7(32'hbbad98cf),
	.w8(32'hbbf38468),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b394c),
	.w1(32'hbb2848fd),
	.w2(32'h3b1897ad),
	.w3(32'h3b724006),
	.w4(32'h3c26a003),
	.w5(32'h3c686f08),
	.w6(32'hbc5caa52),
	.w7(32'hbb0ab8bb),
	.w8(32'h3b8cf020),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1923d),
	.w1(32'hbb915aa4),
	.w2(32'h38d5b00c),
	.w3(32'h3c482278),
	.w4(32'hbc3768d2),
	.w5(32'hbc3ca48e),
	.w6(32'h3c26657e),
	.w7(32'hbc0e31be),
	.w8(32'hbb35eff6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba61e33),
	.w1(32'h3afe34ee),
	.w2(32'h3b3c7588),
	.w3(32'hbc8166c8),
	.w4(32'hbb80fafb),
	.w5(32'h3b82dbbb),
	.w6(32'hbc28376e),
	.w7(32'hba835243),
	.w8(32'h3b08bf9e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b447c3f),
	.w1(32'hbbc11167),
	.w2(32'hbbb4848b),
	.w3(32'hbb03bddd),
	.w4(32'hbc41bc3a),
	.w5(32'hbc24ef9c),
	.w6(32'hbae9a6b6),
	.w7(32'hba877a26),
	.w8(32'hbb671a5e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93bff8),
	.w1(32'hbc4bf274),
	.w2(32'hbbb5f230),
	.w3(32'hbb99e123),
	.w4(32'hbbbfcf06),
	.w5(32'hbbdfb9f6),
	.w6(32'hbaa36dd1),
	.w7(32'hbc1b7c2a),
	.w8(32'hbc481b3b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ef3d4),
	.w1(32'hb9ed9d6a),
	.w2(32'hbbdb40f2),
	.w3(32'hbb8af114),
	.w4(32'hba1e85a5),
	.w5(32'hbc26784c),
	.w6(32'hbc114dc0),
	.w7(32'h3bbe1da4),
	.w8(32'hbc03a935),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a5ebe),
	.w1(32'hbc381405),
	.w2(32'hbb979b10),
	.w3(32'hbc05bbc2),
	.w4(32'h3823414b),
	.w5(32'h3bede703),
	.w6(32'hbba32615),
	.w7(32'hbc202d49),
	.w8(32'hbbe02be8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8af95),
	.w1(32'hbb0f9f62),
	.w2(32'hbbbd9918),
	.w3(32'hbaa2a549),
	.w4(32'hbb2a00e8),
	.w5(32'hba615d23),
	.w6(32'hbb2fbf1b),
	.w7(32'hbb51f2e9),
	.w8(32'hbbf9d762),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3897e37e),
	.w1(32'hb9e0b97a),
	.w2(32'h39ee6d14),
	.w3(32'h3bbb2ab1),
	.w4(32'hba9d9a4c),
	.w5(32'h3c1730be),
	.w6(32'hbb88299e),
	.w7(32'hba1f97bc),
	.w8(32'h39a314f7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77d062),
	.w1(32'hbba91fce),
	.w2(32'hb97e2b98),
	.w3(32'h3b4b7449),
	.w4(32'h3bdbdec6),
	.w5(32'h3bda2ced),
	.w6(32'h3ae8002c),
	.w7(32'h3c46bffd),
	.w8(32'h3c872286),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc1918),
	.w1(32'hbcfede31),
	.w2(32'hbd066f27),
	.w3(32'h3bc217ad),
	.w4(32'h3b56a14a),
	.w5(32'h3b1a59ed),
	.w6(32'h3bd2be1c),
	.w7(32'h3cbfd07f),
	.w8(32'h3cbd503c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce7210f),
	.w1(32'hb99e2121),
	.w2(32'h3bb6643a),
	.w3(32'h3b79bc8e),
	.w4(32'hbb98e4bb),
	.w5(32'hbadcc4de),
	.w6(32'h3cdc4c1f),
	.w7(32'h3a53aad8),
	.w8(32'h3c4fd09b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc3b5b),
	.w1(32'h3c642f2d),
	.w2(32'h3c886f7d),
	.w3(32'hbafc6ea4),
	.w4(32'hbb0ea0f0),
	.w5(32'hbab75d4c),
	.w6(32'h3aca42db),
	.w7(32'hbc0e6428),
	.w8(32'hbb7b4628),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22542d),
	.w1(32'h3c612140),
	.w2(32'h3c8bb36c),
	.w3(32'hbbc2c516),
	.w4(32'hbbdcc00f),
	.w5(32'hbb59c933),
	.w6(32'hba30fefe),
	.w7(32'hba4077eb),
	.w8(32'hbadfe331),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f43e5),
	.w1(32'hbb5b9400),
	.w2(32'hba296875),
	.w3(32'h3a304dc6),
	.w4(32'hbba124c4),
	.w5(32'hba76a028),
	.w6(32'h394ccc52),
	.w7(32'hb98665ce),
	.w8(32'h3ac796a9),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0072f),
	.w1(32'hbb87c067),
	.w2(32'hba369196),
	.w3(32'h39ac3047),
	.w4(32'h3c2d675a),
	.w5(32'h3b5e06d3),
	.w6(32'h3a837060),
	.w7(32'h3a8d9e00),
	.w8(32'hbb1fbb52),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b408e7f),
	.w1(32'hbaf661c7),
	.w2(32'hbc05ce1a),
	.w3(32'h3b04f06c),
	.w4(32'hbba1ea64),
	.w5(32'hbb301162),
	.w6(32'h3b8f9e22),
	.w7(32'hbb3217bb),
	.w8(32'hbc1de72c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d9be0),
	.w1(32'h3a506e09),
	.w2(32'h3b482253),
	.w3(32'h3b26d79e),
	.w4(32'hba9a4252),
	.w5(32'hbaf217ad),
	.w6(32'hbba92587),
	.w7(32'h3a375bde),
	.w8(32'hbadae177),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8866343),
	.w1(32'hba8b6adc),
	.w2(32'h39d8e74a),
	.w3(32'h3b751756),
	.w4(32'h39e86238),
	.w5(32'hbbb9375a),
	.w6(32'hbb6e641c),
	.w7(32'h3a812390),
	.w8(32'h39e94685),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b064140),
	.w1(32'hbb12a0af),
	.w2(32'h386defd1),
	.w3(32'hbbd319f5),
	.w4(32'hbbf111c4),
	.w5(32'hbbd6e1ed),
	.w6(32'h3ab9794f),
	.w7(32'hbc849d0a),
	.w8(32'hbc431587),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7da884),
	.w1(32'h3c1532b9),
	.w2(32'h3c2471bc),
	.w3(32'hbb8269f4),
	.w4(32'hbb0f3823),
	.w5(32'hbc02fa8f),
	.w6(32'hbc1d6ee2),
	.w7(32'hb9fe4240),
	.w8(32'hbbc0c9f0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25eac2),
	.w1(32'hbb80d25b),
	.w2(32'hba8cf071),
	.w3(32'hbbac664c),
	.w4(32'hbc141465),
	.w5(32'hbbba46e3),
	.w6(32'h3a42673e),
	.w7(32'hbbda2ffb),
	.w8(32'hbb7fa14c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2fab4),
	.w1(32'h3a0c4c3a),
	.w2(32'h3c2473c5),
	.w3(32'hbb99e341),
	.w4(32'h3b4644c5),
	.w5(32'h3b5eb205),
	.w6(32'hbc0bd612),
	.w7(32'hbb285dd6),
	.w8(32'h3b74f03b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5a3b4),
	.w1(32'h3c3ed725),
	.w2(32'h3c2bed61),
	.w3(32'h39e5ffe1),
	.w4(32'h3c644636),
	.w5(32'h3c2832ed),
	.w6(32'hbb100da3),
	.w7(32'h3b699923),
	.w8(32'hbb17e70b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c077d08),
	.w1(32'hbb5de505),
	.w2(32'h39f2f980),
	.w3(32'h3c2c9297),
	.w4(32'hbb33847b),
	.w5(32'hbaf94c6c),
	.w6(32'h3b143c12),
	.w7(32'hb8d11e85),
	.w8(32'h3b211abf),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b1a34),
	.w1(32'hbbc6b000),
	.w2(32'h3ac373c6),
	.w3(32'h3b8181f5),
	.w4(32'hba994b59),
	.w5(32'hb9e2fa57),
	.w6(32'h3bc47e0c),
	.w7(32'h3aa014c1),
	.w8(32'h39a4664e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad98a85),
	.w1(32'h3bfc762f),
	.w2(32'h3c48b229),
	.w3(32'hba262e9d),
	.w4(32'h3c2f09f6),
	.w5(32'h3c5ea3a2),
	.w6(32'hbb03d0a9),
	.w7(32'hbb122f6b),
	.w8(32'hbb32d7ee),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f4012),
	.w1(32'h3b0ce7b9),
	.w2(32'h3bc97c63),
	.w3(32'h3ca0110f),
	.w4(32'h3b276eac),
	.w5(32'hbbe5c2dd),
	.w6(32'h3bbc1378),
	.w7(32'h3c23da9b),
	.w8(32'h3b93ab63),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e5c8a),
	.w1(32'h3c67e3bc),
	.w2(32'h3ae224dd),
	.w3(32'hbc16b204),
	.w4(32'h3c099e52),
	.w5(32'h3b960f84),
	.w6(32'h3adb33e5),
	.w7(32'h3c0da08d),
	.w8(32'hb9fb59cb),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22fa4c),
	.w1(32'h3b6df281),
	.w2(32'hbaacbe94),
	.w3(32'hba5a9798),
	.w4(32'hbbefdc22),
	.w5(32'hbc0f1c4d),
	.w6(32'hbb27c656),
	.w7(32'h3a5475c2),
	.w8(32'h3b5a6684),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eaade),
	.w1(32'h3a382710),
	.w2(32'h3b71bbe9),
	.w3(32'hbc201b9c),
	.w4(32'hbb5636b0),
	.w5(32'h39765ca4),
	.w6(32'h3b9134de),
	.w7(32'hbb682424),
	.w8(32'h3b0b08e7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3cf5d),
	.w1(32'hbb00ffca),
	.w2(32'hbb61d83a),
	.w3(32'h3b3f5708),
	.w4(32'hbb3c2231),
	.w5(32'hbc44ef70),
	.w6(32'h3b189174),
	.w7(32'hb7c94eaa),
	.w8(32'h3ac63a87),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00ffa6),
	.w1(32'hbb7463ba),
	.w2(32'hbbaa3cb7),
	.w3(32'hbc0f9b7c),
	.w4(32'hba9e886c),
	.w5(32'hbb563e01),
	.w6(32'hbbcab6b1),
	.w7(32'hb700d28e),
	.w8(32'h392342f0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83d5d8),
	.w1(32'h3993d4a7),
	.w2(32'h3b7598e1),
	.w3(32'hbba8821e),
	.w4(32'hbb409823),
	.w5(32'hbb0cc943),
	.w6(32'h3afc81ad),
	.w7(32'h3994059e),
	.w8(32'h3b7857d9),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77a344),
	.w1(32'hbbd31793),
	.w2(32'hbb5479a4),
	.w3(32'hbb6029f0),
	.w4(32'hba2e342c),
	.w5(32'hbaddfb50),
	.w6(32'h3a0d96f6),
	.w7(32'hbb3bc9d9),
	.w8(32'hba9e9f6f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae753b8),
	.w1(32'hbbb52357),
	.w2(32'hbb3474b4),
	.w3(32'hba67ed7e),
	.w4(32'h3b7555c2),
	.w5(32'h38fe7cdf),
	.w6(32'hbbba7d48),
	.w7(32'h3b7e7303),
	.w8(32'h3c634a5a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbce146),
	.w1(32'hbc3f298e),
	.w2(32'hbc31a6e2),
	.w3(32'h3b860848),
	.w4(32'hbbda3788),
	.w5(32'hbb194670),
	.w6(32'h3bf7c06c),
	.w7(32'h3af8697b),
	.w8(32'h3c4b0bdb),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ee7cd),
	.w1(32'h3bbf62d5),
	.w2(32'h3b4af1f1),
	.w3(32'h3a9a6692),
	.w4(32'h3b3d4e20),
	.w5(32'h3be57a31),
	.w6(32'h3bde9880),
	.w7(32'hbbf52f87),
	.w8(32'hbc47c405),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e44b3),
	.w1(32'h3c16530a),
	.w2(32'h3bd1dc8a),
	.w3(32'h3b5978e5),
	.w4(32'h3c3614bb),
	.w5(32'h3b4b146b),
	.w6(32'hbbce74ab),
	.w7(32'h3bc03893),
	.w8(32'hbb8062f3),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e1c2e),
	.w1(32'h3bd4e594),
	.w2(32'h3ab6f0a4),
	.w3(32'hbad8bbda),
	.w4(32'h3bbc4a2f),
	.w5(32'h3b2106be),
	.w6(32'hbb2b7152),
	.w7(32'h3c0f8317),
	.w8(32'h3bb07b63),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04c242),
	.w1(32'hbaa6018b),
	.w2(32'hbb5983c7),
	.w3(32'h3b6503fc),
	.w4(32'h3bcfccd9),
	.w5(32'hbbb77892),
	.w6(32'h3a1393a1),
	.w7(32'h3bb56724),
	.w8(32'hbb242c54),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad87ba),
	.w1(32'h3c2b793f),
	.w2(32'h3c637837),
	.w3(32'hb94f1c40),
	.w4(32'hbc426498),
	.w5(32'hbabca1b5),
	.w6(32'h3b6e5eb1),
	.w7(32'hbc20e866),
	.w8(32'h3aaf3507),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c705ea1),
	.w1(32'hbba3ac35),
	.w2(32'hbbc461ae),
	.w3(32'h3c5923bb),
	.w4(32'h3b00b92c),
	.w5(32'hbbe0c02b),
	.w6(32'h3b8d0926),
	.w7(32'h3b122f5b),
	.w8(32'hbb25ae1e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdaaa80),
	.w1(32'hbc064a48),
	.w2(32'hbc6df1eb),
	.w3(32'hbbb84c9f),
	.w4(32'h3c0d92ca),
	.w5(32'h3cacffb2),
	.w6(32'hbb9c2b39),
	.w7(32'hbbc7b389),
	.w8(32'hbc6beaa3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13cdc3),
	.w1(32'h3c1cb32b),
	.w2(32'h3b3601e7),
	.w3(32'h3c3bdbb5),
	.w4(32'h3c01a2d8),
	.w5(32'h393fc401),
	.w6(32'hbbd39ff2),
	.w7(32'hb9f4be3c),
	.w8(32'hbc1a2ae4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb070725),
	.w1(32'hbb3919fa),
	.w2(32'h3ba37c8b),
	.w3(32'h3a0a05de),
	.w4(32'h3c10717e),
	.w5(32'h3c5d5a9e),
	.w6(32'hbb8c005b),
	.w7(32'hbb568f04),
	.w8(32'h3aa72e5d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71c0e6),
	.w1(32'hbbcb8c30),
	.w2(32'hbb9860c4),
	.w3(32'h3c28776e),
	.w4(32'hbc063c8f),
	.w5(32'h3a0c8cf6),
	.w6(32'h3bf8106d),
	.w7(32'hbad04858),
	.w8(32'hbb58601d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9ba92),
	.w1(32'hbbe0cddd),
	.w2(32'hbc0496f6),
	.w3(32'hba040f23),
	.w4(32'hbb43e3cf),
	.w5(32'hbc126841),
	.w6(32'hbb033f61),
	.w7(32'hbb1d0a59),
	.w8(32'hbbdd49cf),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcfc58),
	.w1(32'hba68e519),
	.w2(32'h3b391e8e),
	.w3(32'hbb648f68),
	.w4(32'hbbc1e90d),
	.w5(32'hbbfe397f),
	.w6(32'hbbdf4c19),
	.w7(32'hba4858de),
	.w8(32'h3a33cad6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9360184),
	.w1(32'h3c730097),
	.w2(32'h3c52b9bd),
	.w3(32'hbbead7f8),
	.w4(32'h3c5f20cc),
	.w5(32'h3c0c8ce5),
	.w6(32'h3a70f6cc),
	.w7(32'hbb40dfa9),
	.w8(32'hbc170fde),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ea277),
	.w1(32'hb945f75f),
	.w2(32'hbb46b541),
	.w3(32'h3be2144d),
	.w4(32'hbbf2c41b),
	.w5(32'hbc6b8602),
	.w6(32'hbc53cc10),
	.w7(32'h3a1695e8),
	.w8(32'h37a63ff8),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ffe76),
	.w1(32'hbafbc6df),
	.w2(32'h3a3bf5fb),
	.w3(32'hbb603de2),
	.w4(32'h3b346ede),
	.w5(32'h3c637eb1),
	.w6(32'h3b6d160a),
	.w7(32'hbb9831c4),
	.w8(32'h3ae2a750),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91f47e),
	.w1(32'h3b2677a7),
	.w2(32'h3c0076f1),
	.w3(32'h3bad799a),
	.w4(32'h3bbfbed5),
	.w5(32'h3c69acde),
	.w6(32'hbbe25484),
	.w7(32'hbaf9d7dc),
	.w8(32'hbb2809bd),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02562a),
	.w1(32'hbb09bf1f),
	.w2(32'hba586889),
	.w3(32'h3bc3c658),
	.w4(32'hbb20e920),
	.w5(32'h3b4d95a8),
	.w6(32'hbb2edc22),
	.w7(32'hb95842ae),
	.w8(32'h3b1332d3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a615d00),
	.w1(32'h3a149923),
	.w2(32'h3b30dd36),
	.w3(32'h3bc0ba64),
	.w4(32'hbb06ee59),
	.w5(32'hbb75baf3),
	.w6(32'h3b97cc99),
	.w7(32'hbb9cc1a0),
	.w8(32'hbb63c8a6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7e68f),
	.w1(32'hbcb2309a),
	.w2(32'hbccf7cd8),
	.w3(32'hbb83df8e),
	.w4(32'hbbb52afe),
	.w5(32'hbbc10c15),
	.w6(32'hbb2ee1b4),
	.w7(32'h3ca338e5),
	.w8(32'h3cac04fc),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9445ed),
	.w1(32'hbcdbb3eb),
	.w2(32'hbd03fa80),
	.w3(32'h3b1a3e15),
	.w4(32'h3a85a322),
	.w5(32'hbc3c7df4),
	.w6(32'h3cae4f77),
	.w7(32'h3d054159),
	.w8(32'h3cdb0934),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfc2569),
	.w1(32'hbc10b1a8),
	.w2(32'hbb9f458d),
	.w3(32'hbc3957ce),
	.w4(32'hb9d74047),
	.w5(32'hbc39443c),
	.w6(32'h3c9f06d2),
	.w7(32'h39caf11b),
	.w8(32'hbb3a10aa),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b488418),
	.w1(32'h3b02a610),
	.w2(32'h3c332b94),
	.w3(32'hbb88c085),
	.w4(32'h3c54d375),
	.w5(32'h3aa62f1b),
	.w6(32'h3a84ccc2),
	.w7(32'h3b90caea),
	.w8(32'h3a39ccb4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5151c4),
	.w1(32'h39f23e77),
	.w2(32'h3b0a3659),
	.w3(32'h3c4848a6),
	.w4(32'hbb914622),
	.w5(32'hbb12bd1d),
	.w6(32'h3b335bda),
	.w7(32'hbb60ab63),
	.w8(32'h3aeb53cb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c6e81),
	.w1(32'hbb6f9a1c),
	.w2(32'h3c00a6b4),
	.w3(32'hbac72c1e),
	.w4(32'hbb1345f5),
	.w5(32'h3bff665a),
	.w6(32'h3b8b5f82),
	.w7(32'h3b046ba9),
	.w8(32'h3bbca8f1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f8962),
	.w1(32'h3bae6fca),
	.w2(32'h3bf96a64),
	.w3(32'h3b034915),
	.w4(32'h3c07c3b3),
	.w5(32'h3c168efd),
	.w6(32'h3bb59dd0),
	.w7(32'h3b9b6536),
	.w8(32'h3c0fb8c4),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babfdd1),
	.w1(32'h3a783d50),
	.w2(32'hbb33ec4e),
	.w3(32'h3bc77760),
	.w4(32'h3c0530ed),
	.w5(32'hbb719ab3),
	.w6(32'h3b5a8293),
	.w7(32'h3c23c701),
	.w8(32'h3c0324d2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24cc9c),
	.w1(32'h3bd8f928),
	.w2(32'h3c37ed41),
	.w3(32'hbbaaeba2),
	.w4(32'hbbc4c340),
	.w5(32'hbc7c373a),
	.w6(32'h3be01d65),
	.w7(32'h3b56154b),
	.w8(32'h3b0e1739),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5409c),
	.w1(32'h3bd7dc80),
	.w2(32'h3bbd68f8),
	.w3(32'hbbd55ca2),
	.w4(32'h3b8167f3),
	.w5(32'hbafdfcf8),
	.w6(32'hba511656),
	.w7(32'h3b6c44ed),
	.w8(32'hbb189d2b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5317d),
	.w1(32'h3b4a5029),
	.w2(32'hbb1318db),
	.w3(32'h3b9b2b0c),
	.w4(32'h3c0dfad7),
	.w5(32'hbb4b47ac),
	.w6(32'hbbb3ef01),
	.w7(32'hbb330b47),
	.w8(32'hbc5d74aa),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae61dca),
	.w1(32'hbc0a0a06),
	.w2(32'hbbb7af91),
	.w3(32'hb7a7123c),
	.w4(32'hbc193aaf),
	.w5(32'hbbd4e512),
	.w6(32'hbb602331),
	.w7(32'hbadac291),
	.w8(32'h3961808f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb562fa5),
	.w1(32'hbaec296a),
	.w2(32'hbb1755da),
	.w3(32'hbbd94316),
	.w4(32'h3bae91b4),
	.w5(32'h3bd274f1),
	.w6(32'hbb668c9e),
	.w7(32'hbc025b82),
	.w8(32'hbc34f3b3),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b024563),
	.w1(32'hb9d2ccce),
	.w2(32'hb940d546),
	.w3(32'h3b693411),
	.w4(32'hbb6372b2),
	.w5(32'h3b3635b3),
	.w6(32'hbb957e59),
	.w7(32'hbb6a398e),
	.w8(32'h3b3b9134),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ba8db),
	.w1(32'hbbf9e61c),
	.w2(32'hbb855cc4),
	.w3(32'h3c2118eb),
	.w4(32'hbc70e180),
	.w5(32'hbc6eadfd),
	.w6(32'h3b3b74dd),
	.w7(32'h3b1e3632),
	.w8(32'h3c774497),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96287e),
	.w1(32'hbaa795f1),
	.w2(32'h3a97032e),
	.w3(32'hbc060966),
	.w4(32'hbc58bc68),
	.w5(32'hbccf86c8),
	.w6(32'h3c5b8fc9),
	.w7(32'hbbb4d8a3),
	.w8(32'hbc14c954),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe4f0d),
	.w1(32'h3a42d892),
	.w2(32'hbba712f4),
	.w3(32'hbcbdfd9a),
	.w4(32'h3ae5c415),
	.w5(32'hbc13475c),
	.w6(32'hbc45489d),
	.w7(32'hba1acc58),
	.w8(32'hbbc1eaf1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc046e15),
	.w1(32'hbaa47312),
	.w2(32'hbae6fad8),
	.w3(32'hbb123b5b),
	.w4(32'hba201cca),
	.w5(32'h3ab44445),
	.w6(32'hbbf8fefd),
	.w7(32'hba8c09b3),
	.w8(32'h390f863b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33f3e5),
	.w1(32'hbaf0bba5),
	.w2(32'hb9a65d69),
	.w3(32'hbab6db22),
	.w4(32'hbada6396),
	.w5(32'hb8d690fb),
	.w6(32'hbad95fcc),
	.w7(32'hbb13c12b),
	.w8(32'hbabd6add),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07e608),
	.w1(32'hbaa281f8),
	.w2(32'hb980b32c),
	.w3(32'hbab8c42f),
	.w4(32'hba83aecb),
	.w5(32'hbb952b53),
	.w6(32'h3a82a215),
	.w7(32'hba9c29a7),
	.w8(32'hba7182a6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12c653),
	.w1(32'h3988052d),
	.w2(32'hba2fd66f),
	.w3(32'hba9b5080),
	.w4(32'h3b9d1302),
	.w5(32'hb9b6ebae),
	.w6(32'h3a87a90b),
	.w7(32'h3a9c15d4),
	.w8(32'hba92b92b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada0da4),
	.w1(32'hbb0d4c10),
	.w2(32'h396e4704),
	.w3(32'hbb89006a),
	.w4(32'h394bfae3),
	.w5(32'hba50e23f),
	.w6(32'hbb12fc61),
	.w7(32'hba953867),
	.w8(32'hb888710f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94300f7),
	.w1(32'h3b0add95),
	.w2(32'h3b4e903c),
	.w3(32'hbacc424d),
	.w4(32'h3b10da3e),
	.w5(32'h3a738402),
	.w6(32'h3aa5ae6b),
	.w7(32'h39b826d2),
	.w8(32'h3ad05303),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e373f),
	.w1(32'hbb24afd0),
	.w2(32'hbb0301d4),
	.w3(32'hbbbd6919),
	.w4(32'hbb7d0b27),
	.w5(32'hbb75750d),
	.w6(32'hba6d6d89),
	.w7(32'h3aaf187b),
	.w8(32'hb9b65d4c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb292eff),
	.w1(32'hbb4b5df6),
	.w2(32'hbad45c9d),
	.w3(32'hbb22acc4),
	.w4(32'hbb67740d),
	.w5(32'hbb4035d5),
	.w6(32'hb7f8c7d8),
	.w7(32'hbb11b1c8),
	.w8(32'hba7ad693),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51d25c),
	.w1(32'hbb8f38b1),
	.w2(32'hbb3a6f79),
	.w3(32'hbb02840e),
	.w4(32'hbb1b5a91),
	.w5(32'hba451b4f),
	.w6(32'hbb17edc8),
	.w7(32'hbb3cfabe),
	.w8(32'h3aaf195a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64a565),
	.w1(32'hbacb5eaa),
	.w2(32'hbb1af0d9),
	.w3(32'hbb882b9b),
	.w4(32'hba79e40d),
	.w5(32'hbb583aec),
	.w6(32'h3ae7fd3a),
	.w7(32'h3a6309d2),
	.w8(32'hbab4b1a7),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccec9b),
	.w1(32'hbb05f609),
	.w2(32'hbb0a3d18),
	.w3(32'hb91b3bb5),
	.w4(32'hb9ffc88d),
	.w5(32'hbbc42524),
	.w6(32'h3a83c5e1),
	.w7(32'h3903f6a0),
	.w8(32'hbb678fd1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca14c5),
	.w1(32'h3ba18b97),
	.w2(32'h3b34563e),
	.w3(32'hbaa609c1),
	.w4(32'h3b85c97a),
	.w5(32'h3a91d616),
	.w6(32'hbb30a64f),
	.w7(32'h3ba36631),
	.w8(32'h3b45cd0c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fcce0),
	.w1(32'h397ab9e6),
	.w2(32'h39bbc896),
	.w3(32'h3b741a4c),
	.w4(32'h3afb00fa),
	.w5(32'h3ac99694),
	.w6(32'h3b6caf00),
	.w7(32'h3b3b30ad),
	.w8(32'h3b375a86),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e6136),
	.w1(32'hbabf085f),
	.w2(32'h3a847042),
	.w3(32'h3add4e1a),
	.w4(32'hba7f412f),
	.w5(32'hba957231),
	.w6(32'h3aa6f09b),
	.w7(32'hba13b7cd),
	.w8(32'hbaffaa15),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d91ed),
	.w1(32'h3ad12123),
	.w2(32'h3accba69),
	.w3(32'hbbdd78f9),
	.w4(32'hbb061095),
	.w5(32'h3bce4bd5),
	.w6(32'hbb9b29eb),
	.w7(32'hbb1c4539),
	.w8(32'hbba646b4),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfcc05),
	.w1(32'h3b257048),
	.w2(32'h3b990134),
	.w3(32'hba64dfd2),
	.w4(32'h3b9c1fdf),
	.w5(32'h3bc66140),
	.w6(32'h3ac23e5f),
	.w7(32'h3b83a6f0),
	.w8(32'h3b9b21ce),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba557434),
	.w1(32'hbb9cb39d),
	.w2(32'hbb61e2b4),
	.w3(32'hbadc0085),
	.w4(32'hbba9a524),
	.w5(32'hba164b7a),
	.w6(32'h3ab52f8f),
	.w7(32'hbb3f513c),
	.w8(32'hbb320781),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe19696),
	.w1(32'hbbd0ea3f),
	.w2(32'hb8bfccf6),
	.w3(32'hbbc5e36c),
	.w4(32'hbbe93394),
	.w5(32'hbb5126b2),
	.w6(32'hbb7040c4),
	.w7(32'h3b1754a5),
	.w8(32'h3b92d658),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba771300),
	.w1(32'h3b001b67),
	.w2(32'h3aadc1c2),
	.w3(32'h3891378b),
	.w4(32'h3b2989c9),
	.w5(32'h3b26d421),
	.w6(32'hba89e532),
	.w7(32'h3a60a32e),
	.w8(32'h3937e92d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0408aa),
	.w1(32'hb99cd5db),
	.w2(32'hba76ba0a),
	.w3(32'hb9de262e),
	.w4(32'hbae5cd95),
	.w5(32'hbab70294),
	.w6(32'h3a7b715b),
	.w7(32'hbaf007da),
	.w8(32'hbb8b1104),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb68187),
	.w1(32'hbb6cd36e),
	.w2(32'h3bd18237),
	.w3(32'hbbaeffcf),
	.w4(32'hbb150a25),
	.w5(32'h3c51ab59),
	.w6(32'hbbf016e5),
	.w7(32'hbb862953),
	.w8(32'h3bff8755),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cb32cb),
	.w1(32'h39f3a09b),
	.w2(32'h3b276094),
	.w3(32'hba6e478c),
	.w4(32'h3b2bcfc2),
	.w5(32'h3aa81408),
	.w6(32'hbb76ded0),
	.w7(32'h3b1c90b4),
	.w8(32'hbb20299f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2642ad),
	.w1(32'hbb3f2c0f),
	.w2(32'h3911d4c8),
	.w3(32'hbb39e04a),
	.w4(32'hbb1953c3),
	.w5(32'h3b884283),
	.w6(32'hbb6f42c1),
	.w7(32'hbb9287c8),
	.w8(32'h3ac64a9b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c0d42),
	.w1(32'hbaa06fa3),
	.w2(32'hb9c72616),
	.w3(32'hbb070295),
	.w4(32'hbb2080c8),
	.w5(32'h3a2a2a08),
	.w6(32'h398fdf51),
	.w7(32'hbaa54589),
	.w8(32'hba0315a1),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20d662),
	.w1(32'hbaa0433e),
	.w2(32'hba5f21cb),
	.w3(32'hba1e9f6d),
	.w4(32'hbaa63439),
	.w5(32'hbae56ac3),
	.w6(32'h3b14c587),
	.w7(32'hba2777ac),
	.w8(32'hbb252b19),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89f8183),
	.w1(32'h3aca2d14),
	.w2(32'h3a4450a4),
	.w3(32'h39486fca),
	.w4(32'hbb066a46),
	.w5(32'hbaf92b8c),
	.w6(32'hba0a0330),
	.w7(32'hbaddcf67),
	.w8(32'hba81d7d5),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92c28a),
	.w1(32'hbb150d73),
	.w2(32'h39e57c96),
	.w3(32'hbb861a01),
	.w4(32'hbb0bc311),
	.w5(32'hbb45f70a),
	.w6(32'hba1a1c19),
	.w7(32'hbb578ff6),
	.w8(32'hbb88c195),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb150ca),
	.w1(32'hb7192800),
	.w2(32'hb92c0dd1),
	.w3(32'hbbc186d4),
	.w4(32'h38e5fbed),
	.w5(32'h3a62475a),
	.w6(32'hbb4b27ac),
	.w7(32'h3a39cd42),
	.w8(32'hb98f5247),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f2ccf),
	.w1(32'hb921ce72),
	.w2(32'hbb043ae2),
	.w3(32'hbb4458d0),
	.w4(32'hba39bba8),
	.w5(32'hbadcbe5b),
	.w6(32'h3985c549),
	.w7(32'hbac567e0),
	.w8(32'h38d2dd8f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5785b8),
	.w1(32'h3b41353e),
	.w2(32'h3b5d49b5),
	.w3(32'hba312407),
	.w4(32'h3b37378c),
	.w5(32'h3bcebd27),
	.w6(32'hba61062f),
	.w7(32'h3abeaab9),
	.w8(32'h3b6c6946),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbdc93),
	.w1(32'h3acd4247),
	.w2(32'hba272715),
	.w3(32'hb9b11b62),
	.w4(32'hbb163b16),
	.w5(32'hbab4f768),
	.w6(32'hbaa1ab6c),
	.w7(32'hbaaf753c),
	.w8(32'hbb1b6a2a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59cf79),
	.w1(32'hba17bb8c),
	.w2(32'h3a03b7ae),
	.w3(32'hbb59e42e),
	.w4(32'hba2454e7),
	.w5(32'h3a54d1ea),
	.w6(32'hbb631901),
	.w7(32'h39bb0387),
	.w8(32'h39ef6ce9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0775f2),
	.w1(32'h39ed49ed),
	.w2(32'h39d4bd94),
	.w3(32'hbac4e3ac),
	.w4(32'h38b10a73),
	.w5(32'h3b14f21f),
	.w6(32'h3ab1a4a9),
	.w7(32'h39212afc),
	.w8(32'h3b3ff1ae),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ea7aa),
	.w1(32'h39f4668b),
	.w2(32'h3b694db2),
	.w3(32'h3a12b10c),
	.w4(32'hb9efdb2a),
	.w5(32'h3a84a87e),
	.w6(32'h39d8e266),
	.w7(32'h389e4a5b),
	.w8(32'h3ad2983a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9165fd2),
	.w1(32'h3b4ebae8),
	.w2(32'h3b83b289),
	.w3(32'hb99982f6),
	.w4(32'h3b85835a),
	.w5(32'h3b4397e5),
	.w6(32'h3a4fca0f),
	.w7(32'h3b04d668),
	.w8(32'h3bb5a9ab),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2313d5),
	.w1(32'h3b15421d),
	.w2(32'h3b4e7bd4),
	.w3(32'hbb0c68c5),
	.w4(32'hb97f2606),
	.w5(32'hba669b08),
	.w6(32'h3a4ab1a9),
	.w7(32'h3a127c49),
	.w8(32'hba5817ae),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af51569),
	.w1(32'h3b3fa535),
	.w2(32'h3b15c259),
	.w3(32'hbb2acf2f),
	.w4(32'hb7dcc53a),
	.w5(32'h3aab8e1e),
	.w6(32'hbb01ee5e),
	.w7(32'hb968dd68),
	.w8(32'h3aefb5f8),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eafa73),
	.w1(32'h3a84561e),
	.w2(32'h3b03adf7),
	.w3(32'h3a967792),
	.w4(32'h3b1e0fd6),
	.w5(32'hb9d27737),
	.w6(32'hbadd431a),
	.w7(32'h3b173405),
	.w8(32'h3a5a1cf5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40970e),
	.w1(32'hba889017),
	.w2(32'hb6438316),
	.w3(32'h39d49eb2),
	.w4(32'hba42970c),
	.w5(32'h3b47ba1b),
	.w6(32'h3a50336a),
	.w7(32'hb9fdee6a),
	.w8(32'h3a07b23e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9836f1e),
	.w1(32'h3b1b6575),
	.w2(32'h3b5b6cca),
	.w3(32'h3adef3db),
	.w4(32'h39db9455),
	.w5(32'h3b174634),
	.w6(32'h38daa35a),
	.w7(32'h3ab406a2),
	.w8(32'h3aef78be),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba5448),
	.w1(32'hba8c3c93),
	.w2(32'hbb1d0990),
	.w3(32'h39549f7a),
	.w4(32'hbb361113),
	.w5(32'hb8c4773b),
	.w6(32'h3ae9cece),
	.w7(32'hbb2b2d77),
	.w8(32'hba537ff7),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e031c),
	.w1(32'hba02174f),
	.w2(32'hba6feab7),
	.w3(32'hbaf8fab1),
	.w4(32'h3839284f),
	.w5(32'hba555c7d),
	.w6(32'hb89db020),
	.w7(32'hb9f986a1),
	.w8(32'hbafaeb3c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc5f32),
	.w1(32'hbb5513e6),
	.w2(32'hbb0a0a83),
	.w3(32'h3b036aeb),
	.w4(32'hbb1c8d01),
	.w5(32'hbba3772d),
	.w6(32'hba358e38),
	.w7(32'h3a8249f9),
	.w8(32'h391eef4f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb266d0e),
	.w1(32'hba29157a),
	.w2(32'h3b2301f0),
	.w3(32'hbb65c97b),
	.w4(32'h3adb3c65),
	.w5(32'h3a0c6b47),
	.w6(32'hbb7b3557),
	.w7(32'h3a56de95),
	.w8(32'h3b127967),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0f5d7),
	.w1(32'h39c56d25),
	.w2(32'h3aa31fc9),
	.w3(32'hba7c39bd),
	.w4(32'hb9a76b4a),
	.w5(32'h3a5cf7d3),
	.w6(32'hb9e2f642),
	.w7(32'h3ac57072),
	.w8(32'h3b254f5e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9536943),
	.w1(32'h3a12d351),
	.w2(32'h3af92025),
	.w3(32'hbb5358d5),
	.w4(32'hbb00d572),
	.w5(32'h3ae7842b),
	.w6(32'hb970b79e),
	.w7(32'hbb2ab218),
	.w8(32'hb89f791a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef3736),
	.w1(32'hba416467),
	.w2(32'hbab4d2e8),
	.w3(32'h3ae5e811),
	.w4(32'hbb0e2d55),
	.w5(32'hbab25d37),
	.w6(32'h3aeca045),
	.w7(32'hbb069d1d),
	.w8(32'hba7111c2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba410762),
	.w1(32'h3a8555e7),
	.w2(32'hba84d4e1),
	.w3(32'hb98c0025),
	.w4(32'hba05c236),
	.w5(32'h3b072b6d),
	.w6(32'hba572f94),
	.w7(32'h3a082821),
	.w8(32'hb92b2def),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf666d1),
	.w1(32'h3ac62044),
	.w2(32'h3b66a01b),
	.w3(32'hba12ff2d),
	.w4(32'h3a3aecb8),
	.w5(32'h3a3a4197),
	.w6(32'hba73bdf7),
	.w7(32'hbad9a5c3),
	.w8(32'h3a71a7c3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ca2d0),
	.w1(32'h3b128ceb),
	.w2(32'h3ba80069),
	.w3(32'h3ae1e275),
	.w4(32'h3b50872f),
	.w5(32'h3aafd1b5),
	.w6(32'hb9a731d4),
	.w7(32'h3b04cc8c),
	.w8(32'h3b38e3a0),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6110f5),
	.w1(32'hbad8d896),
	.w2(32'hbada7841),
	.w3(32'hb96cf17e),
	.w4(32'hba873e0b),
	.w5(32'hba33ddaa),
	.w6(32'h3b234676),
	.w7(32'hba39ff7e),
	.w8(32'hb8963f67),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade541f),
	.w1(32'hba18439f),
	.w2(32'hbaa2703e),
	.w3(32'hbac9cdc7),
	.w4(32'hba7155e4),
	.w5(32'h3a335db4),
	.w6(32'h3a1b8da1),
	.w7(32'h390a33e7),
	.w8(32'hbae3910e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40a736),
	.w1(32'h3a02379a),
	.w2(32'hbab26d19),
	.w3(32'hbb273f0d),
	.w4(32'hbb6074fd),
	.w5(32'hb9f7803c),
	.w6(32'hbb11b628),
	.w7(32'hbb06052a),
	.w8(32'hbab4106e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96e6c9),
	.w1(32'h3a0b918f),
	.w2(32'hb9b69553),
	.w3(32'hba977db9),
	.w4(32'hba1a732a),
	.w5(32'hbaf5f4ce),
	.w6(32'hba4a9e54),
	.w7(32'hba3fff82),
	.w8(32'hbb441b41),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49e03b),
	.w1(32'h3a0949d1),
	.w2(32'h39a4c165),
	.w3(32'hbb7681fc),
	.w4(32'hbad7f1d0),
	.w5(32'h3a5c0e73),
	.w6(32'hbb608927),
	.w7(32'hba052bab),
	.w8(32'h39d133dc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25f006),
	.w1(32'hb9dc5dd8),
	.w2(32'hba34b349),
	.w3(32'hbb07318d),
	.w4(32'hbb1764ef),
	.w5(32'hbaf63598),
	.w6(32'hba4e86b0),
	.w7(32'hb8953aa1),
	.w8(32'hb8f3955b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0a08a),
	.w1(32'hba45bb7e),
	.w2(32'h3b1beffc),
	.w3(32'hba08f645),
	.w4(32'hba4f83b6),
	.w5(32'hbb4dcf70),
	.w6(32'h3b3eccdd),
	.w7(32'h3b8aed24),
	.w8(32'h3b870dc5),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ded99),
	.w1(32'hbb30c700),
	.w2(32'hbb32e7f5),
	.w3(32'hbafdd8d4),
	.w4(32'hbb1d8ba4),
	.w5(32'hba8d6087),
	.w6(32'hba281eae),
	.w7(32'hbb46c9d4),
	.w8(32'h385e827f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb131a3c),
	.w1(32'hbb33090f),
	.w2(32'hba94cd78),
	.w3(32'hbb822f22),
	.w4(32'hbba4c783),
	.w5(32'h3b0359a5),
	.w6(32'h3a4f68a8),
	.w7(32'hbaf99fd1),
	.w8(32'hbb5e4cbc),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule