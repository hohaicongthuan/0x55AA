module layer_10_featuremap_252(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38930381),
	.w1(32'h3a07eb6a),
	.w2(32'hb9494053),
	.w3(32'hb9afe6d3),
	.w4(32'hbadecb6e),
	.w5(32'h3b03800b),
	.w6(32'h39e412c4),
	.w7(32'hb9be8476),
	.w8(32'h3a2b9f0e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4649c),
	.w1(32'hba0e12ff),
	.w2(32'h385822f6),
	.w3(32'h3a6600b6),
	.w4(32'h3af37878),
	.w5(32'hbaf759db),
	.w6(32'h3adc5482),
	.w7(32'h3a0d958f),
	.w8(32'hbacaebf0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fad618),
	.w1(32'h38d9a70d),
	.w2(32'hbaa08739),
	.w3(32'hbb28d76d),
	.w4(32'hbb1a38c2),
	.w5(32'h39889e73),
	.w6(32'h3ab963f7),
	.w7(32'h3aa29416),
	.w8(32'h3a32ab4b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a059d97),
	.w1(32'h3a04b0cf),
	.w2(32'h396a3cfe),
	.w3(32'h3a2efbb6),
	.w4(32'h398b0585),
	.w5(32'hb89e00f9),
	.w6(32'hb8881863),
	.w7(32'hb88346ed),
	.w8(32'hbb3df377),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9780b2),
	.w1(32'hbabf1541),
	.w2(32'hbac64866),
	.w3(32'h39962e34),
	.w4(32'h3a1010a8),
	.w5(32'h3a92105a),
	.w6(32'hbb0f79b1),
	.w7(32'hba80c671),
	.w8(32'h3a9b449e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25e226),
	.w1(32'h3a387b03),
	.w2(32'h3a124a03),
	.w3(32'h3aa0a3fb),
	.w4(32'h3a4fda0f),
	.w5(32'h3b34ce79),
	.w6(32'h3a72ca03),
	.w7(32'h399f5a2a),
	.w8(32'h3b08f3ab),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf858f),
	.w1(32'hbaac4f15),
	.w2(32'hbb2ee311),
	.w3(32'h3b343d7a),
	.w4(32'hb9d57ac5),
	.w5(32'hba8e5610),
	.w6(32'h3aff0363),
	.w7(32'hbab62393),
	.w8(32'hba63b907),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1470c4),
	.w1(32'h39b0d219),
	.w2(32'h3c00132c),
	.w3(32'hba3c322d),
	.w4(32'h3b074ae5),
	.w5(32'h3b5bcd00),
	.w6(32'h39165c07),
	.w7(32'h3b0eedaa),
	.w8(32'h3ae0d817),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff49d6),
	.w1(32'h3aa1f0fd),
	.w2(32'h3a81c27a),
	.w3(32'h3b08762d),
	.w4(32'h3ad319e9),
	.w5(32'h3a0bd093),
	.w6(32'h3b1458f5),
	.w7(32'h3b13c551),
	.w8(32'h38d0a7f4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba869e9c),
	.w1(32'hbaaa3e69),
	.w2(32'hbb34b06b),
	.w3(32'h3af45423),
	.w4(32'h3aa7568d),
	.w5(32'h3a6a2d6d),
	.w6(32'hbb2b9229),
	.w7(32'hb9d18f90),
	.w8(32'hbb03baa1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5cbb7),
	.w1(32'hba0ea7be),
	.w2(32'hb9935b7d),
	.w3(32'h3a1e73ae),
	.w4(32'hb92d29c0),
	.w5(32'h3a5c1691),
	.w6(32'h3906481c),
	.w7(32'hb88ecdd9),
	.w8(32'h3a00f42b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bcdf3),
	.w1(32'hba31bddc),
	.w2(32'hbb2bdb13),
	.w3(32'h3b59fdee),
	.w4(32'h3a7dd3b6),
	.w5(32'hbb18f4b0),
	.w6(32'h3b854015),
	.w7(32'h3a90b54d),
	.w8(32'hbb545973),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f46ed6),
	.w1(32'hba93c56b),
	.w2(32'hbb4af828),
	.w3(32'h3b082943),
	.w4(32'h3b1a4298),
	.w5(32'hb9604a3a),
	.w6(32'hb9e2867c),
	.w7(32'h3894d069),
	.w8(32'hbb298379),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafded83),
	.w1(32'hba8a959c),
	.w2(32'h3a9ba688),
	.w3(32'h3af79bd3),
	.w4(32'h3b50a00c),
	.w5(32'h3b7449e3),
	.w6(32'h3b34d87d),
	.w7(32'h3b634086),
	.w8(32'h3b5bfa27),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1ad93),
	.w1(32'hb98ff89e),
	.w2(32'hba1b51ab),
	.w3(32'hb8eb3e2b),
	.w4(32'h3ac43c8e),
	.w5(32'hb9e423b0),
	.w6(32'hbab812ec),
	.w7(32'hb9a47f95),
	.w8(32'hbaabbd9a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1d682),
	.w1(32'hba8143cd),
	.w2(32'h3a8490d5),
	.w3(32'hbb20c180),
	.w4(32'h3a8eda2b),
	.w5(32'h3bcc1043),
	.w6(32'hbb84cb31),
	.w7(32'hbae36da1),
	.w8(32'h3b21391a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac50b3c),
	.w1(32'h3abda4c4),
	.w2(32'h3a9d5e5d),
	.w3(32'h3ab44c63),
	.w4(32'h3aa6e9fa),
	.w5(32'hba29b0de),
	.w6(32'h3aedec48),
	.w7(32'h3a8c7b34),
	.w8(32'hba4cf478),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9efa2e),
	.w1(32'hbbaabe65),
	.w2(32'hbacab6d2),
	.w3(32'hbaec0bee),
	.w4(32'hbb193079),
	.w5(32'hbb05044c),
	.w6(32'hbb4dcfa5),
	.w7(32'hbb88a810),
	.w8(32'hbb518d51),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0618ad),
	.w1(32'hbb2a6d2a),
	.w2(32'hbaf286d9),
	.w3(32'hbac8ad4f),
	.w4(32'hbafff0ee),
	.w5(32'hb9ba2064),
	.w6(32'hbb50f53d),
	.w7(32'hbb46128d),
	.w8(32'hbb553d97),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984fdfb),
	.w1(32'hba8f9597),
	.w2(32'hbb035a11),
	.w3(32'h37bbfe23),
	.w4(32'hb7bceaf6),
	.w5(32'h368d2141),
	.w6(32'hba803702),
	.w7(32'hba6c2d16),
	.w8(32'hba43da3c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd6f9f),
	.w1(32'h390fbe13),
	.w2(32'hb9a6101f),
	.w3(32'h38a45ade),
	.w4(32'h39e56806),
	.w5(32'h3b002f04),
	.w6(32'h3a06818a),
	.w7(32'hb9e94e0a),
	.w8(32'h3b063fd4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16ad3d),
	.w1(32'h3b03839f),
	.w2(32'h3ac5a0cf),
	.w3(32'h3b1ae6c7),
	.w4(32'h3b2c0de1),
	.w5(32'h3a9ebead),
	.w6(32'h3af60cc2),
	.w7(32'h3b1e9a4a),
	.w8(32'h3a443638),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8e78f),
	.w1(32'h39ada146),
	.w2(32'hba1ecdee),
	.w3(32'hbb2f45c5),
	.w4(32'h3ab5ed1e),
	.w5(32'h3b073232),
	.w6(32'hbc003456),
	.w7(32'hbb5de119),
	.w8(32'hbbb56bf4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45af86),
	.w1(32'hba2371ad),
	.w2(32'hbb228bbf),
	.w3(32'h39bbc053),
	.w4(32'h39770ef6),
	.w5(32'hbaf371f1),
	.w6(32'hbb5cb4d9),
	.w7(32'hbad71122),
	.w8(32'hbb9269a0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c7884),
	.w1(32'hba537a7a),
	.w2(32'hbb247cc3),
	.w3(32'hbaadb3d6),
	.w4(32'h3a305fc6),
	.w5(32'hba05148d),
	.w6(32'hbaba9e54),
	.w7(32'hb994a121),
	.w8(32'hbb806d92),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ff0fa),
	.w1(32'h3abd23c4),
	.w2(32'h3a96c039),
	.w3(32'h3a8d32cf),
	.w4(32'h3ad298de),
	.w5(32'h3aadf507),
	.w6(32'hba383f91),
	.w7(32'h39990ffb),
	.w8(32'h3a413e93),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ffab9),
	.w1(32'h39b9b27c),
	.w2(32'h3a39b992),
	.w3(32'h39f42388),
	.w4(32'h3a597a50),
	.w5(32'hba3e15bb),
	.w6(32'h3989e207),
	.w7(32'h3a002114),
	.w8(32'hba6218ef),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4597d),
	.w1(32'h3b1d8327),
	.w2(32'hb92a3aee),
	.w3(32'h3aae3d83),
	.w4(32'h3b9ae5f7),
	.w5(32'h3aeff6fd),
	.w6(32'h3b6903d9),
	.w7(32'h3b80e61e),
	.w8(32'h3a2e96e6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c55911),
	.w1(32'hba4e2c1f),
	.w2(32'hba753266),
	.w3(32'h3b3af449),
	.w4(32'h3b017655),
	.w5(32'hb9f50be8),
	.w6(32'h3ae4ad8a),
	.w7(32'h3abdd7c1),
	.w8(32'hb95a9c1d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ee52d),
	.w1(32'h3a897948),
	.w2(32'hb9a9bdd3),
	.w3(32'hbb0b11c7),
	.w4(32'h3b1875d3),
	.w5(32'h3838006e),
	.w6(32'hbb36ef1f),
	.w7(32'h3a2fbe69),
	.w8(32'hbb09f2c0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36f23a),
	.w1(32'hbb1971d5),
	.w2(32'hbafbe48a),
	.w3(32'hbaa0652c),
	.w4(32'hba2a4e2c),
	.w5(32'hba7c7ad5),
	.w6(32'hbadc66d5),
	.w7(32'hbaba79a1),
	.w8(32'h3917beea),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba540d43),
	.w1(32'hbac6ce47),
	.w2(32'hba8aed8d),
	.w3(32'hba405ff8),
	.w4(32'hba2ebf60),
	.w5(32'hba05ad93),
	.w6(32'h3a4109f5),
	.w7(32'h3a2cd414),
	.w8(32'h3a83892c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce7e81),
	.w1(32'hba957ff1),
	.w2(32'hbacb5d7b),
	.w3(32'h3a402cfe),
	.w4(32'hba7a6832),
	.w5(32'hb9e1aaf7),
	.w6(32'hbaa886e2),
	.w7(32'h39b8c323),
	.w8(32'hbb419695),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dcb2a),
	.w1(32'hbb44ea2c),
	.w2(32'hbb186451),
	.w3(32'hbaafe0e6),
	.w4(32'hba336d0b),
	.w5(32'hba4dd0bc),
	.w6(32'hbb03bdcd),
	.w7(32'hbb17dcf1),
	.w8(32'h38a8f860),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95a43f),
	.w1(32'h3a325261),
	.w2(32'h3a5dab98),
	.w3(32'h3a031742),
	.w4(32'h3a01bf5a),
	.w5(32'hbab1b322),
	.w6(32'h3a0c54d2),
	.w7(32'h3a98b389),
	.w8(32'hbabd814b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e4e43),
	.w1(32'hbb2f2ad5),
	.w2(32'hbb38216c),
	.w3(32'hba901e3b),
	.w4(32'hbb1680e2),
	.w5(32'h3a515a88),
	.w6(32'hba6cf0e1),
	.w7(32'hbb3facb9),
	.w8(32'hbb2b3a4f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb842483),
	.w1(32'hbb959d02),
	.w2(32'hba2435fc),
	.w3(32'hbb121ddf),
	.w4(32'hbb584e74),
	.w5(32'hbaee7bd2),
	.w6(32'hbb6a889d),
	.w7(32'hbb670699),
	.w8(32'hbbb95ea3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb820658),
	.w1(32'h3ad42541),
	.w2(32'hbaa9fc8a),
	.w3(32'hbb547538),
	.w4(32'h3b00f360),
	.w5(32'hbaee29eb),
	.w6(32'hbb01e294),
	.w7(32'h391611cf),
	.w8(32'hbb32c7bc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39914c9a),
	.w1(32'hb8c0570a),
	.w2(32'hbb91b7fa),
	.w3(32'h39955d41),
	.w4(32'h3a85c259),
	.w5(32'hbadc28be),
	.w6(32'h3b4ef4f8),
	.w7(32'h3b3bc060),
	.w8(32'h3ab37454),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2269f),
	.w1(32'h39b6cb6d),
	.w2(32'hb9f2f696),
	.w3(32'hba155c98),
	.w4(32'hba27feab),
	.w5(32'hb8bc2a08),
	.w6(32'hb94604da),
	.w7(32'h38ff2a74),
	.w8(32'hb8a3a3a0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2522e),
	.w1(32'hb9db5cde),
	.w2(32'h3a2a0725),
	.w3(32'h39bff166),
	.w4(32'hba816877),
	.w5(32'h3b00a77e),
	.w6(32'hba7b11f1),
	.w7(32'hba0c8e9a),
	.w8(32'h3abfd51d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7a7e4),
	.w1(32'h3aca3f7f),
	.w2(32'h3a9f5272),
	.w3(32'h3af2e017),
	.w4(32'h3acfae7b),
	.w5(32'hbb11ac68),
	.w6(32'h3aae337d),
	.w7(32'h3ab283e3),
	.w8(32'hba62da47),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10e935),
	.w1(32'hba1c7b71),
	.w2(32'hb8e65ddd),
	.w3(32'h3a8f06c0),
	.w4(32'h3aa97df0),
	.w5(32'h3a8868ec),
	.w6(32'hb9d5a296),
	.w7(32'h3a49b1b1),
	.w8(32'h3ada86f1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4649b9),
	.w1(32'hb985ec16),
	.w2(32'h38b9d804),
	.w3(32'hba103ee7),
	.w4(32'h3b87ee47),
	.w5(32'h3ba304ad),
	.w6(32'hbb1beebc),
	.w7(32'hb9b9e201),
	.w8(32'h3af65ccb),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efa334),
	.w1(32'h3b2c666f),
	.w2(32'h39f72657),
	.w3(32'h39d5a2ed),
	.w4(32'h3addbd3f),
	.w5(32'h3ad91184),
	.w6(32'hbb213f69),
	.w7(32'h3a40188d),
	.w8(32'hba8726e5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a585f1),
	.w1(32'h3b09454d),
	.w2(32'h39f4e1f7),
	.w3(32'h3b461905),
	.w4(32'h3b623d51),
	.w5(32'h3973417b),
	.w6(32'hba9d2ec3),
	.w7(32'hb9cc6289),
	.w8(32'hbb67cd62),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68aa5b),
	.w1(32'h3afcccd4),
	.w2(32'hb772de7b),
	.w3(32'hb9e56e45),
	.w4(32'h3aa08780),
	.w5(32'h39f89399),
	.w6(32'hbad8f759),
	.w7(32'hb956f090),
	.w8(32'hbaddeb35),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3207d),
	.w1(32'h3b1e4726),
	.w2(32'h3b43c495),
	.w3(32'h3bb06d3a),
	.w4(32'h3bbb1511),
	.w5(32'h3b441e36),
	.w6(32'h3b3a9c7f),
	.w7(32'h3b86b685),
	.w8(32'h388b2942),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae5a27),
	.w1(32'hbadd6780),
	.w2(32'hbad9d24e),
	.w3(32'hbad188a6),
	.w4(32'hba99c906),
	.w5(32'h3aa4a79f),
	.w6(32'hba9b79ae),
	.w7(32'hb9a32d22),
	.w8(32'h3aac337b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada367c),
	.w1(32'h3a8e1764),
	.w2(32'h3a8af85f),
	.w3(32'h3a47ee57),
	.w4(32'h3a328b25),
	.w5(32'hbaebe711),
	.w6(32'h3a0c0c31),
	.w7(32'h3aae6d1a),
	.w8(32'hbac47490),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a7230),
	.w1(32'h396ec7f1),
	.w2(32'h3a69f472),
	.w3(32'hb91c8cf5),
	.w4(32'h3ab996f5),
	.w5(32'h39859d93),
	.w6(32'h392d4bc9),
	.w7(32'h3a52cecc),
	.w8(32'h3a5e690a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9388d1),
	.w1(32'hbb0d630c),
	.w2(32'hb7d8cda6),
	.w3(32'hb9b69b96),
	.w4(32'h3b29cfd6),
	.w5(32'h39d95d2b),
	.w6(32'hbb2c9536),
	.w7(32'hbad14dc4),
	.w8(32'hbb54d54f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35532d),
	.w1(32'hbacc9126),
	.w2(32'h3a6f8b49),
	.w3(32'hbb008eb9),
	.w4(32'hbaa5a564),
	.w5(32'h3b021f8c),
	.w6(32'hba9f6cde),
	.w7(32'h39f61ee2),
	.w8(32'h3a11620c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed1851),
	.w1(32'hbb08fba7),
	.w2(32'h39f1fcba),
	.w3(32'h397d6d18),
	.w4(32'hb99142b3),
	.w5(32'h3a4e2af2),
	.w6(32'hb9880a9b),
	.w7(32'h389333f3),
	.w8(32'hbaf1d696),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a86d6),
	.w1(32'hba419bf7),
	.w2(32'hba87b4a4),
	.w3(32'hb96886d4),
	.w4(32'h393449eb),
	.w5(32'hbac82268),
	.w6(32'hba3c0f1e),
	.w7(32'hb9e858b4),
	.w8(32'hb9b58c26),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993f160),
	.w1(32'h3a230746),
	.w2(32'h3a00bfea),
	.w3(32'hba02c267),
	.w4(32'h3a4bb27d),
	.w5(32'h39d3aae5),
	.w6(32'hba3424eb),
	.w7(32'h3a1fb536),
	.w8(32'h3a18d7bc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b0a2b),
	.w1(32'h332f993c),
	.w2(32'h38626550),
	.w3(32'h38c6a22a),
	.w4(32'hb9bd3321),
	.w5(32'h39505e8b),
	.w6(32'hba386436),
	.w7(32'hb9b24662),
	.w8(32'hb90fa4cf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb35fbf50),
	.w1(32'h39aaf221),
	.w2(32'hba104fc9),
	.w3(32'h39fda10e),
	.w4(32'hba06f90d),
	.w5(32'h3a9210f2),
	.w6(32'h3a9d1b3b),
	.w7(32'h399acaf3),
	.w8(32'h3a5b0953),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae69204),
	.w1(32'h3ac3c0ae),
	.w2(32'h3a8e641c),
	.w3(32'h3ae3d877),
	.w4(32'h3afc22c3),
	.w5(32'h399e4965),
	.w6(32'h3acfaaa9),
	.w7(32'h3b1a77ab),
	.w8(32'h3afa5780),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92cd72),
	.w1(32'h3af9079c),
	.w2(32'h3b064696),
	.w3(32'hba8305eb),
	.w4(32'h38aa8cee),
	.w5(32'hba016048),
	.w6(32'h3af576cb),
	.w7(32'h3ab40bb4),
	.w8(32'hbaefdc08),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e9de7),
	.w1(32'hbae3e17f),
	.w2(32'hba4b864a),
	.w3(32'h3a243761),
	.w4(32'h3a324dc5),
	.w5(32'h3b178460),
	.w6(32'h398e907c),
	.w7(32'hba4cd081),
	.w8(32'h39b18c91),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ad72f),
	.w1(32'h3884c639),
	.w2(32'h3a3fe47d),
	.w3(32'h39e723c8),
	.w4(32'h3b403b2f),
	.w5(32'h3a590574),
	.w6(32'h392431a6),
	.w7(32'h3b4c6a3c),
	.w8(32'h3a951553),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11160a),
	.w1(32'h39a6d1b2),
	.w2(32'h39df0ee8),
	.w3(32'h38d47d3b),
	.w4(32'h3a4b26f7),
	.w5(32'h39f21321),
	.w6(32'h3a222412),
	.w7(32'h3acbedae),
	.w8(32'h3a076805),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392501b1),
	.w1(32'h38519768),
	.w2(32'h3a396f8e),
	.w3(32'h3a4292c5),
	.w4(32'h3a52daf0),
	.w5(32'h3a0d3512),
	.w6(32'hb9b57062),
	.w7(32'h3a7781b2),
	.w8(32'h3a574e45),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f4196),
	.w1(32'h3a2aad36),
	.w2(32'h39870ca7),
	.w3(32'h3a22d261),
	.w4(32'h3a96c68f),
	.w5(32'hb99fcb99),
	.w6(32'hb892c749),
	.w7(32'h3a84cd0b),
	.w8(32'hbae9313e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22aa2b),
	.w1(32'hba57ca6f),
	.w2(32'hb905e682),
	.w3(32'hb9f21539),
	.w4(32'hb9c39649),
	.w5(32'h3a865ded),
	.w6(32'hba6300d8),
	.w7(32'hb9066b91),
	.w8(32'h39824ac6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96868d7),
	.w1(32'hbafa1986),
	.w2(32'h3a66ebf0),
	.w3(32'hbae26101),
	.w4(32'hbabb740a),
	.w5(32'h3b2bd938),
	.w6(32'hb9d42583),
	.w7(32'hb94c6b6a),
	.w8(32'h3b16769e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d3fac),
	.w1(32'hbb53cf5b),
	.w2(32'h3a9a7970),
	.w3(32'h3b49e37e),
	.w4(32'h3aeb297a),
	.w5(32'hbb034683),
	.w6(32'hbb3a8ddb),
	.w7(32'hbb6ac9fa),
	.w8(32'hbbb0fbfa),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9682be),
	.w1(32'hbb4c955e),
	.w2(32'hbb5e203a),
	.w3(32'hbac57b20),
	.w4(32'hb9d6a319),
	.w5(32'hbb834a82),
	.w6(32'hba9316a1),
	.w7(32'hbb0a38d8),
	.w8(32'hbb801a59),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f8da8),
	.w1(32'hbb74f467),
	.w2(32'hbbc27884),
	.w3(32'hbb4a8805),
	.w4(32'hba8fe027),
	.w5(32'hbb8b014e),
	.w6(32'hbbe12783),
	.w7(32'hbbf2e9e3),
	.w8(32'hbbe2f604),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba377e70),
	.w1(32'hba67d167),
	.w2(32'hb849483a),
	.w3(32'hb9a6d9e2),
	.w4(32'h38e75687),
	.w5(32'h39aea940),
	.w6(32'hba936749),
	.w7(32'h369db459),
	.w8(32'hb9705acf),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374ca955),
	.w1(32'h39b5fe3e),
	.w2(32'h3a73287f),
	.w3(32'h389e8ece),
	.w4(32'h397e3cdd),
	.w5(32'hba9a2c57),
	.w6(32'h3ac3dfde),
	.w7(32'h3a979c5e),
	.w8(32'hb9db033c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c04c48),
	.w1(32'hb9c916a5),
	.w2(32'hba311b61),
	.w3(32'hba2975e6),
	.w4(32'hba9d0420),
	.w5(32'h3acec840),
	.w6(32'h39dba9f5),
	.w7(32'hba17f52f),
	.w8(32'h399ce92b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c3032),
	.w1(32'hbac51ab6),
	.w2(32'hba6ea183),
	.w3(32'h3a50987a),
	.w4(32'h3aa542c6),
	.w5(32'h391dbbfd),
	.w6(32'h3a4d5dc4),
	.w7(32'h39774010),
	.w8(32'h38a1c5c0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dff001),
	.w1(32'h39f4ba83),
	.w2(32'h3a51dc91),
	.w3(32'h3a132279),
	.w4(32'hb9ebb7d0),
	.w5(32'hbb0fe4c3),
	.w6(32'h3a19c9dc),
	.w7(32'h3a0de654),
	.w8(32'hbaceaed1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15dcda),
	.w1(32'hbb6a5e01),
	.w2(32'hbb3f9011),
	.w3(32'hbb1b8de1),
	.w4(32'hbb0834e2),
	.w5(32'h3ad77b6c),
	.w6(32'hbb145ac6),
	.w7(32'hbb3c5667),
	.w8(32'hba78bd10),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d48fb),
	.w1(32'hb99e9292),
	.w2(32'h3b043eb1),
	.w3(32'hbad39167),
	.w4(32'hba605738),
	.w5(32'h3b106bd4),
	.w6(32'hba4ab817),
	.w7(32'hbb1c1498),
	.w8(32'hb9a63e54),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba845b01),
	.w1(32'h3a151f3d),
	.w2(32'h39509249),
	.w3(32'h3ae33e7a),
	.w4(32'h3b3e8f9d),
	.w5(32'h3957ea09),
	.w6(32'hba62d641),
	.w7(32'h39f512cb),
	.w8(32'hba977fcf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf1dbd),
	.w1(32'hba4f9dee),
	.w2(32'hb8f3dc9a),
	.w3(32'hbab557f6),
	.w4(32'hba8cdab9),
	.w5(32'h3b3ef55b),
	.w6(32'hbab25c73),
	.w7(32'hba9b4cd6),
	.w8(32'h3aacd147),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab5147),
	.w1(32'h389f5249),
	.w2(32'hb794f00e),
	.w3(32'h3b1943e4),
	.w4(32'h3a8808ec),
	.w5(32'hbab7e676),
	.w6(32'h3a57fb17),
	.w7(32'hb9a148dd),
	.w8(32'hbb0a9731),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4dbe6),
	.w1(32'hba488480),
	.w2(32'hbaa2aaf6),
	.w3(32'hbb171695),
	.w4(32'h390a441b),
	.w5(32'hba593199),
	.w6(32'hbb6d704d),
	.w7(32'h388b29e2),
	.w8(32'hbb2858cc),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae966ef),
	.w1(32'hbafc28f5),
	.w2(32'hbb189aee),
	.w3(32'hb9ac93f0),
	.w4(32'hb99042a4),
	.w5(32'h3a17182f),
	.w6(32'hbaf427e2),
	.w7(32'hbb0ddc81),
	.w8(32'hbac0a3a5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba370f3b),
	.w1(32'hb8b534cd),
	.w2(32'hba5cf691),
	.w3(32'hba968313),
	.w4(32'hba314aa6),
	.w5(32'hba393722),
	.w6(32'hba5d4bd2),
	.w7(32'hba857412),
	.w8(32'h397f7b1f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a0b6c8),
	.w1(32'hba0b940b),
	.w2(32'hba056f1b),
	.w3(32'hba527cb3),
	.w4(32'hba96dc06),
	.w5(32'h398c1315),
	.w6(32'h38bf4238),
	.w7(32'hb85464df),
	.w8(32'hb9ccac61),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16a1d7),
	.w1(32'h3a6b3978),
	.w2(32'hb9e30202),
	.w3(32'hba12505c),
	.w4(32'hba31bee0),
	.w5(32'h3aa88e26),
	.w6(32'hb95f6d96),
	.w7(32'hb9936c63),
	.w8(32'h3aaf6785),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefc270),
	.w1(32'h3ab29c0a),
	.w2(32'h3aa2ed28),
	.w3(32'h3ab716da),
	.w4(32'h3a9229cc),
	.w5(32'hb9d8956b),
	.w6(32'h3b275c26),
	.w7(32'h3a7b1fd6),
	.w8(32'hb9952b72),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5a03b),
	.w1(32'h3af71a31),
	.w2(32'h39c8e19b),
	.w3(32'hbb0379a6),
	.w4(32'hb967d746),
	.w5(32'hba1e2542),
	.w6(32'hb9bb7faf),
	.w7(32'h3a1a9bbe),
	.w8(32'hbb35c69b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba469f82),
	.w1(32'hba526fcd),
	.w2(32'hbaa575d8),
	.w3(32'h398ff2ea),
	.w4(32'h39b53839),
	.w5(32'h3afe0f80),
	.w6(32'h398b306d),
	.w7(32'h38861116),
	.w8(32'h3b0323e5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86ba03a),
	.w1(32'h3ad78077),
	.w2(32'h3b22cab1),
	.w3(32'h3a538149),
	.w4(32'h3b1ee422),
	.w5(32'h3ae51dce),
	.w6(32'hba9f2723),
	.w7(32'h394cf33d),
	.w8(32'hba92ccad),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac00ba),
	.w1(32'hbbaae276),
	.w2(32'hba35cd8c),
	.w3(32'hbb342c78),
	.w4(32'hba8712be),
	.w5(32'h3b14c69f),
	.w6(32'hbb7b1fc6),
	.w7(32'hbb53b992),
	.w8(32'h39169265),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa8212),
	.w1(32'h3b2359b5),
	.w2(32'hba0d3bd7),
	.w3(32'h3a91ab44),
	.w4(32'h3a5c258e),
	.w5(32'h387799f6),
	.w6(32'h3aa8219a),
	.w7(32'h3ae9647a),
	.w8(32'h3ac1155a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f5658),
	.w1(32'hbb79a141),
	.w2(32'hbbb21eb1),
	.w3(32'hb8e6e786),
	.w4(32'hbaf654cb),
	.w5(32'hba81a2c7),
	.w6(32'hbb1b0156),
	.w7(32'hbb3cdaa3),
	.w8(32'hbaee7ca7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a031051),
	.w1(32'h3a033ff7),
	.w2(32'hbb3de0a9),
	.w3(32'h3aa7751e),
	.w4(32'h3a226b87),
	.w5(32'hbb67a113),
	.w6(32'hba971ffd),
	.w7(32'h3a1e9542),
	.w8(32'hbb8acd99),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8d6af),
	.w1(32'hbbccb95e),
	.w2(32'hbb3eafd1),
	.w3(32'hbb534979),
	.w4(32'hba9c0f0f),
	.w5(32'h3b41eaac),
	.w6(32'hbb9c5bac),
	.w7(32'hbb528cbe),
	.w8(32'hba57c320),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45046e),
	.w1(32'hba936a0b),
	.w2(32'hba455e99),
	.w3(32'hbabbb060),
	.w4(32'hbab407d6),
	.w5(32'hb9c4af20),
	.w6(32'hbb36a9fb),
	.w7(32'hbb211d24),
	.w8(32'hba67cb9e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b261a),
	.w1(32'hbb09f263),
	.w2(32'hbb2985d3),
	.w3(32'hbb895f96),
	.w4(32'hbae4b69e),
	.w5(32'hbae02133),
	.w6(32'hba5a593a),
	.w7(32'hba80dc9c),
	.w8(32'hb94feffa),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7f709),
	.w1(32'h3ae8ffd8),
	.w2(32'h3ac03862),
	.w3(32'h3a74f9f3),
	.w4(32'h39d4177a),
	.w5(32'hba367873),
	.w6(32'h3ad58ea3),
	.w7(32'h3a241a33),
	.w8(32'hb916bc1b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49ec4e),
	.w1(32'hbb1bff08),
	.w2(32'hbad3cf2f),
	.w3(32'hba0ceb98),
	.w4(32'hba7c5dc6),
	.w5(32'hbb45bd90),
	.w6(32'hbb673ba7),
	.w7(32'hbacc80f8),
	.w8(32'hbbbabe08),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16678f),
	.w1(32'hbb7242b3),
	.w2(32'hbbbabd28),
	.w3(32'hbb2efef9),
	.w4(32'hbb98788e),
	.w5(32'hbb99b2cf),
	.w6(32'hbb4d9d05),
	.w7(32'hbb984888),
	.w8(32'hbbe66b1e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b34b5),
	.w1(32'hbc117b4e),
	.w2(32'hba911e3c),
	.w3(32'h39ba90bb),
	.w4(32'h35d01780),
	.w5(32'hb728cb2e),
	.w6(32'h3a00f105),
	.w7(32'hbb1d491d),
	.w8(32'hbbb4179c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb145168),
	.w1(32'h3b18f886),
	.w2(32'hbc0964c3),
	.w3(32'h3a5414e4),
	.w4(32'h3bbbf353),
	.w5(32'hbb068eb2),
	.w6(32'hb8becb69),
	.w7(32'h3b3c5c19),
	.w8(32'hbb7960da),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc68d79),
	.w1(32'h3a2cbaf0),
	.w2(32'h3b68d7ee),
	.w3(32'hb9220709),
	.w4(32'h3ba2987b),
	.w5(32'hba93caf5),
	.w6(32'hbbfa4087),
	.w7(32'hb9ef97b6),
	.w8(32'hbbb4fafe),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c278c),
	.w1(32'hbbbfe136),
	.w2(32'h3a18eab0),
	.w3(32'hbac001c5),
	.w4(32'hb994b9e9),
	.w5(32'hbb802595),
	.w6(32'hbbac2dd7),
	.w7(32'hbafdf61f),
	.w8(32'hbc1d5cb7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26b871),
	.w1(32'hbb8de67a),
	.w2(32'hbbd09773),
	.w3(32'hbaa8d4ea),
	.w4(32'hbb880d6b),
	.w5(32'hbb12cbd6),
	.w6(32'hbb67b311),
	.w7(32'hbb9bd13a),
	.w8(32'h3a37708e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc08d1a),
	.w1(32'hbbd9f56d),
	.w2(32'hbbc41393),
	.w3(32'hbb24ea6d),
	.w4(32'hba3ca9b1),
	.w5(32'hbb238235),
	.w6(32'h3addcdd6),
	.w7(32'hbaada587),
	.w8(32'hbc0f63f9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa089a5),
	.w1(32'hbb296c27),
	.w2(32'hbbb92377),
	.w3(32'hbacbd302),
	.w4(32'hb9dd8bb8),
	.w5(32'hbbfa2752),
	.w6(32'hba85cbb8),
	.w7(32'hb84f35df),
	.w8(32'hbbf747ee),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86968f),
	.w1(32'hbbbcc80c),
	.w2(32'hbb6281f9),
	.w3(32'hbb11bb74),
	.w4(32'hbafbb6fb),
	.w5(32'h3bd3c688),
	.w6(32'hbb723a2c),
	.w7(32'hbb120dd1),
	.w8(32'h3a97720c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b678763),
	.w1(32'h393a40c1),
	.w2(32'h3ad8ffc8),
	.w3(32'h3a376f9a),
	.w4(32'h3b830637),
	.w5(32'hbb7f3a18),
	.w6(32'hbb1e78fa),
	.w7(32'h3b76a900),
	.w8(32'hbbd9a1ed),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56dcf7),
	.w1(32'hbb27b4c0),
	.w2(32'hbb3e036f),
	.w3(32'hbb44fb89),
	.w4(32'hbae31660),
	.w5(32'h3bd5ff6b),
	.w6(32'hbbdd9ba2),
	.w7(32'hbb81160b),
	.w8(32'h3b2b356d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bf420),
	.w1(32'h39aca155),
	.w2(32'hba2348c5),
	.w3(32'hbab74537),
	.w4(32'h3b06d3fd),
	.w5(32'hbbc79fe6),
	.w6(32'hbc0af1eb),
	.w7(32'hbaaf4030),
	.w8(32'hbbb4d2b5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae5e4b),
	.w1(32'hbb19a7f3),
	.w2(32'hbb5f4fea),
	.w3(32'hbbc43e14),
	.w4(32'hbb90afdc),
	.w5(32'hbb720e7a),
	.w6(32'hb953520b),
	.w7(32'h3ace0ba9),
	.w8(32'h39f09efd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6dcdc9),
	.w1(32'h39f77080),
	.w2(32'hb91609b5),
	.w3(32'hbadbd6d3),
	.w4(32'hba4ed598),
	.w5(32'h3b7f47d0),
	.w6(32'hbb3ec25d),
	.w7(32'hbb170e6e),
	.w8(32'h3bc2e502),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55a582),
	.w1(32'h3bb06cd3),
	.w2(32'h3c028f97),
	.w3(32'h3b8f8bf5),
	.w4(32'h3b940efe),
	.w5(32'h3b14c5bc),
	.w6(32'h3b71c209),
	.w7(32'h3b332385),
	.w8(32'hbac56fda),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f136f),
	.w1(32'hbad772fd),
	.w2(32'hba520d68),
	.w3(32'hbadb5ccd),
	.w4(32'h3b0052b4),
	.w5(32'h3b3e2080),
	.w6(32'hb9d749c7),
	.w7(32'h3a56b108),
	.w8(32'hbb4b70bd),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1a5e6),
	.w1(32'hbb0df51a),
	.w2(32'h3b02ed91),
	.w3(32'hba60b892),
	.w4(32'hb9e63e69),
	.w5(32'hbb22420e),
	.w6(32'h3b5e16c7),
	.w7(32'hba4925f5),
	.w8(32'hbb9f3d61),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70a7d8),
	.w1(32'hbab8c749),
	.w2(32'h3957be75),
	.w3(32'hbac21dfc),
	.w4(32'h379a7f8e),
	.w5(32'h3b1da755),
	.w6(32'hbb47a483),
	.w7(32'h3a0a9e7c),
	.w8(32'h3bec48af),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbebb3),
	.w1(32'h3c30c326),
	.w2(32'h3c023d87),
	.w3(32'h3b687036),
	.w4(32'h3b680128),
	.w5(32'hbb83d46e),
	.w6(32'h3c1bd60e),
	.w7(32'h3bdf3a89),
	.w8(32'hbb70ec40),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20df1b),
	.w1(32'hba8e3f78),
	.w2(32'hbb803a45),
	.w3(32'hbb9abf6a),
	.w4(32'hbb97a16c),
	.w5(32'hb994811c),
	.w6(32'hbbc7b42b),
	.w7(32'hbb994498),
	.w8(32'hba60d022),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391ee604),
	.w1(32'hb8af9056),
	.w2(32'h3a9193e4),
	.w3(32'h393b4ab0),
	.w4(32'h39a8fab5),
	.w5(32'hbb4567e5),
	.w6(32'hba4751dd),
	.w7(32'hb9d6df43),
	.w8(32'hbb83f55d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb37082),
	.w1(32'hbbd305f3),
	.w2(32'hbbfa3365),
	.w3(32'hbb9164a5),
	.w4(32'hbb86c396),
	.w5(32'hbb558e2b),
	.w6(32'hbc043b34),
	.w7(32'hbc1035c5),
	.w8(32'hbb0cdd25),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5116b4),
	.w1(32'h386e3dc8),
	.w2(32'hbb30968f),
	.w3(32'hb85b9ac4),
	.w4(32'hba925083),
	.w5(32'h3ba134ca),
	.w6(32'hb9bbe7b7),
	.w7(32'hba4f5012),
	.w8(32'h3bc77759),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc53d5),
	.w1(32'h3b92c5eb),
	.w2(32'hbb66c0af),
	.w3(32'h3bb13bef),
	.w4(32'hbab98061),
	.w5(32'h3c075fa1),
	.w6(32'h3c0476a6),
	.w7(32'hbb0445de),
	.w8(32'hba13a629),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bc667),
	.w1(32'hbb7ffac4),
	.w2(32'hbad86c9c),
	.w3(32'h3b8700bf),
	.w4(32'h3b133ed5),
	.w5(32'h3b735dc7),
	.w6(32'hbb8a2631),
	.w7(32'h3a56c6b9),
	.w8(32'h3ba03d7a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba635aa),
	.w1(32'h3c12bf9e),
	.w2(32'h3b260b39),
	.w3(32'h392ba8bc),
	.w4(32'hbb1483b6),
	.w5(32'h3ad2824a),
	.w6(32'h3b52f388),
	.w7(32'h3b0f5ca7),
	.w8(32'h3acfdaa1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90db90),
	.w1(32'hbb4a579d),
	.w2(32'h3b1ce614),
	.w3(32'hb9b9572b),
	.w4(32'h3ac3afa6),
	.w5(32'h3848988a),
	.w6(32'h3b817df7),
	.w7(32'h3b1c1723),
	.w8(32'h39e93038),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b211fa0),
	.w1(32'h3ac2352d),
	.w2(32'hb9e877d2),
	.w3(32'hbb0937ff),
	.w4(32'hbb66c150),
	.w5(32'h3be71ed1),
	.w6(32'hbac27e57),
	.w7(32'hbb0a9386),
	.w8(32'h3bad6b7d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda685a),
	.w1(32'h3b834311),
	.w2(32'h3aee66c3),
	.w3(32'h392d4ff4),
	.w4(32'h3b161252),
	.w5(32'h39899187),
	.w6(32'h3abb3f3e),
	.w7(32'h3b2f2811),
	.w8(32'hba284cb3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5880ab),
	.w1(32'hbb313496),
	.w2(32'h3a862b76),
	.w3(32'h3a33ca61),
	.w4(32'hba806da0),
	.w5(32'h3b77b5d2),
	.w6(32'h3a56d146),
	.w7(32'hbb816425),
	.w8(32'hbb111b48),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1e165),
	.w1(32'hbc0e4f72),
	.w2(32'hbbaed996),
	.w3(32'h3a170c65),
	.w4(32'hbb4d4990),
	.w5(32'h3b2a1f5f),
	.w6(32'hbc52711b),
	.w7(32'hbc1d0d4c),
	.w8(32'h3ac9a7e7),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb526874),
	.w1(32'hbb65b6f4),
	.w2(32'h3ae45227),
	.w3(32'hbaa952ba),
	.w4(32'hbb401d96),
	.w5(32'hba3e24d8),
	.w6(32'hbb1f7133),
	.w7(32'hbb9013f6),
	.w8(32'hbb41671c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d71e0),
	.w1(32'hbbb61b77),
	.w2(32'hbb6254ad),
	.w3(32'hbb00be13),
	.w4(32'hba33cf76),
	.w5(32'hbb848736),
	.w6(32'hbbbd91aa),
	.w7(32'hbb753245),
	.w8(32'hba5a0c6d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a200c),
	.w1(32'hbab9b3c8),
	.w2(32'hbb30df04),
	.w3(32'hbb98331c),
	.w4(32'hbbd6eb49),
	.w5(32'h3bd7e68a),
	.w6(32'h3a4105c7),
	.w7(32'hbb737c18),
	.w8(32'hba685a03),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b345b26),
	.w1(32'h3b2e999d),
	.w2(32'h3af41777),
	.w3(32'h3ae84686),
	.w4(32'h3a9f4a66),
	.w5(32'h3970de0e),
	.w6(32'hbbabc88b),
	.w7(32'hbb804b91),
	.w8(32'hb9db63fc),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42ef5d),
	.w1(32'hbb85c389),
	.w2(32'hbb0e0a87),
	.w3(32'hbbe5f2db),
	.w4(32'hbb6c4431),
	.w5(32'h3b07125e),
	.w6(32'hbbb78e1d),
	.w7(32'hbb671732),
	.w8(32'h3b1a170b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43eb7d),
	.w1(32'hb9eae12d),
	.w2(32'hbafe213c),
	.w3(32'h3a090e04),
	.w4(32'hb8eb4b93),
	.w5(32'hbc03d250),
	.w6(32'h39fdddf2),
	.w7(32'hbb2bbaf6),
	.w8(32'hbbdf2532),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e816),
	.w1(32'hbb5dd4ab),
	.w2(32'hb9a36a98),
	.w3(32'hbb8937fa),
	.w4(32'hbb2b62c6),
	.w5(32'h3aedc9c7),
	.w6(32'hba638deb),
	.w7(32'hb9ad1aba),
	.w8(32'h3b05717f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11e81d),
	.w1(32'h3b9c3221),
	.w2(32'h3b70a76f),
	.w3(32'hb96e28ee),
	.w4(32'h3b30b70a),
	.w5(32'h3a2d8f1f),
	.w6(32'hba480349),
	.w7(32'h3a884d1c),
	.w8(32'hbaf8f0f8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c27c9),
	.w1(32'hbb27f5c5),
	.w2(32'hbb7b9e02),
	.w3(32'hbb6c59ff),
	.w4(32'hbba71e6f),
	.w5(32'hbaced84e),
	.w6(32'hbbc33fd0),
	.w7(32'hbbce2f9f),
	.w8(32'hba78ae2e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af77631),
	.w1(32'hbae789a8),
	.w2(32'hb862ca7c),
	.w3(32'hbb1047b1),
	.w4(32'hbb2df3d5),
	.w5(32'hba62aca0),
	.w6(32'hbb22b5dc),
	.w7(32'hbb4b3298),
	.w8(32'hbbe6cfbb),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e5ae6),
	.w1(32'hbbed1e54),
	.w2(32'hbc161dbf),
	.w3(32'hbb5cdf02),
	.w4(32'hbad6a1e0),
	.w5(32'h3bca41df),
	.w6(32'hbbfc20aa),
	.w7(32'hbb9d9bc8),
	.w8(32'hba6382c4),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cc058),
	.w1(32'hbbdeac59),
	.w2(32'hbbb42b32),
	.w3(32'h3b78055c),
	.w4(32'h3a6feb6c),
	.w5(32'h3ad01433),
	.w6(32'h3a092a71),
	.w7(32'h3a2fde49),
	.w8(32'hba66b2fe),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb567509),
	.w1(32'hbaafc4e9),
	.w2(32'hbab24c59),
	.w3(32'hbb0f91af),
	.w4(32'hbaff82de),
	.w5(32'hbbe3b125),
	.w6(32'hbbbfde42),
	.w7(32'hbb347155),
	.w8(32'hbba64528),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeed00c),
	.w1(32'hbbcb10a4),
	.w2(32'hbbe94380),
	.w3(32'hbbdecede),
	.w4(32'hbbd3fb87),
	.w5(32'h3aaadce4),
	.w6(32'hbb1dca8e),
	.w7(32'hbb7d4261),
	.w8(32'hb9875903),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6fe31),
	.w1(32'hb9ea9b59),
	.w2(32'h3b419302),
	.w3(32'h3af58c5b),
	.w4(32'h39e80ea0),
	.w5(32'h3b4a584c),
	.w6(32'h3a7c5b36),
	.w7(32'h3aed3a2b),
	.w8(32'hbb3f8aca),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a935241),
	.w1(32'hbb591c3f),
	.w2(32'hba38834b),
	.w3(32'hba35093d),
	.w4(32'h3b2d1756),
	.w5(32'hba9c0aa6),
	.w6(32'hbb7368b3),
	.w7(32'h3ac9f3fc),
	.w8(32'hba086fc4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383b8a93),
	.w1(32'h3a8fe3d1),
	.w2(32'hbaf9be42),
	.w3(32'h39a8ff47),
	.w4(32'hba96fca5),
	.w5(32'hbb892861),
	.w6(32'h3abf0984),
	.w7(32'hbab981d2),
	.w8(32'hbbbb7b99),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7c2a5),
	.w1(32'hbb7d0bff),
	.w2(32'hbbdae63d),
	.w3(32'hbbbf3dd5),
	.w4(32'hbbc28dd3),
	.w5(32'hbbc29e67),
	.w6(32'hbbeb4af6),
	.w7(32'hbc08718f),
	.w8(32'hbb63b4c8),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc704b9),
	.w1(32'h3b6c48fa),
	.w2(32'h3a089c2a),
	.w3(32'h3a210345),
	.w4(32'h3b1e56fe),
	.w5(32'h3be53f64),
	.w6(32'h3afb1052),
	.w7(32'hba130730),
	.w8(32'h3b20b16a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac33318),
	.w1(32'h3b980438),
	.w2(32'h3b39e57c),
	.w3(32'h3bbb03a1),
	.w4(32'h3bb95b26),
	.w5(32'h3a91ae3f),
	.w6(32'h3b982f3a),
	.w7(32'h3b696c79),
	.w8(32'h3b677662),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34445a),
	.w1(32'h3b9f1e58),
	.w2(32'h3ae9ccb3),
	.w3(32'h3b231ea7),
	.w4(32'h3abe8dc0),
	.w5(32'hbb2fb17f),
	.w6(32'h3b91a321),
	.w7(32'h3a814460),
	.w8(32'hbbbb5884),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f80b0),
	.w1(32'hbb6340c3),
	.w2(32'hb98abe49),
	.w3(32'hba19fd03),
	.w4(32'h3a686780),
	.w5(32'h3a90db4c),
	.w6(32'hbbae3e05),
	.w7(32'hbb3e34af),
	.w8(32'hbb9da973),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43da97),
	.w1(32'hbbaff200),
	.w2(32'h3ba301e5),
	.w3(32'h3900a3d1),
	.w4(32'h3b6ad1db),
	.w5(32'hbb149278),
	.w6(32'hbb8763d4),
	.w7(32'h3be95308),
	.w8(32'hbbac011b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96042a),
	.w1(32'h3ad8614c),
	.w2(32'h39027a4d),
	.w3(32'hbb63761c),
	.w4(32'h3b178ecb),
	.w5(32'hbad18eaa),
	.w6(32'hbbbb8825),
	.w7(32'hbad0c585),
	.w8(32'hbb972e0a),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34abbd),
	.w1(32'hbb648f0e),
	.w2(32'hbbe03664),
	.w3(32'hbb0946af),
	.w4(32'hb970cd33),
	.w5(32'hbb1d331d),
	.w6(32'hba9a98a9),
	.w7(32'hb9a08b97),
	.w8(32'hbb4ad388),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9010a5),
	.w1(32'hbaab29f2),
	.w2(32'hbafd2ce7),
	.w3(32'hbb245e2a),
	.w4(32'hbad3029f),
	.w5(32'h3b929e2f),
	.w6(32'hbac0953d),
	.w7(32'hbafd8e81),
	.w8(32'h3b38e408),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b733bc2),
	.w1(32'h3b83179d),
	.w2(32'h3baccf19),
	.w3(32'h39fbb9e9),
	.w4(32'h3b4a2265),
	.w5(32'h3b94889e),
	.w6(32'hbbc8e3b9),
	.w7(32'h3b11d97d),
	.w8(32'h3b2532d6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886ce6b),
	.w1(32'hbb1ff254),
	.w2(32'hbbdbaefb),
	.w3(32'hbb7e35d5),
	.w4(32'hbc03f6ca),
	.w5(32'h3b74f58f),
	.w6(32'hbb9aff8f),
	.w7(32'hbbf59a83),
	.w8(32'h3b2cc986),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab6b25),
	.w1(32'h3a9c798f),
	.w2(32'hbb3ec415),
	.w3(32'h3a2fb592),
	.w4(32'h3af6064c),
	.w5(32'hbb5f2270),
	.w6(32'h38e7a70e),
	.w7(32'hba6536a9),
	.w8(32'hba1a8b5c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cd75a),
	.w1(32'hb988362c),
	.w2(32'hba88c18d),
	.w3(32'hbb949cac),
	.w4(32'hbb19f91c),
	.w5(32'h3b1c92e5),
	.w6(32'hba9b0092),
	.w7(32'h3b34124e),
	.w8(32'h3a86b303),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac01303),
	.w1(32'h3b1232a2),
	.w2(32'h3b7353c1),
	.w3(32'h3b123c20),
	.w4(32'h3b447bab),
	.w5(32'hbb8743b2),
	.w6(32'h3bc32e83),
	.w7(32'h3b34c310),
	.w8(32'hbb7b87dd),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb839689),
	.w1(32'hbaaf8ec2),
	.w2(32'h3aa6a6ec),
	.w3(32'hbadaeaf5),
	.w4(32'hbae98d5e),
	.w5(32'hba49e73b),
	.w6(32'hba50ecc3),
	.w7(32'hbaa5c8a2),
	.w8(32'hbb21f66a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac639e8),
	.w1(32'hba81f2f0),
	.w2(32'hbb0b64be),
	.w3(32'hbb286382),
	.w4(32'hbb36ebac),
	.w5(32'hba812894),
	.w6(32'hba34426b),
	.w7(32'hbad94324),
	.w8(32'h3aa1c2ce),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a694b92),
	.w1(32'h3b490fa4),
	.w2(32'h3ad5bf37),
	.w3(32'hba9b64f8),
	.w4(32'h3a7c0e2e),
	.w5(32'hbba36ec4),
	.w6(32'hbac2c70f),
	.w7(32'h3917ca6a),
	.w8(32'hbbdc816d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb629962),
	.w1(32'hbbb538b0),
	.w2(32'hbb0b23d0),
	.w3(32'hbb08df2b),
	.w4(32'hbac953b8),
	.w5(32'hbb3cc6f2),
	.w6(32'hbb95522a),
	.w7(32'hbb7379b6),
	.w8(32'h3a3361e9),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba684c50),
	.w1(32'hba44e638),
	.w2(32'hbb868d14),
	.w3(32'h3b1db385),
	.w4(32'hba107207),
	.w5(32'h38642956),
	.w6(32'h3b7f9c85),
	.w7(32'h3ad7f190),
	.w8(32'hb9385c11),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd39749),
	.w1(32'h3acdab58),
	.w2(32'hbb1f7d6d),
	.w3(32'h3a3a7e80),
	.w4(32'hbaa43d48),
	.w5(32'hbb14c73b),
	.w6(32'hba6f46ef),
	.w7(32'hbbbe1801),
	.w8(32'h3a1f09e2),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b65e09),
	.w1(32'h3b6ab9f5),
	.w2(32'h3b94ca01),
	.w3(32'hba953cc2),
	.w4(32'hb8741ea7),
	.w5(32'hb9d6e27b),
	.w6(32'hbb112a65),
	.w7(32'h38b09f04),
	.w8(32'h3b0ef01c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967c44),
	.w1(32'h3b4bac65),
	.w2(32'hbb2b6cc8),
	.w3(32'hbb0cd7f6),
	.w4(32'hbb378834),
	.w5(32'h3aa4feb4),
	.w6(32'hbbaf17e0),
	.w7(32'hbbf1ea1a),
	.w8(32'h3a065b2b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb066d5b),
	.w1(32'hbbbc5409),
	.w2(32'hbbc0ed2e),
	.w3(32'hb9984ddc),
	.w4(32'hbb11a522),
	.w5(32'h3bd8b2fa),
	.w6(32'hbc048ac5),
	.w7(32'hbbe8cc54),
	.w8(32'hb9b74142),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba74d7c),
	.w1(32'h3b426b54),
	.w2(32'hbb0f14d1),
	.w3(32'h3b8fed42),
	.w4(32'h3bbf0f54),
	.w5(32'h3a7cd21c),
	.w6(32'h3baa11e0),
	.w7(32'h3b61f150),
	.w8(32'h3b1f3dcb),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3767b),
	.w1(32'h3bfaf039),
	.w2(32'h3bc07644),
	.w3(32'h3b00ebd7),
	.w4(32'h3b9be4c5),
	.w5(32'hbbd85d9a),
	.w6(32'h39d2d00f),
	.w7(32'h3b14479b),
	.w8(32'hbc409284),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc34c7a),
	.w1(32'hbc0578c9),
	.w2(32'hbb88640f),
	.w3(32'hbc348470),
	.w4(32'hbbe40ca9),
	.w5(32'hbab56787),
	.w6(32'hbc27faba),
	.w7(32'hbbd618e1),
	.w8(32'hba7e528c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb11ee3),
	.w1(32'hbba3442c),
	.w2(32'hbc120b17),
	.w3(32'hb9fadd11),
	.w4(32'hbb0c2ca6),
	.w5(32'h3b3e5586),
	.w6(32'h3a04430d),
	.w7(32'hbbaca6f5),
	.w8(32'hba38d465),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a978820),
	.w1(32'hbb7b9299),
	.w2(32'hbb3c8f12),
	.w3(32'h3a9368a8),
	.w4(32'h3c14e7df),
	.w5(32'h3a100f1a),
	.w6(32'hb9c39e83),
	.w7(32'h3c0a59a9),
	.w8(32'hba89f171),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10c778),
	.w1(32'hbb891201),
	.w2(32'hbb24e0c9),
	.w3(32'hbb488847),
	.w4(32'hb88ddb4d),
	.w5(32'h3ba1e241),
	.w6(32'hbbafb2ba),
	.w7(32'hbadd5e4e),
	.w8(32'h3b800fa1),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba726f0),
	.w1(32'h3bb50627),
	.w2(32'h3bbfc1c2),
	.w3(32'h3b80d56e),
	.w4(32'h3b75999f),
	.w5(32'hb9c6007b),
	.w6(32'h3bb3514e),
	.w7(32'h3b9a66ba),
	.w8(32'hbb14fc0e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe46f11),
	.w1(32'hbc1fe1c4),
	.w2(32'hbba9fc19),
	.w3(32'hbb1f8f42),
	.w4(32'hbb227766),
	.w5(32'h3b85c119),
	.w6(32'hbbb66453),
	.w7(32'hbb800fbc),
	.w8(32'h3be7931d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1dc94),
	.w1(32'h3c009d40),
	.w2(32'h3bac8100),
	.w3(32'h3b884a8b),
	.w4(32'h3b26ced9),
	.w5(32'hba072e83),
	.w6(32'h3c211a57),
	.w7(32'h3b8fbb59),
	.w8(32'hbb6f86a3),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb901cee),
	.w1(32'hba0c3294),
	.w2(32'h397a0dfa),
	.w3(32'h3ac5e0bf),
	.w4(32'h3b1002ee),
	.w5(32'hbb8aafb8),
	.w6(32'hba35339c),
	.w7(32'hba9262d7),
	.w8(32'hbbad21a4),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43e807),
	.w1(32'hbb6559ea),
	.w2(32'hbb3800df),
	.w3(32'hbb98ccf2),
	.w4(32'hbb873615),
	.w5(32'hbb359511),
	.w6(32'hbba54765),
	.w7(32'hbb825fb5),
	.w8(32'h39f39c72),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9a395),
	.w1(32'hbbd6e625),
	.w2(32'hbbde784e),
	.w3(32'hba714706),
	.w4(32'hbb18a9c7),
	.w5(32'h3a83ed28),
	.w6(32'hbb0e0af3),
	.w7(32'hbb7de043),
	.w8(32'h3ad5bcee),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa95d9a),
	.w1(32'h3ac5800d),
	.w2(32'hbb7f6bdf),
	.w3(32'hb978c727),
	.w4(32'h3b0639bc),
	.w5(32'hbb0835a8),
	.w6(32'h3a2d6122),
	.w7(32'h39544c76),
	.w8(32'hbae558a7),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa181af),
	.w1(32'hbab71d0b),
	.w2(32'hb9f22604),
	.w3(32'hbb3ba3b8),
	.w4(32'h3a83feb8),
	.w5(32'h3b0f708a),
	.w6(32'hba4352d6),
	.w7(32'h3abb4d47),
	.w8(32'hb96181f7),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcbe99),
	.w1(32'hb657bf92),
	.w2(32'h3ab7c49e),
	.w3(32'h3a93355b),
	.w4(32'h3b103d87),
	.w5(32'hb9aab419),
	.w6(32'hba1d8f35),
	.w7(32'h38f494b0),
	.w8(32'h368df757),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb044b6e),
	.w1(32'hbb00c182),
	.w2(32'h3a0f9e74),
	.w3(32'h3a151902),
	.w4(32'h3a88cb81),
	.w5(32'hba55dba2),
	.w6(32'hbaab195a),
	.w7(32'h3b21099a),
	.w8(32'h3b0ff723),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01c2f7),
	.w1(32'hbafc429a),
	.w2(32'h3ad4dc07),
	.w3(32'hbb25f2d3),
	.w4(32'hb9f5d01b),
	.w5(32'h3b65a773),
	.w6(32'h39c6d1e7),
	.w7(32'hb934842c),
	.w8(32'h3bac4620),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bced1a7),
	.w1(32'h3c0d8fa9),
	.w2(32'h3b85a374),
	.w3(32'h3b919c8f),
	.w4(32'h3b17b38c),
	.w5(32'hbbfbb3f2),
	.w6(32'h3c03b9df),
	.w7(32'h3b84bce5),
	.w8(32'hbbf6b0b3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d6380),
	.w1(32'h3b64b050),
	.w2(32'h3a859c86),
	.w3(32'h3b9167c4),
	.w4(32'h3c1ab1ec),
	.w5(32'hb8f32460),
	.w6(32'h3b9bb0c7),
	.w7(32'h3c1817ef),
	.w8(32'h3b2259c8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7a03a),
	.w1(32'h3bd8d89a),
	.w2(32'h3bbe322f),
	.w3(32'hbb6bfde1),
	.w4(32'h3a37ae4d),
	.w5(32'h3b1da709),
	.w6(32'h38b1cf4b),
	.w7(32'h3b6359b2),
	.w8(32'h3aa88b9b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9810188),
	.w1(32'hbb8f2f2a),
	.w2(32'hbb5d6e97),
	.w3(32'hbb5b017a),
	.w4(32'hbbcfa89b),
	.w5(32'hb9ecf0b3),
	.w6(32'hba9b82fc),
	.w7(32'h3a954d02),
	.w8(32'hbb6907f0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7792ba),
	.w1(32'h3a2e9eea),
	.w2(32'hb7a31fad),
	.w3(32'hb9916a47),
	.w4(32'h3aa28de6),
	.w5(32'hbb1478ae),
	.w6(32'hbb46ebea),
	.w7(32'h38278c96),
	.w8(32'hbae83ce1),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafaed40),
	.w1(32'hbb3d2bba),
	.w2(32'hb9610a26),
	.w3(32'hbaadcbab),
	.w4(32'h394cd8b2),
	.w5(32'hbba614ff),
	.w6(32'hbaae0788),
	.w7(32'hb7826582),
	.w8(32'hba9c9315),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac57526),
	.w1(32'hbb42494f),
	.w2(32'h398a61c9),
	.w3(32'hbbed41b6),
	.w4(32'hbb494023),
	.w5(32'h3a839117),
	.w6(32'hbb7a2447),
	.w7(32'h3ad72e96),
	.w8(32'hbae86465),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab001d),
	.w1(32'hbb779707),
	.w2(32'hbb6fe1c6),
	.w3(32'hbab1570d),
	.w4(32'hba5c772e),
	.w5(32'hbb972222),
	.w6(32'hbbc66235),
	.w7(32'hbb524393),
	.w8(32'hba169e3f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3570a),
	.w1(32'hbbd0084e),
	.w2(32'hbbdbcb19),
	.w3(32'hba778c05),
	.w4(32'hbb32852d),
	.w5(32'hbbcc6051),
	.w6(32'h39f5aa6c),
	.w7(32'hba649ada),
	.w8(32'hbc0a6bb2),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5a966),
	.w1(32'hbbcd2a11),
	.w2(32'hbb96c859),
	.w3(32'hbb605a41),
	.w4(32'h3b0f869a),
	.w5(32'hbbbe392a),
	.w6(32'hbbd82c68),
	.w7(32'hbb0c4bbe),
	.w8(32'hbbefb7d9),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd10601),
	.w1(32'hbb76da93),
	.w2(32'h3bc6c913),
	.w3(32'hbb3ee422),
	.w4(32'h3b60aa23),
	.w5(32'hbb1589a6),
	.w6(32'hbb061ea4),
	.w7(32'h3b8bd39a),
	.w8(32'hbba0be14),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb071e99),
	.w1(32'hbab079c2),
	.w2(32'hbb5c49b7),
	.w3(32'hbaa0a12f),
	.w4(32'h3adde9ce),
	.w5(32'hbaa35866),
	.w6(32'hba918e16),
	.w7(32'hbac541e9),
	.w8(32'hbaaa25a2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9961d3f),
	.w1(32'h3a9d214d),
	.w2(32'hba4cc819),
	.w3(32'h3aa6ab7e),
	.w4(32'hb9c47314),
	.w5(32'hbb274715),
	.w6(32'h3b26b78c),
	.w7(32'hba092a5f),
	.w8(32'hbb0cb5db),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e3ffd),
	.w1(32'hbba0fc63),
	.w2(32'hbb93b110),
	.w3(32'hbb2a7847),
	.w4(32'hbb80543e),
	.w5(32'hbb9aa000),
	.w6(32'hbb9f9c58),
	.w7(32'hbb6ef578),
	.w8(32'hbc066679),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaffda),
	.w1(32'hbb973000),
	.w2(32'h3b7cd7cb),
	.w3(32'hbb2fc15c),
	.w4(32'hbba03c3e),
	.w5(32'h3b5e1319),
	.w6(32'hbbd7e691),
	.w7(32'h3aa18970),
	.w8(32'h3b301310),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa70906),
	.w1(32'h3aa9aa66),
	.w2(32'hb929b004),
	.w3(32'hbb232388),
	.w4(32'hbb78be89),
	.w5(32'h3a3ca38a),
	.w6(32'hb906ebd3),
	.w7(32'hbad30b72),
	.w8(32'h3ac79d5d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69dd1f),
	.w1(32'hbbd4fd58),
	.w2(32'hbb210559),
	.w3(32'hbb5686e0),
	.w4(32'hbb632534),
	.w5(32'hbb2ca238),
	.w6(32'hbbe88b07),
	.w7(32'hbb8d7610),
	.w8(32'hbbd6b137),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac264d),
	.w1(32'hbbc1433a),
	.w2(32'hbbd287fd),
	.w3(32'hba857133),
	.w4(32'h39be97e8),
	.w5(32'hbb3eed97),
	.w6(32'hbb8ad102),
	.w7(32'hbb7ef347),
	.w8(32'hbbae3b71),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88750e),
	.w1(32'hbb8517d8),
	.w2(32'hbb1b2665),
	.w3(32'h3ae5f82d),
	.w4(32'h3afb8992),
	.w5(32'hbb432c9e),
	.w6(32'hbbc7ed07),
	.w7(32'hbb2c8442),
	.w8(32'hbbcfd2ae),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb227d17),
	.w1(32'hbb6201c4),
	.w2(32'hba66ba8a),
	.w3(32'hbad24ff6),
	.w4(32'hbac2a5cb),
	.w5(32'hbba21843),
	.w6(32'hbb0e79f6),
	.w7(32'hbadf3a04),
	.w8(32'hb9f8f789),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb903fbf),
	.w1(32'hbb91ebf9),
	.w2(32'hbb6e3539),
	.w3(32'hba47823a),
	.w4(32'hbbc1b119),
	.w5(32'h3aaaad6a),
	.w6(32'hbb4a4b6e),
	.w7(32'hbb869a77),
	.w8(32'hbb2f08b1),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922f71d),
	.w1(32'hbb866536),
	.w2(32'hbaf15dab),
	.w3(32'hba8fca7e),
	.w4(32'h3af24d48),
	.w5(32'h3b07356c),
	.w6(32'hbba6d869),
	.w7(32'h3b1b3eb7),
	.w8(32'h3afaa7a3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70c925),
	.w1(32'h3b1c42a1),
	.w2(32'hbb87bc78),
	.w3(32'h3b58d0dd),
	.w4(32'h3a239d7e),
	.w5(32'hbb59d0be),
	.w6(32'h3b6e7721),
	.w7(32'hbb1c7251),
	.w8(32'hbbb44991),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89abc2),
	.w1(32'hbb0f5edc),
	.w2(32'hba966d4f),
	.w3(32'hb9b6f932),
	.w4(32'hb9fe71bb),
	.w5(32'hbbf8389f),
	.w6(32'hb9b987f0),
	.w7(32'hba51705b),
	.w8(32'hbbb5c34e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba23a0c),
	.w1(32'hbb6589e6),
	.w2(32'h3bf23706),
	.w3(32'hbb1b3321),
	.w4(32'h39d16509),
	.w5(32'hbb8b96a5),
	.w6(32'hbb775525),
	.w7(32'h3aed8eac),
	.w8(32'hbbeddffa),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92c105),
	.w1(32'hbb8c6ecc),
	.w2(32'hbbcabffa),
	.w3(32'hbaf6e949),
	.w4(32'hbaf4b933),
	.w5(32'hbbdf958d),
	.w6(32'hbbcfcbdf),
	.w7(32'hbbeceda2),
	.w8(32'hbbf79da8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8c2a1),
	.w1(32'hbb57f774),
	.w2(32'h3b08dcf1),
	.w3(32'hbb3602ea),
	.w4(32'h397b3f84),
	.w5(32'h3b6183e8),
	.w6(32'hbbde873e),
	.w7(32'hbb012629),
	.w8(32'hbb1a7d35),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65b7d2),
	.w1(32'h3ad54568),
	.w2(32'h3ba015ef),
	.w3(32'hba08398e),
	.w4(32'h3a8ce904),
	.w5(32'hbba80b0c),
	.w6(32'hbbbfc0f5),
	.w7(32'h3b9d4b2e),
	.w8(32'hbbeee552),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ba462),
	.w1(32'hbbcf6958),
	.w2(32'hbb942c25),
	.w3(32'hbbc31ab1),
	.w4(32'hbb77bbbc),
	.w5(32'hba8ddcf7),
	.w6(32'hbbb85d12),
	.w7(32'hbb7930e1),
	.w8(32'hbb79e0ed),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc322d),
	.w1(32'h3a92000d),
	.w2(32'hba9c6545),
	.w3(32'hba9be51a),
	.w4(32'h3a75c8bb),
	.w5(32'h3b1fb7e9),
	.w6(32'hbb9e13fe),
	.w7(32'hbb4c3ac2),
	.w8(32'h3b6f938a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f3b7c),
	.w1(32'h3ad88b04),
	.w2(32'h3b055453),
	.w3(32'h396af074),
	.w4(32'hba950fb8),
	.w5(32'h3c08288e),
	.w6(32'h3b70cbdc),
	.w7(32'h3aa3fc4e),
	.w8(32'h3bdf0daa),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bbce0),
	.w1(32'hbb9a734e),
	.w2(32'hbbd778b1),
	.w3(32'h39b1da26),
	.w4(32'h39d82916),
	.w5(32'h3b2649e0),
	.w6(32'h3a1cfaaa),
	.w7(32'hbb318d18),
	.w8(32'hba9d214e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3c57f),
	.w1(32'hbb9d55af),
	.w2(32'h3aa5c86a),
	.w3(32'h3bb0a6ce),
	.w4(32'h39123943),
	.w5(32'hbb90d762),
	.w6(32'h3b64a2d9),
	.w7(32'hbab445bc),
	.w8(32'hbbb70e18),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a789d),
	.w1(32'hbb9f9c41),
	.w2(32'hbb6f8d8d),
	.w3(32'hbaecc762),
	.w4(32'hbb8ec7fd),
	.w5(32'h3b1c15c9),
	.w6(32'hbb65cf99),
	.w7(32'hbb497a5a),
	.w8(32'hbb0aee0f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c240d),
	.w1(32'hba9f0166),
	.w2(32'h3b202f11),
	.w3(32'hb9c21e22),
	.w4(32'h3a6ef237),
	.w5(32'h39ba9de1),
	.w6(32'h39af0295),
	.w7(32'hbac95415),
	.w8(32'hba0a0d67),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef86e9),
	.w1(32'hb9cdab58),
	.w2(32'hbab44cbf),
	.w3(32'hb9bef150),
	.w4(32'hb949898a),
	.w5(32'h3a17af5d),
	.w6(32'hbb1beb7a),
	.w7(32'hba407e91),
	.w8(32'hba636c5c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04cb96),
	.w1(32'hbaec611c),
	.w2(32'hbb4ef859),
	.w3(32'h3a7df26f),
	.w4(32'hbab7520d),
	.w5(32'hbb1dff73),
	.w6(32'hbb626ce0),
	.w7(32'hbbec2a8e),
	.w8(32'hba05c123),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46a6f9),
	.w1(32'hba4e5cb0),
	.w2(32'h3b01c21b),
	.w3(32'hba8dabd8),
	.w4(32'h398cc8b6),
	.w5(32'hbacf518b),
	.w6(32'hbae2dc47),
	.w7(32'hbb9d1aa0),
	.w8(32'hb84a0695),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6c8fb),
	.w1(32'h3b438d24),
	.w2(32'h3b442d15),
	.w3(32'h3961c6f5),
	.w4(32'hbad79d4a),
	.w5(32'h3a346544),
	.w6(32'h3ac36783),
	.w7(32'hba97a572),
	.w8(32'hbb48ae8e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c5148),
	.w1(32'h388b0a69),
	.w2(32'h3b55b02f),
	.w3(32'hb9cb83fe),
	.w4(32'h3aecffbf),
	.w5(32'hba7e17d9),
	.w6(32'hb9b57195),
	.w7(32'h3b4e8cc1),
	.w8(32'hba30ba46),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9460a60),
	.w1(32'hbb092ad3),
	.w2(32'hbb35b3b9),
	.w3(32'hb96dff62),
	.w4(32'hb98b1bdd),
	.w5(32'hba368188),
	.w6(32'hbae17c5d),
	.w7(32'hb967ed12),
	.w8(32'hbad2840c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99ee9d),
	.w1(32'hbaec9fc7),
	.w2(32'hbb00b566),
	.w3(32'hbb031cd2),
	.w4(32'h3abb2fab),
	.w5(32'hba35b146),
	.w6(32'hbbbd14eb),
	.w7(32'hbb741967),
	.w8(32'hbb0c1a44),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387038e7),
	.w1(32'hbaac431f),
	.w2(32'hb9a892bd),
	.w3(32'hba9af3e2),
	.w4(32'h3aa7251e),
	.w5(32'hbb2944e7),
	.w6(32'h3a6bf0c9),
	.w7(32'hb90da33d),
	.w8(32'hbae769c5),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe0c45),
	.w1(32'hba0c95a2),
	.w2(32'h3acc791c),
	.w3(32'hb76ca4de),
	.w4(32'h3b12dd3b),
	.w5(32'h381dd1a5),
	.w6(32'h3b5682c8),
	.w7(32'h3b3cb243),
	.w8(32'h39f5cba3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88f29b),
	.w1(32'hbb836f2d),
	.w2(32'hbaf2e61d),
	.w3(32'h39d1bbb0),
	.w4(32'hba29fe63),
	.w5(32'h3a0d1678),
	.w6(32'hbacc2290),
	.w7(32'hbb548a4f),
	.w8(32'hbb2b9270),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f7e40),
	.w1(32'hbaf0651f),
	.w2(32'hbac2d067),
	.w3(32'hba6dbad1),
	.w4(32'hba088144),
	.w5(32'hb9461555),
	.w6(32'hba7938fd),
	.w7(32'hba5c0cf2),
	.w8(32'hb66fd36a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf4027),
	.w1(32'h3aba5d39),
	.w2(32'hba930e5d),
	.w3(32'h3b2bba4b),
	.w4(32'h3b68b456),
	.w5(32'hb98444e9),
	.w6(32'hbaec40f8),
	.w7(32'h3a1d42f5),
	.w8(32'hba59100d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba859de2),
	.w1(32'h3a26e86c),
	.w2(32'hb9931639),
	.w3(32'hbade5b27),
	.w4(32'hb9c2428c),
	.w5(32'h3b08beaf),
	.w6(32'hbb3604f7),
	.w7(32'hb9cc952a),
	.w8(32'hba1445ee),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db284e),
	.w1(32'h3b0582d8),
	.w2(32'h3a21519f),
	.w3(32'h3640c0ed),
	.w4(32'h3a1a396d),
	.w5(32'h3ab749b3),
	.w6(32'hbac11d3a),
	.w7(32'hb9910d41),
	.w8(32'h3aa80291),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4e31f),
	.w1(32'h3a186334),
	.w2(32'hb8d8f8ec),
	.w3(32'h3ab3b7fd),
	.w4(32'h3a89a190),
	.w5(32'hba4861ca),
	.w6(32'h39746435),
	.w7(32'hb96dba14),
	.w8(32'hba358721),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9149976),
	.w1(32'hb9c482cd),
	.w2(32'h39199845),
	.w3(32'h3886ad1c),
	.w4(32'h3a08b913),
	.w5(32'h3abb1814),
	.w6(32'hba49539e),
	.w7(32'hb71fbf28),
	.w8(32'h3a86e900),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb28dc),
	.w1(32'h37bdb12d),
	.w2(32'h391159ad),
	.w3(32'hb97493d0),
	.w4(32'h393d2e83),
	.w5(32'hba10f998),
	.w6(32'h38e8e075),
	.w7(32'h3a8ebca3),
	.w8(32'h3a5abaa0),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bc9a7),
	.w1(32'hb9b963a0),
	.w2(32'h39964624),
	.w3(32'hb86bef2b),
	.w4(32'h3a31a4b0),
	.w5(32'hbb2414b1),
	.w6(32'h3803c827),
	.w7(32'hb96da77f),
	.w8(32'hbb24c40a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ba4f1),
	.w1(32'h3951a559),
	.w2(32'hbb21beaf),
	.w3(32'hbb0b48e2),
	.w4(32'hbb0be63b),
	.w5(32'hb9f99d88),
	.w6(32'hbb96069f),
	.w7(32'hbb467e46),
	.w8(32'hbabb0999),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba673eb2),
	.w1(32'hbb057496),
	.w2(32'hbac14983),
	.w3(32'hbad75d66),
	.w4(32'hbb12086b),
	.w5(32'hba9fa610),
	.w6(32'hbb12f2b7),
	.w7(32'hbaee0e7e),
	.w8(32'hba8e5282),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00d6a2),
	.w1(32'h3a9ed458),
	.w2(32'hba2f1763),
	.w3(32'h3aca01e8),
	.w4(32'h3a08b152),
	.w5(32'h3a1c94ce),
	.w6(32'h39798995),
	.w7(32'hba53d605),
	.w8(32'h3ae09edc),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32477e),
	.w1(32'h3bbdce6c),
	.w2(32'hba177cc2),
	.w3(32'h3b6ddd4d),
	.w4(32'h3af0c83e),
	.w5(32'hbabac4aa),
	.w6(32'h3afb26ab),
	.w7(32'h39b7a0ef),
	.w8(32'hbad7d27d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae42947),
	.w1(32'hba299ca8),
	.w2(32'hb9cee300),
	.w3(32'hba8c6c07),
	.w4(32'hba4d195a),
	.w5(32'h3a59a3f8),
	.w6(32'hba614c14),
	.w7(32'hb98590ae),
	.w8(32'hba13aea3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad185fb),
	.w1(32'hba54d20d),
	.w2(32'hb9a7b4df),
	.w3(32'h3a3b3205),
	.w4(32'hba49e839),
	.w5(32'hba19198e),
	.w6(32'h388db1fa),
	.w7(32'hb8bb3138),
	.w8(32'hb8b528a1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff9097),
	.w1(32'h3aa5df05),
	.w2(32'h3a81aa04),
	.w3(32'hba38894d),
	.w4(32'h3b70e5bb),
	.w5(32'h3882172c),
	.w6(32'hb94fc63d),
	.w7(32'h388f8504),
	.w8(32'hba89021e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e380),
	.w1(32'hbb99344a),
	.w2(32'hbb74247f),
	.w3(32'hbba6a414),
	.w4(32'hbb043250),
	.w5(32'hbb737bf9),
	.w6(32'hbbd506f3),
	.w7(32'hbb7c63d1),
	.w8(32'hbb97289d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac997d8),
	.w1(32'hbb02330f),
	.w2(32'hbb2fdff8),
	.w3(32'hbbb78c31),
	.w4(32'hbb857bef),
	.w5(32'h3aaa45a8),
	.w6(32'hbb4aed47),
	.w7(32'hbb83622b),
	.w8(32'hb980cb7c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f0964),
	.w1(32'h3982416e),
	.w2(32'h39f4d53d),
	.w3(32'h3adec687),
	.w4(32'h3a654ef9),
	.w5(32'hbb072bd6),
	.w6(32'hba6da3fc),
	.w7(32'h3adf6fe2),
	.w8(32'hba01d7c1),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcf1e9),
	.w1(32'h3a6eabdd),
	.w2(32'h3a85d084),
	.w3(32'hbb357771),
	.w4(32'h3aadd680),
	.w5(32'hbaa27891),
	.w6(32'hbabd9de5),
	.w7(32'h3a4f5103),
	.w8(32'h3a8b51d7),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb195109),
	.w1(32'hba296881),
	.w2(32'h3a977a24),
	.w3(32'hb984ae9e),
	.w4(32'hba452f1b),
	.w5(32'h3ada0ab3),
	.w6(32'h3b4c81e1),
	.w7(32'h3aad8132),
	.w8(32'hba9c20da),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a2645),
	.w1(32'h3adfa528),
	.w2(32'h3af19c03),
	.w3(32'h3b7a5510),
	.w4(32'h3a6791c2),
	.w5(32'hbb80b599),
	.w6(32'h3b9cc0c0),
	.w7(32'h3ae6d4e9),
	.w8(32'hbb1ad18a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c4c36),
	.w1(32'h3b0ee65f),
	.w2(32'hb931c9d7),
	.w3(32'h39c4d2ab),
	.w4(32'hba6eb463),
	.w5(32'hba2aaa94),
	.w6(32'h39b59a78),
	.w7(32'h3ab71037),
	.w8(32'h3a009a16),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb406f4c),
	.w1(32'hbb22e093),
	.w2(32'hba6f21cb),
	.w3(32'hbb3bd0b3),
	.w4(32'h3b0ff1a7),
	.w5(32'h3b6938f3),
	.w6(32'h3a5f9128),
	.w7(32'h3af5c459),
	.w8(32'h3a632c61),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380195ea),
	.w1(32'hba6b3cb5),
	.w2(32'hba15e9df),
	.w3(32'h398efb40),
	.w4(32'h39a662ea),
	.w5(32'hba16ddda),
	.w6(32'h389ebd0c),
	.w7(32'h387c5081),
	.w8(32'h38a421bf),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2658f9),
	.w1(32'h3aa48422),
	.w2(32'h3b772c84),
	.w3(32'hb9b13c22),
	.w4(32'h3ad95c96),
	.w5(32'hbb378b17),
	.w6(32'hbb1b2948),
	.w7(32'hbad6a27e),
	.w8(32'hbb514406),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule