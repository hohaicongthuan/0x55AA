module layer_8_featuremap_18(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a707816),
	.w1(32'hbbd68575),
	.w2(32'hbc5c1f86),
	.w3(32'h3c15cc65),
	.w4(32'h3996a3a7),
	.w5(32'hbc2bb161),
	.w6(32'hbb212475),
	.w7(32'hbbcc006f),
	.w8(32'h3b8c21f4),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5075e),
	.w1(32'h3b891503),
	.w2(32'h3c463ef6),
	.w3(32'h3b68479b),
	.w4(32'h3bbae023),
	.w5(32'h37786c46),
	.w6(32'hbb9d7367),
	.w7(32'hbba0026c),
	.w8(32'h3a1ddf4f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25b7c8),
	.w1(32'h3b3f2b49),
	.w2(32'h3c10bbcc),
	.w3(32'h3b80ff82),
	.w4(32'h3bb180d5),
	.w5(32'h3abd130e),
	.w6(32'h3bd3cca3),
	.w7(32'h3af2318c),
	.w8(32'h3b2e2550),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae8eda),
	.w1(32'hbb92eac0),
	.w2(32'h3b988c51),
	.w3(32'hbb85f96a),
	.w4(32'h3af69920),
	.w5(32'hbb2483db),
	.w6(32'h3b63f268),
	.w7(32'h3bb2b0c5),
	.w8(32'hbb8ae8dd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a53de),
	.w1(32'hbad957e1),
	.w2(32'hbb18df63),
	.w3(32'hb9a39deb),
	.w4(32'h3c6c23b2),
	.w5(32'hbad96389),
	.w6(32'h3bc34770),
	.w7(32'h3bb6d9fa),
	.w8(32'hbb547308),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c263113),
	.w1(32'h3affac3f),
	.w2(32'hbad208be),
	.w3(32'h3c4d8b5b),
	.w4(32'h3bd4fbf6),
	.w5(32'h39f0e4c4),
	.w6(32'h3bf21a91),
	.w7(32'h3b45041d),
	.w8(32'hb8c2a2a4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2693f6),
	.w1(32'h3b887d6d),
	.w2(32'h3b3b629f),
	.w3(32'h3ab3c5e2),
	.w4(32'hbb58ad4f),
	.w5(32'hb9a81cfa),
	.w6(32'h3c2d8cc4),
	.w7(32'h3c70b173),
	.w8(32'h3ab12945),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2407f9),
	.w1(32'h3ba17b4c),
	.w2(32'h3c2c96a1),
	.w3(32'h3b0c9c8c),
	.w4(32'h39ad1f14),
	.w5(32'h39f5e713),
	.w6(32'hbb3f795e),
	.w7(32'h3b5b50fc),
	.w8(32'hbb0a84d2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0316da),
	.w1(32'h3bb4cc62),
	.w2(32'h3aae3707),
	.w3(32'h3b04d82b),
	.w4(32'hbafafddd),
	.w5(32'h3a870184),
	.w6(32'hbb8cb0e9),
	.w7(32'hbb8847a8),
	.w8(32'hbbbc3cb2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b6086),
	.w1(32'hbad3f93c),
	.w2(32'hbb586097),
	.w3(32'h3b84a4ce),
	.w4(32'h3a8a2a60),
	.w5(32'hba86d2fa),
	.w6(32'h3b1a354e),
	.w7(32'hba78cbcb),
	.w8(32'h3b543c42),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd38ef1),
	.w1(32'h3add1555),
	.w2(32'h3682fef3),
	.w3(32'h3b8cd74b),
	.w4(32'hbbd8526f),
	.w5(32'hbb90abfc),
	.w6(32'h37abbf4d),
	.w7(32'hbc07092f),
	.w8(32'hbb78901b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5df51),
	.w1(32'h3c9eaddb),
	.w2(32'hbb027d6d),
	.w3(32'h3aa12909),
	.w4(32'hba72f4aa),
	.w5(32'hbba475fe),
	.w6(32'h3b15c95a),
	.w7(32'hbaa65a66),
	.w8(32'hb9217215),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb26d02),
	.w1(32'h3bcda453),
	.w2(32'hbab9622f),
	.w3(32'h3b3a683f),
	.w4(32'h3c69dacf),
	.w5(32'h3c44bc79),
	.w6(32'h3b3672a9),
	.w7(32'h3cbf7fb6),
	.w8(32'h3d644c27),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca549b0),
	.w1(32'hbc38d09c),
	.w2(32'hbc568371),
	.w3(32'hbc5e29f5),
	.w4(32'hbc399202),
	.w5(32'h3bf40445),
	.w6(32'hbc9be2e6),
	.w7(32'hbba0cf94),
	.w8(32'hb8bd8004),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b5f81),
	.w1(32'hbd1fd084),
	.w2(32'h3c6f156f),
	.w3(32'hbc397ab0),
	.w4(32'h3b207cb0),
	.w5(32'h38ed5a26),
	.w6(32'hbc1f7300),
	.w7(32'hbc95bfd3),
	.w8(32'h3d4cbffe),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b95e1),
	.w1(32'hbc0aca6d),
	.w2(32'hbc22fe65),
	.w3(32'hbc1bd25c),
	.w4(32'hbc409aae),
	.w5(32'hbbda5c4c),
	.w6(32'hbc7fa790),
	.w7(32'h3d8adfe5),
	.w8(32'hbbb353e6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d18d8c4),
	.w1(32'hbb7444e6),
	.w2(32'hb901f2f0),
	.w3(32'h3cec8536),
	.w4(32'hbc3acdfa),
	.w5(32'hbc6fc52c),
	.w6(32'hbcce8b84),
	.w7(32'h3c78eb1e),
	.w8(32'hbc39b687),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27c89a),
	.w1(32'hbbe366f4),
	.w2(32'hbc04b2f1),
	.w3(32'h3c76d6cb),
	.w4(32'hbc35606a),
	.w5(32'hbc8eec9e),
	.w6(32'hbc64cbec),
	.w7(32'hbcd4d91a),
	.w8(32'hbb8bac9e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9d853),
	.w1(32'hbcb4b55c),
	.w2(32'hbcac91cf),
	.w3(32'hbce6dca9),
	.w4(32'hbcb21074),
	.w5(32'hbcc890fa),
	.w6(32'h3d4fa1ea),
	.w7(32'hbc777a4e),
	.w8(32'h3becd300),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adca562),
	.w1(32'hbce29afc),
	.w2(32'hbc959e1d),
	.w3(32'h3c3f51e8),
	.w4(32'hbcce8672),
	.w5(32'hbc32ae7b),
	.w6(32'hbc3b19b6),
	.w7(32'hbb744fc9),
	.w8(32'hbc80cba0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb953caf),
	.w1(32'h3a9169ed),
	.w2(32'h3c33c073),
	.w3(32'h3b4109fe),
	.w4(32'h3b9f732e),
	.w5(32'hb92df370),
	.w6(32'hbcb9fca7),
	.w7(32'h3c80b0a3),
	.w8(32'hbbf351c0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fdf89),
	.w1(32'h3b806f05),
	.w2(32'hbc27cba3),
	.w3(32'hb9b6164c),
	.w4(32'hbc2fcf74),
	.w5(32'hbc95600c),
	.w6(32'hbad087b7),
	.w7(32'hbc33ab4b),
	.w8(32'hbb9089ed),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2c7f2a),
	.w1(32'hbd40f9e4),
	.w2(32'h3ccf9d30),
	.w3(32'h3c5a17c2),
	.w4(32'hbba62f47),
	.w5(32'hbc5fada0),
	.w6(32'h3bfdceea),
	.w7(32'h3d385711),
	.w8(32'hbbce5be4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29a835),
	.w1(32'hbcc01477),
	.w2(32'h3d2fbfaf),
	.w3(32'hbccc7458),
	.w4(32'hbb3bdeae),
	.w5(32'h3b6198bf),
	.w6(32'hb91dffe4),
	.w7(32'hbcc15e3f),
	.w8(32'h3c915564),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b2ad3),
	.w1(32'hbaf5ab97),
	.w2(32'hbc8e19fd),
	.w3(32'hbc6c66ba),
	.w4(32'h3abab34c),
	.w5(32'hbc848bd3),
	.w6(32'hbbd02db6),
	.w7(32'hbc1e72fb),
	.w8(32'h3bf3b3f1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c142c39),
	.w1(32'h3bd85834),
	.w2(32'hb9905010),
	.w3(32'h3bc8f7a3),
	.w4(32'hbb9eadba),
	.w5(32'hbd2ba400),
	.w6(32'hbbac942c),
	.w7(32'hbc61ffe6),
	.w8(32'hbc374d60),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbfeedf),
	.w1(32'h3c35d926),
	.w2(32'h3ac0b1e7),
	.w3(32'h3ce814ff),
	.w4(32'hbc83535d),
	.w5(32'hbae09d57),
	.w6(32'h3b726b00),
	.w7(32'hbcba0f9c),
	.w8(32'hba8beaf5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd232c34),
	.w1(32'hbd4751b2),
	.w2(32'hbcf81610),
	.w3(32'hbaeabb9c),
	.w4(32'hbd1a01ab),
	.w5(32'hbdafdfd6),
	.w6(32'h3c229bb8),
	.w7(32'hbd22f704),
	.w8(32'hbd55630d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c100583),
	.w1(32'h3bc63d35),
	.w2(32'hb9f664c1),
	.w3(32'hba6c5141),
	.w4(32'h3b87f603),
	.w5(32'hb92aa352),
	.w6(32'h3bf9c7a0),
	.w7(32'hbaf405fd),
	.w8(32'hba8aa203),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b793fdc),
	.w1(32'h3bede88c),
	.w2(32'h3b9584bc),
	.w3(32'hbb0207f6),
	.w4(32'hbaa2345b),
	.w5(32'h39a01ddd),
	.w6(32'hba424c66),
	.w7(32'h3bae953c),
	.w8(32'hbb46e047),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba67e86),
	.w1(32'h3c0d215c),
	.w2(32'h3b684c06),
	.w3(32'h39105273),
	.w4(32'h3ac87ec4),
	.w5(32'hbc006513),
	.w6(32'hba37f011),
	.w7(32'hbb856634),
	.w8(32'h39da0e08),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc98ff),
	.w1(32'h3aea23e5),
	.w2(32'hbc0951cb),
	.w3(32'hbac0c472),
	.w4(32'hbb581ba4),
	.w5(32'h3c1f22b6),
	.w6(32'hba549acd),
	.w7(32'h3b914c3a),
	.w8(32'hbb448d38),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c083f5e),
	.w1(32'h3bf4b2c1),
	.w2(32'hbb7d2d80),
	.w3(32'hbb767435),
	.w4(32'h3b09bc46),
	.w5(32'hbb245ed3),
	.w6(32'h3b9fd833),
	.w7(32'h3b5842bf),
	.w8(32'hbb07a44d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdeb0a0),
	.w1(32'h3b8af0a8),
	.w2(32'h3be42637),
	.w3(32'h3b52a2d1),
	.w4(32'hbb3550ee),
	.w5(32'hbc351447),
	.w6(32'h3ad448f6),
	.w7(32'h3c71d61b),
	.w8(32'h3b417efe),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb78682),
	.w1(32'hbb8b3675),
	.w2(32'hbad93747),
	.w3(32'hbb2ac328),
	.w4(32'h3c026454),
	.w5(32'h3ace383e),
	.w6(32'h3bcf031b),
	.w7(32'h3c74bd77),
	.w8(32'hbb11d8c3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac97e7),
	.w1(32'hbbf9a209),
	.w2(32'hbb8c15b6),
	.w3(32'hbb97f647),
	.w4(32'h37dd8610),
	.w5(32'hbc293585),
	.w6(32'hbb94c91c),
	.w7(32'h3bb53259),
	.w8(32'hbc0c9fb4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef2219),
	.w1(32'hbb0ca13b),
	.w2(32'hb9c16ca6),
	.w3(32'hbad06182),
	.w4(32'hb93f50a3),
	.w5(32'hbb4ce4cb),
	.w6(32'h3adfe9f7),
	.w7(32'h3bced51e),
	.w8(32'hbbb6b354),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8cac9),
	.w1(32'h3bc4c729),
	.w2(32'h3b8eab7e),
	.w3(32'hbadc333f),
	.w4(32'h3b03b10c),
	.w5(32'hbb757c63),
	.w6(32'h3b2e8f52),
	.w7(32'h3c0ae338),
	.w8(32'h3bc00bb6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e672e),
	.w1(32'h3b2813cd),
	.w2(32'h3c00b292),
	.w3(32'hbb47739f),
	.w4(32'hbb204b9b),
	.w5(32'h3c4e8ace),
	.w6(32'hbb97bcdc),
	.w7(32'hbb3846b9),
	.w8(32'hbb8711a8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e2595),
	.w1(32'hbcb649d2),
	.w2(32'hbaaecdff),
	.w3(32'hbaab0e3f),
	.w4(32'hb9bd41dc),
	.w5(32'hbb028594),
	.w6(32'h3b80d2c6),
	.w7(32'h3a8ab7e2),
	.w8(32'hbc642010),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18944d),
	.w1(32'h3a88d89d),
	.w2(32'hbbd61409),
	.w3(32'hbb913a4a),
	.w4(32'hbbf8eb25),
	.w5(32'hbc952596),
	.w6(32'hbbe1852c),
	.w7(32'hbca69b88),
	.w8(32'h3ac4dff2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a7d4f),
	.w1(32'hba102776),
	.w2(32'hbc64e00d),
	.w3(32'hbbab576e),
	.w4(32'hbc0ae76b),
	.w5(32'h3a69a890),
	.w6(32'hbba545c4),
	.w7(32'h39dc85a3),
	.w8(32'hba49cdc8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c963264),
	.w1(32'hbb7405b5),
	.w2(32'h3c8ccb59),
	.w3(32'h3b96cf31),
	.w4(32'hbbcfa936),
	.w5(32'h3b84f6a2),
	.w6(32'hbc35d97a),
	.w7(32'h3ae7785d),
	.w8(32'hbbd63860),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d8ced),
	.w1(32'hbc27126d),
	.w2(32'hb9c841fb),
	.w3(32'h3b416f62),
	.w4(32'hbbba5939),
	.w5(32'hbaa74af3),
	.w6(32'h3b65a31d),
	.w7(32'h3c4cdfed),
	.w8(32'hbcc4270c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb4640),
	.w1(32'h3b8ea976),
	.w2(32'h3b84aae5),
	.w3(32'h3c345a3e),
	.w4(32'hbc1fa9bf),
	.w5(32'hbca6801b),
	.w6(32'hbc042d4e),
	.w7(32'h3c139add),
	.w8(32'h3c2ef09b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc459d0d),
	.w1(32'hbb231297),
	.w2(32'h38bcc23a),
	.w3(32'hbb6cfd4d),
	.w4(32'hbc3240b5),
	.w5(32'h3a140cc7),
	.w6(32'h3c3e8407),
	.w7(32'hba88e795),
	.w8(32'h3bd9846d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23b76f),
	.w1(32'h3a0cdf77),
	.w2(32'h3c0c8ff4),
	.w3(32'h3af5a02c),
	.w4(32'hba3fc0c7),
	.w5(32'h3baab03b),
	.w6(32'h3d038d8b),
	.w7(32'hbbebc4a7),
	.w8(32'hb9a4418f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7d164),
	.w1(32'h3c31188f),
	.w2(32'hbb0aa80f),
	.w3(32'h3c99042a),
	.w4(32'hbbaa360d),
	.w5(32'hba53c94a),
	.w6(32'h3a47697f),
	.w7(32'h39b58b60),
	.w8(32'hbb97bde0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd1610e),
	.w1(32'hbc3570e9),
	.w2(32'hba06c219),
	.w3(32'h3bc64855),
	.w4(32'hbbb83c39),
	.w5(32'h3c0e0d32),
	.w6(32'hbc1b886a),
	.w7(32'h3bf015ec),
	.w8(32'h3c981df7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18ae4f),
	.w1(32'h3b2082b6),
	.w2(32'h3c05314d),
	.w3(32'hbbd154bd),
	.w4(32'h3a2b4d4d),
	.w5(32'h3c918ee0),
	.w6(32'h3ced36f4),
	.w7(32'hb9c5db22),
	.w8(32'hbb15fb64),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c167ff4),
	.w1(32'h3c698370),
	.w2(32'h3b355ba6),
	.w3(32'h3c1c093f),
	.w4(32'h3cb9b398),
	.w5(32'hbbc42f4d),
	.w6(32'h3d12b0a3),
	.w7(32'h3bc7ae54),
	.w8(32'h3b88dcd7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80ee96),
	.w1(32'hba34c1cc),
	.w2(32'h3bdf9836),
	.w3(32'h38d35e74),
	.w4(32'hbc1830e1),
	.w5(32'hba980b40),
	.w6(32'hba0bfa73),
	.w7(32'hbc84d9c1),
	.w8(32'h3bfbff30),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c078193),
	.w1(32'hbc926392),
	.w2(32'h3ba81586),
	.w3(32'hbc13fb24),
	.w4(32'hbbb7e35e),
	.w5(32'h3aa30ef5),
	.w6(32'hbc0235b3),
	.w7(32'hbb8b14b5),
	.w8(32'h3bff7e80),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11788f),
	.w1(32'hbc7e7b7e),
	.w2(32'hbc56f921),
	.w3(32'hbc916265),
	.w4(32'hbb1ebea0),
	.w5(32'h3aabaaa9),
	.w6(32'hbc8bafaa),
	.w7(32'hbca69557),
	.w8(32'hbc0386b5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eef3b),
	.w1(32'h3a7076f9),
	.w2(32'h3c0d96c4),
	.w3(32'hbc902111),
	.w4(32'hbb86d107),
	.w5(32'hbca994cf),
	.w6(32'h3b861b0d),
	.w7(32'h3c23d927),
	.w8(32'h3bb69191),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a155444),
	.w1(32'hbc463d08),
	.w2(32'hbc57615d),
	.w3(32'h3a9e7d74),
	.w4(32'hb9aea36a),
	.w5(32'hbd31fe3d),
	.w6(32'hbcd7e877),
	.w7(32'h3ba5da53),
	.w8(32'hbc566edf),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3276d),
	.w1(32'hbcd51c2f),
	.w2(32'hbaf5226e),
	.w3(32'h3bf22387),
	.w4(32'hbc2ed9c3),
	.w5(32'hbc5a6354),
	.w6(32'hbb6f123f),
	.w7(32'hbc36fa98),
	.w8(32'h3b850e44),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7cb508),
	.w1(32'h3d025322),
	.w2(32'h3cb3c4cc),
	.w3(32'hbc082164),
	.w4(32'hbcd9cb2a),
	.w5(32'h3dcb346c),
	.w6(32'hbd144314),
	.w7(32'hbd0d4a9f),
	.w8(32'h3be19efe),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c228555),
	.w1(32'hbc37d13c),
	.w2(32'hbcacc3b0),
	.w3(32'hbc009ad1),
	.w4(32'hbd10b0f6),
	.w5(32'h3c4f6431),
	.w6(32'h3ba1169a),
	.w7(32'hbcae163b),
	.w8(32'hbcb7c88b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2804c7),
	.w1(32'hb979d83d),
	.w2(32'hbbe22047),
	.w3(32'hbc61791d),
	.w4(32'hb9b725ce),
	.w5(32'h39f5fa8a),
	.w6(32'hbc8f5a49),
	.w7(32'h3a2e1aa9),
	.w8(32'h3c132bcc),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e39ca),
	.w1(32'hbcae504b),
	.w2(32'h3cee074d),
	.w3(32'hbd1e818d),
	.w4(32'hbcf2b386),
	.w5(32'hbc137c32),
	.w6(32'hbc4b84b3),
	.w7(32'h397b0fe5),
	.w8(32'hbc3f6192),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd9fd3),
	.w1(32'h3c0bf837),
	.w2(32'hb8dc0140),
	.w3(32'hbca3d375),
	.w4(32'hbd2f3e2f),
	.w5(32'hbb0f2483),
	.w6(32'h3b0858fe),
	.w7(32'h3a32f2a4),
	.w8(32'h3c8cbba6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba066b6c),
	.w1(32'hbc2f3c18),
	.w2(32'h3ba07b09),
	.w3(32'h3cadc0ca),
	.w4(32'hbb61589e),
	.w5(32'hbbdc2607),
	.w6(32'hba260575),
	.w7(32'hbc7702ab),
	.w8(32'hbcaa40c0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbeca1f),
	.w1(32'h3c00bab8),
	.w2(32'h3c8e8031),
	.w3(32'h3c80438d),
	.w4(32'hbb800c0a),
	.w5(32'hbb9cf041),
	.w6(32'hbc480b10),
	.w7(32'h3b3e5f3e),
	.w8(32'h3abaad4a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39774010),
	.w1(32'hbc442c3d),
	.w2(32'hbc344f10),
	.w3(32'hbce6a0b9),
	.w4(32'h3cf5dc70),
	.w5(32'hbca3ec51),
	.w6(32'hbc03d5b1),
	.w7(32'h3d803f4a),
	.w8(32'hbb0cf7c0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b8e8b),
	.w1(32'hbc65f0d1),
	.w2(32'h393214fc),
	.w3(32'hbb78e804),
	.w4(32'hbcae10d4),
	.w5(32'hbc86d39b),
	.w6(32'h3cc282d0),
	.w7(32'hbc86ade5),
	.w8(32'hbb6427de),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8bb838),
	.w1(32'h3d2c10ef),
	.w2(32'hbc363265),
	.w3(32'h3ad3512c),
	.w4(32'hbcd4f76f),
	.w5(32'h3a652265),
	.w6(32'hbca2e136),
	.w7(32'hbd02c80b),
	.w8(32'h3d151ac9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62a65a),
	.w1(32'h3addda60),
	.w2(32'hbc8d1b23),
	.w3(32'h37b3c86a),
	.w4(32'hbc0607ae),
	.w5(32'h3b818e20),
	.w6(32'h3c06e1ec),
	.w7(32'hbc977b8c),
	.w8(32'h3c98ccc1),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd40487),
	.w1(32'h3bdc746d),
	.w2(32'hbc98006f),
	.w3(32'hba85c1db),
	.w4(32'hbbb09b3a),
	.w5(32'h3cc2c4c3),
	.w6(32'hbc926f50),
	.w7(32'h3aa86deb),
	.w8(32'hbc0fcb6d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10f3d1),
	.w1(32'hbb906c9d),
	.w2(32'h3ae37cc6),
	.w3(32'hbbe1a476),
	.w4(32'hbcad52ba),
	.w5(32'hbcb6a856),
	.w6(32'h3bf65d03),
	.w7(32'hbc866d97),
	.w8(32'hbc26fcd5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb62051),
	.w1(32'hbb0ce4e1),
	.w2(32'hbb8ed4db),
	.w3(32'hbbc552a0),
	.w4(32'hbc85176d),
	.w5(32'h3ae02034),
	.w6(32'hbb9a7fd5),
	.w7(32'h3ab9f90f),
	.w8(32'hbb152a64),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86e4e2),
	.w1(32'h3ae1160f),
	.w2(32'hbc211464),
	.w3(32'hbbb7e6f5),
	.w4(32'hbbfb5e87),
	.w5(32'hbbbd9c1b),
	.w6(32'hba92e422),
	.w7(32'hbc343f01),
	.w8(32'hbb915be6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb747799),
	.w1(32'hbbaabe79),
	.w2(32'h3cc52930),
	.w3(32'hbba37591),
	.w4(32'hbb8bf438),
	.w5(32'hbb2c586e),
	.w6(32'h3c4b9caa),
	.w7(32'h3b946943),
	.w8(32'h3c442623),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c058c8c),
	.w1(32'hbab7db16),
	.w2(32'hbc1219d3),
	.w3(32'h3c0053c7),
	.w4(32'hbba7e216),
	.w5(32'hbb85b6e4),
	.w6(32'hbc1bc30b),
	.w7(32'h3aa218b9),
	.w8(32'hbbc93a89),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8da2d2),
	.w1(32'hbb506348),
	.w2(32'h3bfca8f4),
	.w3(32'h3c8d0988),
	.w4(32'hbc0b484c),
	.w5(32'hbb2618c5),
	.w6(32'h3c1da6e6),
	.w7(32'hbacf4112),
	.w8(32'hba01d7ea),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd75bf),
	.w1(32'hbc113aac),
	.w2(32'hb9b94086),
	.w3(32'h3c297d1c),
	.w4(32'hbb136278),
	.w5(32'hbbc65a71),
	.w6(32'h3aa25087),
	.w7(32'h3b51daa1),
	.w8(32'hbb605345),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba61ca),
	.w1(32'hbc40fdea),
	.w2(32'h3c9cfdc7),
	.w3(32'hbb02d58f),
	.w4(32'hbabe8bc5),
	.w5(32'hbb1e70b3),
	.w6(32'hbb57fa5a),
	.w7(32'h3cfa87c8),
	.w8(32'hbb8e0a50),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92c040),
	.w1(32'hbc3a5b3a),
	.w2(32'h3a78c9bb),
	.w3(32'hbbffb5ba),
	.w4(32'hbc3e7363),
	.w5(32'hbc31f649),
	.w6(32'h3c1112ee),
	.w7(32'hbc55cbd7),
	.w8(32'h38eafda0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cbc4d6),
	.w1(32'hbc6ab1d5),
	.w2(32'h3c40a391),
	.w3(32'h3ab96acb),
	.w4(32'hbb5f3e7a),
	.w5(32'h3a4b6ded),
	.w6(32'h3bc85d19),
	.w7(32'hbb885f08),
	.w8(32'h3adc860b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba134a9),
	.w1(32'hba9dc0a9),
	.w2(32'hbbac1e7b),
	.w3(32'hba5d80a4),
	.w4(32'hbbe44bb6),
	.w5(32'h3c7a3b6f),
	.w6(32'h3cb66722),
	.w7(32'hb850c81b),
	.w8(32'h3c0b227b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a735060),
	.w1(32'h3bd88b71),
	.w2(32'hbb58b7eb),
	.w3(32'hba485094),
	.w4(32'hbab25df9),
	.w5(32'hbc1ad5fd),
	.w6(32'hbb3f6098),
	.w7(32'hbc659b7c),
	.w8(32'hbbbd9808),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b986d0f),
	.w1(32'h3ba0d36e),
	.w2(32'hbb9189c4),
	.w3(32'h3baf722b),
	.w4(32'h3bd89b88),
	.w5(32'hbb73a4ca),
	.w6(32'hbb157d75),
	.w7(32'hbba76948),
	.w8(32'h3c926a93),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46b18c),
	.w1(32'h3a3c0106),
	.w2(32'hbb7c1732),
	.w3(32'h3ab667c5),
	.w4(32'hbc2afdce),
	.w5(32'hbc0ffc12),
	.w6(32'h3c30a2bc),
	.w7(32'hbc8b5795),
	.w8(32'hbc575e50),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9095b9),
	.w1(32'hbc0adaad),
	.w2(32'hbbd52a06),
	.w3(32'h3c0bb440),
	.w4(32'hbc0fb0c8),
	.w5(32'hbc605a2e),
	.w6(32'hbc9f9170),
	.w7(32'h3ae57fc9),
	.w8(32'hbbd85c36),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5da285),
	.w1(32'hbc25946a),
	.w2(32'h3cb105ee),
	.w3(32'hbc52cf93),
	.w4(32'hbc8e2514),
	.w5(32'hbd0445c1),
	.w6(32'hb91708b2),
	.w7(32'hbbf52bf9),
	.w8(32'hbcb11882),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8fee8),
	.w1(32'h3cd82862),
	.w2(32'h3b4391c7),
	.w3(32'h3a3a3a5b),
	.w4(32'hbbeb060a),
	.w5(32'hbc5e34de),
	.w6(32'h3b189b0d),
	.w7(32'hbc15e204),
	.w8(32'hbbcd8534),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f8feb),
	.w1(32'h3b5a9ab0),
	.w2(32'h3b5c559b),
	.w3(32'hbb02f79c),
	.w4(32'h3b3a891c),
	.w5(32'h3b14817f),
	.w6(32'hbba21b7c),
	.w7(32'hbab57768),
	.w8(32'hbc70303c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb929b808),
	.w1(32'hbb949163),
	.w2(32'hbbc7d057),
	.w3(32'hbc327376),
	.w4(32'h3b85f972),
	.w5(32'h3a703303),
	.w6(32'h3bbe716a),
	.w7(32'hbaa768b1),
	.w8(32'h3cb17859),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb839afb),
	.w1(32'hbc52efa6),
	.w2(32'hbb430dfd),
	.w3(32'h3a13d819),
	.w4(32'h3a9c9fe6),
	.w5(32'hbc8e6e65),
	.w6(32'h3b14fa2e),
	.w7(32'hbad81d63),
	.w8(32'h3c3058d2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b956a6c),
	.w1(32'h3b817395),
	.w2(32'h3bb85004),
	.w3(32'h3b535009),
	.w4(32'hba44d54e),
	.w5(32'h3b712d3f),
	.w6(32'hbae61926),
	.w7(32'hbbe6dc2b),
	.w8(32'hbb050a5f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4084b4),
	.w1(32'hbbcdd54e),
	.w2(32'hbc5de0be),
	.w3(32'h3aa86072),
	.w4(32'hbb6d731b),
	.w5(32'h3b2767e6),
	.w6(32'h3bad3a0f),
	.w7(32'h3c47307b),
	.w8(32'hbc125c54),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6a5a8),
	.w1(32'hbb2ce935),
	.w2(32'h3b03d936),
	.w3(32'hbadc3709),
	.w4(32'hbba5be0f),
	.w5(32'h38207dbf),
	.w6(32'hba8d535e),
	.w7(32'h3c62a93d),
	.w8(32'h3c0a25d5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d9dac),
	.w1(32'h3c22c8ba),
	.w2(32'h3a87719a),
	.w3(32'hbc7b7a53),
	.w4(32'h3c95675e),
	.w5(32'h3c15ceb4),
	.w6(32'h3a80b95c),
	.w7(32'hbbdfea28),
	.w8(32'hbb0ae03e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf21226),
	.w1(32'h3a7945d0),
	.w2(32'hbbe3b2c0),
	.w3(32'hbba7926b),
	.w4(32'hbc27f8b0),
	.w5(32'hbb8cf885),
	.w6(32'hbb5f9b50),
	.w7(32'hba8844ef),
	.w8(32'hbb370093),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23b510),
	.w1(32'h3b07be13),
	.w2(32'h3bdfbeef),
	.w3(32'hbb3b996e),
	.w4(32'h39aed5c5),
	.w5(32'hbae281ad),
	.w6(32'hbc23d5ea),
	.w7(32'hbb969233),
	.w8(32'hbb5ba312),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b081339),
	.w1(32'hbb401616),
	.w2(32'h3c4e988a),
	.w3(32'h3b9ce4ca),
	.w4(32'hbb79725a),
	.w5(32'hbc20cb64),
	.w6(32'h3bf2503a),
	.w7(32'h3c4ebdde),
	.w8(32'hbcb4cc20),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d05a9),
	.w1(32'hbb485b1e),
	.w2(32'hbb2ddea7),
	.w3(32'hbb08e5e1),
	.w4(32'hbbf822e6),
	.w5(32'hbbccff43),
	.w6(32'hb9b94210),
	.w7(32'hbcd51faa),
	.w8(32'hbb6ab1a8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a533a),
	.w1(32'hba82fb69),
	.w2(32'hba1e9022),
	.w3(32'hb7c318f1),
	.w4(32'hba1108d9),
	.w5(32'h3bd4438e),
	.w6(32'h3b8cead8),
	.w7(32'hbb91911c),
	.w8(32'hbd416c2f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b854567),
	.w1(32'h3c224d7c),
	.w2(32'hbc1307a5),
	.w3(32'hbb8b0c64),
	.w4(32'hbc3b031b),
	.w5(32'hbb435e45),
	.w6(32'hbb7d30d5),
	.w7(32'hba2a44d1),
	.w8(32'hbd7f5dcb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84b024a),
	.w1(32'hbb6f9b2c),
	.w2(32'h3c268995),
	.w3(32'h3c894228),
	.w4(32'hbc74bf18),
	.w5(32'h3bb82f0b),
	.w6(32'hbae6aaf7),
	.w7(32'hbd57955c),
	.w8(32'hbb8c8dc2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d4a59),
	.w1(32'hbba0153d),
	.w2(32'h3c0b5375),
	.w3(32'hbcae590a),
	.w4(32'hba473026),
	.w5(32'hbb12c276),
	.w6(32'h3c059261),
	.w7(32'h3b4e2587),
	.w8(32'h3bf4a7b3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6796c),
	.w1(32'h3d012a24),
	.w2(32'h3c1b8d6a),
	.w3(32'h3d8ba170),
	.w4(32'h3d0b28a7),
	.w5(32'hbc170bc7),
	.w6(32'hbbc975e0),
	.w7(32'h3c2d9189),
	.w8(32'hbb2fc750),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cf438),
	.w1(32'h3bcecda1),
	.w2(32'h3c34d191),
	.w3(32'hbd1a30f8),
	.w4(32'h3c229b56),
	.w5(32'hbc0795bb),
	.w6(32'hbba9d069),
	.w7(32'h3d51f5e4),
	.w8(32'h3bbce9b6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b2ec0),
	.w1(32'hbbfc89e6),
	.w2(32'hbc050d45),
	.w3(32'hbc49fde5),
	.w4(32'h3ad06209),
	.w5(32'hbc1c9135),
	.w6(32'hbc0f0a9b),
	.w7(32'h3c3e668a),
	.w8(32'h3b8cdcc4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b0e03),
	.w1(32'hbaa2eb2c),
	.w2(32'h3c08b037),
	.w3(32'hbb024a68),
	.w4(32'h3c267497),
	.w5(32'hbd371e3a),
	.w6(32'hbb4281d4),
	.w7(32'hbb45d22f),
	.w8(32'h3d7b1415),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c76ff),
	.w1(32'h3c296198),
	.w2(32'h3b385363),
	.w3(32'h3c7c4e1a),
	.w4(32'hbbb7f10a),
	.w5(32'hbd88cb8b),
	.w6(32'h3b575e44),
	.w7(32'hbc5021dd),
	.w8(32'hbc5e08bd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4485e0),
	.w1(32'h3c97a393),
	.w2(32'hbc52ebc1),
	.w3(32'hbc2b6da5),
	.w4(32'hbc1267ee),
	.w5(32'hbbfddf2c),
	.w6(32'hbc2714ff),
	.w7(32'hbc5fdcb1),
	.w8(32'hbc03a61b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf396f1),
	.w1(32'hb9e24066),
	.w2(32'h3d7c6ba7),
	.w3(32'h3b200360),
	.w4(32'h3a134ce0),
	.w5(32'hbb2a3eaf),
	.w6(32'h3be24400),
	.w7(32'hbb913e8b),
	.w8(32'hbc185602),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1556a2),
	.w1(32'h3c544c84),
	.w2(32'hbb39ee64),
	.w3(32'h3bdd51e4),
	.w4(32'hb89a8adc),
	.w5(32'hbb54a210),
	.w6(32'h3c965d50),
	.w7(32'hbb07abd1),
	.w8(32'hbb1164b5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb034462),
	.w1(32'hbaad8b54),
	.w2(32'h3bf51c58),
	.w3(32'hbbbb6d21),
	.w4(32'h3a0fa137),
	.w5(32'hbc2a828c),
	.w6(32'h3c441a0d),
	.w7(32'h3b85b1e9),
	.w8(32'hbc4b821b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1213f2),
	.w1(32'h3bcce949),
	.w2(32'h3b1eacc5),
	.w3(32'h3c455c00),
	.w4(32'h3c990e65),
	.w5(32'h3ab1fcf6),
	.w6(32'hbc018e24),
	.w7(32'h3aad44ce),
	.w8(32'h3c28dcc8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b33d3),
	.w1(32'hbbb0d664),
	.w2(32'h3c65d1a1),
	.w3(32'h3b14e343),
	.w4(32'hbc181955),
	.w5(32'h39c1ae7a),
	.w6(32'hbb19e10e),
	.w7(32'h3c41b585),
	.w8(32'hbbea5401),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab1a0a),
	.w1(32'h3bb076a4),
	.w2(32'h3b9acacc),
	.w3(32'hbb9797fe),
	.w4(32'hbb871b55),
	.w5(32'h3a7cdf21),
	.w6(32'hbb26ceae),
	.w7(32'h3aa5c100),
	.w8(32'h3c20fa16),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13325e),
	.w1(32'h3c267479),
	.w2(32'hbaee515e),
	.w3(32'h3c726a17),
	.w4(32'hb98034d5),
	.w5(32'h3bf187c3),
	.w6(32'h3b94106c),
	.w7(32'hbb119abe),
	.w8(32'h3ad3df5a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995a1f1),
	.w1(32'h39ab6b4a),
	.w2(32'hbbcdfd78),
	.w3(32'h3b97d012),
	.w4(32'hbc0c5abc),
	.w5(32'hbb2eb13d),
	.w6(32'h3b9919c9),
	.w7(32'hbc57dac9),
	.w8(32'h3b23cba3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4db861),
	.w1(32'hb81df3d2),
	.w2(32'h3b96ca03),
	.w3(32'h3b3efdf9),
	.w4(32'h3baf8bc2),
	.w5(32'h3c99b16d),
	.w6(32'hbbadb770),
	.w7(32'hbabafc1d),
	.w8(32'hbbb42989),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4aab1),
	.w1(32'h3c0ce0f9),
	.w2(32'hba8c104b),
	.w3(32'h38d1e94f),
	.w4(32'hbb89cdf8),
	.w5(32'h3bb9be34),
	.w6(32'hb9f96ae2),
	.w7(32'hbb5c74ef),
	.w8(32'h3b06193d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc324a50),
	.w1(32'h3b962019),
	.w2(32'hbca34e48),
	.w3(32'hba3b5e7a),
	.w4(32'hbad77e5a),
	.w5(32'hbb851eb1),
	.w6(32'hbb1b4a7a),
	.w7(32'hbc0a8a85),
	.w8(32'hbb5404a1),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ccccc),
	.w1(32'hbc257c5e),
	.w2(32'h3bb0b89b),
	.w3(32'h3a4ca642),
	.w4(32'h3ab99973),
	.w5(32'hbb7524f5),
	.w6(32'h3ba012f9),
	.w7(32'h3ba132ba),
	.w8(32'h3c81d7a7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5e748),
	.w1(32'hbb629ddc),
	.w2(32'hbc313333),
	.w3(32'hba124a4f),
	.w4(32'hba46352d),
	.w5(32'hbbf619d0),
	.w6(32'h3c0cbb29),
	.w7(32'h3be1542a),
	.w8(32'h3b94dd7e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c519530),
	.w1(32'h3ca67e52),
	.w2(32'h3a7df694),
	.w3(32'hbb518c9d),
	.w4(32'h3be180e6),
	.w5(32'h3c8dafae),
	.w6(32'hbb45d5b9),
	.w7(32'h3cda791f),
	.w8(32'h3c5f0483),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb1579),
	.w1(32'h3bbd6842),
	.w2(32'h3ab55d39),
	.w3(32'hbc6d6756),
	.w4(32'h3a89adc6),
	.w5(32'h38c33dfe),
	.w6(32'hbbe8abed),
	.w7(32'hbaff665d),
	.w8(32'h3986a9cc),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad40c74),
	.w1(32'hbbb1be51),
	.w2(32'h3c349265),
	.w3(32'hbc08603b),
	.w4(32'hba97bd1c),
	.w5(32'hb93ae389),
	.w6(32'hbb81c144),
	.w7(32'h3b97ac40),
	.w8(32'h3b19520b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27d5f9),
	.w1(32'hbb8bb7f5),
	.w2(32'hb977918a),
	.w3(32'h3c10b4ff),
	.w4(32'h3c8eb7b7),
	.w5(32'h3ba0c508),
	.w6(32'hbbfca773),
	.w7(32'hbbb6faad),
	.w8(32'h3b1b39cf),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a60bd),
	.w1(32'hbb233f9e),
	.w2(32'hbb8c6e39),
	.w3(32'h3c4e9282),
	.w4(32'hbad76858),
	.w5(32'h3b915f99),
	.w6(32'hbadd0242),
	.w7(32'h3b24cbc7),
	.w8(32'h3b537544),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20a4e6),
	.w1(32'h3ada9f92),
	.w2(32'h3b4b4711),
	.w3(32'hba6a81e4),
	.w4(32'h3aebc759),
	.w5(32'h3bd23615),
	.w6(32'hbbece860),
	.w7(32'hbb9d2489),
	.w8(32'hbab01e00),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87b0f0),
	.w1(32'hbc9722ae),
	.w2(32'h3c6d14ec),
	.w3(32'hbb1ba700),
	.w4(32'hbc5a9cfa),
	.w5(32'hbb105aa0),
	.w6(32'hbb654d65),
	.w7(32'hba0d223f),
	.w8(32'hbbdfd834),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fcc49),
	.w1(32'hbc8e9663),
	.w2(32'h3b2ce388),
	.w3(32'h3bb56e94),
	.w4(32'hbbfb4ef9),
	.w5(32'h3bcabd73),
	.w6(32'hbc4fcb4e),
	.w7(32'h38926796),
	.w8(32'h3bc8446f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule