module layer_6_featuremap_26(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdef3b),
	.w1(32'h3a30bd73),
	.w2(32'h3b9df21c),
	.w3(32'hbbf34003),
	.w4(32'h3c1229d4),
	.w5(32'h3cd054ee),
	.w6(32'hbc06e542),
	.w7(32'hbbef089d),
	.w8(32'hbc2e1b75),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64d429),
	.w1(32'h3c951ad6),
	.w2(32'h3c1cb62e),
	.w3(32'h3ce8b999),
	.w4(32'h3c0dae2c),
	.w5(32'h3a9a71e2),
	.w6(32'h3bec42ea),
	.w7(32'hbb599685),
	.w8(32'hbbc739d4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b923687),
	.w1(32'h3c808496),
	.w2(32'hbb4b46e8),
	.w3(32'h3a5b2a02),
	.w4(32'h3c611ee3),
	.w5(32'hbb682307),
	.w6(32'h3c881c3c),
	.w7(32'h3b5e6fc7),
	.w8(32'hbbdc99b8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4edce2),
	.w1(32'hbc207df2),
	.w2(32'hbc2f45a5),
	.w3(32'hbc299015),
	.w4(32'hbc0ffff6),
	.w5(32'hbc02bda6),
	.w6(32'h3c2404b0),
	.w7(32'h3b2e3557),
	.w8(32'hbb3198d1),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27aaeb),
	.w1(32'hbc02c778),
	.w2(32'h3aba36ed),
	.w3(32'h3bb81d6e),
	.w4(32'hbbad19e9),
	.w5(32'h3b6934ac),
	.w6(32'hbc301186),
	.w7(32'hbb21600f),
	.w8(32'h394ad2be),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d92d0),
	.w1(32'h3c01dbe8),
	.w2(32'hbb7a8cc7),
	.w3(32'h3b8b2470),
	.w4(32'h3b403386),
	.w5(32'hbbd83eba),
	.w6(32'hb8b1e4ea),
	.w7(32'hbbd352ee),
	.w8(32'hbb83c1ba),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb78f12),
	.w1(32'h3b0da351),
	.w2(32'h3af233bf),
	.w3(32'hbc23f0ca),
	.w4(32'h3a81779d),
	.w5(32'h3a3328cb),
	.w6(32'h3b37e36a),
	.w7(32'h3b4e45cc),
	.w8(32'h3bb97430),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba86773),
	.w1(32'h3a9564cb),
	.w2(32'hbaa64f00),
	.w3(32'h3b5666cb),
	.w4(32'h3b38f255),
	.w5(32'h3a2211e7),
	.w6(32'hbb39160e),
	.w7(32'h3b51411e),
	.w8(32'h3c319812),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c049b5b),
	.w1(32'hbb841985),
	.w2(32'hbab1e8a7),
	.w3(32'h3c0de51a),
	.w4(32'hbb5d0ebb),
	.w5(32'hbaa38547),
	.w6(32'hbbaba419),
	.w7(32'hbb1fe6ef),
	.w8(32'hb9833b1e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16af23),
	.w1(32'h3a7f5ccb),
	.w2(32'h3a8498bb),
	.w3(32'hbb0f6c43),
	.w4(32'hb8aaabaf),
	.w5(32'h390fda8e),
	.w6(32'h3b014837),
	.w7(32'h3ad7afe6),
	.w8(32'h3af3e651),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6de771),
	.w1(32'hbb72c52b),
	.w2(32'hbb0b51d0),
	.w3(32'h3b0f781e),
	.w4(32'hbb362b53),
	.w5(32'hbb83bdad),
	.w6(32'h39295566),
	.w7(32'h3ac22261),
	.w8(32'h3b524de2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1aaa0a),
	.w1(32'hbc7b7f85),
	.w2(32'h395abad8),
	.w3(32'hbb2af70f),
	.w4(32'hbc80373f),
	.w5(32'h3b622b9c),
	.w6(32'hbc07889a),
	.w7(32'hbbea0e7c),
	.w8(32'hbb248d11),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13d95d),
	.w1(32'h3c2681f8),
	.w2(32'h3ac14306),
	.w3(32'h3b88f530),
	.w4(32'h3c7d37bf),
	.w5(32'h3abab525),
	.w6(32'h3c324de7),
	.w7(32'h3b81d09a),
	.w8(32'hba82b1c2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87f05e),
	.w1(32'h3c0eabed),
	.w2(32'h3bf437c6),
	.w3(32'hbc003ff8),
	.w4(32'h3b92ea8f),
	.w5(32'h3c08fec3),
	.w6(32'h3bdf9333),
	.w7(32'h3c3e6b6b),
	.w8(32'h3c55f6a4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3331e9),
	.w1(32'h37f88950),
	.w2(32'hbc0ee619),
	.w3(32'h3c0dd25c),
	.w4(32'h3bfb731d),
	.w5(32'hbbae7fa3),
	.w6(32'h3b4853fd),
	.w7(32'hb9d8607e),
	.w8(32'hbc0b9f14),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bf74d),
	.w1(32'h3bbab661),
	.w2(32'hbc7b8b88),
	.w3(32'hbc403113),
	.w4(32'h3b8c4d95),
	.w5(32'hbc4fdc68),
	.w6(32'hb8a5edf5),
	.w7(32'hbc0742aa),
	.w8(32'hbc2b03f1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94add1),
	.w1(32'hbb83fe2a),
	.w2(32'h3bb10285),
	.w3(32'hbc86d475),
	.w4(32'hbc37a8d6),
	.w5(32'h3c18685f),
	.w6(32'hba603f14),
	.w7(32'h3c2204a2),
	.w8(32'h3ba5f624),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5531b6),
	.w1(32'hbc902749),
	.w2(32'hbcfdfb55),
	.w3(32'h3c763614),
	.w4(32'hbc026ca5),
	.w5(32'hbcafddb8),
	.w6(32'hbca31e93),
	.w7(32'hbcd6e470),
	.w8(32'hbcdcdb32),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0f41bc),
	.w1(32'hbc188014),
	.w2(32'hbb854c8c),
	.w3(32'hbce50feb),
	.w4(32'hbc0d6c8b),
	.w5(32'hbb4924e2),
	.w6(32'hbc325ab6),
	.w7(32'hbbae5e7b),
	.w8(32'hbb429524),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec4394),
	.w1(32'h3c5bbd51),
	.w2(32'h3c48b640),
	.w3(32'hbb0183b0),
	.w4(32'h3c7007dd),
	.w5(32'h3c0b6798),
	.w6(32'h3beb17e6),
	.w7(32'h3ac79687),
	.w8(32'h3b36c0fd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c0334),
	.w1(32'hbb9ccef8),
	.w2(32'hbb27d92b),
	.w3(32'h3c6851ce),
	.w4(32'h3ba0f259),
	.w5(32'h3b65232d),
	.w6(32'hbbe405a4),
	.w7(32'h3b04d636),
	.w8(32'h3b49a327),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389c7292),
	.w1(32'hbc2a1ba0),
	.w2(32'hbb56a097),
	.w3(32'h3b3ad945),
	.w4(32'hbbe5cc60),
	.w5(32'hbab56f60),
	.w6(32'hbc4584b0),
	.w7(32'hbbfe03c4),
	.w8(32'hbb3a4cf6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98577b1),
	.w1(32'hb9a01ad6),
	.w2(32'hbb51c6fe),
	.w3(32'h3a664a17),
	.w4(32'h3b27488d),
	.w5(32'hbaa92b74),
	.w6(32'hbb7b35e4),
	.w7(32'h385fd142),
	.w8(32'hb9f12a3e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3972b209),
	.w1(32'h3bb523b6),
	.w2(32'hbb4e3b95),
	.w3(32'h3b29a747),
	.w4(32'h3ad00a38),
	.w5(32'hbbf3a3a1),
	.w6(32'h3a8f3964),
	.w7(32'hbb929a39),
	.w8(32'hbb00f8e8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc98da2),
	.w1(32'hbb794fa4),
	.w2(32'hbba3e8e1),
	.w3(32'hbc83837d),
	.w4(32'h3b21627d),
	.w5(32'hbb422b47),
	.w6(32'hbb9b732c),
	.w7(32'hbb759e4c),
	.w8(32'h3a89bdbd),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde049b),
	.w1(32'h3be8d681),
	.w2(32'h3aa70939),
	.w3(32'h3bb97a85),
	.w4(32'h3c4df10d),
	.w5(32'h3a366493),
	.w6(32'h3c03db22),
	.w7(32'h3c062c4c),
	.w8(32'h394a5af6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb9330),
	.w1(32'h3c1e30e8),
	.w2(32'hbbff876d),
	.w3(32'hbbbebe5e),
	.w4(32'h3bea2876),
	.w5(32'hbbdf55f6),
	.w6(32'h3c91b851),
	.w7(32'h3c056f42),
	.w8(32'hbbe028cb),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f4657),
	.w1(32'h3b4ea1b3),
	.w2(32'hbc37811e),
	.w3(32'hbc58f0c2),
	.w4(32'hbaa1b4a7),
	.w5(32'hbc478217),
	.w6(32'h3bc3ed8c),
	.w7(32'hbb824cae),
	.w8(32'hbc1a32e9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68e098),
	.w1(32'h3c1567aa),
	.w2(32'h39d5261f),
	.w3(32'hbc4e0836),
	.w4(32'hbb0ba9c1),
	.w5(32'hbbf1f46e),
	.w6(32'h3c70c554),
	.w7(32'h3bc0699d),
	.w8(32'h3873f79d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcddd3c),
	.w1(32'h3c21e3c4),
	.w2(32'h3c4b5855),
	.w3(32'hbc0c778e),
	.w4(32'hbab35a94),
	.w5(32'h3c076145),
	.w6(32'h3c8896b8),
	.w7(32'h3bccde46),
	.w8(32'h3bc932cb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1af866),
	.w1(32'hb8531e5b),
	.w2(32'hb8814b02),
	.w3(32'h3b482857),
	.w4(32'hb8b37cdf),
	.w5(32'hb8e3235b),
	.w6(32'hb8976ba9),
	.w7(32'hb877970b),
	.w8(32'hb8b11ceb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01deb2),
	.w1(32'hb9aac1f5),
	.w2(32'hb8dfe739),
	.w3(32'hb9b9ef16),
	.w4(32'hb94d2f6c),
	.w5(32'hb6044a2f),
	.w6(32'hba089ecc),
	.w7(32'hb9f106bc),
	.w8(32'hb9da6106),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91136bd),
	.w1(32'hb8575610),
	.w2(32'hb722b0da),
	.w3(32'h3611bacd),
	.w4(32'hb6ec9ca4),
	.w5(32'h38473aa5),
	.w6(32'hb879d9d9),
	.w7(32'hb85e50ec),
	.w8(32'hb85d125c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38633f32),
	.w1(32'h3908b3ac),
	.w2(32'h3986f91a),
	.w3(32'h38bf2b75),
	.w4(32'h38b50716),
	.w5(32'h39689227),
	.w6(32'h390396d3),
	.w7(32'h39071347),
	.w8(32'h398558bb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9445929),
	.w1(32'hb8b0f0a0),
	.w2(32'h37a3f034),
	.w3(32'hb96796c5),
	.w4(32'hb9078657),
	.w5(32'h38e60f96),
	.w6(32'hb80d9a7d),
	.w7(32'hb90bf52f),
	.w8(32'h3823eb2a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67bfc9),
	.w1(32'hba083bc8),
	.w2(32'hb9e89359),
	.w3(32'hb99b645f),
	.w4(32'hb931d700),
	.w5(32'hb7bfecd0),
	.w6(32'hba05d0a4),
	.w7(32'hba3c290e),
	.w8(32'hba70a209),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379154b8),
	.w1(32'hb90b9dd3),
	.w2(32'hb9bd4dcb),
	.w3(32'h3792256f),
	.w4(32'hb875570e),
	.w5(32'hb98b5fca),
	.w6(32'hb99b322e),
	.w7(32'hb98af694),
	.w8(32'hb9eae542),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba417985),
	.w1(32'hb9b8f8e4),
	.w2(32'hba17dd7a),
	.w3(32'hb81581c0),
	.w4(32'h388b21fe),
	.w5(32'hb938b81c),
	.w6(32'hb9644fb2),
	.w7(32'hb93b0c05),
	.w8(32'hb9b6f51c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9302c1d),
	.w1(32'hb903af7f),
	.w2(32'hb6c2d21e),
	.w3(32'h391054b9),
	.w4(32'h398f4042),
	.w5(32'h39eb7ddb),
	.w6(32'h391cd980),
	.w7(32'h39b8a4c8),
	.w8(32'h3a103353),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9841b7),
	.w1(32'hbb356c63),
	.w2(32'hbb86f340),
	.w3(32'hbb79eb50),
	.w4(32'hbb58140a),
	.w5(32'hbb8615fe),
	.w6(32'hbb98cdbf),
	.w7(32'hbb8e04f8),
	.w8(32'hbb59b2d6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3706722d),
	.w1(32'h38c4f1cd),
	.w2(32'h39a0a7ec),
	.w3(32'h384f886c),
	.w4(32'h39aca284),
	.w5(32'h39d1cbaf),
	.w6(32'hb8f75fc0),
	.w7(32'h37b35eef),
	.w8(32'h3974c19b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b4c6b),
	.w1(32'hb9fad494),
	.w2(32'hba3bacbd),
	.w3(32'h37a7122c),
	.w4(32'hb9146c00),
	.w5(32'hba4c4815),
	.w6(32'h38cc2163),
	.w7(32'hb9ac73e0),
	.w8(32'hba4f06cd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb797f590),
	.w1(32'hb809bd31),
	.w2(32'hb81b3046),
	.w3(32'hb829e16e),
	.w4(32'hb82afbb7),
	.w5(32'hb88c758e),
	.w6(32'hb81155ae),
	.w7(32'hb810545d),
	.w8(32'hb84f08b0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba854c8e),
	.w1(32'hba795a2a),
	.w2(32'hbaa19642),
	.w3(32'hba90cfdd),
	.w4(32'hba4af018),
	.w5(32'hba635a93),
	.w6(32'hba777683),
	.w7(32'hba37c929),
	.w8(32'hba79d446),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0be3b5),
	.w1(32'h3a120d73),
	.w2(32'h3a5946ce),
	.w3(32'h3a5f6b9b),
	.w4(32'h3a78dcd2),
	.w5(32'h3a953b8c),
	.w6(32'h3a4f6b50),
	.w7(32'h3a04c661),
	.w8(32'h3a2403a9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376ec69d),
	.w1(32'h362e930d),
	.w2(32'h37816bb9),
	.w3(32'h36f9e3fc),
	.w4(32'h361c50a0),
	.w5(32'h371e374d),
	.w6(32'h36f513c1),
	.w7(32'hb6a57590),
	.w8(32'hb55c8905),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3751cd89),
	.w1(32'h363c2cb8),
	.w2(32'h37699a23),
	.w3(32'hb77ca2e6),
	.w4(32'hb850e7a7),
	.w5(32'h3754d56b),
	.w6(32'hb79e6aae),
	.w7(32'hb8500491),
	.w8(32'hb6cff514),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29b2fd),
	.w1(32'hb9e15767),
	.w2(32'hba05f42b),
	.w3(32'hb91bee71),
	.w4(32'hb89d02f9),
	.w5(32'hb96249e0),
	.w6(32'h39632079),
	.w7(32'h39e07921),
	.w8(32'h36e05548),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387a9d18),
	.w1(32'h375e0bd6),
	.w2(32'h390c3cd3),
	.w3(32'h39b8da02),
	.w4(32'h39b058c7),
	.w5(32'h39cdcdce),
	.w6(32'h39be2acc),
	.w7(32'h3a229989),
	.w8(32'h3a2835a2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03a085),
	.w1(32'h3a3e3882),
	.w2(32'h3a8f0b01),
	.w3(32'h3a91df33),
	.w4(32'h3ac66871),
	.w5(32'h3aec0e8e),
	.w6(32'h3aafb34d),
	.w7(32'h3addc6bb),
	.w8(32'h3b021695),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba840038),
	.w1(32'hbaa755bc),
	.w2(32'hbab3492d),
	.w3(32'hba52305b),
	.w4(32'hba61ac2b),
	.w5(32'hba7430c1),
	.w6(32'hba966a82),
	.w7(32'hba9f609e),
	.w8(32'hba9f2eef),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a188bdb),
	.w1(32'h39fba723),
	.w2(32'h399e4b97),
	.w3(32'h3a2c7990),
	.w4(32'h3a8be698),
	.w5(32'h3a5536d8),
	.w6(32'h3a48e983),
	.w7(32'h3aa231fb),
	.w8(32'h3abe4027),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9860a6f),
	.w1(32'hb8cd9429),
	.w2(32'h382281ef),
	.w3(32'h38eb8562),
	.w4(32'hb6e814db),
	.w5(32'hb8ad3e7d),
	.w6(32'h39163f91),
	.w7(32'h392d6a5d),
	.w8(32'h39a05998),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f8409),
	.w1(32'h3a0c7b3a),
	.w2(32'h3a25ae3f),
	.w3(32'h3aaab01b),
	.w4(32'h3aee7e11),
	.w5(32'h3b021d61),
	.w6(32'h3a8a3cec),
	.w7(32'h3ab74ab9),
	.w8(32'h3acfff8b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98075bd),
	.w1(32'hb9a6a4f7),
	.w2(32'h39d49bff),
	.w3(32'h39f1be0e),
	.w4(32'h3a60492c),
	.w5(32'h3aa3ad91),
	.w6(32'h39810f19),
	.w7(32'h3a537c42),
	.w8(32'h3ac46952),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7dee1),
	.w1(32'hbbd99d17),
	.w2(32'hbbdfdce3),
	.w3(32'hbbb9da8c),
	.w4(32'hbbc38d00),
	.w5(32'hbbe15d1a),
	.w6(32'hbb9cdfb3),
	.w7(32'hbb764a4c),
	.w8(32'hbb841c22),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60e787),
	.w1(32'h3b3093b9),
	.w2(32'h3b248245),
	.w3(32'h3b842ac4),
	.w4(32'h3b817e71),
	.w5(32'h3b90cebd),
	.w6(32'h3b6cf048),
	.w7(32'h3b2b991a),
	.w8(32'h3b392bac),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc178e71),
	.w1(32'hbc3795f0),
	.w2(32'hbc399630),
	.w3(32'hbc193b87),
	.w4(32'hbc38ee4c),
	.w5(32'hbc49b51d),
	.w6(32'hbc1b7a87),
	.w7(32'hbc47f777),
	.w8(32'hbc415934),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ea4f6),
	.w1(32'hb8cff759),
	.w2(32'h39fdf86a),
	.w3(32'h37482e02),
	.w4(32'h3a4771d1),
	.w5(32'h3a93359f),
	.w6(32'h3a02c94c),
	.w7(32'h39b58609),
	.w8(32'hba0f95e3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d62e8),
	.w1(32'h3ae6298a),
	.w2(32'h3b4f63c9),
	.w3(32'h3b32df8b),
	.w4(32'h3b7f233d),
	.w5(32'h3b95d84c),
	.w6(32'h3b00b2ef),
	.w7(32'h3b2e7c1d),
	.w8(32'h3b740bc6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb1098),
	.w1(32'hbbb5cfb6),
	.w2(32'hbc1c9628),
	.w3(32'hbc0d8191),
	.w4(32'hbc28f997),
	.w5(32'hbc1d593f),
	.w6(32'hbbaf4848),
	.w7(32'hbbeb5af9),
	.w8(32'hbbfbc3b6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf469af),
	.w1(32'hbae86708),
	.w2(32'hb8bff7f2),
	.w3(32'hbaca636f),
	.w4(32'hbaaaf9e9),
	.w5(32'h3a4dc419),
	.w6(32'hba894fcc),
	.w7(32'hba99e618),
	.w8(32'hba9e45cc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35ce2b),
	.w1(32'hbb69ddea),
	.w2(32'hbb41a926),
	.w3(32'hbb6ccfc8),
	.w4(32'hbb95341d),
	.w5(32'hbb87c925),
	.w6(32'hbb6df60e),
	.w7(32'hbb6b5002),
	.w8(32'hbb932d33),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9d5bf),
	.w1(32'h3a35b491),
	.w2(32'h3a598052),
	.w3(32'h3aaf953e),
	.w4(32'h3a84cfa2),
	.w5(32'h3aa1802b),
	.w6(32'h3953f4d8),
	.w7(32'h38524e02),
	.w8(32'h38b9245e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule