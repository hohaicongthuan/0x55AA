module layer_10_featuremap_152(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb620dca6),
	.w1(32'h3727e974),
	.w2(32'h36f9dd8e),
	.w3(32'hb7028740),
	.w4(32'h3764cf74),
	.w5(32'h370825b9),
	.w6(32'hb631e74e),
	.w7(32'h361207ed),
	.w8(32'hb6157933),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394611cc),
	.w1(32'hba4c9406),
	.w2(32'hba2aa476),
	.w3(32'h39fd7ce4),
	.w4(32'hb9de5403),
	.w5(32'hba17d8c8),
	.w6(32'h39855d3e),
	.w7(32'hb9ebf69a),
	.w8(32'hba00ec9a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb523ef46),
	.w1(32'h343de7c9),
	.w2(32'h361f29f0),
	.w3(32'hb5180fac),
	.w4(32'h35c7cbae),
	.w5(32'h367e4afa),
	.w6(32'hb6adf3b3),
	.w7(32'hb614bff6),
	.w8(32'hb5ae2b4a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932ba55),
	.w1(32'h397a1eba),
	.w2(32'h398da432),
	.w3(32'h38d7641f),
	.w4(32'h390d2c30),
	.w5(32'h3974878d),
	.w6(32'h38a3adf0),
	.w7(32'h39230052),
	.w8(32'h39897891),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eba9df),
	.w1(32'h38337055),
	.w2(32'h383dde70),
	.w3(32'h383f3f0b),
	.w4(32'h381be8e9),
	.w5(32'h380acf19),
	.w6(32'h37cfdcd5),
	.w7(32'h3822bdb6),
	.w8(32'h3805c51a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73cbb03),
	.w1(32'hb781c4c3),
	.w2(32'hb7b632c1),
	.w3(32'hb62f5527),
	.w4(32'hb6f50170),
	.w5(32'h36b1da27),
	.w6(32'hb73c42f5),
	.w7(32'hb71e9712),
	.w8(32'h36dc2dd8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acbae5),
	.w1(32'h39922afe),
	.w2(32'h39f62227),
	.w3(32'h39ac2c11),
	.w4(32'h39885d76),
	.w5(32'h3a810909),
	.w6(32'h3a05c260),
	.w7(32'h3a0fffde),
	.w8(32'h3a7fb866),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93cc5c),
	.w1(32'h3ab68e5e),
	.w2(32'h3b2f469f),
	.w3(32'h3b286673),
	.w4(32'h3b1dca93),
	.w5(32'h3ad1dffb),
	.w6(32'h3b78d753),
	.w7(32'h3b8ec2e0),
	.w8(32'h3b4ba55e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb823878e),
	.w1(32'h381c1d9d),
	.w2(32'hb92a9a0d),
	.w3(32'h397493ee),
	.w4(32'h390cd966),
	.w5(32'hb9129c50),
	.w6(32'h39aab108),
	.w7(32'h3932dd87),
	.w8(32'hb98a551d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9301ce7),
	.w1(32'hbb32ff9d),
	.w2(32'hbb856d39),
	.w3(32'hb98a36ff),
	.w4(32'hbb272c0c),
	.w5(32'hbb22ae91),
	.w6(32'h3a0b2ebf),
	.w7(32'hba1dd09b),
	.w8(32'hbab6e68a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36214f70),
	.w1(32'hb851443b),
	.w2(32'h37f74411),
	.w3(32'h38c4e11f),
	.w4(32'hb6a4f0df),
	.w5(32'h383d138d),
	.w6(32'hb8e9899f),
	.w7(32'hb92f9d37),
	.w8(32'hb88edf61),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93efee),
	.w1(32'h3ac1fe05),
	.w2(32'h3abb8273),
	.w3(32'h3a98b458),
	.w4(32'h3ad13b22),
	.w5(32'h3b03052c),
	.w6(32'h3aa76bf8),
	.w7(32'h3a8f51c4),
	.w8(32'h3b0acfc8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98dcae),
	.w1(32'hbb434307),
	.w2(32'hbb865f59),
	.w3(32'hba97eb74),
	.w4(32'hbb391308),
	.w5(32'hbb365e8e),
	.w6(32'hba01e92b),
	.w7(32'hba8d46bd),
	.w8(32'hbb058501),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9221a),
	.w1(32'hba47b6bf),
	.w2(32'h3a1d8ffc),
	.w3(32'h3975217a),
	.w4(32'hb87a38b5),
	.w5(32'h3a2b0d87),
	.w6(32'h396cd9b2),
	.w7(32'hb95034e5),
	.w8(32'h39b9d12b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbdb5f),
	.w1(32'hba6886b3),
	.w2(32'hba27197b),
	.w3(32'hba09371e),
	.w4(32'hba779fcd),
	.w5(32'hb98c65ec),
	.w6(32'h39b32270),
	.w7(32'h39d2b57a),
	.w8(32'h39a8fd44),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72f477),
	.w1(32'hbaaf95af),
	.w2(32'hbb12c2fc),
	.w3(32'h3aa1acfc),
	.w4(32'hba46ea70),
	.w5(32'hbabfb34c),
	.w6(32'h3add2eaa),
	.w7(32'h39d69d5d),
	.w8(32'hb9c43230),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82cc412),
	.w1(32'hb92bac66),
	.w2(32'hb8900f76),
	.w3(32'hb944d29f),
	.w4(32'hb95f0753),
	.w5(32'h37ce4488),
	.w6(32'hb9a7a26b),
	.w7(32'hb9b8d17f),
	.w8(32'h38073663),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b339a2f),
	.w1(32'h3b4eb6df),
	.w2(32'h3b87d6f8),
	.w3(32'h3b871760),
	.w4(32'h3b72a6fd),
	.w5(32'h3b82fc11),
	.w6(32'h3bda400b),
	.w7(32'h3bd0c626),
	.w8(32'h3bd4138d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c844a3),
	.w1(32'hb9ed2a53),
	.w2(32'hba82cf16),
	.w3(32'h3aa03f64),
	.w4(32'hb940d1d3),
	.w5(32'hba4570a6),
	.w6(32'h3b011da3),
	.w7(32'h3ab52074),
	.w8(32'h3a72adc9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5cf1064),
	.w1(32'hb69bcaed),
	.w2(32'hb7201c66),
	.w3(32'hb717e670),
	.w4(32'h363501d2),
	.w5(32'hb6d419a4),
	.w6(32'hb71cdbfb),
	.w7(32'h3722c70f),
	.w8(32'h368cef2e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66ab4d7),
	.w1(32'h37a79b10),
	.w2(32'h37147b95),
	.w3(32'hb7d12c56),
	.w4(32'h37bcb3fe),
	.w5(32'h3609a14a),
	.w6(32'h370e963a),
	.w7(32'h379b1c2f),
	.w8(32'hb790026e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a17bf5),
	.w1(32'hb8ff46e7),
	.w2(32'hb8983f2d),
	.w3(32'hb81f7859),
	.w4(32'hb88ebc23),
	.w5(32'hb8633a44),
	.w6(32'hb8fde180),
	.w7(32'hb99108a2),
	.w8(32'hb975f865),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa8471),
	.w1(32'h3bab66c5),
	.w2(32'h3b9a8820),
	.w3(32'h3bff4d4c),
	.w4(32'h3baf0585),
	.w5(32'h3bd3453c),
	.w6(32'h3c2397fa),
	.w7(32'h3bf6c9bc),
	.w8(32'h3c27b8ac),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec5bde),
	.w1(32'hbb302a2d),
	.w2(32'hbb81eef0),
	.w3(32'hb8264c0f),
	.w4(32'hbb0c5b60),
	.w5(32'hbb177095),
	.w6(32'h3a336747),
	.w7(32'hba41ed67),
	.w8(32'hba963602),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb716e1f4),
	.w1(32'hbb2534da),
	.w2(32'hbb555be5),
	.w3(32'h3a09644c),
	.w4(32'hbae9ed88),
	.w5(32'hbb13385f),
	.w6(32'h3a1e8076),
	.w7(32'hbab3454b),
	.w8(32'hbab821e5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39181720),
	.w1(32'hb8cb1e30),
	.w2(32'hb918fba5),
	.w3(32'hb880533f),
	.w4(32'hb99c55e4),
	.w5(32'hb92c2abc),
	.w6(32'hb9127efc),
	.w7(32'h35b7e229),
	.w8(32'hb923fc27),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7331149),
	.w1(32'h373bf8c8),
	.w2(32'h383bed6e),
	.w3(32'hb5376453),
	.w4(32'h37efc734),
	.w5(32'h386187e1),
	.w6(32'hb7d0c15b),
	.w7(32'hb308c33e),
	.w8(32'h38115337),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2fa97),
	.w1(32'h397efc67),
	.w2(32'h39948bd1),
	.w3(32'hba1d0012),
	.w4(32'hba1df8a7),
	.w5(32'hb80be2a1),
	.w6(32'hbae39774),
	.w7(32'hba827e2a),
	.w8(32'hb8ea9929),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbe1d3),
	.w1(32'h3a4894b7),
	.w2(32'h3a193548),
	.w3(32'h3a03513a),
	.w4(32'h3a99f908),
	.w5(32'h3a3e505d),
	.w6(32'h39da29e6),
	.w7(32'h3a2b10bf),
	.w8(32'h39784855),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9630127),
	.w1(32'hbb224f54),
	.w2(32'hbb377ef1),
	.w3(32'hba533efe),
	.w4(32'hbb2a4f2b),
	.w5(32'hbb1108b9),
	.w6(32'hbab7ce87),
	.w7(32'hbb050bfc),
	.w8(32'hbadec120),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368ed9a8),
	.w1(32'hb745a234),
	.w2(32'hb63accf1),
	.w3(32'h35ea3d96),
	.w4(32'hb7649e2a),
	.w5(32'hb6664863),
	.w6(32'hb7325329),
	.w7(32'hb7ccd26d),
	.w8(32'hb77421a0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b942d9),
	.w1(32'hb80e0cb4),
	.w2(32'h37290384),
	.w3(32'h379a741c),
	.w4(32'hb84aef17),
	.w5(32'hb7ace5a5),
	.w6(32'hb89e0f3e),
	.w7(32'hb8c8233e),
	.w8(32'hb78f2702),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d835d3),
	.w1(32'hba1f2690),
	.w2(32'hba8b3164),
	.w3(32'h3a2285bd),
	.w4(32'hb950cce8),
	.w5(32'hb98c1595),
	.w6(32'h3a833ad9),
	.w7(32'h3a32f8bd),
	.w8(32'h3a0a3a51),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eefb6b),
	.w1(32'hba8653d1),
	.w2(32'hba4767dc),
	.w3(32'hb9c81b10),
	.w4(32'hba4a1af8),
	.w5(32'hba3a37e9),
	.w6(32'hb9842952),
	.w7(32'hba29a951),
	.w8(32'hba179b95),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972e1b3),
	.w1(32'hb808033f),
	.w2(32'hb8c1e9a0),
	.w3(32'hb91a093b),
	.w4(32'hb88cf259),
	.w5(32'hb8e93081),
	.w6(32'hb9ebbdb7),
	.w7(32'hb998fa39),
	.w8(32'hb978a9ae),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d6eb5),
	.w1(32'h399b061f),
	.w2(32'hb7ccc359),
	.w3(32'h39b63944),
	.w4(32'h39e0d68b),
	.w5(32'h39022188),
	.w6(32'h3a25294f),
	.w7(32'h3a095c4a),
	.w8(32'h39fb7678),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ee525),
	.w1(32'h3aee38ce),
	.w2(32'hb920abdf),
	.w3(32'h3a9628c7),
	.w4(32'h3a6e952c),
	.w5(32'hba82e572),
	.w6(32'h3afbc31d),
	.w7(32'h3b18380b),
	.w8(32'h3a9fde65),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacad011),
	.w1(32'hbb2bfb8e),
	.w2(32'hba7d3590),
	.w3(32'hb7127ddf),
	.w4(32'hba360f79),
	.w5(32'hb90b5906),
	.w6(32'hba28e8d7),
	.w7(32'hba0fe29d),
	.w8(32'h3a273d35),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5ff2b),
	.w1(32'hbadf03d7),
	.w2(32'h3aca5c6a),
	.w3(32'hbad5fbc7),
	.w4(32'hba21e62f),
	.w5(32'h3add5b73),
	.w6(32'hbaf2e409),
	.w7(32'hbacc40cb),
	.w8(32'h3a1b02a4),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ccad5),
	.w1(32'hb9b4f898),
	.w2(32'hb99e7d9c),
	.w3(32'hb90eb8da),
	.w4(32'hb935a678),
	.w5(32'h398b1439),
	.w6(32'h38ff5d98),
	.w7(32'h399dde53),
	.w8(32'h3a254368),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73377c8),
	.w1(32'hb8cbcba1),
	.w2(32'hb864fecb),
	.w3(32'hb84b7d51),
	.w4(32'hb8df0ac7),
	.w5(32'hb8bebec1),
	.w6(32'hb8b73bf7),
	.w7(32'hb888462e),
	.w8(32'hb8abf3f6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85feaa1),
	.w1(32'h38591f50),
	.w2(32'h3865cf63),
	.w3(32'hb8310917),
	.w4(32'h38900d60),
	.w5(32'h383a6ecb),
	.w6(32'hb888fdfa),
	.w7(32'h3783f2de),
	.w8(32'h3719d622),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8701d6),
	.w1(32'h3a8bf8df),
	.w2(32'h3a97211d),
	.w3(32'h3a845dbb),
	.w4(32'h3a823ba2),
	.w5(32'h3a97302d),
	.w6(32'h3a1fd9e7),
	.w7(32'h3a175abf),
	.w8(32'h38e57e88),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a588d4),
	.w1(32'hbac6770c),
	.w2(32'hbb0a2857),
	.w3(32'h396d9295),
	.w4(32'h3932a2f7),
	.w5(32'hba5f2c0f),
	.w6(32'h3aed0d47),
	.w7(32'h3ae97905),
	.w8(32'h3a52b3ea),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edc9e5),
	.w1(32'hbb29f0cc),
	.w2(32'hbb64b4cf),
	.w3(32'hb92459c3),
	.w4(32'hbb054079),
	.w5(32'hbb16a38f),
	.w6(32'hb8a3ff72),
	.w7(32'hba83c577),
	.w8(32'hbab9dd82),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90269af),
	.w1(32'hbb4704ea),
	.w2(32'hbb927ec9),
	.w3(32'h39488771),
	.w4(32'hbb170fb6),
	.w5(32'hbb462c66),
	.w6(32'h3a8c78f7),
	.w7(32'hba408f3a),
	.w8(32'hbad0071b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a99bb7),
	.w1(32'hba98e159),
	.w2(32'hbaf54cbe),
	.w3(32'h3a8762e3),
	.w4(32'hb9ae2eb7),
	.w5(32'hba5e21c3),
	.w6(32'h3aea6753),
	.w7(32'h39dd809b),
	.w8(32'h3a52abf9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b998144),
	.w1(32'h3b59c7ac),
	.w2(32'h3b1d4544),
	.w3(32'h3ba7556c),
	.w4(32'h3b3ebb8c),
	.w5(32'h3b2fe692),
	.w6(32'h3bed136b),
	.w7(32'h3bd22ad2),
	.w8(32'h3bc1ea20),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378052d2),
	.w1(32'h38195844),
	.w2(32'hb8312f02),
	.w3(32'hb886723a),
	.w4(32'h38d15525),
	.w5(32'hb76fd88f),
	.w6(32'h38a50114),
	.w7(32'h38c459ce),
	.w8(32'h36846c6d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39374bbe),
	.w1(32'h396eba6e),
	.w2(32'h382565fa),
	.w3(32'h3913f171),
	.w4(32'h3923b8a0),
	.w5(32'hb173d220),
	.w6(32'h3997d2d6),
	.w7(32'h3922bf2e),
	.w8(32'h38881546),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b25a69),
	.w1(32'h39596329),
	.w2(32'h394144fe),
	.w3(32'h39732ee4),
	.w4(32'h396c5c6a),
	.w5(32'h398d347d),
	.w6(32'h39958396),
	.w7(32'h399ff67d),
	.w8(32'h39ae8ff9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dda4ad),
	.w1(32'hba21b363),
	.w2(32'hba9abcc5),
	.w3(32'h39db11d7),
	.w4(32'hb9d50c5f),
	.w5(32'hb9de5381),
	.w6(32'h3a403e94),
	.w7(32'h388aedf8),
	.w8(32'h39459ea6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0225e5),
	.w1(32'h39edd342),
	.w2(32'h39b9cb32),
	.w3(32'h3a3b4a6c),
	.w4(32'h3a149a9d),
	.w5(32'h39b829e4),
	.w6(32'h3a802b12),
	.w7(32'h3a49ace4),
	.w8(32'h3a77c424),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd2d27),
	.w1(32'h3aa3c3dc),
	.w2(32'h39a0ffde),
	.w3(32'h3b363ecd),
	.w4(32'h3b1ed638),
	.w5(32'h3b0aff1b),
	.w6(32'h3ba313bf),
	.w7(32'h3bad0a9c),
	.w8(32'h3b951120),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d66d7),
	.w1(32'h3a1eedd7),
	.w2(32'h3a2acd6f),
	.w3(32'h3a0c31b6),
	.w4(32'h3a34b564),
	.w5(32'h3a3f2b15),
	.w6(32'h3a297b4b),
	.w7(32'h3a6689d5),
	.w8(32'h3a877c18),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3891e892),
	.w1(32'hb823cb1b),
	.w2(32'hb860a640),
	.w3(32'h37a92e8e),
	.w4(32'hb83cfb60),
	.w5(32'hb708358f),
	.w6(32'h3754c3c5),
	.w7(32'hb79bad65),
	.w8(32'hb811b29a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68dea6a),
	.w1(32'hb7e50876),
	.w2(32'hb7f1f262),
	.w3(32'h37ca9fd9),
	.w4(32'hb50fcaf4),
	.w5(32'hb6e99393),
	.w6(32'h37e64308),
	.w7(32'h36aa1b08),
	.w8(32'hb7b403aa),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8850893),
	.w1(32'h3644785e),
	.w2(32'h38ae4f30),
	.w3(32'hb8aceffa),
	.w4(32'hb7b5df4b),
	.w5(32'h39063bc6),
	.w6(32'hb8ea2894),
	.w7(32'hb85deb3c),
	.w8(32'h388e2821),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fa4168),
	.w1(32'h390d81b1),
	.w2(32'h399ad78b),
	.w3(32'h390678ff),
	.w4(32'h399fd0b8),
	.w5(32'h39bf9a21),
	.w6(32'hb85a83e4),
	.w7(32'h3900b8b1),
	.w8(32'h392d692f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8adeac3),
	.w1(32'hb8dd30e4),
	.w2(32'h38bae8be),
	.w3(32'hb8d46c95),
	.w4(32'hb88217a8),
	.w5(32'h3962d971),
	.w6(32'hb959049c),
	.w7(32'hb89ccfe7),
	.w8(32'h3993b2f6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8914874),
	.w1(32'h3a32c0da),
	.w2(32'h3a6bd0a1),
	.w3(32'hb87bf57e),
	.w4(32'h3a0de22d),
	.w5(32'h3a0869e2),
	.w6(32'h3a2404d5),
	.w7(32'h3a83818b),
	.w8(32'h3a9d026c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab48aae),
	.w1(32'h3b00f18d),
	.w2(32'h3add18f3),
	.w3(32'h3b05442b),
	.w4(32'h3ae4f6d4),
	.w5(32'h3b1202e3),
	.w6(32'h3af94ec8),
	.w7(32'h3b1c1186),
	.w8(32'h3b15c84a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a9ca92),
	.w1(32'hb68264a6),
	.w2(32'hb76582eb),
	.w3(32'hb77ec2a1),
	.w4(32'hb793fd27),
	.w5(32'hb70b2090),
	.w6(32'hb76c54fd),
	.w7(32'hb7257c3e),
	.w8(32'h3764e0d5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70c03d5),
	.w1(32'hb5d0cabb),
	.w2(32'h35e31a10),
	.w3(32'hb744e162),
	.w4(32'hb7256a2e),
	.w5(32'h356dc5af),
	.w6(32'hb7212388),
	.w7(32'hb6f4381c),
	.w8(32'hb62293df),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39031eb4),
	.w1(32'h38ca7cd3),
	.w2(32'h387e15cd),
	.w3(32'h391f5053),
	.w4(32'h38f26b7e),
	.w5(32'h385318e7),
	.w6(32'h38cad632),
	.w7(32'h38989edb),
	.w8(32'h388ca95e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75c2fd9),
	.w1(32'hb72dfab6),
	.w2(32'h37ab0c25),
	.w3(32'hb786b48a),
	.w4(32'hb739e10a),
	.w5(32'h375aa053),
	.w6(32'hb7c02426),
	.w7(32'hb7654649),
	.w8(32'hb6cc8a50),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a773117),
	.w1(32'h3a762c7d),
	.w2(32'h3809cba9),
	.w3(32'h3aa3a1c7),
	.w4(32'h3a7fc96d),
	.w5(32'h3a53f0f8),
	.w6(32'h3a8be850),
	.w7(32'h3ad3dec5),
	.w8(32'h3ae6956c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3942af6f),
	.w1(32'hbb096b51),
	.w2(32'hbb3826f8),
	.w3(32'h3aa38dd7),
	.w4(32'hba302e5b),
	.w5(32'hbaf04cfd),
	.w6(32'h3b0060b6),
	.w7(32'hb81728f3),
	.w8(32'h37e3322f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02c4f3),
	.w1(32'h3b55e5ee),
	.w2(32'h3b4cd9e5),
	.w3(32'h3b6ec175),
	.w4(32'h3b84226f),
	.w5(32'h3b6cd8b7),
	.w6(32'h3bc018f0),
	.w7(32'h3bc0d94e),
	.w8(32'h3bbd673d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dde8bb),
	.w1(32'hbb7381bd),
	.w2(32'hbbaf4974),
	.w3(32'h396a3546),
	.w4(32'hbb527879),
	.w5(32'hbb8e793c),
	.w6(32'h3a552a89),
	.w7(32'hbae76f4e),
	.w8(32'hbb30f1c9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364e3132),
	.w1(32'h3716efc3),
	.w2(32'h37961d6e),
	.w3(32'hb7221984),
	.w4(32'hb773f2c6),
	.w5(32'h36be59e3),
	.w6(32'hb78db41e),
	.w7(32'hb7767b1e),
	.w8(32'h36c632d6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d32f6f),
	.w1(32'h3776b825),
	.w2(32'h37dfb5e4),
	.w3(32'hb70f8e9e),
	.w4(32'hb5a570ac),
	.w5(32'h375854ca),
	.w6(32'hb802d62b),
	.w7(32'hb767d25f),
	.w8(32'hb6783831),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bd51b3),
	.w1(32'hb6af0ed9),
	.w2(32'h36e31635),
	.w3(32'hb875b051),
	.w4(32'hb7f4a961),
	.w5(32'hb77e9556),
	.w6(32'hb8747547),
	.w7(32'hb825cb07),
	.w8(32'hb81afb92),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3868b28d),
	.w1(32'h39b65118),
	.w2(32'h39862404),
	.w3(32'h3a0b395d),
	.w4(32'h3a0b10da),
	.w5(32'h3879cffe),
	.w6(32'h39e06ee1),
	.w7(32'h3a2f85dc),
	.w8(32'h39921686),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73d3051),
	.w1(32'h380050eb),
	.w2(32'h37631b04),
	.w3(32'hb79fce40),
	.w4(32'h382ea678),
	.w5(32'h37a584b9),
	.w6(32'hb7bc9cfb),
	.w7(32'h380490b0),
	.w8(32'h37add70a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b731b),
	.w1(32'h3b54842c),
	.w2(32'h3b12726b),
	.w3(32'h3b214192),
	.w4(32'h3b120d6d),
	.w5(32'h3aeb0407),
	.w6(32'h3b460d7f),
	.w7(32'h3b5e7bfb),
	.w8(32'h3b7069a2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f63c2),
	.w1(32'h3b4695ac),
	.w2(32'h3b500019),
	.w3(32'h3b2314e4),
	.w4(32'h3b38f489),
	.w5(32'h3b1127c3),
	.w6(32'h3b83fb85),
	.w7(32'h3b90523d),
	.w8(32'h3b9c2e55),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9975786),
	.w1(32'hbb375315),
	.w2(32'hbb7c70f9),
	.w3(32'hb998f543),
	.w4(32'hbb3832ca),
	.w5(32'hbb54e1f7),
	.w6(32'hba2f0c48),
	.w7(32'hbaf17dc3),
	.w8(32'hbb4483df),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39898e03),
	.w1(32'h3800f385),
	.w2(32'h37cf206f),
	.w3(32'h3a934197),
	.w4(32'h3a44db45),
	.w5(32'h3a1167af),
	.w6(32'h3ae4dc5e),
	.w7(32'h3ae7375f),
	.w8(32'h3a9f9674),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65d35b),
	.w1(32'h38cc6bda),
	.w2(32'hba893bd2),
	.w3(32'h3a82e0b8),
	.w4(32'h382c54c7),
	.w5(32'hb9ddcca6),
	.w6(32'h39e047dd),
	.w7(32'h39b36220),
	.w8(32'h387f321c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921a501),
	.w1(32'hba3eadb3),
	.w2(32'hba7e4ce5),
	.w3(32'hb97b04ae),
	.w4(32'hba34750c),
	.w5(32'hba1d5d0b),
	.w6(32'hb9779466),
	.w7(32'hb99a265e),
	.w8(32'hba029b6d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6b5ed),
	.w1(32'h3aca49bd),
	.w2(32'h3aa8e947),
	.w3(32'h3acd1c3a),
	.w4(32'h3a95c16c),
	.w5(32'h3a94f7e5),
	.w6(32'h3b0cb9ff),
	.w7(32'h3afe97c1),
	.w8(32'h3ada8957),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bac5d7),
	.w1(32'hb64928ed),
	.w2(32'hb60f4dba),
	.w3(32'hb6f6de49),
	.w4(32'hb59444b5),
	.w5(32'hb5a9fce2),
	.w6(32'hb7025723),
	.w7(32'hb6af5b18),
	.w8(32'hb6571898),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37465fe5),
	.w1(32'hb50ebddf),
	.w2(32'hb7199837),
	.w3(32'h36da5950),
	.w4(32'h32c6acba),
	.w5(32'h36485908),
	.w6(32'hb5014755),
	.w7(32'h36446a14),
	.w8(32'h368598b8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe5e27),
	.w1(32'hb98b7d7a),
	.w2(32'hb93aa4d7),
	.w3(32'hb923a8ac),
	.w4(32'hb9865f39),
	.w5(32'hb93baa63),
	.w6(32'hb950a572),
	.w7(32'hb96e3bdf),
	.w8(32'hb946fb52),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84f1141),
	.w1(32'h3814227b),
	.w2(32'h38abb89d),
	.w3(32'hb8881041),
	.w4(32'h37deb095),
	.w5(32'h38bc326b),
	.w6(32'hb8f30b15),
	.w7(32'hb8093124),
	.w8(32'h38000900),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3878ad07),
	.w1(32'hbaa1d100),
	.w2(32'hbb09f754),
	.w3(32'h39d57ad5),
	.w4(32'hba93261f),
	.w5(32'hba9cb742),
	.w6(32'h3a3cd1aa),
	.w7(32'h38c0fe5d),
	.w8(32'h3a050b0b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d7e7b),
	.w1(32'hb91406df),
	.w2(32'h38135ee9),
	.w3(32'hb87bd674),
	.w4(32'h39356749),
	.w5(32'h396fc2e2),
	.w6(32'hb8e3b5fc),
	.w7(32'hb8b8df21),
	.w8(32'h3922252a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a301011),
	.w1(32'hba49b071),
	.w2(32'hbac5cb11),
	.w3(32'h3ab47205),
	.w4(32'hb8d14bbe),
	.w5(32'hb9e7a15b),
	.w6(32'h3ae85651),
	.w7(32'h3a490b38),
	.w8(32'h3a36bfd1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6157d4),
	.w1(32'h3b82bc2f),
	.w2(32'h3ba1f0e8),
	.w3(32'h3b99adc8),
	.w4(32'h3b8af8b6),
	.w5(32'h3bbca4b5),
	.w6(32'h3bd756b6),
	.w7(32'h3be017d9),
	.w8(32'h3bf46792),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba038cd0),
	.w1(32'hb923e059),
	.w2(32'h39c98bb4),
	.w3(32'hba03901a),
	.w4(32'h390df90b),
	.w5(32'h3a297b4e),
	.w6(32'hba3d7cfa),
	.w7(32'hb9f5bf22),
	.w8(32'h399973c1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377a0436),
	.w1(32'hb969a4d1),
	.w2(32'hb98e0b5e),
	.w3(32'h39fd7729),
	.w4(32'hb9134738),
	.w5(32'hb870fb84),
	.w6(32'h3ae56ef7),
	.w7(32'h3a80854e),
	.w8(32'h3b286d0c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f8f6f),
	.w1(32'hb91ad328),
	.w2(32'hba95c2e8),
	.w3(32'h39d55d13),
	.w4(32'h394d4a25),
	.w5(32'hba12bf83),
	.w6(32'h397f9dfc),
	.w7(32'h39e3d1d0),
	.w8(32'h38e2254a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23d75c),
	.w1(32'hba2a4749),
	.w2(32'hba196197),
	.w3(32'h3b125a0c),
	.w4(32'h3a6e4cab),
	.w5(32'h3a2900aa),
	.w6(32'h3b939574),
	.w7(32'h3b54051e),
	.w8(32'h3b2b7e9b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6788c),
	.w1(32'h3a2d0a8d),
	.w2(32'hb93dd0e7),
	.w3(32'h3adad79b),
	.w4(32'h3a44b96b),
	.w5(32'h3a51ca37),
	.w6(32'h3ac6048e),
	.w7(32'h3a9e8c5c),
	.w8(32'h3afeddfd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a531bb),
	.w1(32'hbae53379),
	.w2(32'hba5c8327),
	.w3(32'hb9563816),
	.w4(32'hba9ba4de),
	.w5(32'hb8e9d4a3),
	.w6(32'h38054584),
	.w7(32'hb975a7d2),
	.w8(32'h3a2a6c27),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f9da63),
	.w1(32'h38c98c57),
	.w2(32'hb79dcf5c),
	.w3(32'h3907426f),
	.w4(32'h3800990b),
	.w5(32'hb8f3e188),
	.w6(32'h383f1637),
	.w7(32'hb83e5ed2),
	.w8(32'hb8c8a470),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917d785),
	.w1(32'hba8c49e7),
	.w2(32'hbad82cee),
	.w3(32'h3a9d7c17),
	.w4(32'hb821ac96),
	.w5(32'hba558aeb),
	.w6(32'h3b3dc69b),
	.w7(32'h3afb44b2),
	.w8(32'h3ad34e50),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a84ba),
	.w1(32'h3a72cf3e),
	.w2(32'hb8e8f3b6),
	.w3(32'h3ac34fba),
	.w4(32'h3a550f25),
	.w5(32'h3ad44840),
	.w6(32'h3b46e531),
	.w7(32'h3aecfed7),
	.w8(32'h3b5d0ab5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af44a3d),
	.w1(32'h3b51b0f7),
	.w2(32'h3aab8bee),
	.w3(32'h3b8b2139),
	.w4(32'h3b94a804),
	.w5(32'h3b0f1e28),
	.w6(32'h3bce5ac1),
	.w7(32'h3baa45ab),
	.w8(32'h3b9c7785),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae641d),
	.w1(32'h3aafa441),
	.w2(32'h3b233fa4),
	.w3(32'h3ae901a6),
	.w4(32'h3a2557e6),
	.w5(32'h3b314cc5),
	.w6(32'h3b3372b9),
	.w7(32'h3abdafe8),
	.w8(32'h3b8d585c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f5214f),
	.w1(32'hbb6646ba),
	.w2(32'hbb9ce672),
	.w3(32'hb8af510e),
	.w4(32'hbb40af6f),
	.w5(32'hbb7cb850),
	.w6(32'h3a041444),
	.w7(32'hbaca0522),
	.w8(32'hbb29af5a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa56c58),
	.w1(32'h3a92668e),
	.w2(32'h3a36a673),
	.w3(32'h3af7da30),
	.w4(32'h3ab1b135),
	.w5(32'h3aa64d22),
	.w6(32'h3b625479),
	.w7(32'h3b6de249),
	.w8(32'h3b863b42),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f4151),
	.w1(32'h391c9c36),
	.w2(32'h3792617e),
	.w3(32'hb90f4c6a),
	.w4(32'h38ca2e32),
	.w5(32'hb8ceadff),
	.w6(32'hb90942a7),
	.w7(32'hb93f2d32),
	.w8(32'h36e1803b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ede6c),
	.w1(32'h3bbee6c7),
	.w2(32'h3b9a21d7),
	.w3(32'h3b951e50),
	.w4(32'h3b8bf672),
	.w5(32'h3b3ba368),
	.w6(32'h3b880863),
	.w7(32'h3bc5acf1),
	.w8(32'h3bc1e742),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981bf5a),
	.w1(32'hb7ce640a),
	.w2(32'hba542bee),
	.w3(32'hb9f074ec),
	.w4(32'hba735e22),
	.w5(32'hba0e4920),
	.w6(32'hba20baed),
	.w7(32'hbac79d2a),
	.w8(32'hb9038895),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77fd7f8),
	.w1(32'hb7e2a3fe),
	.w2(32'h3719b8b8),
	.w3(32'hb7c81c3d),
	.w4(32'hb7be9129),
	.w5(32'h379570ec),
	.w6(32'hb81e9b84),
	.w7(32'hb87326ea),
	.w8(32'hb7d9dd56),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a40bb1),
	.w1(32'hb9d65d6d),
	.w2(32'hb93546cf),
	.w3(32'h393d90bb),
	.w4(32'hb9895c68),
	.w5(32'hb88c5669),
	.w6(32'h3a4dab4d),
	.w7(32'h39332a68),
	.w8(32'h392288c7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eeb3ae),
	.w1(32'hbb0472c3),
	.w2(32'hbb3aaf6d),
	.w3(32'h3941263a),
	.w4(32'hbaa9ed9d),
	.w5(32'hbb065212),
	.w6(32'h3a33edec),
	.w7(32'h37a3ea6a),
	.w8(32'hba9e9284),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f7845),
	.w1(32'hbad68664),
	.w2(32'hbb23b8a1),
	.w3(32'h387bb604),
	.w4(32'hbacd2bb0),
	.w5(32'hbb0af283),
	.w6(32'h388b9c6b),
	.w7(32'hba63d2e4),
	.w8(32'hbacd8dc6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c78e1),
	.w1(32'hb989ec5e),
	.w2(32'h3a5f6aef),
	.w3(32'h39d504fc),
	.w4(32'h392219a5),
	.w5(32'h3a6f35e4),
	.w6(32'h39ead72a),
	.w7(32'h3a9c91e8),
	.w8(32'h3b0c449c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04f5a3),
	.w1(32'hbac6e2b2),
	.w2(32'hbaa00954),
	.w3(32'hb8f1a1c6),
	.w4(32'hba66e483),
	.w5(32'hb9e82b3c),
	.w6(32'h3a11229f),
	.w7(32'hba20ac14),
	.w8(32'hb8a49675),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fd7d6),
	.w1(32'hb8250ae6),
	.w2(32'hb9f40f59),
	.w3(32'h3afd914f),
	.w4(32'h3ac39cb3),
	.w5(32'h384cfb42),
	.w6(32'h3ae95476),
	.w7(32'h3aaf1297),
	.w8(32'h3a72d95f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a818dc3),
	.w1(32'h38ae5cdc),
	.w2(32'hb9c36b01),
	.w3(32'h3a7936a1),
	.w4(32'h39ecccb1),
	.w5(32'hb7ee4a00),
	.w6(32'h3a6d4bc6),
	.w7(32'h39f4e644),
	.w8(32'h39b3a62f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9357314),
	.w1(32'hbab53f21),
	.w2(32'hbb06a01f),
	.w3(32'hb93b7486),
	.w4(32'hbaa86023),
	.w5(32'hbab7dc6b),
	.w6(32'h39240911),
	.w7(32'hba21abf8),
	.w8(32'hba440031),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8760068),
	.w1(32'hb8640a62),
	.w2(32'hb7ec5a9d),
	.w3(32'hb8665072),
	.w4(32'hb874c2bc),
	.w5(32'hb75e2787),
	.w6(32'hb8689fb3),
	.w7(32'hb851fcb3),
	.w8(32'hb7ab6a62),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376555c4),
	.w1(32'hb7570c9a),
	.w2(32'hb77aa0f5),
	.w3(32'h382825a4),
	.w4(32'h36b8a2eb),
	.w5(32'hb7a05a18),
	.w6(32'h38243f1d),
	.w7(32'hb817ae53),
	.w8(32'hb6984766),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3797b405),
	.w1(32'hb81012be),
	.w2(32'hb89f8e70),
	.w3(32'h38a0a2aa),
	.w4(32'h3913477b),
	.w5(32'h3889998f),
	.w6(32'h3801e62e),
	.w7(32'h387b77d2),
	.w8(32'h38394cc3),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7894236),
	.w1(32'h3832baec),
	.w2(32'h38f2514b),
	.w3(32'h3857e720),
	.w4(32'h388a698d),
	.w5(32'h38dc811d),
	.w6(32'h3890b063),
	.w7(32'h384b2e24),
	.w8(32'h38d73cd6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e358e),
	.w1(32'hbb06b0a6),
	.w2(32'hbb2ca430),
	.w3(32'hba034222),
	.w4(32'hbae591b2),
	.w5(32'hbaf38d0b),
	.w6(32'hb9c95b28),
	.w7(32'hbaa79c7d),
	.w8(32'hbadbe435),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97cf9c2),
	.w1(32'hb957e159),
	.w2(32'h382cac4c),
	.w3(32'hb936a2b0),
	.w4(32'hb8982a3e),
	.w5(32'h387fee4e),
	.w6(32'hb88cd2b7),
	.w7(32'hb8c07431),
	.w8(32'hb6f8404f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f379b),
	.w1(32'h39808cba),
	.w2(32'h393c78eb),
	.w3(32'h3a3d2d89),
	.w4(32'h39ac2026),
	.w5(32'h39e4824a),
	.w6(32'h3aaa1977),
	.w7(32'h3ab32d20),
	.w8(32'h3abb1749),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6c86f),
	.w1(32'hbb1eeb87),
	.w2(32'hbaf788f4),
	.w3(32'h3796011e),
	.w4(32'hbad99c13),
	.w5(32'hba930313),
	.w6(32'hba3a4b3c),
	.w7(32'hbaf97327),
	.w8(32'hba02a4d3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89397d0),
	.w1(32'hb7fa139c),
	.w2(32'h38109dcd),
	.w3(32'hb86314fb),
	.w4(32'h371b684c),
	.w5(32'h380a0132),
	.w6(32'h38207247),
	.w7(32'h38ae554f),
	.w8(32'h37f81aff),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36513d37),
	.w1(32'h38ad31f0),
	.w2(32'h38e63315),
	.w3(32'h38e98e95),
	.w4(32'h3914b347),
	.w5(32'h38fea1f2),
	.w6(32'h38abd89d),
	.w7(32'h38e93a84),
	.w8(32'h38a43981),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372fcfe2),
	.w1(32'hb5e71c67),
	.w2(32'h37bbb339),
	.w3(32'h36b0f60d),
	.w4(32'hb6cd915b),
	.w5(32'h3736f828),
	.w6(32'hb48d3b1f),
	.w7(32'hb7363541),
	.w8(32'h3727a8b5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d8bdc8),
	.w1(32'hbb8e6817),
	.w2(32'hbb025785),
	.w3(32'h3842fab3),
	.w4(32'hbb594529),
	.w5(32'hbb106ca7),
	.w6(32'hbae82fc4),
	.w7(32'h3b226552),
	.w8(32'h397e390f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00a18c),
	.w1(32'h3b177564),
	.w2(32'h3b6c0f63),
	.w3(32'hbaa50a2a),
	.w4(32'h3a79cf90),
	.w5(32'h3abda258),
	.w6(32'h3aaaa4b3),
	.w7(32'hbb64e701),
	.w8(32'hbaa245ee),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3973509b),
	.w1(32'hbb5cb094),
	.w2(32'hbd2b41a8),
	.w3(32'h3b14cb1f),
	.w4(32'h3c109729),
	.w5(32'h3c858abb),
	.w6(32'hbc476f71),
	.w7(32'hbc3351e1),
	.w8(32'hbaac6794),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc103dc0),
	.w1(32'h3b64f9fd),
	.w2(32'h3b3ed55e),
	.w3(32'hbb258552),
	.w4(32'hbaa0f84b),
	.w5(32'h3b5364f9),
	.w6(32'hba28c73b),
	.w7(32'hbc1ce622),
	.w8(32'hbb7c43a5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ffc28),
	.w1(32'h3b975695),
	.w2(32'hba7a3fbd),
	.w3(32'hbb312b5c),
	.w4(32'h39d4259b),
	.w5(32'hbb40b896),
	.w6(32'hbb00c68c),
	.w7(32'h3a713a4d),
	.w8(32'h3a51ab9e),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ad12e),
	.w1(32'hbbb9acf6),
	.w2(32'h3c43da48),
	.w3(32'hbaf8911e),
	.w4(32'hbaf835b7),
	.w5(32'hbc1139f5),
	.w6(32'hbbf2bf10),
	.w7(32'hbc39f53d),
	.w8(32'hbc183eb9),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2ecae),
	.w1(32'h39718c5e),
	.w2(32'h3c2253fd),
	.w3(32'hbb9e24fc),
	.w4(32'hbbff8c6e),
	.w5(32'h3b3f731b),
	.w6(32'h3b96bea4),
	.w7(32'hbc0c166c),
	.w8(32'hbc4f6e50),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cc9b9),
	.w1(32'h3a0d7e77),
	.w2(32'h3a25f1fd),
	.w3(32'h3c05fc27),
	.w4(32'hbacf92c8),
	.w5(32'h3bee73d9),
	.w6(32'hb90babe1),
	.w7(32'hbc53ea1e),
	.w8(32'hbbda01a5),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e07fb),
	.w1(32'h3b810966),
	.w2(32'h3a3ee9c2),
	.w3(32'h3b9cfdf1),
	.w4(32'hba6fb4a5),
	.w5(32'h3b8b48c7),
	.w6(32'h3becc3be),
	.w7(32'hbb68f9b7),
	.w8(32'h3a4dd720),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1665bf),
	.w1(32'hbb4e720c),
	.w2(32'hbb2e64bd),
	.w3(32'h3aa39523),
	.w4(32'hbb81d501),
	.w5(32'hbc02aaeb),
	.w6(32'h3a8bc160),
	.w7(32'h3b95feb4),
	.w8(32'h39c850cb),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a160652),
	.w1(32'h3b0cc614),
	.w2(32'h3b33534b),
	.w3(32'h38992e7f),
	.w4(32'hbaf823ed),
	.w5(32'h37e9dd6b),
	.w6(32'h39ebb442),
	.w7(32'hba90e8b5),
	.w8(32'h3a55b821),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b579cf0),
	.w1(32'h3af9f71e),
	.w2(32'h3b5480d3),
	.w3(32'hba45550f),
	.w4(32'hbb07588f),
	.w5(32'h3b9915d2),
	.w6(32'h3b45c37a),
	.w7(32'hbb4ea602),
	.w8(32'h3b007242),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed7afa),
	.w1(32'hbb1c895c),
	.w2(32'hba5ccbda),
	.w3(32'hb9c01e66),
	.w4(32'h3bedb5e5),
	.w5(32'h3b2b2895),
	.w6(32'hbb4676cd),
	.w7(32'hb98db425),
	.w8(32'hbab0cdd8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a316f),
	.w1(32'hbc4cefe7),
	.w2(32'hb76e7f23),
	.w3(32'h3c0d60ee),
	.w4(32'hba501cfe),
	.w5(32'h3ba341bd),
	.w6(32'h3c2a92ab),
	.w7(32'h3c853953),
	.w8(32'h3c1145b0),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28d02d),
	.w1(32'hba9da144),
	.w2(32'hba6e2dba),
	.w3(32'h3975b9b2),
	.w4(32'hbab4ff1d),
	.w5(32'h3983732b),
	.w6(32'hbb476bdf),
	.w7(32'h3b4007fd),
	.w8(32'h3b23d849),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7d117),
	.w1(32'hbc34df50),
	.w2(32'hbc0e6a10),
	.w3(32'hb98783dd),
	.w4(32'hbc6b957e),
	.w5(32'hbcf21a3a),
	.w6(32'hbada1a80),
	.w7(32'h3cbbb622),
	.w8(32'h3b9fa9a2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02d230),
	.w1(32'hbcb4e992),
	.w2(32'h3c504e26),
	.w3(32'hbbaf4b89),
	.w4(32'hbc485ced),
	.w5(32'hbca6c833),
	.w6(32'hbc2470d2),
	.w7(32'hbca5e49f),
	.w8(32'hbb6b66b2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd958f),
	.w1(32'h3b90a55b),
	.w2(32'h3bf7a7b6),
	.w3(32'hbc6fbcb1),
	.w4(32'hbafebaa5),
	.w5(32'h3a1730a3),
	.w6(32'hbaade622),
	.w7(32'hbb8455a2),
	.w8(32'hba6379d1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c1960),
	.w1(32'h3b744939),
	.w2(32'h3a4d1816),
	.w3(32'hbb35df02),
	.w4(32'h3b597f4b),
	.w5(32'hba179cb1),
	.w6(32'hbb458f3a),
	.w7(32'hbb799abd),
	.w8(32'hbaac6a05),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a7e93),
	.w1(32'h3b0c8f80),
	.w2(32'hb9e50d85),
	.w3(32'h3b45d32a),
	.w4(32'h3834b05d),
	.w5(32'h3b2c2bb2),
	.w6(32'hbb028992),
	.w7(32'hbc1d3259),
	.w8(32'hbba38958),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2172b0),
	.w1(32'h3b1ddc4e),
	.w2(32'h3a140196),
	.w3(32'h39ebda1d),
	.w4(32'h3a401dcb),
	.w5(32'h3b213515),
	.w6(32'hb9e96da4),
	.w7(32'hbb54ce06),
	.w8(32'hb917c05b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85f0a2c),
	.w1(32'hbb09b6d6),
	.w2(32'hbb541caa),
	.w3(32'h394d7995),
	.w4(32'hbb4abc98),
	.w5(32'hbabf6e8a),
	.w6(32'hbb2642fc),
	.w7(32'hbb8d2073),
	.w8(32'hbb47a1a6),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fc6ca),
	.w1(32'h3858efea),
	.w2(32'hb9aa7b78),
	.w3(32'hba783abd),
	.w4(32'hbacd085f),
	.w5(32'hba958369),
	.w6(32'h39f5f132),
	.w7(32'h3a860d3d),
	.w8(32'h393f19bb),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8ecbd),
	.w1(32'hbc1bdeda),
	.w2(32'hbcac5a35),
	.w3(32'hbaa877bf),
	.w4(32'hbbdae601),
	.w5(32'h3b4181ba),
	.w6(32'hbc47faa9),
	.w7(32'hbb2a63b4),
	.w8(32'hbc5bf1af),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf25023),
	.w1(32'h3b834511),
	.w2(32'h3a959a0c),
	.w3(32'h3aef46c5),
	.w4(32'hbb8834ce),
	.w5(32'hb960ca54),
	.w6(32'hbb2ca101),
	.w7(32'hbbed5489),
	.w8(32'hbc1c474a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b5e2a),
	.w1(32'h3a1cbdc0),
	.w2(32'h39557490),
	.w3(32'hbb6b7ec8),
	.w4(32'hbb2ef5d6),
	.w5(32'hbbb8e869),
	.w6(32'h3af061b1),
	.w7(32'h3bbbef87),
	.w8(32'h3b2af944),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4a231),
	.w1(32'h38c753ff),
	.w2(32'h3bb05ff4),
	.w3(32'hbb013644),
	.w4(32'hbba73541),
	.w5(32'h398c5b6d),
	.w6(32'h3b44f288),
	.w7(32'hbb542711),
	.w8(32'h3ae06869),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa9bfb),
	.w1(32'hbc48104d),
	.w2(32'hbc6fdcf4),
	.w3(32'hbb891946),
	.w4(32'hbb7fbe28),
	.w5(32'hbb96a9d0),
	.w6(32'hbb513d0f),
	.w7(32'hbae3809f),
	.w8(32'h3b4b489d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ef011),
	.w1(32'hbafeed2d),
	.w2(32'hbaa54736),
	.w3(32'hbbbd79f6),
	.w4(32'hbaa6557b),
	.w5(32'hb98882d4),
	.w6(32'hbb08dd48),
	.w7(32'hbb2122ae),
	.w8(32'hb9ee994a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04390f),
	.w1(32'h3b16ef6a),
	.w2(32'h3c357e1a),
	.w3(32'hbaafe9f0),
	.w4(32'hbbd2ac51),
	.w5(32'h3ade405e),
	.w6(32'h3b8bd742),
	.w7(32'hbba030a8),
	.w8(32'hbb9e58cb),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93b217),
	.w1(32'hbbc41e57),
	.w2(32'hbb42801c),
	.w3(32'hbadac992),
	.w4(32'h3a9b81d2),
	.w5(32'h3bc9d88b),
	.w6(32'hb8f9019f),
	.w7(32'h3af6529d),
	.w8(32'hb9989034),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85bf13),
	.w1(32'h3b99b581),
	.w2(32'hba9f2c2f),
	.w3(32'h3afa62e4),
	.w4(32'h3b6f9b7a),
	.w5(32'hba885fdc),
	.w6(32'h3aaba95b),
	.w7(32'hbb801999),
	.w8(32'hbabe3547),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1eeda0),
	.w1(32'h3a248b6f),
	.w2(32'hb83af5b5),
	.w3(32'h3ab1e025),
	.w4(32'hb957bd4f),
	.w5(32'h3a4581f9),
	.w6(32'h3a684b88),
	.w7(32'h3a65c939),
	.w8(32'h3a215175),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba996e73),
	.w1(32'hbb08ce91),
	.w2(32'hba26a667),
	.w3(32'hb9be36b4),
	.w4(32'hba33d068),
	.w5(32'hb9d23277),
	.w6(32'hbb77013f),
	.w7(32'hbb03861f),
	.w8(32'h3a8d77d9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf1783),
	.w1(32'h3b5fe726),
	.w2(32'h3aa784ff),
	.w3(32'h3a21731f),
	.w4(32'h3b9e8100),
	.w5(32'h3bb40217),
	.w6(32'h3b011e86),
	.w7(32'h3a43c178),
	.w8(32'hbb5642ed),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99cad9),
	.w1(32'hbbbd8f03),
	.w2(32'hbb008449),
	.w3(32'h3b648513),
	.w4(32'h3a7ef7b7),
	.w5(32'h3b89e0f0),
	.w6(32'hbbdefb27),
	.w7(32'hbb00bf51),
	.w8(32'h3b69d1f0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12964e),
	.w1(32'hba823cea),
	.w2(32'hba3ea4fd),
	.w3(32'hbafaf799),
	.w4(32'hba7282c9),
	.w5(32'h3bccb19b),
	.w6(32'hbc00be88),
	.w7(32'hbc9c1ac4),
	.w8(32'hbbdd363c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7321e1),
	.w1(32'hbb1645b8),
	.w2(32'hb9b62a77),
	.w3(32'hba8eb4c2),
	.w4(32'hbaebc299),
	.w5(32'hb9b4a2bd),
	.w6(32'h39eb3765),
	.w7(32'h38c4f811),
	.w8(32'h3ae0d9bb),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed344c),
	.w1(32'h3c07865c),
	.w2(32'h3c70de35),
	.w3(32'h3af935c5),
	.w4(32'h3b02a8e1),
	.w5(32'h3c1b807d),
	.w6(32'h3948cd25),
	.w7(32'hbc534fb8),
	.w8(32'hbbf20758),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6e50b),
	.w1(32'h3a444842),
	.w2(32'hbb52c463),
	.w3(32'hb845c1fd),
	.w4(32'hbb838ceb),
	.w5(32'hbaba2c85),
	.w6(32'h39603677),
	.w7(32'hbbc95056),
	.w8(32'hbb820276),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951dad3),
	.w1(32'h3ac9161d),
	.w2(32'h3a9344f1),
	.w3(32'hba62528d),
	.w4(32'hba312f27),
	.w5(32'hba9721db),
	.w6(32'hbaea6ee5),
	.w7(32'hbb2265a1),
	.w8(32'hba1b6f0c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6037c),
	.w1(32'h39b28f83),
	.w2(32'h3b956b0a),
	.w3(32'hba84fa64),
	.w4(32'hb91dba1f),
	.w5(32'h3b5f271f),
	.w6(32'h3b23eb37),
	.w7(32'hbb05ac35),
	.w8(32'h3acb63e3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d85ce),
	.w1(32'h3b5c7d7f),
	.w2(32'hb9747190),
	.w3(32'h3b8ba752),
	.w4(32'h3a535bba),
	.w5(32'hb9b73384),
	.w6(32'h3bffd193),
	.w7(32'h3b8a1297),
	.w8(32'h3b8b1cfa),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b0d67a),
	.w1(32'hbbcbdfa0),
	.w2(32'hbbf8e60b),
	.w3(32'hba16898a),
	.w4(32'hbac30b36),
	.w5(32'hba036137),
	.w6(32'hb994f3d3),
	.w7(32'hbb9abd72),
	.w8(32'hbb942a91),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc458c73),
	.w1(32'hbb1d8f66),
	.w2(32'hbadb4742),
	.w3(32'hba99ff71),
	.w4(32'hbb7789e5),
	.w5(32'hbb9c8c5d),
	.w6(32'hbb0d62cd),
	.w7(32'h3aa4dfe2),
	.w8(32'h3a276db1),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1203e5),
	.w1(32'h3b865f91),
	.w2(32'h3b00a17e),
	.w3(32'hb9ef711a),
	.w4(32'hbb32a637),
	.w5(32'h3ab82caf),
	.w6(32'h3b702b3f),
	.w7(32'hbb2fe2c8),
	.w8(32'h3a6122d8),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fb62f),
	.w1(32'hbc21e0b1),
	.w2(32'hbce161e0),
	.w3(32'hbab45e77),
	.w4(32'hbc3625ad),
	.w5(32'hbc7dd5c2),
	.w6(32'hbb422913),
	.w7(32'h3ca01e89),
	.w8(32'h3bb7ef13),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de2510),
	.w1(32'hbbcfa965),
	.w2(32'hbc6b0573),
	.w3(32'hbbb53603),
	.w4(32'hbbfce50f),
	.w5(32'hbb5f4b71),
	.w6(32'h3b96036a),
	.w7(32'h3c6402f0),
	.w8(32'h3b8228a9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986f07b),
	.w1(32'hbc0f356a),
	.w2(32'h3d27f400),
	.w3(32'h3b79609a),
	.w4(32'h3a9eb543),
	.w5(32'h3b8b6727),
	.w6(32'h3bc5ee2d),
	.w7(32'h3b690de0),
	.w8(32'hbabf4e32),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e00d3),
	.w1(32'hbb6e600a),
	.w2(32'hbbd019d0),
	.w3(32'h3b964f45),
	.w4(32'h3b95bccc),
	.w5(32'h3b1b1e8f),
	.w6(32'hbb262db0),
	.w7(32'hbae12422),
	.w8(32'h3a64d2eb),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0aa2b5),
	.w1(32'hbb085232),
	.w2(32'hbb0eb988),
	.w3(32'h3b49dd77),
	.w4(32'hba03f29b),
	.w5(32'hbac0c331),
	.w6(32'hbb047464),
	.w7(32'h3a4f0099),
	.w8(32'h3aaf2d86),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97bd0b6),
	.w1(32'hbabe6386),
	.w2(32'hbadc7827),
	.w3(32'h38c95b86),
	.w4(32'hbb66ae4b),
	.w5(32'hbc061c16),
	.w6(32'h3ab28d32),
	.w7(32'h3c21dda6),
	.w8(32'h3b1a6223),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b2f68),
	.w1(32'hbbcae443),
	.w2(32'h3b25c814),
	.w3(32'hbad64c30),
	.w4(32'hbbe528b1),
	.w5(32'hbc540cfa),
	.w6(32'h3aeaea7a),
	.w7(32'h3c5a420a),
	.w8(32'hba2e9e81),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdbb17),
	.w1(32'h3c5faa44),
	.w2(32'h3c87a944),
	.w3(32'hbb170c62),
	.w4(32'h3b856fd2),
	.w5(32'h3c00a38a),
	.w6(32'hba39f6fd),
	.w7(32'hbc961cba),
	.w8(32'hbb3b2929),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaa456),
	.w1(32'h3b262163),
	.w2(32'h3ba33023),
	.w3(32'hbc85445a),
	.w4(32'hbae81139),
	.w5(32'h3bbec50a),
	.w6(32'h3a8fdf9b),
	.w7(32'hbc1c9aec),
	.w8(32'h39ab49b1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa93c16),
	.w1(32'hba98f462),
	.w2(32'h3b353038),
	.w3(32'hbb8e402e),
	.w4(32'hbb4225c9),
	.w5(32'h3c2cc904),
	.w6(32'hb89752c1),
	.w7(32'hbc738404),
	.w8(32'hbc0f80f1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4deba),
	.w1(32'h3a7304c1),
	.w2(32'h3ab9bb86),
	.w3(32'h3b92bb52),
	.w4(32'hbb0d2728),
	.w5(32'h3a346796),
	.w6(32'hbb29cb30),
	.w7(32'hbbcadf17),
	.w8(32'h397bf884),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1502bf),
	.w1(32'hbb1bbb9b),
	.w2(32'hbbb93dd5),
	.w3(32'hbb265dd7),
	.w4(32'h3ab77f18),
	.w5(32'h39095f68),
	.w6(32'h3b803cfc),
	.w7(32'hbb5fe079),
	.w8(32'hbb61e5b2),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe7a6f),
	.w1(32'hbb87f758),
	.w2(32'hbbc28254),
	.w3(32'h39fc363d),
	.w4(32'hbbbbd573),
	.w5(32'hbc388572),
	.w6(32'hb98efd8f),
	.w7(32'h3c11d541),
	.w8(32'h3b2c6ad6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86ed50),
	.w1(32'hbbbbbc2b),
	.w2(32'hbc2acfa9),
	.w3(32'hbbc08748),
	.w4(32'hbb4ee7a8),
	.w5(32'hbbb0258c),
	.w6(32'hbb0c5513),
	.w7(32'hbba3d9aa),
	.w8(32'hbb9f905f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f4882),
	.w1(32'h3bbc0046),
	.w2(32'h3b940c93),
	.w3(32'hb926cd32),
	.w4(32'h38d0007e),
	.w5(32'h3b5050eb),
	.w6(32'h3ad4663e),
	.w7(32'hbbd14568),
	.w8(32'h3aa7c2a7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86bd5f),
	.w1(32'h39cc3f79),
	.w2(32'hbba243a8),
	.w3(32'hba907039),
	.w4(32'hba79e816),
	.w5(32'hbb8b5cde),
	.w6(32'hba7e979d),
	.w7(32'h38fbe6e9),
	.w8(32'hbaa158a3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca4d3d),
	.w1(32'hba801729),
	.w2(32'hba61ea6b),
	.w3(32'hba49912b),
	.w4(32'hbb477847),
	.w5(32'hba5eb3a5),
	.w6(32'h3a805bac),
	.w7(32'hbb20cecb),
	.w8(32'hb8b42339),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39847de5),
	.w1(32'hbb240183),
	.w2(32'hbc4fa563),
	.w3(32'hbaa0232f),
	.w4(32'hb934e292),
	.w5(32'hbb23a02e),
	.w6(32'hba8a9469),
	.w7(32'h3b6abeb7),
	.w8(32'hba046e2b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bb7d4),
	.w1(32'h3afdd997),
	.w2(32'h3bb160bf),
	.w3(32'hbae063ed),
	.w4(32'hbac2154f),
	.w5(32'h3c5b5d93),
	.w6(32'hbc0b0068),
	.w7(32'h3a03373e),
	.w8(32'hbc643f92),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b9c2f),
	.w1(32'h3b1d63ea),
	.w2(32'h3b1db311),
	.w3(32'h3b928b37),
	.w4(32'hbb136409),
	.w5(32'h3afcc574),
	.w6(32'h3ac16136),
	.w7(32'hbb8d2f6d),
	.w8(32'h3986ba5d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1497de),
	.w1(32'h3b2fd468),
	.w2(32'h3ac19085),
	.w3(32'hba993c37),
	.w4(32'hb940f135),
	.w5(32'h3b269d2a),
	.w6(32'hba91b62a),
	.w7(32'hbb99eb10),
	.w8(32'hbb71003f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a490c71),
	.w1(32'hbb285923),
	.w2(32'hbbdb1154),
	.w3(32'h3ac1d729),
	.w4(32'h39d5dff8),
	.w5(32'hbb6cda2a),
	.w6(32'h3ba818eb),
	.w7(32'h3b11776f),
	.w8(32'hbbe840f3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a581705),
	.w1(32'hb733d736),
	.w2(32'hbbbef137),
	.w3(32'h3a142dfd),
	.w4(32'h3b62eec5),
	.w5(32'h3b35b267),
	.w6(32'h3ac3217f),
	.w7(32'hbb734065),
	.w8(32'hbad5b308),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf796ea),
	.w1(32'hba679603),
	.w2(32'hbb522f39),
	.w3(32'hbb08f5e4),
	.w4(32'hbb24cf33),
	.w5(32'hbb9aabd0),
	.w6(32'hbb27adc7),
	.w7(32'hbb9b20da),
	.w8(32'hbb1a16b1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b0204),
	.w1(32'h3ad0ba3d),
	.w2(32'h3bc18599),
	.w3(32'hb98d1711),
	.w4(32'hbb2577e3),
	.w5(32'hbad2111f),
	.w6(32'h3a43aac7),
	.w7(32'hbb2c803b),
	.w8(32'h3abe3cd1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f1260),
	.w1(32'hbc0cc587),
	.w2(32'hbab0cd00),
	.w3(32'hbb83b07d),
	.w4(32'hbc753a55),
	.w5(32'hbc9aebf3),
	.w6(32'h3c32c285),
	.w7(32'h3cdf294e),
	.w8(32'h3b23ee0e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba00e95),
	.w1(32'h3a55b94a),
	.w2(32'hbb2db9fa),
	.w3(32'hb9833065),
	.w4(32'hbafaddd2),
	.w5(32'h3b11cbdd),
	.w6(32'hbbade462),
	.w7(32'hbc43b317),
	.w8(32'hbbad7462),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ec14c),
	.w1(32'h38a43857),
	.w2(32'h3b02c7e5),
	.w3(32'hbb32c0bf),
	.w4(32'hba5747a8),
	.w5(32'hbaf83b3f),
	.w6(32'hbae9b88c),
	.w7(32'hbaed4a8f),
	.w8(32'hbad589e1),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e0198),
	.w1(32'h3b7047ac),
	.w2(32'h3b378fd3),
	.w3(32'h3a90509b),
	.w4(32'h3a77a134),
	.w5(32'hba162a56),
	.w6(32'hba034c6f),
	.w7(32'hba9087e3),
	.w8(32'h3a4ebadd),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2c8e6),
	.w1(32'hba28d622),
	.w2(32'hb9e96137),
	.w3(32'hbab59f7a),
	.w4(32'hb997275f),
	.w5(32'h392b6056),
	.w6(32'hbb04160b),
	.w7(32'hbaa186b9),
	.w8(32'h3b1265c9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db533b),
	.w1(32'h3bc57b3e),
	.w2(32'h3c241a9f),
	.w3(32'h3ac084b8),
	.w4(32'h3ae07545),
	.w5(32'h3bb44acc),
	.w6(32'h3b2dd183),
	.w7(32'hbb4707aa),
	.w8(32'h3bc7b46d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec5593),
	.w1(32'hbcedd107),
	.w2(32'hbb7a60b5),
	.w3(32'h3b8d0efc),
	.w4(32'hbc4ddc6f),
	.w5(32'hbc7f6f83),
	.w6(32'h3a035c0f),
	.w7(32'hbbb4a4ff),
	.w8(32'hbc80be0b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfc66d8),
	.w1(32'hbae96863),
	.w2(32'hbbafc2a8),
	.w3(32'hbc0bb976),
	.w4(32'hbb3d1f04),
	.w5(32'hbc039a1e),
	.w6(32'h3b27c6f7),
	.w7(32'h3c2811af),
	.w8(32'h3a271a90),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03f0d9),
	.w1(32'h3b0210a3),
	.w2(32'h3a5addf9),
	.w3(32'h3a76983f),
	.w4(32'h3a1e03f6),
	.w5(32'h3af047b5),
	.w6(32'hbb1f2752),
	.w7(32'hb97e244d),
	.w8(32'hbb905d23),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac00b17),
	.w1(32'hb9e7ffb1),
	.w2(32'h3ac9f9e9),
	.w3(32'h3a18c7e1),
	.w4(32'hbb96a7ab),
	.w5(32'hbbe8ff2e),
	.w6(32'hbb59158d),
	.w7(32'hbb339a6c),
	.w8(32'hba7edae4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0cc31),
	.w1(32'h3a0231ab),
	.w2(32'hb9413e18),
	.w3(32'hbbc85d7e),
	.w4(32'hb9c4e3a4),
	.w5(32'hba94eddb),
	.w6(32'h3a921c88),
	.w7(32'h3ac3c4c2),
	.w8(32'hba28fa9d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdf15d),
	.w1(32'hbb878895),
	.w2(32'hbbc58cc2),
	.w3(32'hbafd49e3),
	.w4(32'hbaa79fb8),
	.w5(32'hba806d84),
	.w6(32'hba56bb19),
	.w7(32'hbbd1d9ae),
	.w8(32'hbb94ab9d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebde15),
	.w1(32'h3b76a9b2),
	.w2(32'h3c112b71),
	.w3(32'h3aa343ea),
	.w4(32'hbb83cd18),
	.w5(32'h3bef7829),
	.w6(32'h3b606618),
	.w7(32'hba9a09c6),
	.w8(32'h3b536c81),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebce5e),
	.w1(32'hbb307356),
	.w2(32'hbbc32dc5),
	.w3(32'h3b3533a9),
	.w4(32'hbabf1daa),
	.w5(32'hbaea28c3),
	.w6(32'h3b0cf2fb),
	.w7(32'hbb894ff0),
	.w8(32'hba5b43f6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d9d8d),
	.w1(32'h3b71c692),
	.w2(32'hbb05eb44),
	.w3(32'hbb6156da),
	.w4(32'h3a62bf08),
	.w5(32'h3bbd407c),
	.w6(32'h3aab708b),
	.w7(32'hbb2476f5),
	.w8(32'h3b853fa9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd44554),
	.w1(32'h3bd2bc87),
	.w2(32'h3a897f4f),
	.w3(32'h3b2553ad),
	.w4(32'h3bea4331),
	.w5(32'h3b9642e7),
	.w6(32'h3b5ff844),
	.w7(32'h3b6f3f64),
	.w8(32'h3b9e6e47),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba95b32),
	.w1(32'h3ac9a6aa),
	.w2(32'hb93b8fbf),
	.w3(32'h3bfbfad9),
	.w4(32'h3a3bfac4),
	.w5(32'hb913bd85),
	.w6(32'h3b3dff68),
	.w7(32'hb9853090),
	.w8(32'hbb1cb87c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23a52a),
	.w1(32'hbc3bc7af),
	.w2(32'hbbcb00b5),
	.w3(32'h39be7b62),
	.w4(32'hbc269e94),
	.w5(32'hbc0bb46c),
	.w6(32'hbbe3d94b),
	.w7(32'h3b95e924),
	.w8(32'hbb4b6844),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3826b),
	.w1(32'hb92d93a2),
	.w2(32'hb90b578b),
	.w3(32'hbbc751cc),
	.w4(32'hba80993e),
	.w5(32'hb6de2330),
	.w6(32'hb8b61474),
	.w7(32'hb6e4c1f2),
	.w8(32'h38afeb18),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf9c1c),
	.w1(32'h3ada96bf),
	.w2(32'h3a429b71),
	.w3(32'hba1008bb),
	.w4(32'hba6df7f7),
	.w5(32'h3a4745eb),
	.w6(32'hbb811517),
	.w7(32'hbc1fc855),
	.w8(32'hbb2fab79),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95207b),
	.w1(32'hba461256),
	.w2(32'h3aae1704),
	.w3(32'hba62f35c),
	.w4(32'hbab1e2d3),
	.w5(32'hb9350fa9),
	.w6(32'h394c28b7),
	.w7(32'h3a8fd114),
	.w8(32'h3ac5aaeb),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8fd19),
	.w1(32'h3a44aaaf),
	.w2(32'hbab80676),
	.w3(32'hbad43464),
	.w4(32'h3a0c8a15),
	.w5(32'h3b0a42fd),
	.w6(32'hba471b03),
	.w7(32'hb993871e),
	.w8(32'h3aa34de8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b134b50),
	.w1(32'h3b451a75),
	.w2(32'h38ff7392),
	.w3(32'h3b957616),
	.w4(32'hbaa437b8),
	.w5(32'hb8564700),
	.w6(32'h3bcea845),
	.w7(32'h3ba3b767),
	.w8(32'h3ac9f048),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a97e3),
	.w1(32'h3bd20983),
	.w2(32'h3b1309ea),
	.w3(32'h3a6286a5),
	.w4(32'h3bce8f25),
	.w5(32'h3c8f6b42),
	.w6(32'hbbbfb06e),
	.w7(32'hbc800653),
	.w8(32'hbba20e8e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d240c),
	.w1(32'hbb86bf9f),
	.w2(32'hbbc6abb0),
	.w3(32'h3a6b337f),
	.w4(32'hbaa69906),
	.w5(32'hba4c4041),
	.w6(32'hba9c9b64),
	.w7(32'hbbb6c2e6),
	.w8(32'hbb1e74e4),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b14ff),
	.w1(32'hb9c86066),
	.w2(32'hbb76ad0f),
	.w3(32'hb979ea68),
	.w4(32'h37566a13),
	.w5(32'h38f9e3f0),
	.w6(32'hbb6b9d1e),
	.w7(32'hbb601174),
	.w8(32'hbb27f1fe),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a5f8f),
	.w1(32'hbb5a8954),
	.w2(32'hbc825c6d),
	.w3(32'hba3459a1),
	.w4(32'hba815b32),
	.w5(32'h3cd71c82),
	.w6(32'hbbdab2c5),
	.w7(32'hbbdf7413),
	.w8(32'hbc1cccc7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ee6e3),
	.w1(32'hb8c37578),
	.w2(32'h3b29300e),
	.w3(32'h3b9bdea3),
	.w4(32'hbb76047b),
	.w5(32'h3a8df400),
	.w6(32'hba59bc27),
	.w7(32'hba226071),
	.w8(32'hbbc64c59),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbef795),
	.w1(32'h3b99aac9),
	.w2(32'hbb57178f),
	.w3(32'hbbb15819),
	.w4(32'h3b41a7c9),
	.w5(32'h3c5c5f6f),
	.w6(32'hbba58e0e),
	.w7(32'hbc729f2a),
	.w8(32'hbbdb6032),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb015f63),
	.w1(32'h3ab3a12b),
	.w2(32'h3b8e042e),
	.w3(32'h3a183060),
	.w4(32'hba7b0dcd),
	.w5(32'h3bfdd8fe),
	.w6(32'hba8188d0),
	.w7(32'hbbd559e9),
	.w8(32'hbb58adf2),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34ac3b),
	.w1(32'h3bfa6d1b),
	.w2(32'h3c3df0d8),
	.w3(32'h3b8b2c86),
	.w4(32'h3b9f284d),
	.w5(32'h3c77fd5b),
	.w6(32'hb9173969),
	.w7(32'hbc53cbe7),
	.w8(32'hba86b7bd),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaada004),
	.w1(32'hbc12caa2),
	.w2(32'hbc85a491),
	.w3(32'hbaa5217b),
	.w4(32'hbb8f6e58),
	.w5(32'hbc98bd66),
	.w6(32'hba71d745),
	.w7(32'hbc0d26cc),
	.w8(32'hbbc93746),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b20b4),
	.w1(32'hbb3921e9),
	.w2(32'hbc82eb4c),
	.w3(32'hbb6a62f1),
	.w4(32'hbad6fee9),
	.w5(32'h3c475738),
	.w6(32'h3b4509bd),
	.w7(32'hbb8c4342),
	.w8(32'hbc1203ff),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19051d),
	.w1(32'h39a581dc),
	.w2(32'hbb875609),
	.w3(32'h3be13c29),
	.w4(32'hba9b31f9),
	.w5(32'hbc124e51),
	.w6(32'h3bfa959b),
	.w7(32'h3ca3ea1e),
	.w8(32'h3bbea4ee),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa79b85),
	.w1(32'hbb054f83),
	.w2(32'h3b2a8522),
	.w3(32'h3afb2e35),
	.w4(32'hbb0a63a5),
	.w5(32'hbb12f2c7),
	.w6(32'hbad0bd34),
	.w7(32'hbb1d289d),
	.w8(32'hba8a07c0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39858ef7),
	.w1(32'h3977bc86),
	.w2(32'hbad36a02),
	.w3(32'h3a1c6b90),
	.w4(32'hba801f39),
	.w5(32'hbb87514d),
	.w6(32'h3a9e3345),
	.w7(32'h3be10ae9),
	.w8(32'h3a3ffe8b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3b5f6),
	.w1(32'h398e41ec),
	.w2(32'hb99db39f),
	.w3(32'h3ae296d7),
	.w4(32'hbaa12fd5),
	.w5(32'h399e9be7),
	.w6(32'h3a7a5daa),
	.w7(32'h3abd1435),
	.w8(32'h3a25f319),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f773d),
	.w1(32'h3bb8638a),
	.w2(32'h3aa7b3a5),
	.w3(32'hbae2431b),
	.w4(32'h398ffbd7),
	.w5(32'h39d3e669),
	.w6(32'hbb1606f2),
	.w7(32'hbb101b7e),
	.w8(32'hbb9d34d8),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b633a),
	.w1(32'h3a443493),
	.w2(32'hba195356),
	.w3(32'h3a34d57b),
	.w4(32'hba649df8),
	.w5(32'h3a1e1627),
	.w6(32'hba2f25ed),
	.w7(32'hba3e6de7),
	.w8(32'hba95bfd2),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3f860),
	.w1(32'hba04dcd1),
	.w2(32'hbb501997),
	.w3(32'h39d47c07),
	.w4(32'hbab23cb7),
	.w5(32'hbbb4038f),
	.w6(32'h3b04b119),
	.w7(32'h3c184c27),
	.w8(32'h3a96bd85),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988e5a7),
	.w1(32'h39dd8bc7),
	.w2(32'hbbbc3d5a),
	.w3(32'h3a4bfd66),
	.w4(32'hbb5dc5a6),
	.w5(32'hbc2eee01),
	.w6(32'h3a7aa866),
	.w7(32'h3c40b0d6),
	.w8(32'h3b0e5996),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b605711),
	.w1(32'h3b48c2ba),
	.w2(32'h3b82faf4),
	.w3(32'hba3fbae1),
	.w4(32'hba02e109),
	.w5(32'hba3e3be0),
	.w6(32'hba100406),
	.w7(32'hbb462720),
	.w8(32'h3b10335e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7e364),
	.w1(32'h3acfe5a6),
	.w2(32'hbc857742),
	.w3(32'hbb214ae8),
	.w4(32'hbb2594a4),
	.w5(32'hbc1d69fb),
	.w6(32'hbc34edc6),
	.w7(32'h3ab90670),
	.w8(32'hbc47ee45),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc138dc),
	.w1(32'h3b54c649),
	.w2(32'h3c1fa5a9),
	.w3(32'hbc7b2a10),
	.w4(32'hba456742),
	.w5(32'hba86920f),
	.w6(32'h3af0e8ff),
	.w7(32'hbbb0662c),
	.w8(32'h3ae91c3c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ecca1),
	.w1(32'hbbd09ce3),
	.w2(32'hbc444035),
	.w3(32'hbb349765),
	.w4(32'hbb2be04c),
	.w5(32'hbc00c2de),
	.w6(32'hb9d9075f),
	.w7(32'hb9c0816c),
	.w8(32'hbb01152c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc045089),
	.w1(32'hbc064edb),
	.w2(32'hbb954615),
	.w3(32'hbb0dec18),
	.w4(32'hbc2beb83),
	.w5(32'hbc7224d9),
	.w6(32'hbba631f4),
	.w7(32'h3bfa6385),
	.w8(32'hbbbb2736),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdab324),
	.w1(32'hb98299cd),
	.w2(32'hbb6148cb),
	.w3(32'hbbd1f0ac),
	.w4(32'hbae7815f),
	.w5(32'hbbee2f3c),
	.w6(32'h3b27cd96),
	.w7(32'h3c47ae1e),
	.w8(32'h3ac36b07),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a210483),
	.w1(32'h3a74b5d6),
	.w2(32'hba50a7db),
	.w3(32'h3a7a06e4),
	.w4(32'hba00dfe7),
	.w5(32'hbac38380),
	.w6(32'h3a1f71fa),
	.w7(32'h3ac9cda9),
	.w8(32'hba834cdc),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6218fc),
	.w1(32'h3b097c97),
	.w2(32'hba2e5951),
	.w3(32'h3b0f9389),
	.w4(32'h3a81998a),
	.w5(32'h3a3edc20),
	.w6(32'h39c29161),
	.w7(32'hba226f02),
	.w8(32'hbb16c2bf),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45e728),
	.w1(32'hbc4238d5),
	.w2(32'hbcac9ddd),
	.w3(32'h3b5e3f5e),
	.w4(32'hbc4ee969),
	.w5(32'hbc51be85),
	.w6(32'hbc1a79df),
	.w7(32'hba055c8f),
	.w8(32'hbb80014f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf57238),
	.w1(32'h3b028134),
	.w2(32'hbbc2a8e6),
	.w3(32'hbbd8e30a),
	.w4(32'hba4aea46),
	.w5(32'hbb99e6e8),
	.w6(32'h3b349b18),
	.w7(32'h3a2b9dcc),
	.w8(32'hbab16d44),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39851e18),
	.w1(32'hbbab89b4),
	.w2(32'hbb16a293),
	.w3(32'hba9074ec),
	.w4(32'hbb2c22ac),
	.w5(32'h3a191c91),
	.w6(32'hbb85aa50),
	.w7(32'hbbe9a2e0),
	.w8(32'hbaf1dcd9),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80922b0),
	.w1(32'h3b9bcdf7),
	.w2(32'h3acd9b9b),
	.w3(32'h3af4ca7d),
	.w4(32'h3b078434),
	.w5(32'h3c1425fc),
	.w6(32'hbbb2052f),
	.w7(32'hbc184edd),
	.w8(32'hbb95b12b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7c056),
	.w1(32'hb81971cd),
	.w2(32'hbb16bed7),
	.w3(32'h3a55c3fe),
	.w4(32'hbae2ca13),
	.w5(32'hbb8289a3),
	.w6(32'hba82e5c4),
	.w7(32'h3b59a9b7),
	.w8(32'h3a0d1eb3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa79322),
	.w1(32'hbce9c1b4),
	.w2(32'hbd0e9fc7),
	.w3(32'hbac0003d),
	.w4(32'hbc71fa57),
	.w5(32'hbba1c5af),
	.w6(32'hbc108b14),
	.w7(32'hbc4022a3),
	.w8(32'hbc81a698),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83f407),
	.w1(32'h3aa79bff),
	.w2(32'h3ba7f2b1),
	.w3(32'hba2a391e),
	.w4(32'hba8e25ae),
	.w5(32'h3c917f09),
	.w6(32'hbb726d42),
	.w7(32'hbc837b9d),
	.w8(32'hbbd4de4c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0167c4),
	.w1(32'h3b0bdfab),
	.w2(32'h3ac307a9),
	.w3(32'h3bb658fc),
	.w4(32'h3aca53f0),
	.w5(32'h3b82dc9b),
	.w6(32'h3b6f483f),
	.w7(32'h3ae9dce9),
	.w8(32'h3b14a428),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4eaca8),
	.w1(32'h3741239e),
	.w2(32'h38191d88),
	.w3(32'h3a3f3fec),
	.w4(32'h37ac3637),
	.w5(32'h378ed11e),
	.w6(32'h37011bcc),
	.w7(32'h3818b1e4),
	.w8(32'h380128de),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c9c00),
	.w1(32'hba13f067),
	.w2(32'hba928999),
	.w3(32'h3a8669dd),
	.w4(32'h3a1927f8),
	.w5(32'h3783d9d9),
	.w6(32'h3b3ead04),
	.w7(32'h3b42fba1),
	.w8(32'h3b376698),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule