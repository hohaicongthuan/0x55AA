module layer_8_featuremap_90(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81b950),
	.w1(32'h3c55afc0),
	.w2(32'h3d0e268a),
	.w3(32'h3caf3685),
	.w4(32'hbcdf627a),
	.w5(32'hbb98cb9e),
	.w6(32'h3c861183),
	.w7(32'hbc4ce00c),
	.w8(32'hbc17019d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbbb540),
	.w1(32'hbc43cbe3),
	.w2(32'hbc4a5e7e),
	.w3(32'h3b9cde75),
	.w4(32'hbba042ec),
	.w5(32'h3cb43491),
	.w6(32'hbcf25950),
	.w7(32'h3acc7831),
	.w8(32'h3d16f48a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e5f70),
	.w1(32'hbbd72924),
	.w2(32'h3a9b8e32),
	.w3(32'hbc1c80e6),
	.w4(32'h3ba670c5),
	.w5(32'h3c2c620b),
	.w6(32'h3c1b4c05),
	.w7(32'h3c4aafc2),
	.w8(32'hbbeeb987),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ca37e),
	.w1(32'h3b9cadcb),
	.w2(32'hb97a66b2),
	.w3(32'h3c5e7b1d),
	.w4(32'hbca22ab9),
	.w5(32'hbc87508f),
	.w6(32'hbcb113d5),
	.w7(32'h3c899e55),
	.w8(32'h3c25040e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fe401),
	.w1(32'hbcbcd124),
	.w2(32'h3d710381),
	.w3(32'hbcdb6d07),
	.w4(32'hba61723c),
	.w5(32'h3c0cf108),
	.w6(32'hbc3edf40),
	.w7(32'hbba8b1b3),
	.w8(32'h3bcf136d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be21847),
	.w1(32'h3c1f4935),
	.w2(32'h3c57a475),
	.w3(32'hbd6a395b),
	.w4(32'hbc24a5ba),
	.w5(32'h3c02a16f),
	.w6(32'hbc61e502),
	.w7(32'h3b478423),
	.w8(32'h3c4b1224),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc678106),
	.w1(32'h396f11ce),
	.w2(32'h3caa5e9f),
	.w3(32'h3bca6006),
	.w4(32'hbc02af7e),
	.w5(32'hbcc83614),
	.w6(32'hbc0a7403),
	.w7(32'h3d5ee0ab),
	.w8(32'h3cbf81ad),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc720c11),
	.w1(32'h3d026c0f),
	.w2(32'hbb74fa37),
	.w3(32'hbcb8d6b3),
	.w4(32'h3bb53d54),
	.w5(32'hbc1fbd62),
	.w6(32'hbd07210f),
	.w7(32'hbcb83cf6),
	.w8(32'h3bd3ef7a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb935aa),
	.w1(32'h3c236f13),
	.w2(32'hbc1f6860),
	.w3(32'hbab44f02),
	.w4(32'h3b6ccdf1),
	.w5(32'h3b62544a),
	.w6(32'hbc36d198),
	.w7(32'h3c422a51),
	.w8(32'h3d00f9b5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd26f31f),
	.w1(32'h3c8336e8),
	.w2(32'hbdbcb379),
	.w3(32'hbd3445a7),
	.w4(32'hbc887d77),
	.w5(32'hbb847a9b),
	.w6(32'hbcd56042),
	.w7(32'hbcf47bdf),
	.w8(32'hbb93b864),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac65c0),
	.w1(32'hbcccd531),
	.w2(32'hbb5ef618),
	.w3(32'hbc34b3f7),
	.w4(32'h3c507383),
	.w5(32'h3ac4546a),
	.w6(32'h3ae51ec8),
	.w7(32'hbc8af38e),
	.w8(32'h3b788be5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7dff7),
	.w1(32'hbc8176e8),
	.w2(32'h3ca2c87a),
	.w3(32'h3bd9d299),
	.w4(32'hbbc5e717),
	.w5(32'hbcc1dfe0),
	.w6(32'hbcc30eec),
	.w7(32'hbd5b85b6),
	.w8(32'hbcaade18),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfccf5c),
	.w1(32'hbb7a8841),
	.w2(32'hbbd99231),
	.w3(32'h3babe84f),
	.w4(32'h3b90c347),
	.w5(32'hbb97460a),
	.w6(32'hbd63b81d),
	.w7(32'hbbfe7cb1),
	.w8(32'hb9d32049),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0317e5),
	.w1(32'h3b248ab5),
	.w2(32'h3c3c808a),
	.w3(32'h3b7ec389),
	.w4(32'hbb98d3a8),
	.w5(32'h3b2f0f1e),
	.w6(32'h3bceb6a1),
	.w7(32'hbb61ac4b),
	.w8(32'h3c1a469a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd31bb),
	.w1(32'h3b2ff0eb),
	.w2(32'hbc4863d6),
	.w3(32'h3bb1f54f),
	.w4(32'h3acb6a1b),
	.w5(32'hbb594974),
	.w6(32'h3b179850),
	.w7(32'h3b1890a0),
	.w8(32'h3bf24735),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h358dae96),
	.w1(32'hba162ad0),
	.w2(32'h3c794d7d),
	.w3(32'hbb626c6b),
	.w4(32'h3b911ed4),
	.w5(32'hbbafbef2),
	.w6(32'h3b3e5f88),
	.w7(32'h3b73981c),
	.w8(32'h3cedb7e4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b243fd5),
	.w1(32'hbaa05efe),
	.w2(32'hb9f89e38),
	.w3(32'h3b9a8a29),
	.w4(32'hbb3a57ab),
	.w5(32'hbb09ccc3),
	.w6(32'h3b90facd),
	.w7(32'hbbb2ff4b),
	.w8(32'hbb84c6e6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cf805),
	.w1(32'hbb0b3638),
	.w2(32'hbc0013b3),
	.w3(32'hbbee889d),
	.w4(32'hbc533397),
	.w5(32'hbb9b5994),
	.w6(32'hbc235fe0),
	.w7(32'hbb3792a7),
	.w8(32'hbbd4bfa9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cf934),
	.w1(32'h3bed1157),
	.w2(32'h3c9ba9eb),
	.w3(32'hbc86a48c),
	.w4(32'hbc149fb3),
	.w5(32'hbc24f473),
	.w6(32'hbb10afc3),
	.w7(32'hbc7d2f0e),
	.w8(32'hbc248bcd),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc588e05),
	.w1(32'hbb38c935),
	.w2(32'h3c6cca04),
	.w3(32'hbbcd08a5),
	.w4(32'h3b02fb3d),
	.w5(32'hbbd400d6),
	.w6(32'hbc9587f8),
	.w7(32'h3bce6651),
	.w8(32'hbc6855e9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d307d),
	.w1(32'h3c5c946c),
	.w2(32'hbc26a5e8),
	.w3(32'hbbd18013),
	.w4(32'hbb92a26c),
	.w5(32'h3bacf2b5),
	.w6(32'h3abec678),
	.w7(32'h3c2a189e),
	.w8(32'hba7d7e11),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80e96f),
	.w1(32'h3bbb8842),
	.w2(32'hbaca2c86),
	.w3(32'h3be3c795),
	.w4(32'h3bccc675),
	.w5(32'h3c2260cb),
	.w6(32'hbb999c6f),
	.w7(32'h3c163b56),
	.w8(32'h3b148267),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c379f44),
	.w1(32'hbb98080c),
	.w2(32'h3c81efde),
	.w3(32'hbb4e41ea),
	.w4(32'hbb77a38b),
	.w5(32'h3b4ab7c7),
	.w6(32'hbc285a82),
	.w7(32'hbaa811a4),
	.w8(32'hbc6e74f4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5138cd),
	.w1(32'h3b059045),
	.w2(32'h3b1af7cd),
	.w3(32'h3bb50d3b),
	.w4(32'hbc43a696),
	.w5(32'h3bdee26c),
	.w6(32'hbb9d3e57),
	.w7(32'hba51ee53),
	.w8(32'hbbdfc6e5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e5b1b),
	.w1(32'hbc08958e),
	.w2(32'hba63272a),
	.w3(32'h3c5564b2),
	.w4(32'hbb881048),
	.w5(32'hbb60dd86),
	.w6(32'hbaaaebc0),
	.w7(32'h3bee400c),
	.w8(32'hbb1f601b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe04faf),
	.w1(32'hbb6d3914),
	.w2(32'h39bcac7d),
	.w3(32'hbb7f762a),
	.w4(32'hbb44645b),
	.w5(32'h3b03b5b9),
	.w6(32'hbb65f693),
	.w7(32'hbcebaa19),
	.w8(32'hbb921710),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06297f),
	.w1(32'hbad7ceab),
	.w2(32'h3aec6ca0),
	.w3(32'hba70d78f),
	.w4(32'h3bda25d7),
	.w5(32'h3bcb18ef),
	.w6(32'hbb0887df),
	.w7(32'hbb500633),
	.w8(32'hbbe89e5e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd066583),
	.w1(32'h3ca1fd17),
	.w2(32'h3d545abf),
	.w3(32'hbc1dba06),
	.w4(32'h3d502979),
	.w5(32'h3d05d981),
	.w6(32'hbd5d3ee6),
	.w7(32'h3c926ace),
	.w8(32'hbd33da42),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c232da9),
	.w1(32'h3d79bc5c),
	.w2(32'hbc7e63b9),
	.w3(32'hbca3103b),
	.w4(32'h3b8f16a1),
	.w5(32'h3baf73af),
	.w6(32'hbbcf25dd),
	.w7(32'hbd0fbaca),
	.w8(32'hbb40b327),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d8ba4),
	.w1(32'hbd87ab72),
	.w2(32'h3d0c966a),
	.w3(32'hbc4393ec),
	.w4(32'hbb2a52c0),
	.w5(32'hbb4898c4),
	.w6(32'hbc8b5f92),
	.w7(32'h3ce5d8ae),
	.w8(32'hbc6e8385),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb50370),
	.w1(32'h3c9211c4),
	.w2(32'hbcaab9fe),
	.w3(32'h3c3d34b8),
	.w4(32'hbc80134e),
	.w5(32'h3ac330f7),
	.w6(32'hbaf1a9d3),
	.w7(32'hba9af8d2),
	.w8(32'hbb946763),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9d014),
	.w1(32'hbc298421),
	.w2(32'h3a4deee2),
	.w3(32'hbbac8abd),
	.w4(32'h3b3d6ed5),
	.w5(32'h3cbe80f8),
	.w6(32'hbc88e6e7),
	.w7(32'h3c9879c8),
	.w8(32'h3b30a060),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada8233),
	.w1(32'h3a6e3cac),
	.w2(32'hbc049c22),
	.w3(32'hbcad34cd),
	.w4(32'h3c828a56),
	.w5(32'hbc6c5579),
	.w6(32'hbca98b42),
	.w7(32'hbbd46977),
	.w8(32'hbc823439),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f3edd),
	.w1(32'hbc48ade1),
	.w2(32'h3ba9bb9a),
	.w3(32'hbc95f8c8),
	.w4(32'h3b8bed2e),
	.w5(32'h3cbaf7bb),
	.w6(32'h3c207aa1),
	.w7(32'h3d23f43e),
	.w8(32'hbc24c4ad),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0bd37),
	.w1(32'hbd28dc83),
	.w2(32'hbb4eae81),
	.w3(32'hbc49d1f5),
	.w4(32'h3d28ea28),
	.w5(32'hba717125),
	.w6(32'h3c408a8d),
	.w7(32'hbb15943d),
	.w8(32'hbccfa4a0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd432b58),
	.w1(32'hbc48638f),
	.w2(32'hbc545b70),
	.w3(32'hb8896edc),
	.w4(32'hbc487bc3),
	.w5(32'hbd599de7),
	.w6(32'hbca958ef),
	.w7(32'h3bbeabd4),
	.w8(32'h3d2732cc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9a2fd),
	.w1(32'h3c369917),
	.w2(32'h3b807648),
	.w3(32'hbb33765a),
	.w4(32'h3ba568d7),
	.w5(32'hbd14fcc0),
	.w6(32'hbcc39f63),
	.w7(32'hbc0772ad),
	.w8(32'h3c89b052),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c814bd9),
	.w1(32'hbbf3c1d3),
	.w2(32'hbbe005c6),
	.w3(32'hbc0f212c),
	.w4(32'hbbf975be),
	.w5(32'hbca0efe2),
	.w6(32'hba623a47),
	.w7(32'hbcbd49ea),
	.w8(32'hbd0f7efb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9cafab),
	.w1(32'hbc88e359),
	.w2(32'h3bcc7d01),
	.w3(32'h3d5a0415),
	.w4(32'hbcc9ca6d),
	.w5(32'h3c90b0e6),
	.w6(32'h3c35195d),
	.w7(32'hbb12b015),
	.w8(32'h3c8a8b50),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07306b),
	.w1(32'h3c17c326),
	.w2(32'h3a9a9c14),
	.w3(32'hbc1d2ae8),
	.w4(32'h396dccf6),
	.w5(32'h3bcf37a9),
	.w6(32'h3b600e6d),
	.w7(32'h3bd218bd),
	.w8(32'h3bf26497),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2e24c7),
	.w1(32'hbd263d38),
	.w2(32'h3c80db87),
	.w3(32'hbd43211a),
	.w4(32'hbba2a4aa),
	.w5(32'hbd1aca5f),
	.w6(32'hbd42586b),
	.w7(32'hbc421c4c),
	.w8(32'hbccd21b3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd58c34),
	.w1(32'hbb63de30),
	.w2(32'hbcb8293d),
	.w3(32'hbcf72c34),
	.w4(32'h3c3ef29c),
	.w5(32'h39d70ffb),
	.w6(32'hbbd81fc3),
	.w7(32'h3b269745),
	.w8(32'h3c763162),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b221e),
	.w1(32'h3c0c2612),
	.w2(32'h3c03a13b),
	.w3(32'hbc1cdb29),
	.w4(32'h3cf2ab99),
	.w5(32'hbbd9094f),
	.w6(32'h3d1b8b79),
	.w7(32'h3c8a04a2),
	.w8(32'h3bd58fb0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75dde0),
	.w1(32'h3bc8681a),
	.w2(32'h3c410bae),
	.w3(32'hbd5652ce),
	.w4(32'h3bdbec56),
	.w5(32'hba77fb73),
	.w6(32'hbbe5779a),
	.w7(32'hbc856aea),
	.w8(32'h3c37686a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b961183),
	.w1(32'h3d317590),
	.w2(32'hbc77ed7f),
	.w3(32'hbc6cb89e),
	.w4(32'h3c864c8c),
	.w5(32'h3b37da34),
	.w6(32'hbc8eb382),
	.w7(32'h3d3df3f6),
	.w8(32'hbc2f33ed),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7458e9),
	.w1(32'h3bfac3f4),
	.w2(32'hbb4bb6b7),
	.w3(32'hbc7fdd98),
	.w4(32'hba8d4336),
	.w5(32'h3c89597a),
	.w6(32'hbbfc0b4e),
	.w7(32'hbcff0111),
	.w8(32'hbbb40dde),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce98aba),
	.w1(32'hbc490b14),
	.w2(32'hbb75e26e),
	.w3(32'hbc68a6d5),
	.w4(32'h3c49bdcd),
	.w5(32'h3ac6e3ba),
	.w6(32'h3c58c1f0),
	.w7(32'hbcaf8f1a),
	.w8(32'hbc2dd96a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdccb47),
	.w1(32'h3bfab380),
	.w2(32'h3c3d1cdf),
	.w3(32'hbcdee2d0),
	.w4(32'hbc063d08),
	.w5(32'h3c607876),
	.w6(32'h3c01cd8a),
	.w7(32'hbc564bd3),
	.w8(32'hbc323540),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eb757),
	.w1(32'hbb70fd85),
	.w2(32'h3c5fceb7),
	.w3(32'hbc247613),
	.w4(32'h3c7c26f7),
	.w5(32'h3c977700),
	.w6(32'hba7e1d1a),
	.w7(32'h3b5003bd),
	.w8(32'hbb31c202),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5471c3),
	.w1(32'hbca0212c),
	.w2(32'h3b18fb77),
	.w3(32'h3a41d4e6),
	.w4(32'hbbc1785d),
	.w5(32'hbc6afa82),
	.w6(32'hbc74ee8c),
	.w7(32'h3cbbab81),
	.w8(32'hbb5c6b78),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba389ef3),
	.w1(32'hbc206285),
	.w2(32'hbbfe6a1e),
	.w3(32'h3b345839),
	.w4(32'hbb86a370),
	.w5(32'h3c13e6f8),
	.w6(32'hbd873a3c),
	.w7(32'h3b826984),
	.w8(32'h396391fa),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc662e8),
	.w1(32'hbc5cae90),
	.w2(32'hbc33ddc7),
	.w3(32'hbcdf905b),
	.w4(32'h3c6995af),
	.w5(32'h3c9e405a),
	.w6(32'hbcbfd90a),
	.w7(32'hbbe66740),
	.w8(32'hbc3e1c89),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68501f),
	.w1(32'hbd4961ab),
	.w2(32'hbcad4ada),
	.w3(32'h3d264bd5),
	.w4(32'hbc0e0422),
	.w5(32'hbb949707),
	.w6(32'h3c578c3f),
	.w7(32'h3c53b7fb),
	.w8(32'hbc8cd021),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3010f6),
	.w1(32'hbba9eddb),
	.w2(32'hbc3d35cd),
	.w3(32'h3b8beb05),
	.w4(32'h3c300e90),
	.w5(32'hbbf8aacd),
	.w6(32'hbc22e7e3),
	.w7(32'h3bdfec6e),
	.w8(32'hbc3a3ba9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b3449),
	.w1(32'hbc27a46c),
	.w2(32'h3c3f1c31),
	.w3(32'h3c1a1ea3),
	.w4(32'h3b13293d),
	.w5(32'h3c6c32d7),
	.w6(32'hb8757640),
	.w7(32'h3c881f30),
	.w8(32'hbb613053),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddf328),
	.w1(32'hb9a69365),
	.w2(32'hbc859f9e),
	.w3(32'hbaffca11),
	.w4(32'hbbfef2b6),
	.w5(32'hbc54fea3),
	.w6(32'hbc4b7cc6),
	.w7(32'hbc02d747),
	.w8(32'hbc500b33),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ef769),
	.w1(32'hbc4d0dab),
	.w2(32'hbb33cecf),
	.w3(32'h3b24b26b),
	.w4(32'h3bda8571),
	.w5(32'hbbd323a5),
	.w6(32'hbc355a57),
	.w7(32'hbb6501cd),
	.w8(32'hba830b9f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc034cf8),
	.w1(32'hbbd4da1f),
	.w2(32'h3bb5a43f),
	.w3(32'hbc85cd12),
	.w4(32'hbb01057d),
	.w5(32'h3c585714),
	.w6(32'hbcd94a5d),
	.w7(32'h3c05785a),
	.w8(32'hbbbdd3a8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d409a32),
	.w1(32'h3be0c895),
	.w2(32'hbbd8edaa),
	.w3(32'h3c9296de),
	.w4(32'hbcc3c315),
	.w5(32'hbb8dc73e),
	.w6(32'hbb794d85),
	.w7(32'hbcb36eed),
	.w8(32'hbcea6870),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc572dbd),
	.w1(32'hba2e3dd3),
	.w2(32'hba0db04f),
	.w3(32'h3b9dc23c),
	.w4(32'hbb060dc5),
	.w5(32'h3b788489),
	.w6(32'hbc86604c),
	.w7(32'hbbbcb175),
	.w8(32'h3c0a7967),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf142c),
	.w1(32'hb9d0d09d),
	.w2(32'hbb0ad5cc),
	.w3(32'hbc497f0d),
	.w4(32'hbc432b0c),
	.w5(32'hbb272cc7),
	.w6(32'h3cb3ce5c),
	.w7(32'hbbeab712),
	.w8(32'h3bd1fba3),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36fcbd),
	.w1(32'hbb9521bb),
	.w2(32'h3a940072),
	.w3(32'hbc16c852),
	.w4(32'hbc890190),
	.w5(32'h3b80e5f3),
	.w6(32'h3aa852b7),
	.w7(32'hba7a95de),
	.w8(32'h3b81205a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e38c1),
	.w1(32'h3cbc1515),
	.w2(32'h3a1e483e),
	.w3(32'h3c6b11b7),
	.w4(32'h3afed379),
	.w5(32'h3c23282b),
	.w6(32'hbca01578),
	.w7(32'hbbcfb30b),
	.w8(32'hbcb6c29c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dadc1),
	.w1(32'hbc50de13),
	.w2(32'hba90df09),
	.w3(32'h3c839db4),
	.w4(32'h3bf4820c),
	.w5(32'h3b15abcf),
	.w6(32'hbc34c3fc),
	.w7(32'h3d2eab20),
	.w8(32'hbbf15c11),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a214155),
	.w1(32'hbbad14ad),
	.w2(32'hbc51ba2e),
	.w3(32'hbb33eca0),
	.w4(32'h3c9c2c52),
	.w5(32'hbb637d86),
	.w6(32'h3a060b78),
	.w7(32'hbac0137b),
	.w8(32'h3c4b65bd),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d06a963),
	.w1(32'hbbdd1e75),
	.w2(32'hbb51b07a),
	.w3(32'h3bc15024),
	.w4(32'hbbf0d0f4),
	.w5(32'hbb6f48f6),
	.w6(32'hbc48705f),
	.w7(32'hb90b54b7),
	.w8(32'h3c06a469),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3abca4),
	.w1(32'hbbf9e222),
	.w2(32'hbbac3503),
	.w3(32'hbccdb71d),
	.w4(32'h3b832f3b),
	.w5(32'h3c3331aa),
	.w6(32'hbcc499f6),
	.w7(32'h3bf11fa3),
	.w8(32'h3cc6f7f3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ced07),
	.w1(32'hbba8efa3),
	.w2(32'hbbfc7d2a),
	.w3(32'h3bf0a492),
	.w4(32'hbbbd2ee3),
	.w5(32'hbc5703a6),
	.w6(32'h3c00c087),
	.w7(32'hbb51ffbb),
	.w8(32'h3aa13547),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89a5b1),
	.w1(32'hbb8776a0),
	.w2(32'hbc02e04d),
	.w3(32'hbbae44ef),
	.w4(32'hbbf9ae5a),
	.w5(32'hbb6e4491),
	.w6(32'hbbf337a6),
	.w7(32'h3c557073),
	.w8(32'hbabd2e8f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18d6ef),
	.w1(32'h3c20357c),
	.w2(32'h3b99aa53),
	.w3(32'hbae01dc0),
	.w4(32'hbbe89575),
	.w5(32'hbdaed390),
	.w6(32'hbb501b93),
	.w7(32'h3a31e778),
	.w8(32'hbcd077b7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb51a1),
	.w1(32'hbc20d056),
	.w2(32'h3cd27c1f),
	.w3(32'hbb960a63),
	.w4(32'h3c8dbb91),
	.w5(32'hbbd0c4e5),
	.w6(32'hba1f7a1e),
	.w7(32'hbcc0ea18),
	.w8(32'hbcbca79c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd842867),
	.w1(32'hbc50bb18),
	.w2(32'hb96d7b2e),
	.w3(32'hbc5b9e9c),
	.w4(32'hbb061a99),
	.w5(32'hbce6db58),
	.w6(32'hbb402016),
	.w7(32'h399f1044),
	.w8(32'hbc4cb003),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a9a3a),
	.w1(32'hbcba1406),
	.w2(32'h3bd73b78),
	.w3(32'h3bb3d2e8),
	.w4(32'hbc808ecf),
	.w5(32'h3cd1ec26),
	.w6(32'hbc4e0049),
	.w7(32'hb9ccd601),
	.w8(32'hbdbe4fc5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd14c0),
	.w1(32'hbb50af26),
	.w2(32'hbbf4af48),
	.w3(32'hbc45fa8d),
	.w4(32'hbd189450),
	.w5(32'hbb3f581b),
	.w6(32'h38bc4927),
	.w7(32'h3c2db214),
	.w8(32'hbc2aeb85),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01a8e0),
	.w1(32'h3c9cec3e),
	.w2(32'hbc81dd21),
	.w3(32'hbd07946f),
	.w4(32'hbce6a5be),
	.w5(32'hbb09e276),
	.w6(32'hbbfe9fa5),
	.w7(32'h3beb3b62),
	.w8(32'hbcce7cad),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccf303b),
	.w1(32'h3bd65cb2),
	.w2(32'hbc4023e4),
	.w3(32'hbc816579),
	.w4(32'h3c03e74c),
	.w5(32'hbca1dd53),
	.w6(32'hbc5ce1e6),
	.w7(32'hbc70506b),
	.w8(32'hbb87daba),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb097077),
	.w1(32'h3ccce969),
	.w2(32'h3b1da3d0),
	.w3(32'h3c1039cd),
	.w4(32'h3c2ed4d9),
	.w5(32'h3c09aadf),
	.w6(32'hbc9a97a0),
	.w7(32'h3c0ebcb5),
	.w8(32'hbcfff227),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc737bc2),
	.w1(32'hbc3855ab),
	.w2(32'hbd061c15),
	.w3(32'hbb454032),
	.w4(32'hbd121bb0),
	.w5(32'h3c36fd0c),
	.w6(32'hbd4d56bc),
	.w7(32'hbd43e669),
	.w8(32'hbc733159),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd73de1d),
	.w1(32'h3c894532),
	.w2(32'hbcb51735),
	.w3(32'hba2b67b7),
	.w4(32'hbce9a3f7),
	.w5(32'h3ac9910f),
	.w6(32'hbda46562),
	.w7(32'hbcf16c2d),
	.w8(32'hbc60d450),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddcd4d),
	.w1(32'hbd78a92f),
	.w2(32'h3b49593a),
	.w3(32'hbcff4e2a),
	.w4(32'hbd7f5b82),
	.w5(32'h3b6014c7),
	.w6(32'h3d1fa5cb),
	.w7(32'hbd05292d),
	.w8(32'h3c20bf7c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e5bb3),
	.w1(32'h3b9ce171),
	.w2(32'hbcd748bf),
	.w3(32'hbcdfd461),
	.w4(32'h3bf7b2d5),
	.w5(32'h3d022c07),
	.w6(32'h3cd34648),
	.w7(32'hbd056a6e),
	.w8(32'hbb9b23f0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ecd9e),
	.w1(32'hbda4225e),
	.w2(32'hbc244879),
	.w3(32'hbc4f3b41),
	.w4(32'h3c3c86de),
	.w5(32'hbcf1cd10),
	.w6(32'h3c2e4e50),
	.w7(32'hbba7ef62),
	.w8(32'h3c74c64d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99dc9d),
	.w1(32'h3c3d9b74),
	.w2(32'hbcc34366),
	.w3(32'hbce5eda5),
	.w4(32'h3b897c7c),
	.w5(32'h3af56761),
	.w6(32'hbd9077e3),
	.w7(32'hbc34bf4c),
	.w8(32'h3a94f46b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd895533),
	.w1(32'hbd2bcecc),
	.w2(32'hbd184100),
	.w3(32'hbcdbbd18),
	.w4(32'hbc0be551),
	.w5(32'hbcee3241),
	.w6(32'hbd1ea672),
	.w7(32'hbbff6bf9),
	.w8(32'hbcef185f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f9eb9),
	.w1(32'h3ac64985),
	.w2(32'hbbaeb3a4),
	.w3(32'hbcc404c0),
	.w4(32'hbbad4b70),
	.w5(32'hb973a11b),
	.w6(32'hbcc29301),
	.w7(32'hbc41d1ee),
	.w8(32'hbc305f6d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf32dde),
	.w1(32'hbb05ea13),
	.w2(32'hbba51c6f),
	.w3(32'hbba85dbe),
	.w4(32'h3bcc1309),
	.w5(32'hbc7d2735),
	.w6(32'h3acedee7),
	.w7(32'hba4d7abb),
	.w8(32'hbbcd8f99),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8937a8),
	.w1(32'h3baeaaf7),
	.w2(32'h3b8a5c07),
	.w3(32'hbb891946),
	.w4(32'h37e87442),
	.w5(32'h3c0df421),
	.w6(32'hbc0083cd),
	.w7(32'h3ba4806d),
	.w8(32'hbb647a84),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d29e4b4),
	.w1(32'hbbbc12a6),
	.w2(32'hbaf96f20),
	.w3(32'h3b1729c2),
	.w4(32'hbaff17d6),
	.w5(32'hba3d809e),
	.w6(32'h3bb42ac5),
	.w7(32'hb9e1e170),
	.w8(32'hbbcfddf2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba641296),
	.w1(32'h3b74e223),
	.w2(32'hba8f0c1b),
	.w3(32'hbb60bdda),
	.w4(32'hba2f3811),
	.w5(32'hbc33c3a9),
	.w6(32'hba083838),
	.w7(32'hbc02ee0e),
	.w8(32'hba8ca2e9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71e373),
	.w1(32'h3c9f63be),
	.w2(32'hbb8dd61d),
	.w3(32'h3b7b7917),
	.w4(32'h3ba387c5),
	.w5(32'h3b582505),
	.w6(32'h3b1d37c6),
	.w7(32'hbb923ca5),
	.w8(32'hba46e438),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69d44f),
	.w1(32'hbc46f541),
	.w2(32'hbb07ac9e),
	.w3(32'hbb9cfcd7),
	.w4(32'hbc03f584),
	.w5(32'h3cc2e8da),
	.w6(32'hbbd0e82f),
	.w7(32'hbb8ebe7b),
	.w8(32'hbaeb1bcb),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc455ced),
	.w1(32'hb912d4d3),
	.w2(32'h3c0c3f62),
	.w3(32'hbb9ab261),
	.w4(32'h3ba2cfe4),
	.w5(32'hbc1683ee),
	.w6(32'hbbe70a13),
	.w7(32'hbbf22673),
	.w8(32'hbaab2415),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc03f),
	.w1(32'h3b315059),
	.w2(32'hbbb751b9),
	.w3(32'h3c103be7),
	.w4(32'h3c1b986c),
	.w5(32'hbbb4db17),
	.w6(32'h3b1192b5),
	.w7(32'hba0091ec),
	.w8(32'h3a75fe1c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f9699),
	.w1(32'hbb233652),
	.w2(32'h3baaf6e2),
	.w3(32'hba7fc92d),
	.w4(32'hb9042d58),
	.w5(32'h3b7de424),
	.w6(32'hbc0177ef),
	.w7(32'h3a8078c8),
	.w8(32'hbbcca0f3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31ccf3),
	.w1(32'h3a64a00f),
	.w2(32'hbb58d74a),
	.w3(32'hba72e72c),
	.w4(32'h3ab6c194),
	.w5(32'hbb0ed1f7),
	.w6(32'h3bfd608b),
	.w7(32'hbc7a67f1),
	.w8(32'h3b0f4d2f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58be59),
	.w1(32'h3b8dd2da),
	.w2(32'h3c8065ae),
	.w3(32'hbb00ded3),
	.w4(32'hbbad9b05),
	.w5(32'hbb455fc7),
	.w6(32'h3c034acd),
	.w7(32'hbb0740ad),
	.w8(32'hbb5bb697),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc292862),
	.w1(32'hba67e1a9),
	.w2(32'hbd3783d0),
	.w3(32'hbc31ec62),
	.w4(32'h3a4987fe),
	.w5(32'hbb3e110d),
	.w6(32'hbbf5160a),
	.w7(32'h3b28e595),
	.w8(32'h39461bc7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb388c93),
	.w1(32'hbb63c2b5),
	.w2(32'hbb9ce506),
	.w3(32'h3a9a9a5c),
	.w4(32'hbad5e127),
	.w5(32'h3b84434b),
	.w6(32'hbacce0f1),
	.w7(32'h3b891688),
	.w8(32'h3cb4a9e0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdf14d2),
	.w1(32'h3b29c80f),
	.w2(32'hbb62d1d7),
	.w3(32'hbbace98c),
	.w4(32'h3bb86233),
	.w5(32'hbbf113d9),
	.w6(32'h3c2962fa),
	.w7(32'hbc5f77f4),
	.w8(32'h39f7e172),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6e9b0),
	.w1(32'h3d9296d5),
	.w2(32'hbbd0bf33),
	.w3(32'h3cde0b40),
	.w4(32'hbc2b0c86),
	.w5(32'h3c6ca3df),
	.w6(32'hbc0e6a8a),
	.w7(32'hbb887b2d),
	.w8(32'h3b0744ab),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d60ca69),
	.w1(32'hbcaffdb2),
	.w2(32'h3caebcb8),
	.w3(32'h3c99ee44),
	.w4(32'h3d7368d7),
	.w5(32'hbcd3a32a),
	.w6(32'h3c1a1c47),
	.w7(32'hbba1e2cc),
	.w8(32'hbc9c24e7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9aa98e),
	.w1(32'h3ca47b5a),
	.w2(32'h3b9a06c0),
	.w3(32'h3bc45e8e),
	.w4(32'h3df1b58c),
	.w5(32'h3cbd35a3),
	.w6(32'h3c8c92ba),
	.w7(32'hbc0c93f6),
	.w8(32'hbcb36548),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4365cb),
	.w1(32'hbc9b11b4),
	.w2(32'h3b5019af),
	.w3(32'hbbfa4c84),
	.w4(32'hbba45dff),
	.w5(32'hbca1be98),
	.w6(32'hbca3b93e),
	.w7(32'hbab63fed),
	.w8(32'hbba70422),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbb6f48),
	.w1(32'hbcc288ba),
	.w2(32'hbc8bac4e),
	.w3(32'h3bb2b951),
	.w4(32'hbc43b2d0),
	.w5(32'hbb9d5d99),
	.w6(32'hbccdb02c),
	.w7(32'hbcc079cf),
	.w8(32'hbc43a694),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb71224),
	.w1(32'h3cc663d2),
	.w2(32'hbd483752),
	.w3(32'hbbb10d04),
	.w4(32'hbc0bc342),
	.w5(32'h3c8f7fe0),
	.w6(32'hbc8f3fc5),
	.w7(32'hbba533ae),
	.w8(32'h3cf49dd5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb876b77),
	.w1(32'h3b4b9923),
	.w2(32'hbe04b9db),
	.w3(32'h3c5cf118),
	.w4(32'hbc260a09),
	.w5(32'h3c857b5a),
	.w6(32'hbc8f66aa),
	.w7(32'hbc099783),
	.w8(32'hbc9df054),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc806c88),
	.w1(32'hbc988117),
	.w2(32'hbcc6b53d),
	.w3(32'h3c0c5c43),
	.w4(32'h3b36aa41),
	.w5(32'h3c0f6d39),
	.w6(32'h3c80fd67),
	.w7(32'hbc78ad6e),
	.w8(32'hbdc3aba7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34b2af),
	.w1(32'h3ad02e03),
	.w2(32'h3c892d27),
	.w3(32'hbce3b31b),
	.w4(32'h3cd14dbe),
	.w5(32'h3caf255b),
	.w6(32'hbd236107),
	.w7(32'h3c78d777),
	.w8(32'h3cb2dac1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca1a4),
	.w1(32'hbc8c0b05),
	.w2(32'hbc5caf7d),
	.w3(32'h3bc4ff49),
	.w4(32'h3d0a1b39),
	.w5(32'hbcdb197e),
	.w6(32'hbc987f5b),
	.w7(32'h3b94871c),
	.w8(32'hbb201538),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3db77011),
	.w1(32'h3c01000e),
	.w2(32'hba90f1a6),
	.w3(32'hbc60a59e),
	.w4(32'hbccedb06),
	.w5(32'hbc147d22),
	.w6(32'h3c09eafe),
	.w7(32'hbca309ac),
	.w8(32'hbbc642a0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccaa969),
	.w1(32'h3bdaec90),
	.w2(32'h3be225ef),
	.w3(32'h3875ddec),
	.w4(32'h3c0ecce4),
	.w5(32'h3870ffdd),
	.w6(32'hbc9bbddb),
	.w7(32'hbcc3612b),
	.w8(32'h3d0309ae),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb491c),
	.w1(32'h3b876b31),
	.w2(32'hba8f3c17),
	.w3(32'hbc604185),
	.w4(32'h3c944cf6),
	.w5(32'h3ae886ce),
	.w6(32'hbc9a0bb5),
	.w7(32'hbbcd6cb9),
	.w8(32'hbc3cde23),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c506705),
	.w1(32'hbbdff448),
	.w2(32'h3be77fd2),
	.w3(32'h3af1bb44),
	.w4(32'h3b071f1c),
	.w5(32'hbc6860ad),
	.w6(32'hbc15335f),
	.w7(32'hbba80168),
	.w8(32'h3bb56186),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0b481b),
	.w1(32'h3c1a6fd6),
	.w2(32'hbce53ce3),
	.w3(32'h3ac9289b),
	.w4(32'hbb9b54af),
	.w5(32'hbacc4de7),
	.w6(32'hbb864820),
	.w7(32'h3cc72afb),
	.w8(32'h3be95244),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ba3a0),
	.w1(32'hbb8bdbbc),
	.w2(32'h3d0840c3),
	.w3(32'hbdbc84f9),
	.w4(32'hbca925c8),
	.w5(32'h3c6c2158),
	.w6(32'hbe1b512d),
	.w7(32'h3b16e00b),
	.w8(32'h3c6a7649),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae315bc),
	.w1(32'hbc396647),
	.w2(32'hbc3f33fe),
	.w3(32'hbb2a14ce),
	.w4(32'h3d073a2a),
	.w5(32'h3d6f9fec),
	.w6(32'hbc0cedaf),
	.w7(32'hb9f7f57f),
	.w8(32'hbc866386),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c275482),
	.w1(32'hbbd7502d),
	.w2(32'hbca5e478),
	.w3(32'hbae7e48c),
	.w4(32'h3bca707c),
	.w5(32'h3bece005),
	.w6(32'h3bb2087b),
	.w7(32'h3c4236b1),
	.w8(32'h3c90a207),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1cb0a1),
	.w1(32'h3c35580e),
	.w2(32'hbcd9b2ea),
	.w3(32'h3cbc65a3),
	.w4(32'h3c040dda),
	.w5(32'hbc0d1d8f),
	.w6(32'hbc56f668),
	.w7(32'h3be5ec9c),
	.w8(32'h3c592f27),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27ad1b),
	.w1(32'hbd3357e0),
	.w2(32'h39ef69e3),
	.w3(32'h3b033f46),
	.w4(32'h3d818ef6),
	.w5(32'h3b1b704c),
	.w6(32'hbd037f38),
	.w7(32'hba2f3436),
	.w8(32'hbcd68ac4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62b7be),
	.w1(32'hbb5006c2),
	.w2(32'hbcf3face),
	.w3(32'hbc0a9874),
	.w4(32'h3c8f8b52),
	.w5(32'hbcc535e2),
	.w6(32'h3c809eae),
	.w7(32'hbb8ff567),
	.w8(32'hbc79ff12),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16be45),
	.w1(32'h3d10e204),
	.w2(32'h3c7bef24),
	.w3(32'hbc0c9473),
	.w4(32'h3c0fd140),
	.w5(32'h3d16978e),
	.w6(32'h3970cf3f),
	.w7(32'h3d068e2b),
	.w8(32'hbd5bba35),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca567de),
	.w1(32'hbd132263),
	.w2(32'hbc7ed81c),
	.w3(32'hbd21f408),
	.w4(32'hbd07c7c0),
	.w5(32'hbb26e798),
	.w6(32'hbcd108a6),
	.w7(32'hbce249fa),
	.w8(32'hbb958910),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8991bf),
	.w1(32'hbc059f04),
	.w2(32'h3cca6323),
	.w3(32'h3c1a268a),
	.w4(32'hbba06960),
	.w5(32'h3bbbf9d5),
	.w6(32'hb6a674de),
	.w7(32'hbc06b738),
	.w8(32'h3caf07f7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c2916),
	.w1(32'hbd0b8b2d),
	.w2(32'h3ce15d50),
	.w3(32'hbc15ad8b),
	.w4(32'hbd80e9b5),
	.w5(32'h3c150160),
	.w6(32'hbb9ae4c2),
	.w7(32'hbc7b2cf8),
	.w8(32'hbaf94632),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0ff35),
	.w1(32'hbbf5b55b),
	.w2(32'hb9711737),
	.w3(32'h3cb67baa),
	.w4(32'hbc6b6b7c),
	.w5(32'h3c6098c7),
	.w6(32'h3d1d3989),
	.w7(32'h3c8718f0),
	.w8(32'hbc827461),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb360a86),
	.w1(32'hbd022596),
	.w2(32'hbd926f80),
	.w3(32'h3cb82f37),
	.w4(32'h3bc83088),
	.w5(32'h3ab76fec),
	.w6(32'hbb4d7789),
	.w7(32'hbc9cb99c),
	.w8(32'h3b206f5a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca85805),
	.w1(32'h3b24e98b),
	.w2(32'hbbb2c02f),
	.w3(32'h3c3f1ef4),
	.w4(32'h3c600e1b),
	.w5(32'h3c122703),
	.w6(32'hbb955715),
	.w7(32'hbb603655),
	.w8(32'hbc309cbe),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b996db9),
	.w1(32'h3a48ecc4),
	.w2(32'h3aba062e),
	.w3(32'hbba059f6),
	.w4(32'h3b431165),
	.w5(32'h3b12bb0b),
	.w6(32'h39de3e57),
	.w7(32'h3c3266b6),
	.w8(32'hbb11e375),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule