module layer_10_featuremap_196(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cea0b5),
	.w1(32'h3a5dd07b),
	.w2(32'hb94c6c44),
	.w3(32'h39ecf41f),
	.w4(32'h39a5e0d3),
	.w5(32'hb9d4e8b7),
	.w6(32'h3a505bb2),
	.w7(32'h3a2ab35e),
	.w8(32'h39c18da1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36ea09),
	.w1(32'h3b0ba395),
	.w2(32'h3ad545da),
	.w3(32'h3a8390c5),
	.w4(32'hb9d46513),
	.w5(32'hb962ecb5),
	.w6(32'h3aa25424),
	.w7(32'hba8a4d1c),
	.w8(32'hb991b4c6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9095c36),
	.w1(32'hb87083b6),
	.w2(32'hb9e2edac),
	.w3(32'hb8d4a74b),
	.w4(32'h3858367d),
	.w5(32'hb8dcf80f),
	.w6(32'h388e0d68),
	.w7(32'hb8bbfaa4),
	.w8(32'hb8986572),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f0f98b),
	.w1(32'h39294e41),
	.w2(32'hb81d9063),
	.w3(32'h38bd0182),
	.w4(32'h3a41e9c4),
	.w5(32'h3a71106d),
	.w6(32'hba269708),
	.w7(32'hba2909d4),
	.w8(32'h377d4fbe),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb7769),
	.w1(32'h38819877),
	.w2(32'hba1c0bb8),
	.w3(32'h3a912fc4),
	.w4(32'h393aa425),
	.w5(32'hb9a2d9f5),
	.w6(32'h3a332784),
	.w7(32'h3a1eb3d8),
	.w8(32'h391370a3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f7eb7),
	.w1(32'h3a0d5b13),
	.w2(32'h3a65b59c),
	.w3(32'hb91cc9d0),
	.w4(32'h3a085504),
	.w5(32'h3a6a6107),
	.w6(32'h3a2da4d1),
	.w7(32'h3a7be753),
	.w8(32'h3a5087db),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6b3b6),
	.w1(32'h3a838de2),
	.w2(32'hba250e08),
	.w3(32'h3b3463a1),
	.w4(32'h3a41c564),
	.w5(32'h3a58f754),
	.w6(32'hbb7915bb),
	.w7(32'hba9f7fb1),
	.w8(32'h3a80491d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb225bca),
	.w1(32'hbc23d0fe),
	.w2(32'hbad00592),
	.w3(32'hbad4687d),
	.w4(32'h3b6d4ae3),
	.w5(32'h3aeca607),
	.w6(32'hbbd86eca),
	.w7(32'hbb9bbe89),
	.w8(32'h3a692233),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac5366),
	.w1(32'hb999beb4),
	.w2(32'hba050ca5),
	.w3(32'h3a3b3c20),
	.w4(32'h3976903d),
	.w5(32'hb8b63d3e),
	.w6(32'h3a3abfb0),
	.w7(32'h3a80aeb9),
	.w8(32'h3960a427),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabff586),
	.w1(32'hbaab41f8),
	.w2(32'h3927cffc),
	.w3(32'h3a64031d),
	.w4(32'hbad216c9),
	.w5(32'h395aec5c),
	.w6(32'hbb2683fc),
	.w7(32'hba558960),
	.w8(32'h3a3202c8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f18e1),
	.w1(32'hb9a9420e),
	.w2(32'hba2aeeaf),
	.w3(32'hba48066f),
	.w4(32'hb7c8f9fd),
	.w5(32'hb9f30e71),
	.w6(32'h3a672b09),
	.w7(32'h39a9e2a1),
	.w8(32'hba089927),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61dd9d),
	.w1(32'h3a64de71),
	.w2(32'hba3f9824),
	.w3(32'h3baaa294),
	.w4(32'h3b381f7f),
	.w5(32'h3b235a88),
	.w6(32'hbb28f0ba),
	.w7(32'hb98f599a),
	.w8(32'h3b14814f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a181cad),
	.w1(32'h37e8f7c7),
	.w2(32'hba3bc207),
	.w3(32'h3b2545ee),
	.w4(32'h3aad53f9),
	.w5(32'h3a89d39f),
	.w6(32'h39f07098),
	.w7(32'h3b0522b6),
	.w8(32'h3b037065),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6944e),
	.w1(32'h3a9f66c3),
	.w2(32'h3b250043),
	.w3(32'h3aca4f64),
	.w4(32'h3a1ef55c),
	.w5(32'h3a842060),
	.w6(32'hba21c76c),
	.w7(32'h389fbb7b),
	.w8(32'h3a33f573),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3850ffc0),
	.w1(32'hb99cbc98),
	.w2(32'h3a0bf0e4),
	.w3(32'h3a6c45ac),
	.w4(32'hb9d348bc),
	.w5(32'h36f80f52),
	.w6(32'hba68f12f),
	.w7(32'hbabe6478),
	.w8(32'hb825a051),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba648a8),
	.w1(32'h37b22d56),
	.w2(32'h387d326b),
	.w3(32'hbaa8b35c),
	.w4(32'hbad21e8d),
	.w5(32'h3aa518f9),
	.w6(32'hba829ad9),
	.w7(32'h38a5719f),
	.w8(32'h3a870a25),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a092e54),
	.w1(32'h389c31cc),
	.w2(32'h37231165),
	.w3(32'h39d59dab),
	.w4(32'hb99b98ac),
	.w5(32'hb9d7e1d7),
	.w6(32'hb990236f),
	.w7(32'hb89ed83f),
	.w8(32'hb9285a41),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5eef4),
	.w1(32'hbc1b3b9b),
	.w2(32'hbbe7ea8f),
	.w3(32'hbb8f083b),
	.w4(32'hbba6d9a9),
	.w5(32'hbb1de6cb),
	.w6(32'hbb80bc52),
	.w7(32'hba9a3375),
	.w8(32'hb7e341c4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16ff0b),
	.w1(32'hbb26572d),
	.w2(32'hbae3d3f3),
	.w3(32'hbad8f14a),
	.w4(32'hba95a0cf),
	.w5(32'hb7d692dc),
	.w6(32'hbb1e6aec),
	.w7(32'h3849dd55),
	.w8(32'h3a74d332),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc1f77),
	.w1(32'h384cbf2a),
	.w2(32'hb851a8ff),
	.w3(32'hb8c6030d),
	.w4(32'h38bd7c02),
	.w5(32'h38928235),
	.w6(32'h393ba469),
	.w7(32'h389c4871),
	.w8(32'h3802502a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383a165d),
	.w1(32'h3971b886),
	.w2(32'h39d8ed24),
	.w3(32'h389f1a70),
	.w4(32'h399fa517),
	.w5(32'h39f28f28),
	.w6(32'h3960d769),
	.w7(32'h39adb584),
	.w8(32'h399146ea),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8ac1d),
	.w1(32'h3b03150b),
	.w2(32'h3a6299f0),
	.w3(32'h3af5149c),
	.w4(32'h3aaaf8b7),
	.w5(32'h3988a48d),
	.w6(32'h3b206e30),
	.w7(32'h3a12f13a),
	.w8(32'h389b1f50),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e636c),
	.w1(32'hbbe8a5dc),
	.w2(32'hbbd96a1d),
	.w3(32'hbc1017bf),
	.w4(32'hbbd0c9fe),
	.w5(32'h39bb093f),
	.w6(32'hbc17f6f2),
	.w7(32'hba87fd77),
	.w8(32'h3b1606bf),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ad5ce),
	.w1(32'h39e7e6bf),
	.w2(32'h3b378b1a),
	.w3(32'h39dc92fc),
	.w4(32'h3a94a61f),
	.w5(32'h3b5e8c3d),
	.w6(32'hb95d8e32),
	.w7(32'h3a4be5ff),
	.w8(32'h3b30cc7d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae36422),
	.w1(32'h3b80de51),
	.w2(32'h3b2edbf6),
	.w3(32'h3b3dadc0),
	.w4(32'h3ad6aa45),
	.w5(32'h3a4e4027),
	.w6(32'h3aed8c91),
	.w7(32'hbb552ccf),
	.w8(32'hbb457d0d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e07085),
	.w1(32'h39844221),
	.w2(32'h39a8ba27),
	.w3(32'hb969f645),
	.w4(32'h3972eb5c),
	.w5(32'h3946229f),
	.w6(32'hb7faded1),
	.w7(32'h39994de9),
	.w8(32'h397f076b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d82f4),
	.w1(32'h387dc2cc),
	.w2(32'hb898817d),
	.w3(32'h3984499e),
	.w4(32'hb72315f5),
	.w5(32'h37379b35),
	.w6(32'h39451d1d),
	.w7(32'h38b96824),
	.w8(32'h37d7b6fa),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17365e),
	.w1(32'h3a7d6fe9),
	.w2(32'hbab2ed75),
	.w3(32'h3a371e2b),
	.w4(32'hbb2b8e71),
	.w5(32'hbb895438),
	.w6(32'h3bdbf668),
	.w7(32'h3b8a9579),
	.w8(32'hbaa38a25),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a047a5a),
	.w1(32'h385d636d),
	.w2(32'h39a36c9f),
	.w3(32'h3a527a2e),
	.w4(32'h3a688547),
	.w5(32'h3a14668d),
	.w6(32'h3a8020ab),
	.w7(32'h3a253280),
	.w8(32'h3a32a4a4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add0e8d),
	.w1(32'h3b9d74a9),
	.w2(32'h3b19aac1),
	.w3(32'h395e6bcf),
	.w4(32'hba846729),
	.w5(32'hbb076bf9),
	.w6(32'h3bb4d0e9),
	.w7(32'h39d83e3e),
	.w8(32'hbaa090bc),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3912ef3e),
	.w1(32'h399fc76a),
	.w2(32'h399698e1),
	.w3(32'hb8ce37db),
	.w4(32'h395e9780),
	.w5(32'h399b6553),
	.w6(32'h3964b5f3),
	.w7(32'h399af776),
	.w8(32'h3980d51a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915961f),
	.w1(32'h38e0b871),
	.w2(32'h38faf1cf),
	.w3(32'h3946a885),
	.w4(32'h38bb7db0),
	.w5(32'h38bf02c8),
	.w6(32'h38eb3de3),
	.w7(32'h399d0d89),
	.w8(32'h398a6562),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2aca4),
	.w1(32'h38a01b50),
	.w2(32'h3a1e1309),
	.w3(32'h3a113e55),
	.w4(32'h3a5d8dce),
	.w5(32'h3ad2e622),
	.w6(32'hba955ac4),
	.w7(32'h39c95ed4),
	.w8(32'h3acb9356),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c2443),
	.w1(32'h3a776b81),
	.w2(32'h3937b440),
	.w3(32'h391b463f),
	.w4(32'hb98a47e6),
	.w5(32'hb9c71b72),
	.w6(32'hb8a3af53),
	.w7(32'hbab3ad0a),
	.w8(32'hba8575a2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d47633),
	.w1(32'hb9093b4e),
	.w2(32'hba216945),
	.w3(32'h391322fb),
	.w4(32'hb9f92246),
	.w5(32'hb9233a85),
	.w6(32'hba019575),
	.w7(32'hba11ca87),
	.w8(32'hb9852268),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc98f7),
	.w1(32'hb9c79016),
	.w2(32'hb89b5de9),
	.w3(32'hba6a787b),
	.w4(32'h3a053cf9),
	.w5(32'h3b05d64a),
	.w6(32'hbaf32a61),
	.w7(32'hba0f3cf6),
	.w8(32'h3abceb1f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e87dc),
	.w1(32'hbbfe4835),
	.w2(32'h394ed4bc),
	.w3(32'h3ad26e84),
	.w4(32'hbbc5d0bb),
	.w5(32'h3af9940a),
	.w6(32'hbc09b49b),
	.w7(32'hbbe63ac2),
	.w8(32'h3b9fdce7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de14d8),
	.w1(32'h3b6090c1),
	.w2(32'h3ac07893),
	.w3(32'h3b6e5dad),
	.w4(32'hba060ccc),
	.w5(32'hbb0d99b1),
	.w6(32'h3b962e85),
	.w7(32'hbb6bca23),
	.w8(32'hbb0b8801),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4abff9),
	.w1(32'h3bc84c9a),
	.w2(32'h39b25169),
	.w3(32'h3bd34228),
	.w4(32'h3a08fdae),
	.w5(32'hbb7104d4),
	.w6(32'h3c478aae),
	.w7(32'h3aefb951),
	.w8(32'hbb2f1102),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a919f81),
	.w1(32'h39f04595),
	.w2(32'h3a1aff81),
	.w3(32'h3a602d1d),
	.w4(32'hba16d20a),
	.w5(32'hb981c812),
	.w6(32'h3a0ea9b3),
	.w7(32'hba616d0e),
	.w8(32'h37db9d82),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca7b52),
	.w1(32'hb9b165a1),
	.w2(32'hb88c9a98),
	.w3(32'hb9a43850),
	.w4(32'hb9cbb809),
	.w5(32'hb908a405),
	.w6(32'hba0f8626),
	.w7(32'hb97d4b3f),
	.w8(32'hb8d8ffa0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992edce),
	.w1(32'h39569ff5),
	.w2(32'h37269d9a),
	.w3(32'h392aebd9),
	.w4(32'h38bdb5b0),
	.w5(32'hb91416d1),
	.w6(32'h39912dde),
	.w7(32'hb8a72fbc),
	.w8(32'hb916db92),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17ba51),
	.w1(32'h38ca276d),
	.w2(32'h38b05796),
	.w3(32'hba1d1ce3),
	.w4(32'h396034a8),
	.w5(32'h385e8957),
	.w6(32'hb9b98336),
	.w7(32'h39082323),
	.w8(32'h393d2627),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe52d3c),
	.w1(32'hbb81a52c),
	.w2(32'hbae28c30),
	.w3(32'hbb69a84d),
	.w4(32'hbad09c6d),
	.w5(32'h3b18ba86),
	.w6(32'hb9891811),
	.w7(32'h3b1afb01),
	.w8(32'h3b5e9a95),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cbf2c),
	.w1(32'hb900619c),
	.w2(32'h381d1b3c),
	.w3(32'hbaa54929),
	.w4(32'hb996f935),
	.w5(32'h3a157cd1),
	.w6(32'h38967a3a),
	.w7(32'hba25319a),
	.w8(32'h399a5bd4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e08223),
	.w1(32'h3921e2ba),
	.w2(32'h3ad2164b),
	.w3(32'h38641b70),
	.w4(32'h3ae4b671),
	.w5(32'h3b700a9e),
	.w6(32'h380ec63f),
	.w7(32'hb99f107c),
	.w8(32'h3b1dfb49),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04504f),
	.w1(32'hbb10d987),
	.w2(32'h3a1909ab),
	.w3(32'hba2fe0f7),
	.w4(32'hbab7b800),
	.w5(32'h3a6b3c5f),
	.w6(32'hbb1ef81c),
	.w7(32'hbaa8194b),
	.w8(32'h3a1cee28),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6974f5),
	.w1(32'hbc0ac506),
	.w2(32'hbbda8146),
	.w3(32'hbacdec31),
	.w4(32'hbaec6117),
	.w5(32'hba0768b3),
	.w6(32'hbb74ef0b),
	.w7(32'h3aaa539d),
	.w8(32'h3b5c896d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c576c5),
	.w1(32'hb75f15d2),
	.w2(32'h387d57d1),
	.w3(32'h38befbff),
	.w4(32'h38ff6e2b),
	.w5(32'h39430a5d),
	.w6(32'h3985e7f1),
	.w7(32'h39873f97),
	.w8(32'h392483ba),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba198e24),
	.w1(32'h3937e25b),
	.w2(32'h388ab7c7),
	.w3(32'hba93aa2b),
	.w4(32'hb9d52355),
	.w5(32'hb8adab13),
	.w6(32'hba0b38f9),
	.w7(32'hb9edc165),
	.w8(32'hb989364a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ea1bc),
	.w1(32'hb97c4a59),
	.w2(32'hba21668b),
	.w3(32'h3a803ea4),
	.w4(32'hb809c281),
	.w5(32'hba11146a),
	.w6(32'hb967598d),
	.w7(32'hba0bc05d),
	.w8(32'hba252a2c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5b0d8),
	.w1(32'h3916b659),
	.w2(32'h38b562ec),
	.w3(32'hb9ba7b82),
	.w4(32'h3a0472ed),
	.w5(32'h3a7831a3),
	.w6(32'hb9464ef8),
	.w7(32'hb97e4c8d),
	.w8(32'hb9bf73e9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39667cec),
	.w1(32'hba477d48),
	.w2(32'hb9ce373a),
	.w3(32'hba094a56),
	.w4(32'hb8b1c164),
	.w5(32'h39f3e241),
	.w6(32'hb9ed6eb1),
	.w7(32'h39399653),
	.w8(32'h3a292149),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8348b7),
	.w1(32'hbbd571a7),
	.w2(32'hbb34a984),
	.w3(32'hbb0582ef),
	.w4(32'hbb6c0e11),
	.w5(32'h3982584f),
	.w6(32'hbb7d73b3),
	.w7(32'h3a61b046),
	.w8(32'h3b3c3c08),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae79553),
	.w1(32'hbac1ade8),
	.w2(32'hbac719f5),
	.w3(32'hba1342d5),
	.w4(32'hb95c09ba),
	.w5(32'hb9810e1c),
	.w6(32'h3a440746),
	.w7(32'h3a1e052b),
	.w8(32'hb9973858),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ad8154),
	.w1(32'h399f167f),
	.w2(32'h38f10ca9),
	.w3(32'hb8c5f258),
	.w4(32'hb9025f26),
	.w5(32'hb9605bfa),
	.w6(32'hb86058ff),
	.w7(32'hb9af0db3),
	.w8(32'hb9928b12),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3948f191),
	.w1(32'hb62070fc),
	.w2(32'hb9439267),
	.w3(32'h381fbc29),
	.w4(32'h38332506),
	.w5(32'hb8100a99),
	.w6(32'h36b97c41),
	.w7(32'hb9513603),
	.w8(32'hb85055ba),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb962220a),
	.w1(32'hba056bbe),
	.w2(32'hba2b5a32),
	.w3(32'hb9acc7c1),
	.w4(32'hba17e0ea),
	.w5(32'hba30959c),
	.w6(32'hb8b60116),
	.w7(32'hb9f54008),
	.w8(32'hb948c546),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c02c2),
	.w1(32'h39bebdb8),
	.w2(32'hb8b7dd21),
	.w3(32'h39c66c00),
	.w4(32'h394acc31),
	.w5(32'hb986e1e8),
	.w6(32'h39b9a855),
	.w7(32'hb84876eb),
	.w8(32'h36e37f70),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e8f56),
	.w1(32'h3822f61c),
	.w2(32'h39c59c15),
	.w3(32'hb99c5357),
	.w4(32'h39011119),
	.w5(32'h39ecbac3),
	.w6(32'h3a623d98),
	.w7(32'h3a129cba),
	.w8(32'h39d73f15),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad33c32),
	.w1(32'hbb0870d3),
	.w2(32'hbacd0088),
	.w3(32'hba565a7e),
	.w4(32'hba3e2fdf),
	.w5(32'h39473b5c),
	.w6(32'hba68e70c),
	.w7(32'h39bfc3bc),
	.w8(32'h3a4ce9d7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb73211),
	.w1(32'hba5f8a9b),
	.w2(32'hbac01f92),
	.w3(32'hbb58ff4e),
	.w4(32'hba347b8d),
	.w5(32'hba9ee026),
	.w6(32'h3a4a22ce),
	.w7(32'h3a9707e6),
	.w8(32'hba8d7352),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a022022),
	.w1(32'hb8c5f57b),
	.w2(32'hba2c8355),
	.w3(32'h3a26474f),
	.w4(32'hb8bdb8f4),
	.w5(32'hb9b43bb4),
	.w6(32'hb901835d),
	.w7(32'hb9848d09),
	.w8(32'h393184e7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb924ba38),
	.w1(32'hba0d128f),
	.w2(32'hba38d283),
	.w3(32'hb99de5a6),
	.w4(32'hb9c7656f),
	.w5(32'hba1aa76f),
	.w6(32'hb9e266e1),
	.w7(32'hba2687ad),
	.w8(32'hba05b83a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba381e86),
	.w1(32'hb8372b85),
	.w2(32'hb90e322a),
	.w3(32'hba0970aa),
	.w4(32'h37e5676c),
	.w5(32'hb8e85780),
	.w6(32'hb898168a),
	.w7(32'hb96cf3ae),
	.w8(32'hb8a76291),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4dbad),
	.w1(32'hba025794),
	.w2(32'hb99a60de),
	.w3(32'hb96c8307),
	.w4(32'hb9ce17f9),
	.w5(32'hb94ae6c9),
	.w6(32'hb9a7ac81),
	.w7(32'hb98cef58),
	.w8(32'h398e038d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fd1b3),
	.w1(32'hb98dbb07),
	.w2(32'h3b6e2b0c),
	.w3(32'h3be456ef),
	.w4(32'hb9bee949),
	.w5(32'h390307e8),
	.w6(32'hbab36b05),
	.w7(32'h3b5e6cc4),
	.w8(32'h3b3ee07c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fb674),
	.w1(32'h3762d5c2),
	.w2(32'h36a6250a),
	.w3(32'h3a907b8c),
	.w4(32'h3b8dd828),
	.w5(32'h3b948d97),
	.w6(32'hbb1d9244),
	.w7(32'h3a8ce666),
	.w8(32'h3b2957a9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c38df),
	.w1(32'hbb17147c),
	.w2(32'hbb2adcfc),
	.w3(32'hb9e2d33d),
	.w4(32'h393e4998),
	.w5(32'h39f7a896),
	.w6(32'h38dbc400),
	.w7(32'h3a09c08f),
	.w8(32'hbad2716a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe2f78),
	.w1(32'h3b7fa23e),
	.w2(32'h3ab69d79),
	.w3(32'h3af3171a),
	.w4(32'hba29ad24),
	.w5(32'hb8e87a1c),
	.w6(32'hb9a4d6ec),
	.w7(32'hbbc461be),
	.w8(32'hbb42967c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2da74e),
	.w1(32'hb9851dec),
	.w2(32'hba063e8f),
	.w3(32'hb9bd746b),
	.w4(32'hb96ae911),
	.w5(32'hb9d3f974),
	.w6(32'hb9409834),
	.w7(32'hb9b4e6cd),
	.w8(32'hb978a65a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba048cfc),
	.w1(32'h38de9ac1),
	.w2(32'h393b02cd),
	.w3(32'hb9ba7fce),
	.w4(32'h38b159de),
	.w5(32'h395c9141),
	.w6(32'h38937b3f),
	.w7(32'h38f7ea45),
	.w8(32'h394aa077),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996027d),
	.w1(32'h38f19cea),
	.w2(32'h3953891d),
	.w3(32'h399fe697),
	.w4(32'h39105eee),
	.w5(32'h39853f1b),
	.w6(32'h390ff05a),
	.w7(32'h393bd9e6),
	.w8(32'h39831c7c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9657e34),
	.w1(32'hba6ebfa2),
	.w2(32'hba4a7029),
	.w3(32'h3a0c687e),
	.w4(32'h39408545),
	.w5(32'h3900c381),
	.w6(32'h393c1990),
	.w7(32'h3a1e4a27),
	.w8(32'h3a17a248),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f7c498),
	.w1(32'h394f9b1e),
	.w2(32'h386b0ded),
	.w3(32'h397cf57b),
	.w4(32'h393b63e8),
	.w5(32'hb7ff099a),
	.w6(32'h396475c7),
	.w7(32'h392f2584),
	.w8(32'h38ee8b08),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb129d22),
	.w1(32'hbba0100b),
	.w2(32'hba0f102b),
	.w3(32'hb977e099),
	.w4(32'hbaee2e7e),
	.w5(32'hb99c644c),
	.w6(32'hbb4de2c7),
	.w7(32'hbafbaff9),
	.w8(32'h3ab9b3ca),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2da69f),
	.w1(32'hbbeebeac),
	.w2(32'hbae6b1d0),
	.w3(32'hbabc554c),
	.w4(32'hbb2233ce),
	.w5(32'h3af7dc59),
	.w6(32'hbbaca78f),
	.w7(32'hbb38d673),
	.w8(32'h3aea1fde),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8df4dd),
	.w1(32'h3b15b4ff),
	.w2(32'h3aaf4e4b),
	.w3(32'h3b3d6273),
	.w4(32'h3a78665a),
	.w5(32'h39eea554),
	.w6(32'h3adc8ca5),
	.w7(32'hb9396c61),
	.w8(32'h39de45a5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb191eae),
	.w1(32'hbb03d7cb),
	.w2(32'hba375960),
	.w3(32'hba4f4a24),
	.w4(32'hba272ec4),
	.w5(32'hb998f769),
	.w6(32'hba05aa93),
	.w7(32'h39c7aefd),
	.w8(32'hb930decb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38222b4d),
	.w1(32'hbaee20ae),
	.w2(32'h3a88a0e1),
	.w3(32'h3b71df00),
	.w4(32'hb8961c50),
	.w5(32'h3a9418ad),
	.w6(32'hbaacb561),
	.w7(32'hb8253067),
	.w8(32'h3ae6c2b7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3fd40),
	.w1(32'hba5aaff1),
	.w2(32'hba057a2b),
	.w3(32'hb90378cf),
	.w4(32'hba4c6921),
	.w5(32'hba11ae92),
	.w6(32'h38ccff36),
	.w7(32'hb9846da5),
	.w8(32'hba57ef61),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97a671),
	.w1(32'hbb2a65f1),
	.w2(32'hbaf22929),
	.w3(32'hb8b063f0),
	.w4(32'hba587a31),
	.w5(32'hb78bd9ed),
	.w6(32'hbad99cb4),
	.w7(32'h3921a33a),
	.w8(32'h3a84749a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39398c99),
	.w1(32'h38c1b27a),
	.w2(32'hb885a39b),
	.w3(32'h39348190),
	.w4(32'h38045602),
	.w5(32'hb868bdf7),
	.w6(32'h3813f509),
	.w7(32'h379571c8),
	.w8(32'h37a1af0d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb893b767),
	.w1(32'h393983db),
	.w2(32'h38a437cf),
	.w3(32'hb8a91c88),
	.w4(32'h394b68ef),
	.w5(32'h38c3c96a),
	.w6(32'h38e42f77),
	.w7(32'h391d1039),
	.w8(32'h38e367e8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64dd5a6),
	.w1(32'hba1327c8),
	.w2(32'hb99246c4),
	.w3(32'h3966cec8),
	.w4(32'h37356fa7),
	.w5(32'h3984b5f5),
	.w6(32'hb983340b),
	.w7(32'h3898069d),
	.w8(32'hb897f64d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9810f55),
	.w1(32'hb945609b),
	.w2(32'hb9af90e2),
	.w3(32'h3981af45),
	.w4(32'hb9d0a9d6),
	.w5(32'hb9f18388),
	.w6(32'h3980b099),
	.w7(32'hb9ce2f7b),
	.w8(32'hb9e2258d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d998c8),
	.w1(32'h3b1175d3),
	.w2(32'h3b0ae1ac),
	.w3(32'h3a497fa4),
	.w4(32'hb9291593),
	.w5(32'h3a113691),
	.w6(32'hb9434be8),
	.w7(32'hbade4d78),
	.w8(32'hba13c940),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37390c94),
	.w1(32'h39e9c8cd),
	.w2(32'h3a094a2b),
	.w3(32'h38187ab4),
	.w4(32'h39b9ab8a),
	.w5(32'h39fe4a8d),
	.w6(32'h397e4e63),
	.w7(32'h398e9d47),
	.w8(32'h39c0a56f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85015e),
	.w1(32'h39997728),
	.w2(32'hb9ec4a71),
	.w3(32'hba841f70),
	.w4(32'hba67b515),
	.w5(32'h3a579440),
	.w6(32'hbb0e5082),
	.w7(32'hbaab1c4e),
	.w8(32'h38c14bea),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba063fd),
	.w1(32'hbbc6d180),
	.w2(32'hbb6b8950),
	.w3(32'hbb9e79c0),
	.w4(32'hbb856a19),
	.w5(32'h39b6462a),
	.w6(32'hbbce41db),
	.w7(32'hbb15ef6c),
	.w8(32'h39ad856b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dc3392),
	.w1(32'h3ad0b4f7),
	.w2(32'hb9efe5d8),
	.w3(32'h3ab7ef08),
	.w4(32'hb9e38e64),
	.w5(32'hbadd8865),
	.w6(32'h3b82400f),
	.w7(32'h3a9cf1ee),
	.w8(32'hb9c8aa8f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a292b7e),
	.w1(32'h3a394638),
	.w2(32'hb91cfab8),
	.w3(32'h3bc87525),
	.w4(32'hba9c7a4c),
	.w5(32'hba80fec9),
	.w6(32'h3a4f3056),
	.w7(32'h3b77ba0a),
	.w8(32'h3bb0109c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c7323),
	.w1(32'hb90bfa46),
	.w2(32'h399826c7),
	.w3(32'h3927cd9c),
	.w4(32'hb868a597),
	.w5(32'h3a3e3751),
	.w6(32'h3a9e6ee9),
	.w7(32'hba56b3f5),
	.w8(32'h38875921),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60f390),
	.w1(32'hbb311496),
	.w2(32'h3a05d16f),
	.w3(32'hb9f71231),
	.w4(32'hbab70954),
	.w5(32'h3a9362fa),
	.w6(32'hbb1705ec),
	.w7(32'hb9f26e5e),
	.w8(32'h3a6d6918),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb002777),
	.w1(32'h3a80f743),
	.w2(32'h3ade0086),
	.w3(32'h3a58f378),
	.w4(32'hba2f9195),
	.w5(32'hb8bd9ecb),
	.w6(32'hba317311),
	.w7(32'h3a14e5bd),
	.w8(32'h3a801a6e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393870a0),
	.w1(32'h3b17cb87),
	.w2(32'h3a5c5b9c),
	.w3(32'h3a247de0),
	.w4(32'hbaaa9450),
	.w5(32'hba63f011),
	.w6(32'h3b35e9fa),
	.w7(32'h3a016755),
	.w8(32'hb8b7252e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fa379),
	.w1(32'hb8c593c8),
	.w2(32'hba24958b),
	.w3(32'h3a8396d8),
	.w4(32'h38f41fd7),
	.w5(32'hb9bd1d73),
	.w6(32'hb981a4de),
	.w7(32'h395cb5e7),
	.w8(32'hb8fa7fdf),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa47437),
	.w1(32'hbb26c784),
	.w2(32'hba00b7be),
	.w3(32'hba8af40f),
	.w4(32'hb905b2a7),
	.w5(32'h3b0a184b),
	.w6(32'hbb1bf3f0),
	.w7(32'h3a3ebbca),
	.w8(32'h3b269931),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13f0e6),
	.w1(32'h39d68504),
	.w2(32'h3aa0c3ed),
	.w3(32'h3bc550b9),
	.w4(32'h3b0c9929),
	.w5(32'h3a8d1da6),
	.w6(32'hba06b106),
	.w7(32'h3989fb8e),
	.w8(32'h3af44a74),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b068886),
	.w1(32'hbbd579aa),
	.w2(32'hbaf6e4a9),
	.w3(32'hbbf9c40c),
	.w4(32'hbc00da07),
	.w5(32'h3b707303),
	.w6(32'hbc3908f4),
	.w7(32'hbbeaf6f2),
	.w8(32'h3b345cc5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae46425),
	.w1(32'h3a9334c7),
	.w2(32'hbb32d43f),
	.w3(32'h39868851),
	.w4(32'hbb146c32),
	.w5(32'hbb80181e),
	.w6(32'h3b7ad7b5),
	.w7(32'hba0527cc),
	.w8(32'h3a96c66f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984c7cf),
	.w1(32'h3aaab7d8),
	.w2(32'h3b55a73f),
	.w3(32'hb9d64110),
	.w4(32'hb80e8d0f),
	.w5(32'h3b3190d0),
	.w6(32'hba8c91dd),
	.w7(32'hbb07518b),
	.w8(32'hba0042ad),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d3d27),
	.w1(32'hbba5e89f),
	.w2(32'h38ade93f),
	.w3(32'h3bc19ed0),
	.w4(32'hba8a323c),
	.w5(32'h3b19c7cf),
	.w6(32'hb97dbd00),
	.w7(32'h39c3e9c1),
	.w8(32'h3bba0de4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcdf6c),
	.w1(32'h3a30f12d),
	.w2(32'h3a8b0a31),
	.w3(32'h3aadc233),
	.w4(32'h3a71d31a),
	.w5(32'h3ac56e04),
	.w6(32'h3a158a7b),
	.w7(32'h3abf6c53),
	.w8(32'h3ad4d95e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb169695),
	.w1(32'hbc18cbd5),
	.w2(32'hbbfdd46d),
	.w3(32'hbb4cbf04),
	.w4(32'hbbe81d11),
	.w5(32'hbb560bd0),
	.w6(32'hbc13048e),
	.w7(32'hbc19919b),
	.w8(32'hb8d54244),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f185c),
	.w1(32'h3b0c0156),
	.w2(32'hba8bba54),
	.w3(32'h3b3c8de2),
	.w4(32'h3b262ede),
	.w5(32'h3921e8bc),
	.w6(32'h3ab34a28),
	.w7(32'h3ab56af0),
	.w8(32'h3a304528),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397aa2fe),
	.w1(32'h395408c8),
	.w2(32'hb9948556),
	.w3(32'h3999bc55),
	.w4(32'h394ea33f),
	.w5(32'hb88f54f5),
	.w6(32'h39e5b421),
	.w7(32'h39646ae4),
	.w8(32'h393b0fe2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9aed49),
	.w1(32'h3a7de604),
	.w2(32'h38b99441),
	.w3(32'hba524bf5),
	.w4(32'h38037ca2),
	.w5(32'h398c0ca1),
	.w6(32'hba34db88),
	.w7(32'hb9e5b993),
	.w8(32'hba46b248),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d1cda),
	.w1(32'h3aa059f7),
	.w2(32'h3b056c38),
	.w3(32'h3ac9a94a),
	.w4(32'h3acc7e54),
	.w5(32'h3b440780),
	.w6(32'hb9eda380),
	.w7(32'h3af35628),
	.w8(32'h3b4fc0b4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a607dee),
	.w1(32'h3a2633a0),
	.w2(32'h3a822919),
	.w3(32'h3aba34ee),
	.w4(32'h3a096f10),
	.w5(32'h3a07a1bc),
	.w6(32'h3a53346b),
	.w7(32'hba418486),
	.w8(32'hb93e3029),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e6ebd),
	.w1(32'h39d71231),
	.w2(32'hbab2306c),
	.w3(32'hba18c3f6),
	.w4(32'hbadd50c5),
	.w5(32'hba87b939),
	.w6(32'h3b259c88),
	.w7(32'h3a1e1790),
	.w8(32'hb9f4d369),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d2037),
	.w1(32'h38669f6b),
	.w2(32'hb957d0cf),
	.w3(32'hb7beba0b),
	.w4(32'hbadb1355),
	.w5(32'hba9b0c23),
	.w6(32'hba3b67d4),
	.w7(32'hbb005497),
	.w8(32'hba763c3c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1225c1),
	.w1(32'h3b115ad5),
	.w2(32'h3a5a1869),
	.w3(32'hbb1e17b8),
	.w4(32'h3a51d90d),
	.w5(32'h3b8d8c9d),
	.w6(32'hb9f823e4),
	.w7(32'hb9510271),
	.w8(32'h3b6de3d5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64f6b5),
	.w1(32'hbae30a0f),
	.w2(32'hb9877aba),
	.w3(32'hb9acf315),
	.w4(32'hbb44bbbf),
	.w5(32'hbaa4aa42),
	.w6(32'hbac2f3e6),
	.w7(32'hba62e8c8),
	.w8(32'hb9ecf8a9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c6d5f),
	.w1(32'h3a161e60),
	.w2(32'h3a97223f),
	.w3(32'h39f72df7),
	.w4(32'h3a6aa74d),
	.w5(32'h3a9d8c2e),
	.w6(32'h3abad7df),
	.w7(32'h3a0e1d5a),
	.w8(32'h39fba7cc),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b9381),
	.w1(32'h39b6ced9),
	.w2(32'h3a304e6e),
	.w3(32'h3980c4c2),
	.w4(32'h39f14c69),
	.w5(32'h3a3fff9f),
	.w6(32'h398e3448),
	.w7(32'h3a1c8d61),
	.w8(32'h3a4c6e08),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ba2ec),
	.w1(32'h390fa6d8),
	.w2(32'h39adee3c),
	.w3(32'h3aa8abd9),
	.w4(32'h36841708),
	.w5(32'h3a08b6ce),
	.w6(32'h3a1f4598),
	.w7(32'h3a02be0c),
	.w8(32'h39ede927),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a213445),
	.w1(32'h39e75a4b),
	.w2(32'h3a225856),
	.w3(32'h3a2ca73e),
	.w4(32'h39ddabde),
	.w5(32'h3a232778),
	.w6(32'h39f36157),
	.w7(32'h3a2f9922),
	.w8(32'h3a2c4156),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42dc1f),
	.w1(32'h3a94cb54),
	.w2(32'h3a92cd0c),
	.w3(32'h3a9930e7),
	.w4(32'h3a3e2502),
	.w5(32'h3a7ce1b0),
	.w6(32'h39b9292d),
	.w7(32'h3a23bc4a),
	.w8(32'h39363af8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b3c1e6),
	.w1(32'h3a84ac86),
	.w2(32'h3aab6ec3),
	.w3(32'h39eaf93a),
	.w4(32'h3a3e3b52),
	.w5(32'h3aef2bd4),
	.w6(32'h3a092bf5),
	.w7(32'h3920327c),
	.w8(32'h3ad103b3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f78325),
	.w1(32'h399e8656),
	.w2(32'hba357912),
	.w3(32'h3a373900),
	.w4(32'h3a5f4d89),
	.w5(32'h399fd498),
	.w6(32'h3aa69113),
	.w7(32'h3aa3d3b5),
	.w8(32'h3a0afee8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba732318),
	.w1(32'hbb340d5b),
	.w2(32'hba51d367),
	.w3(32'h3a33aa81),
	.w4(32'hb99ce107),
	.w5(32'h3a01b8b4),
	.w6(32'hbaeec49d),
	.w7(32'h398cd1b1),
	.w8(32'h3ac57dd7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae71b08),
	.w1(32'h3b9d5652),
	.w2(32'h3b103fee),
	.w3(32'h3b138ed1),
	.w4(32'h39454326),
	.w5(32'hba253796),
	.w6(32'h3b3aa639),
	.w7(32'hbb00d1e0),
	.w8(32'hbb052889),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a152719),
	.w1(32'hb7f118fe),
	.w2(32'h3805c387),
	.w3(32'h3a2159e5),
	.w4(32'hb9b6f675),
	.w5(32'hb9b0fe30),
	.w6(32'h39c8ec08),
	.w7(32'h388a2c30),
	.w8(32'hb9d31bbf),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9668697),
	.w1(32'h3a15205a),
	.w2(32'h3a668d7c),
	.w3(32'hb830d338),
	.w4(32'h3a2dc0b9),
	.w5(32'h3a668d8a),
	.w6(32'h3a4fa198),
	.w7(32'h3a8caf72),
	.w8(32'h3a584313),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9df3d3),
	.w1(32'h397f55c7),
	.w2(32'h39c72a64),
	.w3(32'h3a98c126),
	.w4(32'h3986b92e),
	.w5(32'h39e6d157),
	.w6(32'h396b8322),
	.w7(32'h39cd5dc8),
	.w8(32'h3987d20d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d9e5b),
	.w1(32'hba05a764),
	.w2(32'h3a8c0dec),
	.w3(32'h3a858f16),
	.w4(32'h392024bc),
	.w5(32'hbb147f01),
	.w6(32'h3abc1cc9),
	.w7(32'h3ae0803c),
	.w8(32'h3b4ccd9d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79c57f),
	.w1(32'h3b849f39),
	.w2(32'h3c2d5532),
	.w3(32'h3b15cf11),
	.w4(32'h3b0b96a5),
	.w5(32'h3bfbc856),
	.w6(32'hbaf88879),
	.w7(32'h3ab2d6cb),
	.w8(32'h3a0fed21),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ba7f9),
	.w1(32'hbb7ef24d),
	.w2(32'hbc0ceb29),
	.w3(32'hbadeb11c),
	.w4(32'hbb91cad2),
	.w5(32'hbacfdf72),
	.w6(32'hb8bc7129),
	.w7(32'hbc13d5fb),
	.w8(32'h3bcaef18),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b612298),
	.w1(32'hbafd4479),
	.w2(32'hbae28e87),
	.w3(32'hbc813e33),
	.w4(32'hbb364afa),
	.w5(32'h3a120ed1),
	.w6(32'hba33565f),
	.w7(32'hba996dbb),
	.w8(32'hbb0231a4),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad8bfd),
	.w1(32'hbb4f6d9f),
	.w2(32'hbadf3436),
	.w3(32'hbb0dc6cd),
	.w4(32'h3a088f35),
	.w5(32'hba811105),
	.w6(32'hb88e17ef),
	.w7(32'h3a417b33),
	.w8(32'h3b67077b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd4f88),
	.w1(32'h3b54eb84),
	.w2(32'h3c35b101),
	.w3(32'hba50eb9b),
	.w4(32'h38d62af0),
	.w5(32'hbaa77b0a),
	.w6(32'h3c146db9),
	.w7(32'h3bcd91ee),
	.w8(32'hbc4c70c0),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12dfc0),
	.w1(32'hbc114b71),
	.w2(32'h3c50cd20),
	.w3(32'h3b3004c4),
	.w4(32'h3b596995),
	.w5(32'h3c15516d),
	.w6(32'h3b91819e),
	.w7(32'h3be356c6),
	.w8(32'hbb3c1097),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7b5ba),
	.w1(32'h3c5d403a),
	.w2(32'h3c818153),
	.w3(32'h3c27ebaa),
	.w4(32'h3c612126),
	.w5(32'h3c4d9ca4),
	.w6(32'h3c728343),
	.w7(32'h3bf650f3),
	.w8(32'hbb77a901),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdac218),
	.w1(32'hbc243229),
	.w2(32'hbb3afc25),
	.w3(32'hbb0d6b85),
	.w4(32'hbb42948a),
	.w5(32'h3b50da8e),
	.w6(32'hbb21a091),
	.w7(32'h3aff84b6),
	.w8(32'h3bd47861),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2779c3),
	.w1(32'hbb89cfc0),
	.w2(32'h3ab2efb2),
	.w3(32'h3b8b3d0d),
	.w4(32'hbb66ea80),
	.w5(32'hbb253863),
	.w6(32'hbb8cbe97),
	.w7(32'hbb3c0f87),
	.w8(32'hba450cc9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f3df63),
	.w1(32'hb8a80b84),
	.w2(32'hbae62560),
	.w3(32'h3ae439a1),
	.w4(32'hbb22aab2),
	.w5(32'hbb5fa8f2),
	.w6(32'hba0a4ab4),
	.w7(32'hbb06a1f9),
	.w8(32'h398c194b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb292d3c),
	.w1(32'hba9330eb),
	.w2(32'hbbdb8c8f),
	.w3(32'h3a940a13),
	.w4(32'hbadcb177),
	.w5(32'hbb51ebb1),
	.w6(32'hb96c10ca),
	.w7(32'h38b96b19),
	.w8(32'hb98060c5),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ec93d),
	.w1(32'hbb08ea8f),
	.w2(32'h3b5ae356),
	.w3(32'hbbe62635),
	.w4(32'hbbfba3ab),
	.w5(32'hbadd46e6),
	.w6(32'h3b0ebb05),
	.w7(32'h3b5987d3),
	.w8(32'hba25bf62),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09450d),
	.w1(32'hbc0f0a67),
	.w2(32'hba452b85),
	.w3(32'h3b6e9c5f),
	.w4(32'hbbcf5506),
	.w5(32'hbbd8ebb1),
	.w6(32'hbbd93041),
	.w7(32'h3bdbc9ae),
	.w8(32'hbb07402d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2be3f1),
	.w1(32'hbac83f3b),
	.w2(32'h3a9ae482),
	.w3(32'h3c372c36),
	.w4(32'h38d46b2e),
	.w5(32'h3ae42e2e),
	.w6(32'hba7d3823),
	.w7(32'hbaf3f1bd),
	.w8(32'h3bbd06e9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1214a6),
	.w1(32'hbcc68059),
	.w2(32'hbc6c4a3c),
	.w3(32'h3b8079df),
	.w4(32'hbcbac4c9),
	.w5(32'hbc6dc56b),
	.w6(32'hbc84b550),
	.w7(32'hbc123d0b),
	.w8(32'h3c2c16b9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6927de),
	.w1(32'hbcb0aaec),
	.w2(32'h3cabf394),
	.w3(32'h3c6a7a58),
	.w4(32'hbca24df4),
	.w5(32'hbc56043d),
	.w6(32'h3a0ede21),
	.w7(32'h3c9a3032),
	.w8(32'hbc8b7f77),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1be482),
	.w1(32'hbaa0756c),
	.w2(32'h3b429355),
	.w3(32'h3caf178f),
	.w4(32'hba416346),
	.w5(32'h39aac42a),
	.w6(32'h39ce12f1),
	.w7(32'h3aef81c8),
	.w8(32'hbb47902a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ff00f),
	.w1(32'h3a57df35),
	.w2(32'h3b229713),
	.w3(32'h3804bc28),
	.w4(32'h3b545c8a),
	.w5(32'hbb89caef),
	.w6(32'hbad2fde2),
	.w7(32'hbb54933f),
	.w8(32'h3a6eb57c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f9e10),
	.w1(32'h3bad3726),
	.w2(32'h3b168f9b),
	.w3(32'hba92bd1b),
	.w4(32'h3a6935f5),
	.w5(32'h3b6c0071),
	.w6(32'h3bae1f76),
	.w7(32'h3bf17ecc),
	.w8(32'h3b6d93f7),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be832f3),
	.w1(32'hbb1bb522),
	.w2(32'hbab0629c),
	.w3(32'hb9ea22f2),
	.w4(32'hbbe81ae9),
	.w5(32'hbb5ac750),
	.w6(32'hbb03f5e1),
	.w7(32'hbb650d1b),
	.w8(32'hbb6179c4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30af41),
	.w1(32'h3a645bc6),
	.w2(32'h3951cd40),
	.w3(32'hb8191d80),
	.w4(32'h39b1f316),
	.w5(32'hbaddd67a),
	.w6(32'h3aea2c8d),
	.w7(32'hba721219),
	.w8(32'h3a26f42d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed9a00),
	.w1(32'hbb5372ab),
	.w2(32'hbbc6d53e),
	.w3(32'h3a2a2e16),
	.w4(32'hba7dbd2e),
	.w5(32'hbb55da0e),
	.w6(32'hbb75b12a),
	.w7(32'hbb05db9e),
	.w8(32'hbadd5c80),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb740334),
	.w1(32'hbcc48c5b),
	.w2(32'hbc8251ad),
	.w3(32'h3b13dc41),
	.w4(32'hbb1e2e96),
	.w5(32'h3c2f16e9),
	.w6(32'hbc780035),
	.w7(32'hbc867a1f),
	.w8(32'h3ca675ae),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4187e4),
	.w1(32'hbacae7d7),
	.w2(32'hbb44e590),
	.w3(32'hbc170490),
	.w4(32'hbb80f9dd),
	.w5(32'hbb27a895),
	.w6(32'hbafe7cd7),
	.w7(32'hbb8d6461),
	.w8(32'hba91cf81),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb7af7),
	.w1(32'hbc0d9126),
	.w2(32'hbb45d84d),
	.w3(32'h3b1177a1),
	.w4(32'hbbd6c259),
	.w5(32'hbb9d5bf7),
	.w6(32'hbbde95fb),
	.w7(32'hbb6a88d3),
	.w8(32'hbae5f5a8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaf982),
	.w1(32'h3b127ab8),
	.w2(32'h3b53af27),
	.w3(32'hba64d7e6),
	.w4(32'hbc23daa9),
	.w5(32'h3ac41c2a),
	.w6(32'h3b5d78b5),
	.w7(32'h3b374341),
	.w8(32'hbc201b9c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c7d7f),
	.w1(32'hbabf24b3),
	.w2(32'hb91faaa9),
	.w3(32'hbaf0151e),
	.w4(32'hb8ebf162),
	.w5(32'hbbf30fc7),
	.w6(32'h3b4e972e),
	.w7(32'h3b9d60e0),
	.w8(32'hbb97f3f8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b815c91),
	.w1(32'hb88967c3),
	.w2(32'hbb1d7a88),
	.w3(32'hbb84831a),
	.w4(32'hba9856f7),
	.w5(32'hbb8c0379),
	.w6(32'h37d6dcc5),
	.w7(32'hbaf6e597),
	.w8(32'h39b82c7e),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba913063),
	.w1(32'h3c0a21aa),
	.w2(32'h3b3a7e67),
	.w3(32'hba0658dc),
	.w4(32'h3a8faf0c),
	.w5(32'h38c6de3a),
	.w6(32'h3b6cb407),
	.w7(32'hbb8304ce),
	.w8(32'hbc5b82e2),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc123a49),
	.w1(32'h3b9c77f8),
	.w2(32'hbc07ab02),
	.w3(32'hbc23573c),
	.w4(32'h3b7b40bd),
	.w5(32'hbc265469),
	.w6(32'h3bd7c7df),
	.w7(32'hbc1b7d77),
	.w8(32'hbb632578),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2da893),
	.w1(32'hbad950f1),
	.w2(32'h3a4d4db5),
	.w3(32'hbb030ca5),
	.w4(32'hbb58af69),
	.w5(32'hba072538),
	.w6(32'h38ed350d),
	.w7(32'h3a153b54),
	.w8(32'h3ad072ba),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff50ee),
	.w1(32'hbb6180dd),
	.w2(32'hbb9e90fc),
	.w3(32'hba5a9685),
	.w4(32'hbabcfc0e),
	.w5(32'hbb86b808),
	.w6(32'hbb33d42e),
	.w7(32'hbb55f2aa),
	.w8(32'h3a0674df),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8993a),
	.w1(32'hba4a6b97),
	.w2(32'h39c0ae24),
	.w3(32'hb9ea7140),
	.w4(32'h3a60e481),
	.w5(32'hbab57267),
	.w6(32'hba0ce104),
	.w7(32'hba0a058b),
	.w8(32'hb7e62d38),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17a1b6),
	.w1(32'hbc0f54f1),
	.w2(32'h3aa30027),
	.w3(32'hba108f01),
	.w4(32'hbc1acaa6),
	.w5(32'hbbb9dc9e),
	.w6(32'hbbbdc401),
	.w7(32'hbc40b2c0),
	.w8(32'hba99c765),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff9a4f),
	.w1(32'hbaf6f093),
	.w2(32'h3bbed405),
	.w3(32'h3a3537e4),
	.w4(32'hbaa7b001),
	.w5(32'hbc378d7e),
	.w6(32'hbbc8fb6b),
	.w7(32'hbb529b58),
	.w8(32'h3bb67ebc),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c681fd3),
	.w1(32'h3bb68301),
	.w2(32'hbc04fa5e),
	.w3(32'h3bab9c27),
	.w4(32'h3af2c472),
	.w5(32'hbb10a58c),
	.w6(32'h3b048cf5),
	.w7(32'hbb1092e5),
	.w8(32'hbbf0e065),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6cd9d),
	.w1(32'hba936e91),
	.w2(32'hba9d325f),
	.w3(32'hbc1a5719),
	.w4(32'hbb0440e4),
	.w5(32'hbb55ab7f),
	.w6(32'hbb36f9bd),
	.w7(32'hba91a22f),
	.w8(32'hbab0e169),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ed00e),
	.w1(32'h3bbce5df),
	.w2(32'h3c1f7e45),
	.w3(32'h3b77f3bd),
	.w4(32'h3b14c576),
	.w5(32'h3b52d601),
	.w6(32'h3bafa4c7),
	.w7(32'h3bb843bd),
	.w8(32'hbbcc5f1d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3738e0),
	.w1(32'hbb37a242),
	.w2(32'hba476922),
	.w3(32'hbb33f04b),
	.w4(32'hba6d2966),
	.w5(32'h3a9e68c7),
	.w6(32'h3956c7db),
	.w7(32'h3ae99c75),
	.w8(32'h3aef4f41),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2699d),
	.w1(32'hb9c32736),
	.w2(32'h3b252cef),
	.w3(32'h3ad92f30),
	.w4(32'hb9cc592d),
	.w5(32'hba889cae),
	.w6(32'h3add90b3),
	.w7(32'h3ab597f7),
	.w8(32'hbb675045),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb917927),
	.w1(32'hbbf4f38d),
	.w2(32'hbb3929e5),
	.w3(32'hbb01652e),
	.w4(32'hbbe90824),
	.w5(32'hbbcb6b36),
	.w6(32'hbb4f6dd8),
	.w7(32'hbae8e1c0),
	.w8(32'hbb0fc2ea),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b54576),
	.w1(32'hbbbb9ff5),
	.w2(32'hb9134e39),
	.w3(32'hbbc60ee0),
	.w4(32'hbb34f19c),
	.w5(32'h3b774d92),
	.w6(32'hbc00c8e9),
	.w7(32'hb9b014a3),
	.w8(32'h3b968a66),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92ab54),
	.w1(32'hbb6eaa08),
	.w2(32'hb97a58a4),
	.w3(32'h3ae1f290),
	.w4(32'hbbdd982d),
	.w5(32'hbbfaeb18),
	.w6(32'hbab2858e),
	.w7(32'h3b70cd40),
	.w8(32'hbb24eb84),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28563c),
	.w1(32'h3a651c3e),
	.w2(32'h3a5dc82b),
	.w3(32'h3b523219),
	.w4(32'h3a7a2dfa),
	.w5(32'hbb18f5c5),
	.w6(32'h3b525f85),
	.w7(32'hbaa39ef1),
	.w8(32'hbb039c01),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8653b7d),
	.w1(32'hba22be56),
	.w2(32'hbb958da2),
	.w3(32'hba577787),
	.w4(32'hbbbcb65f),
	.w5(32'hbb96a7e2),
	.w6(32'hbb2d3fcb),
	.w7(32'hba986f97),
	.w8(32'h3ac1b100),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22b7e9),
	.w1(32'hbd00ac6d),
	.w2(32'hbccf2c37),
	.w3(32'hbb27a490),
	.w4(32'hbcd00b8a),
	.w5(32'hbc5178c8),
	.w6(32'hbc9258c8),
	.w7(32'hbc2fb7d6),
	.w8(32'h3c9e84a2),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c942a9c),
	.w1(32'hbc64837e),
	.w2(32'hbc07bdd7),
	.w3(32'h3c14db01),
	.w4(32'hbb870609),
	.w5(32'h3a9ac95e),
	.w6(32'hbbf50c51),
	.w7(32'hbba6e1a4),
	.w8(32'h3c868ac5),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbcd8c0),
	.w1(32'hbc6c7b4c),
	.w2(32'hbba8a158),
	.w3(32'h3bdd511e),
	.w4(32'h3b6584d6),
	.w5(32'hbc18dd70),
	.w6(32'hbc5d069c),
	.w7(32'h3b2519b6),
	.w8(32'hbad7a45b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf895fa),
	.w1(32'h39e546ba),
	.w2(32'hbb88a4bf),
	.w3(32'h3c8e1033),
	.w4(32'hb94fbccb),
	.w5(32'hbb87e363),
	.w6(32'h3abccde0),
	.w7(32'hbb48678e),
	.w8(32'hba8ac6c6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4302e),
	.w1(32'h3a3546d9),
	.w2(32'h3b619fdb),
	.w3(32'hbb4cf6d7),
	.w4(32'h39a23615),
	.w5(32'hba457965),
	.w6(32'h3adf489a),
	.w7(32'h38aa6c02),
	.w8(32'h3a84648a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b80da),
	.w1(32'hbc2ae151),
	.w2(32'hbb5734ac),
	.w3(32'h3a18eb4c),
	.w4(32'hbc0a2297),
	.w5(32'hbbb03696),
	.w6(32'hbc0dc8e2),
	.w7(32'hbb85b072),
	.w8(32'h39ba8f26),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e3f79),
	.w1(32'hbc85edb5),
	.w2(32'hbc1a5a56),
	.w3(32'h3b2efa55),
	.w4(32'hbc7cf128),
	.w5(32'hbbf26bcd),
	.w6(32'hbc3f02ed),
	.w7(32'h3aaf94d8),
	.w8(32'h3c517b1e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cafbdb5),
	.w1(32'hba8e5996),
	.w2(32'hbb349a2b),
	.w3(32'h3c5baa59),
	.w4(32'hbc1cdcfe),
	.w5(32'hbc278d8c),
	.w6(32'hbb57e5f8),
	.w7(32'hbbf91470),
	.w8(32'hbc59a3ae),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86c234),
	.w1(32'h39c6e998),
	.w2(32'h3bec316b),
	.w3(32'h3bde7e31),
	.w4(32'hbb063a2f),
	.w5(32'h3b80c870),
	.w6(32'h3ae91cbd),
	.w7(32'h3b775810),
	.w8(32'hbbbd22ed),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4cd3e),
	.w1(32'hbbd77afe),
	.w2(32'h3c72c19e),
	.w3(32'hbac99a0b),
	.w4(32'h3c048758),
	.w5(32'h3c006eb4),
	.w6(32'h39dcff12),
	.w7(32'h3ba1a2f5),
	.w8(32'hbc1eeb32),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc556ef1),
	.w1(32'hba4d60e3),
	.w2(32'hbadae253),
	.w3(32'hbc2f4d78),
	.w4(32'hbb49167f),
	.w5(32'hbb07b4e5),
	.w6(32'hba0a151f),
	.w7(32'hbad1201f),
	.w8(32'hbba489a9),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb133327),
	.w1(32'hba19cf55),
	.w2(32'hbb383673),
	.w3(32'hbabffe56),
	.w4(32'hbb1d92f9),
	.w5(32'hb97a3c9f),
	.w6(32'hb9c56db9),
	.w7(32'hba5e809b),
	.w8(32'hbaf7d161),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae79bd),
	.w1(32'h39d12168),
	.w2(32'hbc2d6c5b),
	.w3(32'h3b374db5),
	.w4(32'h3b013c4c),
	.w5(32'hbae37f0d),
	.w6(32'h3a8fd969),
	.w7(32'h3a35032c),
	.w8(32'h3c2b7676),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8293d8),
	.w1(32'hbcbdccdb),
	.w2(32'h3c136b52),
	.w3(32'h3bf4d96b),
	.w4(32'hbb4e904c),
	.w5(32'h3b34711c),
	.w6(32'hbbef6218),
	.w7(32'h3ba90745),
	.w8(32'h3c5a8deb),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1b3a6),
	.w1(32'hbbecdef1),
	.w2(32'hbbc9e84f),
	.w3(32'h3ca468c9),
	.w4(32'hbbf917b7),
	.w5(32'hbb706d61),
	.w6(32'hbb620c8b),
	.w7(32'hba816172),
	.w8(32'h390eda08),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25d2ac),
	.w1(32'hbb9cb4f3),
	.w2(32'hbad3abdd),
	.w3(32'h39bbf2db),
	.w4(32'hb98f58f3),
	.w5(32'hb9378b88),
	.w6(32'hbb92947e),
	.w7(32'h3953248f),
	.w8(32'h389369ec),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0cad0),
	.w1(32'hbb8fdc21),
	.w2(32'hbb0c4d8b),
	.w3(32'hb99da141),
	.w4(32'hbbedf568),
	.w5(32'hbba6ef5b),
	.w6(32'h3a26c2ff),
	.w7(32'h3a5fc7ec),
	.w8(32'h3b3993a5),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8023b6),
	.w1(32'hbc193204),
	.w2(32'hbbba0fdb),
	.w3(32'hb9a0444d),
	.w4(32'hbbdaaa33),
	.w5(32'hbbbd4a89),
	.w6(32'hbb9f7087),
	.w7(32'hbbce02ba),
	.w8(32'h3b677c81),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba87df4),
	.w1(32'hbc411fba),
	.w2(32'h3b8c382c),
	.w3(32'hbb054f2f),
	.w4(32'hbc0de7b0),
	.w5(32'hbbbe16ee),
	.w6(32'hbc104414),
	.w7(32'hbc2ada3d),
	.w8(32'h3c22f85f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5f34b),
	.w1(32'h3a20cfe1),
	.w2(32'hbb3b9171),
	.w3(32'h3c2f07e9),
	.w4(32'hbb107689),
	.w5(32'hbb1b5e56),
	.w6(32'hba8ffb68),
	.w7(32'hbaa4b918),
	.w8(32'hba87a79a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b121684),
	.w1(32'hba4c6bbb),
	.w2(32'h3b908c19),
	.w3(32'hbb80edc1),
	.w4(32'hbaf2efe2),
	.w5(32'h3ae6a1c4),
	.w6(32'h3b560740),
	.w7(32'h3a3d099e),
	.w8(32'h3b2e5adb),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a9cf9),
	.w1(32'hbcb4e5ab),
	.w2(32'h3bfc262b),
	.w3(32'h3a9f60e0),
	.w4(32'hbbe0a4c4),
	.w5(32'h3bf14e12),
	.w6(32'hbc2f2fe9),
	.w7(32'hbab1c82b),
	.w8(32'h3c9e739a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05132c),
	.w1(32'hbb3cfaa8),
	.w2(32'h39fcb06f),
	.w3(32'h3ca836d1),
	.w4(32'h3a9f4425),
	.w5(32'h3aa4a47a),
	.w6(32'h39a13fb5),
	.w7(32'h3ac94a74),
	.w8(32'hbb245463),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e8b47),
	.w1(32'hbb2aba16),
	.w2(32'hbb4cabc1),
	.w3(32'hbb747fd5),
	.w4(32'hbb0dce59),
	.w5(32'hbab041a2),
	.w6(32'hbb168250),
	.w7(32'hbb827c8f),
	.w8(32'h3a71575f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a677b),
	.w1(32'hbb1daff9),
	.w2(32'h3b590acc),
	.w3(32'h3b0a5d7c),
	.w4(32'h3a3faec5),
	.w5(32'h3b026be7),
	.w6(32'hbb190f69),
	.w7(32'h3afb00d5),
	.w8(32'hbbb116a2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb482d20),
	.w1(32'hbc8ce4f4),
	.w2(32'h3b9895a6),
	.w3(32'h3b286749),
	.w4(32'hbbeea4b9),
	.w5(32'h3ba77940),
	.w6(32'hbc284f33),
	.w7(32'h3c49a588),
	.w8(32'h3cce4460),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d17a48a),
	.w1(32'h3b24d772),
	.w2(32'hbb974d46),
	.w3(32'h3cce9081),
	.w4(32'h394deb66),
	.w5(32'hbaaba739),
	.w6(32'h3b444e0a),
	.w7(32'h3a50b65c),
	.w8(32'hbb2db82b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4ef4a),
	.w1(32'hbb302f24),
	.w2(32'hb9ccaf35),
	.w3(32'hbb45c3d9),
	.w4(32'hbae097bd),
	.w5(32'hba8ea749),
	.w6(32'hbb2aa609),
	.w7(32'hbb077663),
	.w8(32'hba89c44e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a4c8f),
	.w1(32'hbb105944),
	.w2(32'hb9f33ef8),
	.w3(32'h3b18dfe8),
	.w4(32'hbacc298e),
	.w5(32'hbb14773e),
	.w6(32'h3a27ad8f),
	.w7(32'h3aa49269),
	.w8(32'hbb61aa7d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb804f4f),
	.w1(32'hbb0c1467),
	.w2(32'hbae4077c),
	.w3(32'hbabc896d),
	.w4(32'hba3a2d17),
	.w5(32'hbb29edb3),
	.w6(32'hbb4360b0),
	.w7(32'hbb358f88),
	.w8(32'hbb73d1b9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a08cd),
	.w1(32'hbacd7437),
	.w2(32'hbb2c9592),
	.w3(32'hba452e67),
	.w4(32'hbbbd7305),
	.w5(32'hbb20eb90),
	.w6(32'hbb48f562),
	.w7(32'hb94a0b30),
	.w8(32'hbb95aed5),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb333f5f),
	.w1(32'hbc3b3af2),
	.w2(32'hbb1992b2),
	.w3(32'hb92f339d),
	.w4(32'hbc9efa2c),
	.w5(32'hbc388354),
	.w6(32'hbbc016a4),
	.w7(32'hbb587bf2),
	.w8(32'h39fcb469),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73a20f),
	.w1(32'hbb8c3e06),
	.w2(32'h3b2fcaad),
	.w3(32'h3cef3f6d),
	.w4(32'hbb0dd0c8),
	.w5(32'hba35033e),
	.w6(32'hbb6ea73f),
	.w7(32'hbad87181),
	.w8(32'h3b80d7ef),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcc309),
	.w1(32'hbb8146b6),
	.w2(32'hbbe71f01),
	.w3(32'h3bb9269a),
	.w4(32'hbbe2c457),
	.w5(32'hbba7f9c2),
	.w6(32'hbba95fde),
	.w7(32'hbbbaeff3),
	.w8(32'h3bb53f71),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b995c),
	.w1(32'h3bbcabe7),
	.w2(32'h3a815bf3),
	.w3(32'h3b42fafe),
	.w4(32'h38c86e54),
	.w5(32'hba8b9afa),
	.w6(32'h3bb90845),
	.w7(32'hbad704a1),
	.w8(32'hbc0260d9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88213e),
	.w1(32'hbb78f493),
	.w2(32'hbb96f9f6),
	.w3(32'hba43f1a3),
	.w4(32'hbb2d710f),
	.w5(32'hbb9cb736),
	.w6(32'hbb6c27e7),
	.w7(32'hbb5919f2),
	.w8(32'h3928546c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dcaad),
	.w1(32'hbab181f3),
	.w2(32'hbb2452a7),
	.w3(32'h38ed426e),
	.w4(32'hba4c565c),
	.w5(32'hba48bfc5),
	.w6(32'hbb8fcd8f),
	.w7(32'hbb79f26a),
	.w8(32'hbb158ce3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd48b5),
	.w1(32'hbbe984dd),
	.w2(32'hbbdaff6b),
	.w3(32'hbb28389a),
	.w4(32'hbc12876f),
	.w5(32'hbb735511),
	.w6(32'hbbaf65e9),
	.w7(32'hbb70d6ff),
	.w8(32'h3a4c38fd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c7873),
	.w1(32'h3b381f6f),
	.w2(32'h3b014fce),
	.w3(32'hba2cc124),
	.w4(32'hbb84f7cb),
	.w5(32'hbb36e2f0),
	.w6(32'h3aa61fe1),
	.w7(32'h3addc208),
	.w8(32'hbb4f2359),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba024e6e),
	.w1(32'hbbc45567),
	.w2(32'hbbb6228f),
	.w3(32'h3a789a80),
	.w4(32'hbbb91379),
	.w5(32'h3a7bf1e0),
	.w6(32'hbbaa6c3d),
	.w7(32'hbbb309bd),
	.w8(32'h3b8eb00f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5b0f8),
	.w1(32'hbb81a2c4),
	.w2(32'h3ad2d524),
	.w3(32'hbbb9b527),
	.w4(32'hba8429d8),
	.w5(32'h3ba78f9a),
	.w6(32'hbbc918b7),
	.w7(32'hbaa792f6),
	.w8(32'hbaacb198),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb05016),
	.w1(32'h3b1ab48c),
	.w2(32'h3a3be8e3),
	.w3(32'hbb1367c9),
	.w4(32'h3b6d314a),
	.w5(32'h3be14cf3),
	.w6(32'h3b13f386),
	.w7(32'h3b38a4c7),
	.w8(32'h3baab8b2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ab042),
	.w1(32'hbc917b12),
	.w2(32'hbc2c69f6),
	.w3(32'h3c38ef29),
	.w4(32'hbc822303),
	.w5(32'hbc3793a9),
	.w6(32'hbc3c2fa1),
	.w7(32'h3b31b81a),
	.w8(32'h3c4d5519),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c019ee1),
	.w1(32'hbacc7615),
	.w2(32'hbb7d2a54),
	.w3(32'h3b9a5816),
	.w4(32'hba45a8cf),
	.w5(32'hbb422a61),
	.w6(32'hbb12ea66),
	.w7(32'hbb2ae516),
	.w8(32'hba7e5b85),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14d34d),
	.w1(32'hbb864678),
	.w2(32'hbb4bcff2),
	.w3(32'hba206469),
	.w4(32'hbbc1397d),
	.w5(32'hbb5aa017),
	.w6(32'hbb73b0fb),
	.w7(32'hbb4b4e07),
	.w8(32'hbbbe6df0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6695e6),
	.w1(32'hbb54a3bd),
	.w2(32'hbb992df3),
	.w3(32'hbbab9876),
	.w4(32'hbaac5d70),
	.w5(32'hba8b6645),
	.w6(32'hbc16c18c),
	.w7(32'hbbc16bf5),
	.w8(32'h3b3f4b6e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb844d55),
	.w1(32'hbbdc1172),
	.w2(32'hbb8b524d),
	.w3(32'hbb011208),
	.w4(32'hbb061b77),
	.w5(32'hbaac899f),
	.w6(32'hbb9c1e58),
	.w7(32'hba8488db),
	.w8(32'h3b2ca1bf),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa35878),
	.w1(32'hbbfdc4bc),
	.w2(32'hbbe2186b),
	.w3(32'hbad9fdd6),
	.w4(32'hbbb50d1c),
	.w5(32'h3a6e8f91),
	.w6(32'hbbf64a03),
	.w7(32'hbad5b92c),
	.w8(32'h3c2b23da),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25758a),
	.w1(32'h3af83664),
	.w2(32'hbb8d27f7),
	.w3(32'h3be78453),
	.w4(32'hbb313fdb),
	.w5(32'hba964a75),
	.w6(32'hbb3dbbaf),
	.w7(32'hbb9fffae),
	.w8(32'hbc1d9f22),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fd2b3),
	.w1(32'h39316d37),
	.w2(32'hbbd3ea93),
	.w3(32'hbc2e8548),
	.w4(32'hbae90c1f),
	.w5(32'hbbbf39d1),
	.w6(32'hba282e7a),
	.w7(32'hbbc77705),
	.w8(32'hbb313eb4),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83c395),
	.w1(32'hbba44064),
	.w2(32'hbaf794f7),
	.w3(32'hba3927c6),
	.w4(32'hbb33f919),
	.w5(32'hbb0d3714),
	.w6(32'hb9e723c5),
	.w7(32'hb5b3edda),
	.w8(32'h3ac34655),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50a917),
	.w1(32'hbbef6619),
	.w2(32'h3bca1d26),
	.w3(32'hbaf32e6a),
	.w4(32'h3b111fd1),
	.w5(32'h3c3071ed),
	.w6(32'hbb37607c),
	.w7(32'h3845f6e4),
	.w8(32'h3b3fecb2),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7ac85),
	.w1(32'hba3b8315),
	.w2(32'h3a993cc2),
	.w3(32'hbc8dc286),
	.w4(32'hbad5230e),
	.w5(32'h3af00686),
	.w6(32'hbb386276),
	.w7(32'h3a2643bf),
	.w8(32'hb9fd1055),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc053972),
	.w1(32'hbb242eb0),
	.w2(32'h3c8140fb),
	.w3(32'hbbb9c304),
	.w4(32'h3aa5b20c),
	.w5(32'h3b918a79),
	.w6(32'h39ade8db),
	.w7(32'h3b20aadd),
	.w8(32'hbc1a3c05),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb976194),
	.w1(32'hbc34d76c),
	.w2(32'hbc06df3f),
	.w3(32'hbb2f8beb),
	.w4(32'hbc469c68),
	.w5(32'hbbcd4870),
	.w6(32'hbc157745),
	.w7(32'hbba147d1),
	.w8(32'hbaa07745),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90efd1),
	.w1(32'h3b902871),
	.w2(32'h3b9b956a),
	.w3(32'hbb9ee498),
	.w4(32'hb78bae54),
	.w5(32'h3ba4a8de),
	.w6(32'hbb85a92c),
	.w7(32'h3945280d),
	.w8(32'hbc2d3c70),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4de5f3),
	.w1(32'hbc95c76c),
	.w2(32'hbc938fbf),
	.w3(32'hbbf5c30a),
	.w4(32'hbbc4ad27),
	.w5(32'hbcd1db1a),
	.w6(32'h3a2f2e59),
	.w7(32'hbc9c1522),
	.w8(32'hbb6d3cd3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c854529),
	.w1(32'hbbe34e13),
	.w2(32'hba4771fc),
	.w3(32'h3ace3a89),
	.w4(32'h3bb4a28f),
	.w5(32'h3c4d3462),
	.w6(32'h3b8d415e),
	.w7(32'hbbe80147),
	.w8(32'h3cb6f45d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd75d32),
	.w1(32'hbc8096d3),
	.w2(32'h3a88b02d),
	.w3(32'h3b168762),
	.w4(32'hbba6adc8),
	.w5(32'h3a949f57),
	.w6(32'hbc5fb1ba),
	.w7(32'hbba746f3),
	.w8(32'h3c2f27f2),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36345e),
	.w1(32'hbb27e87f),
	.w2(32'h3aadb688),
	.w3(32'h3bf117ed),
	.w4(32'hba70e35b),
	.w5(32'h381ced77),
	.w6(32'hbac67efd),
	.w7(32'h39c19c3d),
	.w8(32'h3ac39642),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b878273),
	.w1(32'hbb4daaa6),
	.w2(32'h3ad58166),
	.w3(32'h3b64d8b4),
	.w4(32'hbafe10c0),
	.w5(32'hbab1b27e),
	.w6(32'hbb551d47),
	.w7(32'hbad60c3b),
	.w8(32'h3ab716d6),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5de08f),
	.w1(32'hbabc0610),
	.w2(32'hbb052ca2),
	.w3(32'h3b1d39ac),
	.w4(32'hbb2344e7),
	.w5(32'hbb8e00d7),
	.w6(32'hba78dea7),
	.w7(32'hbaef559e),
	.w8(32'h3a9b6f9c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1af427),
	.w1(32'hbb4f5a8b),
	.w2(32'hbb8867fb),
	.w3(32'h3a1c2602),
	.w4(32'hba715f73),
	.w5(32'h3961cced),
	.w6(32'h3a797a1c),
	.w7(32'hb9e3178d),
	.w8(32'h3bbec278),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa0b8a),
	.w1(32'hbb385c8a),
	.w2(32'hbbbb4208),
	.w3(32'h3a1f5e6c),
	.w4(32'hbaedda52),
	.w5(32'hbb88e908),
	.w6(32'hbb5fc786),
	.w7(32'hbb55b601),
	.w8(32'hbabd3efb),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc15bb),
	.w1(32'hbb95c18a),
	.w2(32'h3acbfd6d),
	.w3(32'hbaf11646),
	.w4(32'hbb068294),
	.w5(32'hba112eea),
	.w6(32'hbb8cc110),
	.w7(32'hba9e38dc),
	.w8(32'h3b85e13d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7eccf),
	.w1(32'hbc905971),
	.w2(32'hbc6d72e6),
	.w3(32'h3b99c291),
	.w4(32'hbc9234a6),
	.w5(32'hbc289b09),
	.w6(32'hbc2ff257),
	.w7(32'hbc01b983),
	.w8(32'h3c490554),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ea09d),
	.w1(32'h3ac664a3),
	.w2(32'h3ae3624f),
	.w3(32'h3c365faa),
	.w4(32'hba7d5982),
	.w5(32'hbab0eb07),
	.w6(32'h3af66d4c),
	.w7(32'h39e4d361),
	.w8(32'hbbcbfc06),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26d334),
	.w1(32'hbc7704f6),
	.w2(32'hbc378619),
	.w3(32'hba399fef),
	.w4(32'hbc90709e),
	.w5(32'hbc968b32),
	.w6(32'hbc5a77d7),
	.w7(32'hbc9c5119),
	.w8(32'h3c0cd46e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affb4b8),
	.w1(32'h3ab92fd7),
	.w2(32'h3bbd50b1),
	.w3(32'h3b0c52a9),
	.w4(32'h3aee272b),
	.w5(32'h3b40789b),
	.w6(32'h3b3f048d),
	.w7(32'h3b9d411e),
	.w8(32'hbbb075bd),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f39e9),
	.w1(32'hbb37a3db),
	.w2(32'hbaabdcb6),
	.w3(32'hba34e712),
	.w4(32'hbba81e6b),
	.w5(32'hbb4dbacd),
	.w6(32'h3a522199),
	.w7(32'h3b97e8ba),
	.w8(32'h3a206dd4),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1c673),
	.w1(32'hbb9cb1b8),
	.w2(32'hbb9b8f69),
	.w3(32'h3b2591ae),
	.w4(32'hbbb8a849),
	.w5(32'hbb49324e),
	.w6(32'hbbde9c66),
	.w7(32'hbbd98c50),
	.w8(32'h3b81eeb3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb06dc),
	.w1(32'hbbb997a6),
	.w2(32'h3b23bb98),
	.w3(32'h3bab2403),
	.w4(32'hbb47eb3d),
	.w5(32'hbaa9620d),
	.w6(32'hbbc5292d),
	.w7(32'hbb077800),
	.w8(32'h3b898070),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c091960),
	.w1(32'h3a2cf1fa),
	.w2(32'h3b4574a5),
	.w3(32'h3bb5609c),
	.w4(32'h3a7a4d24),
	.w5(32'h3ab93a3e),
	.w6(32'h39a07e07),
	.w7(32'h3a832daf),
	.w8(32'hbaac9b44),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83ac5d),
	.w1(32'h3b5689f2),
	.w2(32'h3b989a70),
	.w3(32'h3b2582ab),
	.w4(32'h3b21cef4),
	.w5(32'h3b04181d),
	.w6(32'h3aed2f01),
	.w7(32'h3aadd278),
	.w8(32'hbb00a449),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8426f6),
	.w1(32'hbc8b3b63),
	.w2(32'hbc55c834),
	.w3(32'h3aa6970a),
	.w4(32'hb9942915),
	.w5(32'h3bb1c066),
	.w6(32'hbc16c0c0),
	.w7(32'hbc7799fa),
	.w8(32'h3c0abe7f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cde7ee6),
	.w1(32'hbbd65ef8),
	.w2(32'h3bfa60e4),
	.w3(32'h3ad97c98),
	.w4(32'hb970dd65),
	.w5(32'h39cd7709),
	.w6(32'hb9655679),
	.w7(32'h3b8c838c),
	.w8(32'h398c6c58),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f8fd8),
	.w1(32'hbc012c74),
	.w2(32'hbaec96f9),
	.w3(32'h3a452cc0),
	.w4(32'hbbbd468e),
	.w5(32'hbbe915e5),
	.w6(32'hbbd82689),
	.w7(32'hbb8d7998),
	.w8(32'hbb172097),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a6057),
	.w1(32'hba9d70ed),
	.w2(32'h3a81bacc),
	.w3(32'hbb501e6e),
	.w4(32'hbb674ac5),
	.w5(32'hbac2f9c9),
	.w6(32'hbaa15818),
	.w7(32'hbaabdce2),
	.w8(32'hbb083054),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83e831),
	.w1(32'hbb9b9bdb),
	.w2(32'hbabe8eb8),
	.w3(32'hbb7e7c9d),
	.w4(32'hbb7256c6),
	.w5(32'hbb776347),
	.w6(32'hbb5f6d51),
	.w7(32'hbb4e59d9),
	.w8(32'hbb56b6b0),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8bb19),
	.w1(32'hbc24cf64),
	.w2(32'hbcb81eb8),
	.w3(32'hba1e7bcf),
	.w4(32'hb9505940),
	.w5(32'h3bbaeb43),
	.w6(32'h3b07ef66),
	.w7(32'hbc138aeb),
	.w8(32'h3c90c11f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb63438),
	.w1(32'h3c10fc27),
	.w2(32'h3c803f9f),
	.w3(32'h3b1eaec1),
	.w4(32'h3bbf0f7e),
	.w5(32'h3c3b1895),
	.w6(32'h3c1dc03f),
	.w7(32'h3bf32a3d),
	.w8(32'hbc0ec9d2),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f63bd),
	.w1(32'hbb8636f4),
	.w2(32'hbbef6c12),
	.w3(32'hbc47b06c),
	.w4(32'hbb89c998),
	.w5(32'hbbeed82c),
	.w6(32'hbb2817e8),
	.w7(32'hbb315fc0),
	.w8(32'h39cfb2fe),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8dba6),
	.w1(32'hb9cbaa25),
	.w2(32'hba062e46),
	.w3(32'h3a211ab9),
	.w4(32'hba055871),
	.w5(32'hb88b8adc),
	.w6(32'hb9cb19f2),
	.w7(32'hba2b4659),
	.w8(32'hba3cbdd8),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e1e27),
	.w1(32'hbae7a38d),
	.w2(32'hbb1af9f7),
	.w3(32'hbb0698c7),
	.w4(32'h3ab22f25),
	.w5(32'h3b3dc078),
	.w6(32'hba3594fb),
	.w7(32'h3981ba67),
	.w8(32'h39631253),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule