module layer_8_featuremap_94(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1fb8a),
	.w1(32'h3a59188e),
	.w2(32'h379c1fb7),
	.w3(32'hbc17dee6),
	.w4(32'h39f69461),
	.w5(32'hbbb10830),
	.w6(32'hbc582dd5),
	.w7(32'hbbb54a6f),
	.w8(32'hbc31cfbf),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e08942),
	.w1(32'h3b49b2ff),
	.w2(32'hb8cae5a1),
	.w3(32'h3c1dcc05),
	.w4(32'h3b8228a1),
	.w5(32'h3c180e98),
	.w6(32'h3bb483ba),
	.w7(32'h3b27aba2),
	.w8(32'h3c6966be),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f787e),
	.w1(32'h3ca9c997),
	.w2(32'h3b966fcd),
	.w3(32'h3ca21eeb),
	.w4(32'h3c070d2a),
	.w5(32'h3c1ec906),
	.w6(32'h3ccc15c0),
	.w7(32'h3c96e915),
	.w8(32'h3c8c0dbf),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c020043),
	.w1(32'h3cf80296),
	.w2(32'hbb59d123),
	.w3(32'h3c85945f),
	.w4(32'h39a1f268),
	.w5(32'hbb595e28),
	.w6(32'h3c7aa32a),
	.w7(32'hba8d6902),
	.w8(32'hbb7de613),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d7747),
	.w1(32'h3b5a119a),
	.w2(32'h3c22bf4c),
	.w3(32'h3b61f794),
	.w4(32'hbb5355a7),
	.w5(32'hbac1ef48),
	.w6(32'hbb92d216),
	.w7(32'h3aec744e),
	.w8(32'h3b075160),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3715c3),
	.w1(32'h3a9aac5f),
	.w2(32'hbaba72e5),
	.w3(32'h3be57885),
	.w4(32'h3c0a888d),
	.w5(32'h3c18cbd1),
	.w6(32'h3a99dc95),
	.w7(32'h3b45af74),
	.w8(32'h3bd8ecb7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2d747),
	.w1(32'hbaf955e6),
	.w2(32'hbb4d7f08),
	.w3(32'h3bf5fb76),
	.w4(32'hbb18847b),
	.w5(32'h3b07663c),
	.w6(32'h3b6bfc91),
	.w7(32'hbacf7128),
	.w8(32'h3bb89e35),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd69a17),
	.w1(32'h3acfb91d),
	.w2(32'h3bc47a37),
	.w3(32'h3ccb9434),
	.w4(32'h3c8be0d3),
	.w5(32'h3bcd94e0),
	.w6(32'h3c81364b),
	.w7(32'h3bc53814),
	.w8(32'hba94e9b8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c975774),
	.w1(32'h3bcdc558),
	.w2(32'h3b101202),
	.w3(32'h3c3d75de),
	.w4(32'h3bcb77fd),
	.w5(32'hba28e920),
	.w6(32'h3c3d98d9),
	.w7(32'h3b82c9b7),
	.w8(32'h38e11af0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8f092),
	.w1(32'h3b962abd),
	.w2(32'h3c5ce520),
	.w3(32'h3be9b858),
	.w4(32'h3c4c5f2f),
	.w5(32'h3b4c5171),
	.w6(32'h3bb508ec),
	.w7(32'h3c2e6f0f),
	.w8(32'h3c5be7b4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf62093),
	.w1(32'hbae2ef37),
	.w2(32'hb9f7ef07),
	.w3(32'hbc1d3aba),
	.w4(32'h3ac5dc32),
	.w5(32'h3b86f7d9),
	.w6(32'hbb505ce9),
	.w7(32'hbc029b07),
	.w8(32'hbba0f545),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b5985),
	.w1(32'h3b74f7f6),
	.w2(32'h3c6dc3ad),
	.w3(32'hbb8c4c95),
	.w4(32'h3c1d7718),
	.w5(32'h3c01aec7),
	.w6(32'hbbb16d1c),
	.w7(32'h3c061184),
	.w8(32'h3bbb2d0d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbdd302),
	.w1(32'h3ba78bbe),
	.w2(32'hbba63dc0),
	.w3(32'h3c5390ff),
	.w4(32'h3bdd2408),
	.w5(32'h3c23f95a),
	.w6(32'h3c358462),
	.w7(32'h3bfe17c6),
	.w8(32'h3c7ba980),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37851604),
	.w1(32'hbb8445db),
	.w2(32'hbb8579fb),
	.w3(32'h3b3c09a7),
	.w4(32'hbaea31de),
	.w5(32'h3b70e4f6),
	.w6(32'h3a95a03d),
	.w7(32'hbb69831c),
	.w8(32'h3aa170f9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80cc57),
	.w1(32'hbc12b821),
	.w2(32'hbb77305a),
	.w3(32'h3c228960),
	.w4(32'hb9a27638),
	.w5(32'hbaecf6fe),
	.w6(32'h3a3a3e9f),
	.w7(32'hb98550b5),
	.w8(32'hbb40fcb3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd38c4),
	.w1(32'hbba73373),
	.w2(32'hbca9804b),
	.w3(32'h3b63d3cd),
	.w4(32'h3b63fcd1),
	.w5(32'hbc3ace24),
	.w6(32'h3a8d6604),
	.w7(32'h3c553192),
	.w8(32'h3cdf3118),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43dd37),
	.w1(32'hbc199fd8),
	.w2(32'h3c2f3aa0),
	.w3(32'hbbc02c1f),
	.w4(32'hbcc72cee),
	.w5(32'hbc96e2ed),
	.w6(32'hbcb7ff92),
	.w7(32'hbbdae006),
	.w8(32'hbb9f2040),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf364d),
	.w1(32'h3c501516),
	.w2(32'hbb2c9859),
	.w3(32'h3903bf3c),
	.w4(32'hbb69110d),
	.w5(32'hbc4069d8),
	.w6(32'h3c3b79ee),
	.w7(32'h3c5b7ed4),
	.w8(32'h3d82e155),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c799a3a),
	.w1(32'h3c66e540),
	.w2(32'h3c046d7f),
	.w3(32'hbcae95a6),
	.w4(32'h3b1836c3),
	.w5(32'hbc98149d),
	.w6(32'hbd14a59d),
	.w7(32'hbc7b704a),
	.w8(32'h3cccbef6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79eae2),
	.w1(32'h3cc4710d),
	.w2(32'h3a9d91d8),
	.w3(32'hbccd1cb3),
	.w4(32'h3c091485),
	.w5(32'hbc97c04f),
	.w6(32'h3b024d98),
	.w7(32'hbca9d3d4),
	.w8(32'h3d3c0eed),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb266c71),
	.w1(32'h3c4e7f58),
	.w2(32'hbb2dc59a),
	.w3(32'hbd5ca4c0),
	.w4(32'h3b19063c),
	.w5(32'h3cd139bd),
	.w6(32'h3b2bf98a),
	.w7(32'hbbfcf77d),
	.w8(32'hbc789546),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aef90),
	.w1(32'hbc645ab2),
	.w2(32'h3ca1f016),
	.w3(32'h3d2ad21f),
	.w4(32'hbc592b0a),
	.w5(32'h3c9f8321),
	.w6(32'h3c828e33),
	.w7(32'h3c62a67f),
	.w8(32'h3c0b2ecf),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86e150),
	.w1(32'h3bfbcffe),
	.w2(32'hbb2eb6b3),
	.w3(32'hba6d3c65),
	.w4(32'h3c33ff76),
	.w5(32'h3bb9e235),
	.w6(32'h3b9f8ca0),
	.w7(32'hbc51e989),
	.w8(32'hbca1b28c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5b6d4),
	.w1(32'hbca790fe),
	.w2(32'h3b2e18a1),
	.w3(32'hbbdab668),
	.w4(32'h3c3bc785),
	.w5(32'h3a470956),
	.w6(32'hbcd0b00a),
	.w7(32'h3c83f8ab),
	.w8(32'h3c5630fd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05562f),
	.w1(32'h3c3660f0),
	.w2(32'h3a286add),
	.w3(32'hbc18feee),
	.w4(32'h3bce08cd),
	.w5(32'h3bb4a7b9),
	.w6(32'h3ac73977),
	.w7(32'h3b6ca44a),
	.w8(32'h3bcd5952),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc13a5),
	.w1(32'h3bfc5f51),
	.w2(32'h3baac09b),
	.w3(32'h3a347b29),
	.w4(32'hbc6fd447),
	.w5(32'h3ce3fbf5),
	.w6(32'hbb986a2f),
	.w7(32'hbcfca0fb),
	.w8(32'hbb6a811f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7169ea),
	.w1(32'h3c1a5f06),
	.w2(32'hbcaa73bf),
	.w3(32'h3c65b645),
	.w4(32'h3c0914fe),
	.w5(32'hbc4f43cb),
	.w6(32'h3d0c9455),
	.w7(32'hbc832736),
	.w8(32'h3c169496),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd6afe6),
	.w1(32'hbcdca05e),
	.w2(32'h3cff9227),
	.w3(32'hbd0de9ed),
	.w4(32'h3c564474),
	.w5(32'h3d190f03),
	.w6(32'hbd223921),
	.w7(32'hbcd261b6),
	.w8(32'hbd2889f7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3735f6),
	.w1(32'h3a3986ca),
	.w2(32'h3c736c04),
	.w3(32'h3cbd58de),
	.w4(32'h3c0fcdfc),
	.w5(32'h3cc5dc4a),
	.w6(32'hbb841e9b),
	.w7(32'hbd3fd04b),
	.w8(32'hbcc15d54),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc2dce2),
	.w1(32'h3b169701),
	.w2(32'hbc2a8c54),
	.w3(32'h3c3e7e77),
	.w4(32'h3b8b585c),
	.w5(32'h3b53665a),
	.w6(32'h3d016b04),
	.w7(32'h3c166c98),
	.w8(32'hb9a42e41),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11684d),
	.w1(32'hbb21942a),
	.w2(32'hba392612),
	.w3(32'h3bf79cb9),
	.w4(32'h3a870337),
	.w5(32'h3a883b2d),
	.w6(32'hbaace090),
	.w7(32'h3b93e67f),
	.w8(32'h3b84d372),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b282dd6),
	.w1(32'h3ba126c5),
	.w2(32'h39a2d99f),
	.w3(32'h3c084a74),
	.w4(32'hba0a2459),
	.w5(32'hbc1e6210),
	.w6(32'h3c2d002c),
	.w7(32'hbc189d0a),
	.w8(32'hbab7eaf8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc75996),
	.w1(32'hbcb60c3a),
	.w2(32'hbb5caa33),
	.w3(32'hbb93318e),
	.w4(32'hbabac967),
	.w5(32'h3c8530ab),
	.w6(32'hbd4484cc),
	.w7(32'h3b6beaae),
	.w8(32'h3c06eeda),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9600ed),
	.w1(32'h3c909f1b),
	.w2(32'hbc23859a),
	.w3(32'hbaa315e0),
	.w4(32'hbc3b6d77),
	.w5(32'hbcff001b),
	.w6(32'h3cb6ff96),
	.w7(32'h3c536ec2),
	.w8(32'h3c70a538),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3a72f),
	.w1(32'h3c1f2bfb),
	.w2(32'hbc267b04),
	.w3(32'hbcdf5a7b),
	.w4(32'h3c6882f7),
	.w5(32'h3cab2e7c),
	.w6(32'h3c8e726e),
	.w7(32'h3bc84eaa),
	.w8(32'h3bbaeeee),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc496964),
	.w1(32'h3a6823bb),
	.w2(32'h3c805853),
	.w3(32'h3c41f47f),
	.w4(32'h3cb18dd1),
	.w5(32'h3cd01bb5),
	.w6(32'h3c0bde6f),
	.w7(32'hbc6ad242),
	.w8(32'hbd1dd3fd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbcaf5d),
	.w1(32'hbd07382d),
	.w2(32'hbbcc3b77),
	.w3(32'h3c7240e6),
	.w4(32'h3c1a100f),
	.w5(32'h3cb12c60),
	.w6(32'h3bc659ad),
	.w7(32'hbcd0a8c5),
	.w8(32'h3c4e8e76),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f8a51),
	.w1(32'hbc85d0f9),
	.w2(32'h3c564333),
	.w3(32'h3c566af2),
	.w4(32'hbc33ce7a),
	.w5(32'hbc71e162),
	.w6(32'h3c3dc8d5),
	.w7(32'h3cca89f6),
	.w8(32'h3b12389e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e80b4),
	.w1(32'h3c7e78de),
	.w2(32'hbb2eae4e),
	.w3(32'hbc093c0b),
	.w4(32'hbb88ce30),
	.w5(32'hbc810d1b),
	.w6(32'h3c459c6f),
	.w7(32'hbc4ec8a7),
	.w8(32'h3ca540aa),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb25faf),
	.w1(32'h3a06ff68),
	.w2(32'h3b2eafe5),
	.w3(32'hbc91966f),
	.w4(32'hbbb77384),
	.w5(32'hba8a6a0b),
	.w6(32'hbaeefb8c),
	.w7(32'hbc39e4e5),
	.w8(32'hbb612ffd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c692eb7),
	.w1(32'h3c73272d),
	.w2(32'hb972fa87),
	.w3(32'h3b6813e7),
	.w4(32'h3c95330c),
	.w5(32'hbcd3492d),
	.w6(32'h3c25be8e),
	.w7(32'h3c895084),
	.w8(32'h3d0edcca),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9691aa),
	.w1(32'h3c2930bc),
	.w2(32'hbc900318),
	.w3(32'hbc560c76),
	.w4(32'h3c9c18ce),
	.w5(32'h3cc41f41),
	.w6(32'hbc815e57),
	.w7(32'h3b5f3d23),
	.w8(32'hbc3536d2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad71217),
	.w1(32'hbc76e08a),
	.w2(32'hbbd6895f),
	.w3(32'h3c455acc),
	.w4(32'hbb19b185),
	.w5(32'h3cb73855),
	.w6(32'hbc2d8011),
	.w7(32'h3baae0ee),
	.w8(32'hbae86b7b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e92cc),
	.w1(32'hbba6df54),
	.w2(32'hbb3b6bdd),
	.w3(32'hbab19958),
	.w4(32'h3b0ca42b),
	.w5(32'h3b8c35d1),
	.w6(32'h3c2e976b),
	.w7(32'hbae3930c),
	.w8(32'h3bbea17b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cd064),
	.w1(32'h3b7e2835),
	.w2(32'h3d04a22d),
	.w3(32'h3b8da7d4),
	.w4(32'hbb202971),
	.w5(32'h3cd211e0),
	.w6(32'hbb74ac70),
	.w7(32'hbce91386),
	.w8(32'hbd1d936c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae95db),
	.w1(32'hbbcb31d8),
	.w2(32'hbb57bfd4),
	.w3(32'h3c8c0ca0),
	.w4(32'h3c309262),
	.w5(32'h3c3c24a2),
	.w6(32'h3c181d48),
	.w7(32'h3a768d3d),
	.w8(32'hbc5db484),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ecf13),
	.w1(32'hbbbfc2c7),
	.w2(32'hbb7eba0b),
	.w3(32'h3bae3bbf),
	.w4(32'h3cfaec51),
	.w5(32'h3cfdfcc1),
	.w6(32'hbc2bac19),
	.w7(32'hbcf1bc9b),
	.w8(32'h3c102f26),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce8e4ff),
	.w1(32'hbc1630d1),
	.w2(32'h3b991818),
	.w3(32'h3b18091a),
	.w4(32'hbb47f81a),
	.w5(32'h3d29869d),
	.w6(32'h3cb3d9da),
	.w7(32'hbcd9cbbb),
	.w8(32'h3c7dfc8e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66bc6d),
	.w1(32'h3c1dedaa),
	.w2(32'hbbf606e9),
	.w3(32'h3c188d6f),
	.w4(32'hbb9e8a65),
	.w5(32'hbc849e08),
	.w6(32'h3d2b0a64),
	.w7(32'h3bcc0f06),
	.w8(32'hbbdc82d4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3d9f21),
	.w1(32'hbbf1f46d),
	.w2(32'h3baaedfc),
	.w3(32'h3a7dd447),
	.w4(32'hbcc94c2d),
	.w5(32'hbd5082c8),
	.w6(32'hbd369112),
	.w7(32'h3c42847e),
	.w8(32'h3cc5a16b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d615309),
	.w1(32'h3c268c4c),
	.w2(32'h3c18f154),
	.w3(32'hbce52f71),
	.w4(32'h3bba2263),
	.w5(32'hbcc3b24e),
	.w6(32'hbd0f43b3),
	.w7(32'h3d170214),
	.w8(32'hbc3415fc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64ea3b),
	.w1(32'h3c25eca2),
	.w2(32'hbc3f83bf),
	.w3(32'h3bd2fdca),
	.w4(32'h3d0962e6),
	.w5(32'h3d2cdb75),
	.w6(32'hbcd40d68),
	.w7(32'hbd336907),
	.w8(32'hbcf23a3d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdcdd4),
	.w1(32'hbc1cb4c7),
	.w2(32'hbc766fd9),
	.w3(32'h3c99ae31),
	.w4(32'h3b148a90),
	.w5(32'hbcb18907),
	.w6(32'h3c3427d6),
	.w7(32'h3ac29c6a),
	.w8(32'hbbc51fc9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78d5da),
	.w1(32'h3c7fd157),
	.w2(32'h3a477c3d),
	.w3(32'h3c08b099),
	.w4(32'h3ad04c9f),
	.w5(32'h3b7702b2),
	.w6(32'h3b491c13),
	.w7(32'h3bec5768),
	.w8(32'h3c40af1b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7be45e),
	.w1(32'hbb93e82f),
	.w2(32'h3bb19203),
	.w3(32'h3b90d8fd),
	.w4(32'h3c57bed4),
	.w5(32'h3d133032),
	.w6(32'h3b0820ff),
	.w7(32'hbce42a39),
	.w8(32'h3b0d8cec),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69a8d1),
	.w1(32'h3c16eeeb),
	.w2(32'h3c74d289),
	.w3(32'h39268a42),
	.w4(32'hbc7c64cf),
	.w5(32'hbcaa6559),
	.w6(32'h3d0c7e75),
	.w7(32'h3ca63865),
	.w8(32'h3c8c6ef2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c562f74),
	.w1(32'h3c37fe25),
	.w2(32'h3bd46cc6),
	.w3(32'hbc0afb32),
	.w4(32'h3c0a8ac0),
	.w5(32'h3bf81d5a),
	.w6(32'h3ac705fa),
	.w7(32'h3c080188),
	.w8(32'hb99cc5bc),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c426bbf),
	.w1(32'h3af43590),
	.w2(32'h3cb21747),
	.w3(32'h3c0e1a7b),
	.w4(32'hb97e9a71),
	.w5(32'h3c839879),
	.w6(32'hbb78ec4d),
	.w7(32'hbc3f14a4),
	.w8(32'hbcf4ed0b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4bb78c),
	.w1(32'h3cc48329),
	.w2(32'hbb48956c),
	.w3(32'h3c093485),
	.w4(32'h3af5811b),
	.w5(32'h3b05d438),
	.w6(32'h3c81e746),
	.w7(32'hbb66fbd7),
	.w8(32'h3ac3e25e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b689d24),
	.w1(32'h3b16669f),
	.w2(32'hbaf4f0ba),
	.w3(32'h3bee4968),
	.w4(32'h3b317b2a),
	.w5(32'h3ba83cfe),
	.w6(32'h3bcb323c),
	.w7(32'h3ae02468),
	.w8(32'h3c6921e2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacc144),
	.w1(32'hba2793f6),
	.w2(32'hbbbbc29d),
	.w3(32'h3b7e2d53),
	.w4(32'hbca63ff0),
	.w5(32'hbc94e61a),
	.w6(32'h3b0279ec),
	.w7(32'h3c1d57ef),
	.w8(32'hbc8bb1a9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ab5b2),
	.w1(32'hbb3c3760),
	.w2(32'h3b9e6d2c),
	.w3(32'h3bd46051),
	.w4(32'hbc04f7f1),
	.w5(32'h3974c85a),
	.w6(32'hbb12494d),
	.w7(32'hbc130335),
	.w8(32'hbc986fba),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5847d2),
	.w1(32'h3bc7793a),
	.w2(32'h3d1442ed),
	.w3(32'h3bd0052b),
	.w4(32'hbce87bc9),
	.w5(32'hba81e794),
	.w6(32'hb785d45e),
	.w7(32'h3c87e322),
	.w8(32'hbb05e60f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47175c),
	.w1(32'hbc19609f),
	.w2(32'h3b8c559f),
	.w3(32'h3c23ea92),
	.w4(32'h3c6828c2),
	.w5(32'h3c1ff4df),
	.w6(32'hbb35d1d0),
	.w7(32'h3c0d6f39),
	.w8(32'hbc5cf6f4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc26933),
	.w1(32'h3c1cbb39),
	.w2(32'h3b4f2f2c),
	.w3(32'h3c8d9988),
	.w4(32'h3c19f158),
	.w5(32'h3ccf18ad),
	.w6(32'hbc10e0e2),
	.w7(32'hbc1c23ef),
	.w8(32'hbc4b5a55),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b540ff3),
	.w1(32'h3b391a38),
	.w2(32'h3ca19543),
	.w3(32'h3cb92302),
	.w4(32'h3aa7cc70),
	.w5(32'hbcc07adc),
	.w6(32'h3bbd5868),
	.w7(32'h3cb24143),
	.w8(32'hbc17f771),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d01b98a),
	.w1(32'h3ced2051),
	.w2(32'h3b6cf6bd),
	.w3(32'h3be94b31),
	.w4(32'h3c87a841),
	.w5(32'hbb353a8c),
	.w6(32'h3c82c281),
	.w7(32'hbbaa24ad),
	.w8(32'h3cfb2c58),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ac8d3),
	.w1(32'h3c8eeb8e),
	.w2(32'hbb28d774),
	.w3(32'hbd436728),
	.w4(32'hbb1dce8c),
	.w5(32'hbb9dcb59),
	.w6(32'h3c7d2dee),
	.w7(32'h3a32ab9f),
	.w8(32'hbc1255e3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62ab47),
	.w1(32'hbbeab25c),
	.w2(32'hbb881c55),
	.w3(32'hbb0dca3f),
	.w4(32'hbada389d),
	.w5(32'hbbec1ac9),
	.w6(32'hbca3a7cb),
	.w7(32'h3c71b2a0),
	.w8(32'h3cab243f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb42176),
	.w1(32'hbbb6959f),
	.w2(32'h3c1dbd81),
	.w3(32'h3b2bdad0),
	.w4(32'h3c094744),
	.w5(32'h3c4dae4a),
	.w6(32'hbd1d2f65),
	.w7(32'hbc1ced70),
	.w8(32'hbca207f7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b2357),
	.w1(32'hbb18f18a),
	.w2(32'h3ce0fc27),
	.w3(32'hbc41707e),
	.w4(32'h3ced376b),
	.w5(32'h3c3b1ec5),
	.w6(32'hbc8e89f4),
	.w7(32'h3c86ee3f),
	.w8(32'hbc30db07),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c877389),
	.w1(32'h3bdbffbc),
	.w2(32'hbbdd9ac6),
	.w3(32'hbb5fb08d),
	.w4(32'hb9de2ce1),
	.w5(32'hbc4dfd4e),
	.w6(32'hbc9478a7),
	.w7(32'h3ce6a675),
	.w8(32'hbc555b68),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ee2e6),
	.w1(32'h3bf23ff0),
	.w2(32'h3c8365b5),
	.w3(32'h3c18236a),
	.w4(32'h3b7c86d1),
	.w5(32'h3bf667fb),
	.w6(32'hbb7da3a3),
	.w7(32'hbc205022),
	.w8(32'hbca8ac1f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cebea3f),
	.w1(32'h3c3fd583),
	.w2(32'h3b67873e),
	.w3(32'h3c34d5c3),
	.w4(32'h3c86a991),
	.w5(32'hbbbcb9b3),
	.w6(32'hbb996d95),
	.w7(32'h3cf72d21),
	.w8(32'h3c16d65c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cabf51f),
	.w1(32'hbadd96e0),
	.w2(32'hbc92a810),
	.w3(32'h3b32835c),
	.w4(32'hbbaa4647),
	.w5(32'hbbd9a318),
	.w6(32'hbd1226c5),
	.w7(32'hbcc275f1),
	.w8(32'h3cfaf8fc),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e7c66),
	.w1(32'hbc09d9b5),
	.w2(32'hbb7a1c99),
	.w3(32'hbcc642ca),
	.w4(32'hbc7e4409),
	.w5(32'hbc55c586),
	.w6(32'h3b9f3b46),
	.w7(32'h3c91e8bd),
	.w8(32'hbb67bd8a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd314af),
	.w1(32'hbb4514e1),
	.w2(32'h386e6185),
	.w3(32'h3bf30f02),
	.w4(32'hb7ac63e3),
	.w5(32'hb5bbb1b4),
	.w6(32'hbb3cb0b1),
	.w7(32'hb883d4d9),
	.w8(32'h3743d95e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ad06a),
	.w1(32'h3bdf3c0b),
	.w2(32'h3bc753e3),
	.w3(32'hba9c306c),
	.w4(32'h3ae2eeb5),
	.w5(32'h3afbf4c8),
	.w6(32'hbc066661),
	.w7(32'hbc3aca84),
	.w8(32'hbc047d96),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bd7a2),
	.w1(32'h3a145f27),
	.w2(32'h3b1da1c5),
	.w3(32'hbac3ff50),
	.w4(32'hbaf2dd7c),
	.w5(32'hb9d04aa7),
	.w6(32'h3b7d83b8),
	.w7(32'h3bb57f83),
	.w8(32'h3bcc5d83),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90593b6),
	.w1(32'hb9dc6bb4),
	.w2(32'hb7ab1f44),
	.w3(32'h3991b9cf),
	.w4(32'h38d89fdb),
	.w5(32'h395ca231),
	.w6(32'h3964080d),
	.w7(32'h38389389),
	.w8(32'h39bcdbea),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35bdb631),
	.w1(32'hb63f7858),
	.w2(32'hb8908544),
	.w3(32'hb8cab6c7),
	.w4(32'hb79ffcd6),
	.w5(32'hb8f837d8),
	.w6(32'hb595f1dd),
	.w7(32'hb7247813),
	.w8(32'hb8ccbe8d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1d9ea),
	.w1(32'h3b3d1a27),
	.w2(32'h3b4eccac),
	.w3(32'h3b1d096d),
	.w4(32'h3bcbc720),
	.w5(32'h3bbbfad0),
	.w6(32'h3b55def9),
	.w7(32'h3b3eca8c),
	.w8(32'h3b08b4ca),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29ae6d),
	.w1(32'h3bac96e7),
	.w2(32'h3ba99926),
	.w3(32'hbaa66661),
	.w4(32'hbaa50d43),
	.w5(32'h3a520bb0),
	.w6(32'hbc07483c),
	.w7(32'hbc19aa0a),
	.w8(32'hbbc00f08),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd8974f),
	.w1(32'h3c7cd440),
	.w2(32'h3c9b9de3),
	.w3(32'h3c8f17cb),
	.w4(32'h3ba7000a),
	.w5(32'h3c29f978),
	.w6(32'hbbf4de50),
	.w7(32'hbb6f62e1),
	.w8(32'h3bd141e2),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30627d),
	.w1(32'h3c8eeb18),
	.w2(32'h3c569681),
	.w3(32'h3bb44b61),
	.w4(32'h3b84f34a),
	.w5(32'h3bea3e39),
	.w6(32'hbc03e09f),
	.w7(32'hbc2f5ab1),
	.w8(32'hbb8b87d1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00ea0d),
	.w1(32'h3c1aea26),
	.w2(32'h3b68efc4),
	.w3(32'h3b70e866),
	.w4(32'h3bdb17c0),
	.w5(32'h3bb364be),
	.w6(32'hbabc3ff7),
	.w7(32'hbb0fb93d),
	.w8(32'hba570b3d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953a036),
	.w1(32'hb8dc56d3),
	.w2(32'hb9c10c5b),
	.w3(32'hb998b25b),
	.w4(32'hb9067c75),
	.w5(32'hb972dc6e),
	.w6(32'hb9037143),
	.w7(32'h39c71b35),
	.w8(32'h39220626),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ca1934),
	.w1(32'h37975015),
	.w2(32'hb82a5ed6),
	.w3(32'hb89bf33c),
	.w4(32'h37a935b9),
	.w5(32'hb80487d9),
	.w6(32'hb7f0bcdc),
	.w7(32'h3836ac36),
	.w8(32'h380d439b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e3842),
	.w1(32'h38ea6fb9),
	.w2(32'hb8a3eeb9),
	.w3(32'hb815c610),
	.w4(32'h38d0eeb8),
	.w5(32'hb8a34d4a),
	.w6(32'h3803d1ec),
	.w7(32'h3924760d),
	.w8(32'hb504be4d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9443d),
	.w1(32'h3b2c3164),
	.w2(32'h39c2a609),
	.w3(32'hba7ae90e),
	.w4(32'h3a3f43a1),
	.w5(32'hba2e373e),
	.w6(32'hbb6057c0),
	.w7(32'hbb6c1913),
	.w8(32'hbb4291e5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9401f9),
	.w1(32'h3b632223),
	.w2(32'h3b71853e),
	.w3(32'h3b257fb6),
	.w4(32'h3b5c57d5),
	.w5(32'h3ba90099),
	.w6(32'h3add3aa1),
	.w7(32'h3b18c28d),
	.w8(32'h3b0e22b9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a4f79),
	.w1(32'h3a03852b),
	.w2(32'h39e99a23),
	.w3(32'h3a82333b),
	.w4(32'h3a150da0),
	.w5(32'h3a5b6902),
	.w6(32'h3afe2c45),
	.w7(32'h3a948100),
	.w8(32'h3a7ce59c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39112a5c),
	.w1(32'hbae087b9),
	.w2(32'h399adb4a),
	.w3(32'h3b728bc1),
	.w4(32'h3b8c60cb),
	.w5(32'h3b917a43),
	.w6(32'h3a9a8c9c),
	.w7(32'hba995fe6),
	.w8(32'hbac861be),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce89e1),
	.w1(32'h3bc6ad48),
	.w2(32'h3b90ddb7),
	.w3(32'h3b76599f),
	.w4(32'h3b4b6305),
	.w5(32'h3b20ef33),
	.w6(32'h3aac3e86),
	.w7(32'hb8aaf635),
	.w8(32'h3a771a56),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0817f5),
	.w1(32'h3a2c5702),
	.w2(32'h3aafd276),
	.w3(32'h3a30ac7f),
	.w4(32'hb94b1e67),
	.w5(32'h3a134553),
	.w6(32'h3badf187),
	.w7(32'h3bc43c7b),
	.w8(32'h3bbe3bb4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a837f0c),
	.w1(32'h3b95e47a),
	.w2(32'h3b82205d),
	.w3(32'h39ca1331),
	.w4(32'h3b024e18),
	.w5(32'h3a6ea514),
	.w6(32'hb928b3f9),
	.w7(32'h39d7c058),
	.w8(32'h3ac5296d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c294bb0),
	.w1(32'h3c04ee77),
	.w2(32'h3a4cbb5a),
	.w3(32'hbb0285e1),
	.w4(32'hbb1dc927),
	.w5(32'hbb3fda14),
	.w6(32'hbc258ba8),
	.w7(32'hbbf2d0d2),
	.w8(32'hbb451097),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f303bb),
	.w1(32'h3893f590),
	.w2(32'h38357af4),
	.w3(32'h378d76ea),
	.w4(32'hb71544a6),
	.w5(32'h37597627),
	.w6(32'h388bc0a3),
	.w7(32'h3943caf4),
	.w8(32'h37fca39c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984b7a1),
	.w1(32'hb8cfdf79),
	.w2(32'hb91f34bf),
	.w3(32'hb899c06c),
	.w4(32'h38f93616),
	.w5(32'hb73297af),
	.w6(32'h3734f3ca),
	.w7(32'h3951b213),
	.w8(32'h37291edc),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97cdde0),
	.w1(32'hb8fa5700),
	.w2(32'hb944fc11),
	.w3(32'hb9429ca9),
	.w4(32'hb7d4c47c),
	.w5(32'hb90dc8ea),
	.w6(32'hb6b171d8),
	.w7(32'h38731793),
	.w8(32'hb6887e65),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ea13a),
	.w1(32'h39191dcd),
	.w2(32'h39475a82),
	.w3(32'h39d075b8),
	.w4(32'h3a0dd454),
	.w5(32'h39d5c764),
	.w6(32'h39a82489),
	.w7(32'h39de11d3),
	.w8(32'h38e4d13a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76386a),
	.w1(32'h3b47aebb),
	.w2(32'h3a27e2a4),
	.w3(32'h3b71b408),
	.w4(32'h3b4e1ce9),
	.w5(32'h3b02c6e2),
	.w6(32'h3b34abba),
	.w7(32'h3b3f60e7),
	.w8(32'h3b41b22c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae57159),
	.w1(32'h3b007f9a),
	.w2(32'h3aad28c2),
	.w3(32'h368dd602),
	.w4(32'h3a78cf5f),
	.w5(32'h3a1f4c80),
	.w6(32'hb9586aef),
	.w7(32'h3ab2a05b),
	.w8(32'h39a537d2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5010e6),
	.w1(32'h3b035136),
	.w2(32'h3b15595d),
	.w3(32'h3b414495),
	.w4(32'h3b93eb6f),
	.w5(32'h3b87e03f),
	.w6(32'h3b7506b9),
	.w7(32'h3b9b595c),
	.w8(32'h3b8750e2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cda9b1),
	.w1(32'hba9dd054),
	.w2(32'hba219ab0),
	.w3(32'h3a109c3a),
	.w4(32'h3a41d1c3),
	.w5(32'h39f87e1d),
	.w6(32'h3b072233),
	.w7(32'h3aeeab32),
	.w8(32'h3aaf18a9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b38f7),
	.w1(32'h3b903390),
	.w2(32'h3b30435a),
	.w3(32'h39964f68),
	.w4(32'h39a7bb57),
	.w5(32'h3abea464),
	.w6(32'hbbe040c6),
	.w7(32'hbc18f14c),
	.w8(32'hbbd6ae57),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cfd2bf),
	.w1(32'h383f21d7),
	.w2(32'hbad18a46),
	.w3(32'hbb87e375),
	.w4(32'hbb4c39c6),
	.w5(32'hbb75a6c0),
	.w6(32'hbbe335fc),
	.w7(32'hbbce1b4e),
	.w8(32'hbb819465),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaced3ed),
	.w1(32'hbad52598),
	.w2(32'hbaa09a5c),
	.w3(32'hba9baf28),
	.w4(32'h382e0cab),
	.w5(32'hb71a2251),
	.w6(32'hbae26757),
	.w7(32'hba846af0),
	.w8(32'h39090ab7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17f51e),
	.w1(32'h3a605585),
	.w2(32'h3b11d429),
	.w3(32'h3b88861f),
	.w4(32'h3b3abf2b),
	.w5(32'h3b3c8513),
	.w6(32'h3ba66535),
	.w7(32'h3b7b5d90),
	.w8(32'h3b587c93),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38fb46),
	.w1(32'h3c153196),
	.w2(32'h3b0386a1),
	.w3(32'h3bb044e4),
	.w4(32'h3bac769b),
	.w5(32'h3b3a4607),
	.w6(32'h3b55fe86),
	.w7(32'h3b9d5e77),
	.w8(32'h3b809d1b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8ff96),
	.w1(32'hbb023482),
	.w2(32'h39731ed0),
	.w3(32'hbb963992),
	.w4(32'hbba6e095),
	.w5(32'hb9a85e80),
	.w6(32'h39c06ad6),
	.w7(32'hb902733c),
	.w8(32'h3b65cb50),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb10bbb),
	.w1(32'h3ac76415),
	.w2(32'h3ba92ed8),
	.w3(32'h3b374936),
	.w4(32'hb979f114),
	.w5(32'h3b92232d),
	.w6(32'h3b913992),
	.w7(32'h390ec8cb),
	.w8(32'h3b69d622),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a290246),
	.w1(32'hba3cae02),
	.w2(32'h3a886156),
	.w3(32'h3b69b9bb),
	.w4(32'h3b4fe7a0),
	.w5(32'h3b67a557),
	.w6(32'h3bc5967f),
	.w7(32'h3bbfe167),
	.w8(32'h3b96e551),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f7656a),
	.w1(32'h3a08feae),
	.w2(32'h384579b4),
	.w3(32'h393ef8cd),
	.w4(32'h3a14a4cf),
	.w5(32'h39686470),
	.w6(32'h37f70c9a),
	.w7(32'h3a255938),
	.w8(32'h39a544f7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a18b9),
	.w1(32'h3abada9b),
	.w2(32'hba768eab),
	.w3(32'h3a4e2784),
	.w4(32'hb9aeba83),
	.w5(32'h39edb577),
	.w6(32'hba3e9bfc),
	.w7(32'hba12b470),
	.w8(32'hba2d37f2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbdb34),
	.w1(32'h3b0a4f64),
	.w2(32'h3aa9c152),
	.w3(32'hb8e37266),
	.w4(32'hb8b4be71),
	.w5(32'hba369205),
	.w6(32'hba08bd49),
	.w7(32'hb92f2528),
	.w8(32'hbac0630e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c59cf),
	.w1(32'hba9edc59),
	.w2(32'h3aa1ace7),
	.w3(32'h39ac7c4c),
	.w4(32'hba17e80f),
	.w5(32'h3b078d17),
	.w6(32'h3a88782c),
	.w7(32'h39f0523c),
	.w8(32'h3b08f41e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dc13c),
	.w1(32'h3b82e1fa),
	.w2(32'h3bc48eff),
	.w3(32'h3ae628c6),
	.w4(32'h3b018fe1),
	.w5(32'h3b889651),
	.w6(32'hbadc2505),
	.w7(32'hbb970c7c),
	.w8(32'hbad9fc64),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885e344),
	.w1(32'hb81327f5),
	.w2(32'hb8798a70),
	.w3(32'hb8128fcd),
	.w4(32'h378d19d1),
	.w5(32'hb8cba88e),
	.w6(32'h37950080),
	.w7(32'h358487c2),
	.w8(32'h375310bf),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22beb8),
	.w1(32'hb8dce618),
	.w2(32'hb90532f9),
	.w3(32'hb97040d5),
	.w4(32'hb9d537cd),
	.w5(32'hb81c571b),
	.w6(32'h39cd692a),
	.w7(32'h3a2de304),
	.w8(32'h39dad10c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf83e3),
	.w1(32'h3b7f6975),
	.w2(32'h3b604f0e),
	.w3(32'h3c024e5d),
	.w4(32'h3c2998fa),
	.w5(32'h3c0dd20c),
	.w6(32'h3c1d0c7d),
	.w7(32'h3c052072),
	.w8(32'h3bbd12b8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c8785),
	.w1(32'h3b1fecdb),
	.w2(32'hb8d21c3a),
	.w3(32'hbbaf6399),
	.w4(32'hbb51b942),
	.w5(32'hbadf5794),
	.w6(32'h3a1651d3),
	.w7(32'h3b7cbaa5),
	.w8(32'h3bb4189a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a256a48),
	.w1(32'h3a9640d2),
	.w2(32'h38dea393),
	.w3(32'h3a8adbaa),
	.w4(32'h3aa45d48),
	.w5(32'h3a596e5a),
	.w6(32'h3ae39ad8),
	.w7(32'h3b145bb7),
	.w8(32'h3ae06d8a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a6be9),
	.w1(32'hbb059906),
	.w2(32'hbad185a4),
	.w3(32'h3ad9b566),
	.w4(32'h3ab1a799),
	.w5(32'h3b14c6bc),
	.w6(32'h3b36c619),
	.w7(32'h3ae923c1),
	.w8(32'h3af091b4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80f118),
	.w1(32'h3adae026),
	.w2(32'h393656f2),
	.w3(32'h3b25b3cd),
	.w4(32'h3ab47d6a),
	.w5(32'h3af7cf76),
	.w6(32'h3ad6daf2),
	.w7(32'h3afba634),
	.w8(32'h3b0d4f64),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54c905),
	.w1(32'h3ba27a16),
	.w2(32'h3b1f0d67),
	.w3(32'h3b92ec25),
	.w4(32'h3ba9f86c),
	.w5(32'h3b3713b5),
	.w6(32'h3bc694da),
	.w7(32'h3b8fc788),
	.w8(32'h3b51cc55),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a79421),
	.w1(32'hb9e92924),
	.w2(32'hbacecd08),
	.w3(32'hbad598bc),
	.w4(32'hba64349d),
	.w5(32'hba8707d0),
	.w6(32'h3ab45ee0),
	.w7(32'h3afeea83),
	.w8(32'h3adc09aa),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74dc7d),
	.w1(32'hbabcd9e7),
	.w2(32'h396e1668),
	.w3(32'hbac0930a),
	.w4(32'h3a1df0a2),
	.w5(32'h3a973071),
	.w6(32'hba9a38cc),
	.w7(32'hbab1a448),
	.w8(32'hba377f79),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule