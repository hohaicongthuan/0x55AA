module layer_10_featuremap_34(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74ba79),
	.w1(32'h3b43d7c3),
	.w2(32'hbb9896c2),
	.w3(32'h3a2de6d5),
	.w4(32'hb994d82b),
	.w5(32'hbbc79ed2),
	.w6(32'hbc260752),
	.w7(32'hbbcd2a71),
	.w8(32'h3bb2627e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91da67),
	.w1(32'hb8ea4a2a),
	.w2(32'hb983d222),
	.w3(32'hbb88b611),
	.w4(32'hbabe2d3f),
	.w5(32'hbb1cca3a),
	.w6(32'hb9e3177a),
	.w7(32'hb889b5e9),
	.w8(32'hbb0ff561),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb5f62),
	.w1(32'h3bb5f51a),
	.w2(32'hbad49fa0),
	.w3(32'h3b872a94),
	.w4(32'h3b63707d),
	.w5(32'hbb26d735),
	.w6(32'h3a6e3331),
	.w7(32'h3b27746f),
	.w8(32'h3a279b2c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ca87e),
	.w1(32'hbb031cfd),
	.w2(32'h3c39ac20),
	.w3(32'hbb30a8a5),
	.w4(32'hbbbc89c0),
	.w5(32'h3bcf0900),
	.w6(32'hbbd23e90),
	.w7(32'h3a9c0da3),
	.w8(32'h3a215b2b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18ae04),
	.w1(32'h3b004e6d),
	.w2(32'h3a93312d),
	.w3(32'h3b063853),
	.w4(32'h3ade76b4),
	.w5(32'h3a060e25),
	.w6(32'h3aad9e2d),
	.w7(32'h3b1aa240),
	.w8(32'hbbcb76d7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9691d8),
	.w1(32'hbbd52ae8),
	.w2(32'hbca0b308),
	.w3(32'hbbbdde41),
	.w4(32'hbc0691fb),
	.w5(32'hbd0762a7),
	.w6(32'hbbed911d),
	.w7(32'hbc45c8c8),
	.w8(32'hbce7a985),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0b97f),
	.w1(32'hbcb07b5c),
	.w2(32'h3b032758),
	.w3(32'hbd631265),
	.w4(32'hbd38cde2),
	.w5(32'h3b23a9d3),
	.w6(32'hbd43d88b),
	.w7(32'hbd13115e),
	.w8(32'h3b615b13),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba70888),
	.w1(32'h3b789188),
	.w2(32'h3aa85f38),
	.w3(32'h3bb5ed4d),
	.w4(32'h3b6d685a),
	.w5(32'h38c6dda8),
	.w6(32'h3b9d108e),
	.w7(32'h3ba14cec),
	.w8(32'hba58a302),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f10f8),
	.w1(32'hb9a54f91),
	.w2(32'h3b3339a2),
	.w3(32'h3a9427fb),
	.w4(32'hbb492949),
	.w5(32'h3c11ce37),
	.w6(32'hb94d37f1),
	.w7(32'hbbb06a89),
	.w8(32'h3ba0d07b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40839c),
	.w1(32'h3c424227),
	.w2(32'hb82f2d01),
	.w3(32'h3c6cd5d0),
	.w4(32'h3c77a8fe),
	.w5(32'h399ea3da),
	.w6(32'h3c56006b),
	.w7(32'h3c2ed144),
	.w8(32'hbb835021),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec6481),
	.w1(32'hb82a1b42),
	.w2(32'hbb1b24b5),
	.w3(32'hba949ee6),
	.w4(32'hbae1fcb7),
	.w5(32'h3b2b9631),
	.w6(32'hbba1eca5),
	.w7(32'hbbe1570f),
	.w8(32'hbab68f25),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b0cfa),
	.w1(32'h3a9c191b),
	.w2(32'h3b038fb3),
	.w3(32'h398f95b3),
	.w4(32'h3b0562e6),
	.w5(32'h3b8a4096),
	.w6(32'hba039b12),
	.w7(32'h3a799143),
	.w8(32'h3b91b562),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d32a3),
	.w1(32'h3ba39a21),
	.w2(32'hbc1bca69),
	.w3(32'h3bceca0e),
	.w4(32'h3bcd568c),
	.w5(32'hbc212c05),
	.w6(32'h3c007157),
	.w7(32'h3c0b50b9),
	.w8(32'hbc3e128f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4a983),
	.w1(32'hbbb4c9a2),
	.w2(32'h3bbabc4c),
	.w3(32'hbc4c95cb),
	.w4(32'hbca2ccb4),
	.w5(32'h3af23115),
	.w6(32'hbc143d9c),
	.w7(32'hbc23525f),
	.w8(32'hbb72f678),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84ba20),
	.w1(32'h3bb47a28),
	.w2(32'hba196a72),
	.w3(32'hba50533b),
	.w4(32'hbb8b74d5),
	.w5(32'h3ace44c7),
	.w6(32'hba6c6b68),
	.w7(32'hba0d7c0f),
	.w8(32'h3bfed28e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f3362),
	.w1(32'hba758867),
	.w2(32'h3b5d3429),
	.w3(32'h3b958285),
	.w4(32'h39cdfd5a),
	.w5(32'hbac2dff8),
	.w6(32'h3be21c11),
	.w7(32'h3bb311e7),
	.w8(32'hbb4130a2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac40668),
	.w1(32'h3b1bce30),
	.w2(32'h3ac1d72c),
	.w3(32'hbc15c2b7),
	.w4(32'hbbd38d1b),
	.w5(32'h3b058f44),
	.w6(32'hbc2a1828),
	.w7(32'hbbd181d6),
	.w8(32'hbb85fe56),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b220419),
	.w1(32'hbb6a3efd),
	.w2(32'hbc13bb5a),
	.w3(32'h3b9078b4),
	.w4(32'hbb6f007d),
	.w5(32'hbc27cbc6),
	.w6(32'hbbe547c9),
	.w7(32'hbc2c1529),
	.w8(32'hbbf5b74f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe13d9d),
	.w1(32'hbbd685da),
	.w2(32'h3be0ea2f),
	.w3(32'hbbf27f63),
	.w4(32'hbc0d7e13),
	.w5(32'hbae172e4),
	.w6(32'hbc0e49e1),
	.w7(32'hbbd087e7),
	.w8(32'h3b969a3f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24696c),
	.w1(32'h3bcdc7d8),
	.w2(32'h3bc8eeee),
	.w3(32'h3bb66a4f),
	.w4(32'hba7bea27),
	.w5(32'h3ba726ad),
	.w6(32'h3a41df65),
	.w7(32'h3b683488),
	.w8(32'h3b5e8ba6),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4a9c5),
	.w1(32'h3902b04b),
	.w2(32'h3b5352e2),
	.w3(32'h3bab93fa),
	.w4(32'h3b318e0a),
	.w5(32'hbb6bf2fc),
	.w6(32'h3afbf8d2),
	.w7(32'hbaacd62a),
	.w8(32'hb9ea9dc8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77d7b4),
	.w1(32'h3b9a79a5),
	.w2(32'h3b7cedf2),
	.w3(32'hbae59870),
	.w4(32'h3a896159),
	.w5(32'hba34b30e),
	.w6(32'hbad682b0),
	.w7(32'hb89edbe9),
	.w8(32'h3949b27b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc23cb2),
	.w1(32'h3c15f6b9),
	.w2(32'hbcbf2c5b),
	.w3(32'h3ba2bf52),
	.w4(32'h3ba0352c),
	.w5(32'hbc841156),
	.w6(32'h3bd7f3d3),
	.w7(32'h3ba0c2f2),
	.w8(32'hbcaecbb1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89ca7f),
	.w1(32'hbc98b87c),
	.w2(32'hbc07f515),
	.w3(32'hbaa93455),
	.w4(32'hbc159451),
	.w5(32'hbc441e64),
	.w6(32'hbc026878),
	.w7(32'hbc65ad36),
	.w8(32'hbc0010c7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2db7a6),
	.w1(32'hbbdd30d2),
	.w2(32'h3ba62568),
	.w3(32'hbc43ff00),
	.w4(32'hbc444732),
	.w5(32'h3c091d54),
	.w6(32'hbc6bbe2b),
	.w7(32'hbc119c44),
	.w8(32'h3b22ddad),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8479e),
	.w1(32'h3c1df396),
	.w2(32'hbb25b29f),
	.w3(32'h3bc1fca4),
	.w4(32'h3c401ff8),
	.w5(32'hbadbe658),
	.w6(32'h3bb7a422),
	.w7(32'h3a322d28),
	.w8(32'hba4be4ff),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb279a88),
	.w1(32'h3b02b3fc),
	.w2(32'hb9429f4c),
	.w3(32'hbb167589),
	.w4(32'h3bdd0c48),
	.w5(32'hbafe7cff),
	.w6(32'h3a4b340d),
	.w7(32'h3b4e03d2),
	.w8(32'h39ca57bb),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ed806),
	.w1(32'h3a398452),
	.w2(32'h3a154f09),
	.w3(32'hbb2699b2),
	.w4(32'hbaa53c7e),
	.w5(32'hbb415170),
	.w6(32'hb9abdec0),
	.w7(32'h3a4ab491),
	.w8(32'h3a67e3a1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca69ae),
	.w1(32'h3bfa193d),
	.w2(32'h3bb01905),
	.w3(32'h3bda22b8),
	.w4(32'h3b294d59),
	.w5(32'h3aac514c),
	.w6(32'h3c175b85),
	.w7(32'h3afd5ce2),
	.w8(32'h3ab59aa6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41f8d8),
	.w1(32'hba7beedc),
	.w2(32'hbb45d07b),
	.w3(32'hb78aba95),
	.w4(32'hbb7739ad),
	.w5(32'hbba38be7),
	.w6(32'hba9f5d11),
	.w7(32'hbbbe971d),
	.w8(32'hbb62198a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c02c1),
	.w1(32'hb9d96a61),
	.w2(32'h3b8d2f3b),
	.w3(32'hbbd64831),
	.w4(32'hbb6c695d),
	.w5(32'h3cd7a572),
	.w6(32'hbbba6bd9),
	.w7(32'hbb6bc9a8),
	.w8(32'h3cfb80e7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcb8d1),
	.w1(32'h3ba1b081),
	.w2(32'h3b8e8788),
	.w3(32'h3d2451c2),
	.w4(32'h3cdd8cd4),
	.w5(32'h3bdf248f),
	.w6(32'h3d3a0190),
	.w7(32'h3cff9a2e),
	.w8(32'h3b59a4d8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f50ce),
	.w1(32'h391bd843),
	.w2(32'hba796818),
	.w3(32'h3c7159e6),
	.w4(32'h3c46b401),
	.w5(32'h3a8e9ae1),
	.w6(32'h3bb8ae7b),
	.w7(32'hb99f677d),
	.w8(32'h3ac6c2f5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a902a00),
	.w1(32'h3a902aef),
	.w2(32'h3c2392aa),
	.w3(32'h3a630bfa),
	.w4(32'h3aa7c52c),
	.w5(32'h3ba20f94),
	.w6(32'h3ac57354),
	.w7(32'hba792ff8),
	.w8(32'h39f15db3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc96c3d),
	.w1(32'hbb8566c5),
	.w2(32'hba84a840),
	.w3(32'hbb89351b),
	.w4(32'hbb39de79),
	.w5(32'h3aecadd8),
	.w6(32'hba86f7b7),
	.w7(32'hbaa82536),
	.w8(32'hba6231d4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfdded),
	.w1(32'hbb6611af),
	.w2(32'h3be2871e),
	.w3(32'h3b00b862),
	.w4(32'h3ab304ff),
	.w5(32'h3ae4844b),
	.w6(32'h3b298a71),
	.w7(32'hba8d167f),
	.w8(32'h3aa9ba5f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd9454),
	.w1(32'h3bb65b8e),
	.w2(32'hbb8a9fb1),
	.w3(32'h3b36cfa2),
	.w4(32'h38b1f76a),
	.w5(32'hbb94dc60),
	.w6(32'hbba7aa57),
	.w7(32'hbb9baaf6),
	.w8(32'hb9cd5ce9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeced9b),
	.w1(32'hbbc6de66),
	.w2(32'h3ac71313),
	.w3(32'hbbcc8877),
	.w4(32'hbbd70e4a),
	.w5(32'h3c462e49),
	.w6(32'hbb502cd9),
	.w7(32'hbc0119cd),
	.w8(32'h3b18ac62),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cc4b9),
	.w1(32'h3b718fac),
	.w2(32'h3b067ab9),
	.w3(32'h3cac16ad),
	.w4(32'h3c8e1b18),
	.w5(32'h3ac14b73),
	.w6(32'h3c374808),
	.w7(32'h3bba21a8),
	.w8(32'hbb2d7ea8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98c984),
	.w1(32'h3b1f9934),
	.w2(32'hbb28f8e0),
	.w3(32'hbb12d229),
	.w4(32'h39da87eb),
	.w5(32'hba6343e6),
	.w6(32'h3a86420d),
	.w7(32'h3b58bfcb),
	.w8(32'hbb1021c5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a369aed),
	.w1(32'hbb26d177),
	.w2(32'hbb081e08),
	.w3(32'hbb1d9eef),
	.w4(32'hba5842a2),
	.w5(32'h3b871ae2),
	.w6(32'hbb3c4ca1),
	.w7(32'hbbb0663c),
	.w8(32'hbbd82c77),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7e544),
	.w1(32'hb9f3611a),
	.w2(32'hba6eb9b8),
	.w3(32'h3c43108c),
	.w4(32'h3c1ff1ba),
	.w5(32'h382441f3),
	.w6(32'hbb4d4291),
	.w7(32'hbb4509c3),
	.w8(32'h3b4ec537),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dcf00),
	.w1(32'hbb3a5eae),
	.w2(32'hba0681d8),
	.w3(32'h3b7500e6),
	.w4(32'h3b2ac58b),
	.w5(32'hbb25fcc1),
	.w6(32'h3c0604c7),
	.w7(32'h3bc471b5),
	.w8(32'hbb53637a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba858647),
	.w1(32'hbb37f65d),
	.w2(32'hb9c1626d),
	.w3(32'hbb0837d9),
	.w4(32'hbae7e5cd),
	.w5(32'h3c089f61),
	.w6(32'hbaeea7e2),
	.w7(32'hbb1ed323),
	.w8(32'h3be9bb8f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a316c2d),
	.w1(32'h3b8f6124),
	.w2(32'h3ba0e846),
	.w3(32'h3bfc7d89),
	.w4(32'h3b59676e),
	.w5(32'h3b8c33f8),
	.w6(32'h3c2135bf),
	.w7(32'h3bda8008),
	.w8(32'h3b463544),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf91fea),
	.w1(32'h3ba74b1d),
	.w2(32'hbba308f9),
	.w3(32'hbb86bec5),
	.w4(32'h3ae893f5),
	.w5(32'hbc1649f4),
	.w6(32'h3b9f892f),
	.w7(32'h3c363d3f),
	.w8(32'hbc0a1f99),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5f304),
	.w1(32'hb88372aa),
	.w2(32'h3baefe0d),
	.w3(32'hbbfd714e),
	.w4(32'hbb7d8d02),
	.w5(32'h3b6aa29e),
	.w6(32'hbc1b2bbe),
	.w7(32'hbb568c43),
	.w8(32'h3c72cec4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b908765),
	.w1(32'h3bfcc278),
	.w2(32'h3b31bdff),
	.w3(32'hba86c4c2),
	.w4(32'h3ba4a9cc),
	.w5(32'h3ac4acd9),
	.w6(32'h3ba89219),
	.w7(32'h3b0dbf35),
	.w8(32'h3af8ebc8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ddeb9),
	.w1(32'hbb17e56b),
	.w2(32'h388ec82b),
	.w3(32'h3ab6f6e3),
	.w4(32'hba4867da),
	.w5(32'hbbcab857),
	.w6(32'h3ab99395),
	.w7(32'hb944d2c4),
	.w8(32'hbc07d038),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce6df8),
	.w1(32'hbb6b8c8f),
	.w2(32'h3bc79a24),
	.w3(32'hbc8a250d),
	.w4(32'hbc135e73),
	.w5(32'h37cb3612),
	.w6(32'hbc06af5e),
	.w7(32'hbb7278da),
	.w8(32'h3b0988ac),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad60fb0),
	.w1(32'h381fe6aa),
	.w2(32'h3bb8d811),
	.w3(32'hbb994182),
	.w4(32'hbbbc9b65),
	.w5(32'hbac68244),
	.w6(32'h3aabc14f),
	.w7(32'h3bdbbdc1),
	.w8(32'h3b15a935),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6f29e),
	.w1(32'h3a89f211),
	.w2(32'h3b81388a),
	.w3(32'hbbad1ffc),
	.w4(32'hbb1218e8),
	.w5(32'h3b6b9357),
	.w6(32'hbb818dab),
	.w7(32'h3be3912a),
	.w8(32'hbad03eb0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a8953),
	.w1(32'h3abf718b),
	.w2(32'hbc26d35f),
	.w3(32'h3a84bb02),
	.w4(32'h3acdea18),
	.w5(32'hbc0dbd02),
	.w6(32'h3b323c7d),
	.w7(32'h3ac18fa0),
	.w8(32'hb77a8859),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb520a),
	.w1(32'hbc51f321),
	.w2(32'h3b977ee9),
	.w3(32'hbc090565),
	.w4(32'hbc266c4a),
	.w5(32'h3b902b6a),
	.w6(32'h3a1648f5),
	.w7(32'hbbd2d3e7),
	.w8(32'h3b38622a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be49e4a),
	.w1(32'h3bd05dea),
	.w2(32'h3a891c8a),
	.w3(32'h38fd626f),
	.w4(32'h3b824fc3),
	.w5(32'h3bd5c680),
	.w6(32'h3bf980a5),
	.w7(32'h3c1f3c1c),
	.w8(32'h3bfc5586),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38c570),
	.w1(32'h3a8c6180),
	.w2(32'h3b715d66),
	.w3(32'h3b9a88d0),
	.w4(32'h3a9c21f3),
	.w5(32'hbc41aa8c),
	.w6(32'h3b8e8c26),
	.w7(32'hbb46c7d0),
	.w8(32'hbbbe4d75),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb45bb2),
	.w1(32'h3a834d9e),
	.w2(32'h3b84313c),
	.w3(32'hbbfd2539),
	.w4(32'hba2b1656),
	.w5(32'h39ff05b8),
	.w6(32'hbb17db9d),
	.w7(32'hb7836d0d),
	.w8(32'h3ad093f4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf54f2),
	.w1(32'hb9d3b2f4),
	.w2(32'h3a049322),
	.w3(32'hbb3c7219),
	.w4(32'hbb943c99),
	.w5(32'h3ba4a2e8),
	.w6(32'hbb8e53aa),
	.w7(32'hbb02c372),
	.w8(32'h3c075856),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b063f51),
	.w1(32'hbbf5061b),
	.w2(32'h39eb2f35),
	.w3(32'h3babd7e8),
	.w4(32'hbb3764d1),
	.w5(32'hbbcf1c23),
	.w6(32'h3c3001ae),
	.w7(32'h3af24372),
	.w8(32'hbbfbe177),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2df146),
	.w1(32'hbad2bd03),
	.w2(32'hbc15815f),
	.w3(32'hbbc56092),
	.w4(32'hbbb2d499),
	.w5(32'hbafb6df3),
	.w6(32'hbbed94b2),
	.w7(32'hbc1aff80),
	.w8(32'hbc154f96),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58918e),
	.w1(32'hbbd6771a),
	.w2(32'hbb0329c6),
	.w3(32'hba5ba8fe),
	.w4(32'hb944f9b8),
	.w5(32'hbc5e1240),
	.w6(32'hbc208972),
	.w7(32'hbbdd7aa2),
	.w8(32'hbb239e6a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c4cc7),
	.w1(32'hbbe6a93e),
	.w2(32'h3c28de51),
	.w3(32'hbca145a4),
	.w4(32'hbbb6526e),
	.w5(32'h3c4eb9a2),
	.w6(32'hbc89f08e),
	.w7(32'hbbd4fd4a),
	.w8(32'h3c4e22ce),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98e1b5),
	.w1(32'h3c592fde),
	.w2(32'hbab31522),
	.w3(32'h3cbba792),
	.w4(32'h3c8bd80e),
	.w5(32'h3ad2c46b),
	.w6(32'h3c0b3024),
	.w7(32'h3c092d65),
	.w8(32'hbb58507f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea9cb7),
	.w1(32'hbab78cdd),
	.w2(32'hbbb4a4a2),
	.w3(32'h3b007951),
	.w4(32'h3b92a5fa),
	.w5(32'hbb5b3c1f),
	.w6(32'hbb9ecedb),
	.w7(32'hbbcb9b7f),
	.w8(32'hbb2c3f4a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07f23e),
	.w1(32'hbbd77c29),
	.w2(32'h3b02984f),
	.w3(32'hbbb68109),
	.w4(32'hbbddae84),
	.w5(32'h3b3c8bc3),
	.w6(32'hbadc5645),
	.w7(32'hbba9429e),
	.w8(32'h3ba5f3eb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b111545),
	.w1(32'h3ab4961f),
	.w2(32'hb9ecf4ce),
	.w3(32'h3b320607),
	.w4(32'h3b733f52),
	.w5(32'h37372ae8),
	.w6(32'h3bc01e99),
	.w7(32'h3bd66f8a),
	.w8(32'hba66e62f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bcc670),
	.w1(32'hb9fb48ba),
	.w2(32'h3ad65a24),
	.w3(32'h3a993eaa),
	.w4(32'h3aebb5f2),
	.w5(32'hba4b9ca9),
	.w6(32'h3a11c216),
	.w7(32'hb9f79922),
	.w8(32'h3b59ede7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6401a8),
	.w1(32'hbb1a2d49),
	.w2(32'h3c422858),
	.w3(32'hba73af72),
	.w4(32'hbaa258aa),
	.w5(32'h3c66a17c),
	.w6(32'hbb56c8c2),
	.w7(32'h3b8c3b60),
	.w8(32'h3c476731),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89fc92),
	.w1(32'h3c1b512b),
	.w2(32'hbb6d03fc),
	.w3(32'h3c2df10b),
	.w4(32'h3c57d97a),
	.w5(32'hbb945e38),
	.w6(32'h3c38ac50),
	.w7(32'h3c1baf09),
	.w8(32'hbb88902d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb793c82),
	.w1(32'hbbb51acc),
	.w2(32'h3b3c4e98),
	.w3(32'hbba3feaf),
	.w4(32'hbbcd9aef),
	.w5(32'h3b5a3303),
	.w6(32'hbb94a4bb),
	.w7(32'hbbb51912),
	.w8(32'h3a8bdbba),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f79bd9),
	.w1(32'h3abe0176),
	.w2(32'h3b344c2f),
	.w3(32'h3ab98bf7),
	.w4(32'h3b92e36b),
	.w5(32'h3a982515),
	.w6(32'h3ad271f9),
	.w7(32'h3b5840c7),
	.w8(32'h3a2c68fc),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfd306),
	.w1(32'h3a5bed68),
	.w2(32'hbb92d397),
	.w3(32'hbac6750b),
	.w4(32'h3a19959d),
	.w5(32'hbb8821b4),
	.w6(32'hb9ef3022),
	.w7(32'h3b842fa7),
	.w8(32'h3985981f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31ccd1),
	.w1(32'hba8ba0ff),
	.w2(32'hba9d53f5),
	.w3(32'hbaf7ba59),
	.w4(32'h3b3db259),
	.w5(32'hbcbfd931),
	.w6(32'hbbfb126c),
	.w7(32'h39cd6634),
	.w8(32'hbcafebe3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc061857),
	.w1(32'hbbc8ec73),
	.w2(32'hbaacb195),
	.w3(32'hbd187169),
	.w4(32'hbd0b9635),
	.w5(32'hbb1da765),
	.w6(32'hbcff8824),
	.w7(32'hbcd7c93c),
	.w8(32'hbb32751f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dbd5e),
	.w1(32'hbb98c7e0),
	.w2(32'h3b460b41),
	.w3(32'hbb9fa64a),
	.w4(32'hbba69545),
	.w5(32'h388d857c),
	.w6(32'hbb8f00b4),
	.w7(32'hbb645593),
	.w8(32'hbb9f8d49),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02eebb),
	.w1(32'h3bbb405c),
	.w2(32'h3b7ee994),
	.w3(32'h3b51f0ee),
	.w4(32'h3b6e537c),
	.w5(32'hbabe3d11),
	.w6(32'hbb16c677),
	.w7(32'h3adc8808),
	.w8(32'hbbc36cfd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b2147),
	.w1(32'h38d06612),
	.w2(32'hbb9856b4),
	.w3(32'hbc0cfb5f),
	.w4(32'hbb6fee6d),
	.w5(32'h3b2ed439),
	.w6(32'hbc47e06a),
	.w7(32'hbb341a57),
	.w8(32'hbbaf1e13),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98437c2),
	.w1(32'h3a0b8e06),
	.w2(32'hbb28f5f5),
	.w3(32'h3bc54629),
	.w4(32'h3b8f0a2d),
	.w5(32'hbb4d572e),
	.w6(32'hbb766495),
	.w7(32'hbb3be07a),
	.w8(32'h3a309f71),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadcae3),
	.w1(32'hb7a6df36),
	.w2(32'hb9f1e83c),
	.w3(32'hbc7e49d2),
	.w4(32'hbb835744),
	.w5(32'hbb9037cb),
	.w6(32'hbba900f9),
	.w7(32'hbb9818ab),
	.w8(32'h3a2ea3f1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86fc2c6),
	.w1(32'h3a29035b),
	.w2(32'h3b2ffa0a),
	.w3(32'hbb83f5b9),
	.w4(32'hbb9e4566),
	.w5(32'h3a820a42),
	.w6(32'h3a55ff70),
	.w7(32'h3ae86f05),
	.w8(32'h3b80adea),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb871a80),
	.w1(32'hbbad100d),
	.w2(32'hbad7c4d2),
	.w3(32'hba70083b),
	.w4(32'hba103f51),
	.w5(32'hbad33dc5),
	.w6(32'h3aee7fa3),
	.w7(32'h394f611a),
	.w8(32'hbae62184),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7f63e),
	.w1(32'h3ae05f5b),
	.w2(32'hba387659),
	.w3(32'hb88ba9dd),
	.w4(32'h3aa6ee01),
	.w5(32'hb9be81f5),
	.w6(32'hb97af18d),
	.w7(32'h3a850cbc),
	.w8(32'h3b5760bb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb56b7c),
	.w1(32'h3a8b8323),
	.w2(32'h3b9ce324),
	.w3(32'hbb813de1),
	.w4(32'h3b427d46),
	.w5(32'hbb438704),
	.w6(32'hbb981e53),
	.w7(32'h3ad178f3),
	.w8(32'h3c29e809),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb082c81),
	.w1(32'h3c0d5bcf),
	.w2(32'h39e36aec),
	.w3(32'hbc2577f8),
	.w4(32'hbb417129),
	.w5(32'hbb296f35),
	.w6(32'hbbaa6413),
	.w7(32'hbbba1c5a),
	.w8(32'h3b17c727),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a485083),
	.w1(32'h3b8cac96),
	.w2(32'h3bd80c34),
	.w3(32'h3bcedd9c),
	.w4(32'h3b059674),
	.w5(32'h3921cfe1),
	.w6(32'h3b2c8cc1),
	.w7(32'h3b306101),
	.w8(32'hbadf5642),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b6aa4),
	.w1(32'h3bbc4fe7),
	.w2(32'h3a998620),
	.w3(32'hbba01496),
	.w4(32'h3bddfa2b),
	.w5(32'h3b36c7d4),
	.w6(32'h3b2a8e2a),
	.w7(32'h3c33ec83),
	.w8(32'h3b69f43f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5312d0),
	.w1(32'h3a5f2346),
	.w2(32'hb8abee6e),
	.w3(32'h3b895f5a),
	.w4(32'h3b5a36d9),
	.w5(32'hbb0b402d),
	.w6(32'h3b316769),
	.w7(32'h3b5b40aa),
	.w8(32'hbb5043c6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aad621),
	.w1(32'hba6a1c20),
	.w2(32'h3c0bb912),
	.w3(32'hbb5cfbcc),
	.w4(32'hbb1b9fd5),
	.w5(32'hbb0dfe85),
	.w6(32'hbb0701d3),
	.w7(32'hbb175520),
	.w8(32'hbb0374d5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99dba5),
	.w1(32'hba4d96f7),
	.w2(32'hbbd976e6),
	.w3(32'hbbf234e1),
	.w4(32'hbbfdee6c),
	.w5(32'h3c1532ae),
	.w6(32'hbb06ea61),
	.w7(32'hbb727e7f),
	.w8(32'h3b568266),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a220e75),
	.w1(32'hbc33c90e),
	.w2(32'h3b3173e1),
	.w3(32'h3c8421d5),
	.w4(32'h3bbb8de9),
	.w5(32'h3bcbedfb),
	.w6(32'h3c93a706),
	.w7(32'h3c0ab1b8),
	.w8(32'h3ba8cc61),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98c238),
	.w1(32'hbb2d7a3b),
	.w2(32'hbbb24041),
	.w3(32'h3bff2c2b),
	.w4(32'hba33968f),
	.w5(32'h3b935c0c),
	.w6(32'h3be7a328),
	.w7(32'hba7a453c),
	.w8(32'h3bc6bd97),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01a1a4),
	.w1(32'hbb227443),
	.w2(32'h3b1d49ed),
	.w3(32'h3c596152),
	.w4(32'h3bfee000),
	.w5(32'hb7a03e51),
	.w6(32'h3c215709),
	.w7(32'h3b2194bf),
	.w8(32'hbb09eb9d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986288d),
	.w1(32'h3b044f09),
	.w2(32'hbaa5ed40),
	.w3(32'hba58a291),
	.w4(32'h3aafb604),
	.w5(32'hbb7a04d4),
	.w6(32'hbb01e410),
	.w7(32'hb9271e15),
	.w8(32'hbba17613),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f4b98),
	.w1(32'hbad86fa4),
	.w2(32'h3c898ad0),
	.w3(32'hbbb2b9df),
	.w4(32'hbb6edef9),
	.w5(32'h3c5cc163),
	.w6(32'hbbc7f1a3),
	.w7(32'hbb81e8f9),
	.w8(32'h3c29008c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f8445),
	.w1(32'h3c2007fa),
	.w2(32'hbba54be8),
	.w3(32'h3c870908),
	.w4(32'h3c84b5d0),
	.w5(32'h3b66f6f0),
	.w6(32'h3c7b6ffc),
	.w7(32'h3c85d499),
	.w8(32'h3b073650),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cf55b),
	.w1(32'h3b6d053e),
	.w2(32'h3b9eec51),
	.w3(32'h3ac2638d),
	.w4(32'h3b80d3b7),
	.w5(32'hbb98b65e),
	.w6(32'h3b7181d7),
	.w7(32'h3ab8c406),
	.w8(32'hbba1f241),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b962b1e),
	.w1(32'h3bfcab97),
	.w2(32'hbb0dc084),
	.w3(32'hbb9bfbce),
	.w4(32'hbb0a5690),
	.w5(32'hbbfcb68c),
	.w6(32'hbb3066b0),
	.w7(32'h3bab6733),
	.w8(32'hbb59d2e6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26e9da),
	.w1(32'h3c33ca0c),
	.w2(32'hbbaf9443),
	.w3(32'hbbca2a65),
	.w4(32'h3b182c89),
	.w5(32'h3b377456),
	.w6(32'hbb17ccdd),
	.w7(32'h3aaa39c3),
	.w8(32'h3c08ba49),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcd7ec),
	.w1(32'hbc01ebb8),
	.w2(32'h3b98f15f),
	.w3(32'h3c829b7d),
	.w4(32'h3c0d63f6),
	.w5(32'h3bf71d14),
	.w6(32'h3c87ae65),
	.w7(32'h3c2335cd),
	.w8(32'h3b85fbf3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b723b),
	.w1(32'hba2d61e6),
	.w2(32'h3b235dae),
	.w3(32'h3becee04),
	.w4(32'h3a0c5309),
	.w5(32'h3bd8786b),
	.w6(32'h3bc94b61),
	.w7(32'hba9c0b9f),
	.w8(32'h3ba043cd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcf632),
	.w1(32'h3859b88d),
	.w2(32'hb9ed4247),
	.w3(32'h3ca6b2f6),
	.w4(32'h3c4f88fe),
	.w5(32'h3c124f2f),
	.w6(32'h3c397448),
	.w7(32'h39b724d3),
	.w8(32'h3c5cce14),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab72e91),
	.w1(32'hbbbc246a),
	.w2(32'h38fe4b97),
	.w3(32'h3c41af0b),
	.w4(32'h3a25d4cd),
	.w5(32'hbb4b572b),
	.w6(32'h3c816959),
	.w7(32'h3c1abd96),
	.w8(32'hbae80bd2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8beea),
	.w1(32'hb9c2746a),
	.w2(32'h3b6b036d),
	.w3(32'hbb449e0d),
	.w4(32'hbb4c66fd),
	.w5(32'h3b8be5ca),
	.w6(32'hbbe18176),
	.w7(32'hbbfa3ed0),
	.w8(32'h3bc75fb9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f3ecb),
	.w1(32'h3a39d97f),
	.w2(32'h3b46c292),
	.w3(32'h3b14370b),
	.w4(32'h392d1e1c),
	.w5(32'h3a3ec932),
	.w6(32'h3ba1f3c8),
	.w7(32'h39a9f0de),
	.w8(32'h3b7b1538),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba903e3b),
	.w1(32'h3b08599f),
	.w2(32'h3b7d3c79),
	.w3(32'hba676f47),
	.w4(32'hbae177ff),
	.w5(32'h3b854193),
	.w6(32'h3bead329),
	.w7(32'h3ab0dbe6),
	.w8(32'h3b995c6c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20ecd8),
	.w1(32'h3b0cf6b6),
	.w2(32'h3baca8a5),
	.w3(32'h3b1240b0),
	.w4(32'h3b02db11),
	.w5(32'h3ba6dbbe),
	.w6(32'h3b88b7ba),
	.w7(32'h3b555bed),
	.w8(32'h3bbcd5ec),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e1cc9),
	.w1(32'h3b86b1c6),
	.w2(32'h3aef518c),
	.w3(32'h3b7266f6),
	.w4(32'h3bb7c9f0),
	.w5(32'hbb1a7044),
	.w6(32'h3ba77615),
	.w7(32'h3bd4050a),
	.w8(32'hbb4fe557),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba523329),
	.w1(32'hbb537d84),
	.w2(32'h3acb3204),
	.w3(32'hbb91fc2f),
	.w4(32'hbbe4e125),
	.w5(32'h3ab28283),
	.w6(32'hbb0b792e),
	.w7(32'hbab52842),
	.w8(32'h3af3612b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06f635),
	.w1(32'h3ba81174),
	.w2(32'h3bcebae1),
	.w3(32'h3aba09af),
	.w4(32'hbb308d8a),
	.w5(32'h3c71305f),
	.w6(32'h3be4b37a),
	.w7(32'h3a3161fb),
	.w8(32'h3c516582),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9c350),
	.w1(32'h3b79fcea),
	.w2(32'h3ac2e97e),
	.w3(32'h3ca0e1e8),
	.w4(32'h3c69eda7),
	.w5(32'hbbcfaaaf),
	.w6(32'h3c868af9),
	.w7(32'h3c8d94d6),
	.w8(32'hbb52177a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52a68e),
	.w1(32'h3b9e50ef),
	.w2(32'hbabda963),
	.w3(32'hbc3f1f50),
	.w4(32'hbb0003bd),
	.w5(32'hbc1fda9d),
	.w6(32'hbc169e27),
	.w7(32'hbbf855ff),
	.w8(32'hbbbef8c6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a088d),
	.w1(32'hbb5ead52),
	.w2(32'h3b5a07df),
	.w3(32'hbc802d76),
	.w4(32'hbbd3dc12),
	.w5(32'h3aae0dce),
	.w6(32'hbc23dc7e),
	.w7(32'hbb9918e6),
	.w8(32'hbb71603f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdbfaa),
	.w1(32'h3ad8a7b6),
	.w2(32'hbad43bdb),
	.w3(32'hbbbe8669),
	.w4(32'hbaf7c12c),
	.w5(32'h3c1318b6),
	.w6(32'hbbd9c74a),
	.w7(32'hbb26b09c),
	.w8(32'h3c2e77a5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb268498),
	.w1(32'hbab1f8a2),
	.w2(32'h3baf67d8),
	.w3(32'h3c427afc),
	.w4(32'h3b82399e),
	.w5(32'h3bb5e516),
	.w6(32'h3ca00389),
	.w7(32'h3c8a5fce),
	.w8(32'h39eef39b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2adca),
	.w1(32'h3b87e3fc),
	.w2(32'h3b176ebc),
	.w3(32'h3c44c634),
	.w4(32'h3c00dadd),
	.w5(32'hbb3833e5),
	.w6(32'h39216bc4),
	.w7(32'hbb3fcfb9),
	.w8(32'hbb0b65b4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abffdea),
	.w1(32'h3b05b08c),
	.w2(32'hbbecec32),
	.w3(32'hbb94cefd),
	.w4(32'hbbb4c37d),
	.w5(32'h3b549958),
	.w6(32'hbb04c616),
	.w7(32'hbb858527),
	.w8(32'h3c07d8eb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0716ee),
	.w1(32'hbbd06188),
	.w2(32'h3aa62323),
	.w3(32'hbb0cf19b),
	.w4(32'hbb79b0c8),
	.w5(32'hbb28a886),
	.w6(32'h3ba4349b),
	.w7(32'h3b871c72),
	.w8(32'hbb9d2761),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bbb8f),
	.w1(32'h398ec65e),
	.w2(32'h3c19e881),
	.w3(32'hb9c1f069),
	.w4(32'hb9cd35de),
	.w5(32'h3ca5e66f),
	.w6(32'hbb7f2c8f),
	.w7(32'hbbd3785b),
	.w8(32'h3ccf4824),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73497e),
	.w1(32'h3c058215),
	.w2(32'h3ac18258),
	.w3(32'h3d0de58d),
	.w4(32'h3c8844a1),
	.w5(32'h3b8d10d3),
	.w6(32'h3d02763c),
	.w7(32'h3cd21b7a),
	.w8(32'h3b05c221),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e37ef),
	.w1(32'hbb8d729f),
	.w2(32'h3c096a71),
	.w3(32'h3b2538b3),
	.w4(32'hbbae542d),
	.w5(32'h3c567f64),
	.w6(32'h3bfd1662),
	.w7(32'hbb47d56e),
	.w8(32'h3bdad9f7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e98c9),
	.w1(32'h3c17113b),
	.w2(32'hbadc84cd),
	.w3(32'h3c26d300),
	.w4(32'h3c4e02f9),
	.w5(32'hbb1a6f33),
	.w6(32'h3bdf3a75),
	.w7(32'h3c2a918f),
	.w8(32'hbb8249a6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d3ecf),
	.w1(32'hbb2313c7),
	.w2(32'hba92349b),
	.w3(32'hbb5ff904),
	.w4(32'hbb6420fe),
	.w5(32'hba79824c),
	.w6(32'hbbab4757),
	.w7(32'hbba6456e),
	.w8(32'hba73daad),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39858aa0),
	.w1(32'h3b020014),
	.w2(32'h3baea47b),
	.w3(32'hbabd7180),
	.w4(32'h3a178a0d),
	.w5(32'h3b65d349),
	.w6(32'hbab3c67d),
	.w7(32'h3adf791f),
	.w8(32'h3c184434),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c101c75),
	.w1(32'h3c7af603),
	.w2(32'h39bb2d5a),
	.w3(32'hbbf8820b),
	.w4(32'hbb2da1ed),
	.w5(32'hbb17d6ba),
	.w6(32'hbb9ce9c6),
	.w7(32'hbb434efe),
	.w8(32'hb8f61808),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac21a28),
	.w1(32'h3b21d21e),
	.w2(32'h3b97baaa),
	.w3(32'hb9919726),
	.w4(32'hb800d7ba),
	.w5(32'hbb2092fb),
	.w6(32'hba3b6da4),
	.w7(32'hbaeef5ea),
	.w8(32'h3979a7d4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e7f14),
	.w1(32'hbb0f323a),
	.w2(32'hbabbe876),
	.w3(32'hbbae3ec4),
	.w4(32'hbbcc1e81),
	.w5(32'hbba42de2),
	.w6(32'h3a4bc376),
	.w7(32'h3c0bbff6),
	.w8(32'hba5d89f1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed4450),
	.w1(32'hbaccd779),
	.w2(32'hbb850817),
	.w3(32'hbc0ea09e),
	.w4(32'hbc088190),
	.w5(32'h37676d80),
	.w6(32'hbaee7615),
	.w7(32'hba461b23),
	.w8(32'h3b07326e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05c2f3),
	.w1(32'hbbd7fc59),
	.w2(32'h3bcf21b8),
	.w3(32'hba58b0a2),
	.w4(32'hbb4f4c91),
	.w5(32'h3b622674),
	.w6(32'hbb84ca17),
	.w7(32'h3b57beaa),
	.w8(32'h3c00c91b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dc51d),
	.w1(32'h3bbf286e),
	.w2(32'h3c2bb2b8),
	.w3(32'h3c0f7b01),
	.w4(32'h3c1f0d49),
	.w5(32'h3b564529),
	.w6(32'h3b4be3e9),
	.w7(32'h3c0a552f),
	.w8(32'h3bce9a7d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c378650),
	.w1(32'h3c20f29e),
	.w2(32'hbb7ee9af),
	.w3(32'h39d55087),
	.w4(32'h3c113d40),
	.w5(32'hbaf3a606),
	.w6(32'h3b8e21ee),
	.w7(32'h3b1b26ac),
	.w8(32'hbbab4e50),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe97973),
	.w1(32'h3ac1d8fd),
	.w2(32'hba3d957e),
	.w3(32'hbbfc45fb),
	.w4(32'hbb846480),
	.w5(32'hbba4b3c0),
	.w6(32'hbb103695),
	.w7(32'hbbb68896),
	.w8(32'h3ac54622),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2f797),
	.w1(32'h3a31faa0),
	.w2(32'h3b0788df),
	.w3(32'hbbd07517),
	.w4(32'hbb921de1),
	.w5(32'hb9080eed),
	.w6(32'hbbfa6999),
	.w7(32'hbbd5ce16),
	.w8(32'h3b2be280),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba32586),
	.w1(32'hbbab7124),
	.w2(32'hbc315c1a),
	.w3(32'h3b81194e),
	.w4(32'h3b8e46f6),
	.w5(32'hbc13a89e),
	.w6(32'h3c0d62fa),
	.w7(32'h3c0f57f6),
	.w8(32'hbc05ee6a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfc223),
	.w1(32'hba40de15),
	.w2(32'hbac44e83),
	.w3(32'hbc24bdcf),
	.w4(32'hbc1bdd0d),
	.w5(32'hbb71aaff),
	.w6(32'hbb98a29a),
	.w7(32'hba99712e),
	.w8(32'hbb9f8597),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9efea1),
	.w1(32'h37b0ac1d),
	.w2(32'hbb1102fe),
	.w3(32'hbb9ac342),
	.w4(32'hbb51879b),
	.w5(32'hbbcae2c1),
	.w6(32'hbbacf52a),
	.w7(32'hbb06b5cf),
	.w8(32'h3925e9d8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ddf5c),
	.w1(32'hbb9002a4),
	.w2(32'h3aacdcd4),
	.w3(32'hbb74d7fe),
	.w4(32'hbb9323f0),
	.w5(32'hbb73faee),
	.w6(32'h3a3f2263),
	.w7(32'hbb2ba49b),
	.w8(32'hbbccaf99),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a894901),
	.w1(32'hbb3dd064),
	.w2(32'hbaa2d751),
	.w3(32'hbb9050dc),
	.w4(32'hbb14eaff),
	.w5(32'h3bcc5c59),
	.w6(32'hb98ba1a6),
	.w7(32'hbb0846f7),
	.w8(32'h3b43ca52),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c366079),
	.w1(32'h3ba21677),
	.w2(32'hb904cc12),
	.w3(32'h3c8f59e8),
	.w4(32'h3c208e2b),
	.w5(32'h3ae06649),
	.w6(32'h3c61c478),
	.w7(32'h3b6f4e46),
	.w8(32'h3b02bd94),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f60ff),
	.w1(32'h3b3756dc),
	.w2(32'hbc0d1a0b),
	.w3(32'h3b4e3a30),
	.w4(32'h3b4e406d),
	.w5(32'hbc146fbf),
	.w6(32'h3b1b5538),
	.w7(32'h3b3d56de),
	.w8(32'hbb83ec96),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d90ce),
	.w1(32'hbb80fcdc),
	.w2(32'h3addc272),
	.w3(32'hbc186602),
	.w4(32'hbbe58a9f),
	.w5(32'h3b2e569a),
	.w6(32'hbc2f1c8c),
	.w7(32'hbc23a5c7),
	.w8(32'h3a3ada9a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc172a),
	.w1(32'h3a84538b),
	.w2(32'h3bb53f63),
	.w3(32'h3a3df490),
	.w4(32'h3a98b279),
	.w5(32'hbbebe5d3),
	.w6(32'hba83ed96),
	.w7(32'h38cac65b),
	.w8(32'hbacb89f6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b61287),
	.w1(32'h3b9faa8d),
	.w2(32'hbb114481),
	.w3(32'hbb1c2f33),
	.w4(32'h3b771c8c),
	.w5(32'hbb8b5451),
	.w6(32'h3ab08e2f),
	.w7(32'h3bdd1ede),
	.w8(32'hbb015c1c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cb41a),
	.w1(32'hbbddb3a5),
	.w2(32'hbb288020),
	.w3(32'hbba68fc6),
	.w4(32'hbba0a3d6),
	.w5(32'hba761dfa),
	.w6(32'hba69424e),
	.w7(32'h3aa9e748),
	.w8(32'hbc040d5c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2c9c4),
	.w1(32'hbbae5403),
	.w2(32'hb9ad298d),
	.w3(32'hbad485c3),
	.w4(32'hbb0caadc),
	.w5(32'h3a201504),
	.w6(32'hbc003d20),
	.w7(32'hbc122491),
	.w8(32'h3814b8d6),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e12c4),
	.w1(32'h3a9b66aa),
	.w2(32'hbb8f7375),
	.w3(32'h3a724f60),
	.w4(32'h3a897c68),
	.w5(32'hba3111e2),
	.w6(32'h39415fc3),
	.w7(32'h3a5ceddc),
	.w8(32'h3b301539),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb860cc9),
	.w1(32'hbc0da9b3),
	.w2(32'hb97f5438),
	.w3(32'hba66b8cc),
	.w4(32'hbbf21ef0),
	.w5(32'hbb058b03),
	.w6(32'h3b980d33),
	.w7(32'h3a33ed71),
	.w8(32'h3b56c552),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa243c9),
	.w1(32'h3a84fc66),
	.w2(32'hbb006254),
	.w3(32'h3b29f392),
	.w4(32'hbae16389),
	.w5(32'hbbe82eb9),
	.w6(32'hba1dfa14),
	.w7(32'h3b09518b),
	.w8(32'hbb360cb3),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81f44e),
	.w1(32'h3b9f180b),
	.w2(32'hba434aa0),
	.w3(32'hbbd8881f),
	.w4(32'hb8248319),
	.w5(32'h3b513930),
	.w6(32'hbbbdb0df),
	.w7(32'hbb9e5d32),
	.w8(32'h3b862043),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a031190),
	.w1(32'hba8a7da4),
	.w2(32'h3b70d287),
	.w3(32'h3b3b1692),
	.w4(32'h3b0a288d),
	.w5(32'hbb4d6ee8),
	.w6(32'h3b5c752e),
	.w7(32'h3ab7d00a),
	.w8(32'h3bbd3d2d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02631f),
	.w1(32'h3bce41c5),
	.w2(32'hbc03fcc6),
	.w3(32'h3b8f7ace),
	.w4(32'h3c4db5e0),
	.w5(32'hbc25b10e),
	.w6(32'h39a58988),
	.w7(32'hba8d650a),
	.w8(32'hbc183da2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae65f3),
	.w1(32'hbb88e77d),
	.w2(32'hbb376654),
	.w3(32'hbc69dc38),
	.w4(32'hbc24927c),
	.w5(32'hbb01f30a),
	.w6(32'hbc3ff957),
	.w7(32'hbb67e67d),
	.w8(32'hbb5a5cfe),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b9026),
	.w1(32'hbad105e5),
	.w2(32'h3bc0b9aa),
	.w3(32'hbb58fb45),
	.w4(32'hbb0dcb45),
	.w5(32'h3b0ed5aa),
	.w6(32'hbba059b4),
	.w7(32'hbb53f66d),
	.w8(32'h3b436e09),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2d543),
	.w1(32'hbaf80eb3),
	.w2(32'h3bac72c1),
	.w3(32'hbb3909bc),
	.w4(32'hbb4cf040),
	.w5(32'h3b9981b5),
	.w6(32'h39c95a08),
	.w7(32'h3b701fef),
	.w8(32'h3c0b4426),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0ce9f),
	.w1(32'h39509f2d),
	.w2(32'hba04a4ed),
	.w3(32'h3b246bde),
	.w4(32'h3b49b581),
	.w5(32'hbb1495ed),
	.w6(32'h3b9ca7dc),
	.w7(32'h3b364f4c),
	.w8(32'h38e08445),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3ad88),
	.w1(32'h3ab4f945),
	.w2(32'h39f0025a),
	.w3(32'hbc011ef9),
	.w4(32'hbbd8e6ae),
	.w5(32'h3b6bb194),
	.w6(32'hbc22d4ef),
	.w7(32'hbba7d72b),
	.w8(32'h3a9faf13),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7c608),
	.w1(32'h3a5e68c5),
	.w2(32'hbb15d75c),
	.w3(32'h3bca59b0),
	.w4(32'h3b7c144a),
	.w5(32'hbc27b983),
	.w6(32'h3b72cc56),
	.w7(32'h3ac7af04),
	.w8(32'hbc1c5f3c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6bc0f),
	.w1(32'hba236221),
	.w2(32'h39e63795),
	.w3(32'hbc1bbbdd),
	.w4(32'h3a521c4d),
	.w5(32'h3bef07ac),
	.w6(32'hbba3c244),
	.w7(32'h3c0d1923),
	.w8(32'h3c10c000),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad58241),
	.w1(32'h3c7968da),
	.w2(32'h3b2a5e8a),
	.w3(32'hbbccf304),
	.w4(32'h3b9ab96a),
	.w5(32'h3af2ec3b),
	.w6(32'hbb7cfbea),
	.w7(32'hbb94ddd8),
	.w8(32'h384a8c62),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99bbf49),
	.w1(32'hbb2525ca),
	.w2(32'h3a4f398f),
	.w3(32'h395e03a3),
	.w4(32'hbada3a66),
	.w5(32'h3c4c1a28),
	.w6(32'hba81dd34),
	.w7(32'hbb27f32e),
	.w8(32'h3b2cdd83),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9f81a),
	.w1(32'hba3d6a5e),
	.w2(32'h3b673deb),
	.w3(32'h3caa7fa3),
	.w4(32'h3c3cc8c1),
	.w5(32'h3c322784),
	.w6(32'h3c21e9cf),
	.w7(32'h3bbc8f74),
	.w8(32'h3c79e6eb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af25781),
	.w1(32'hb9976924),
	.w2(32'h3be8e5c9),
	.w3(32'h3c06d697),
	.w4(32'hbb205b65),
	.w5(32'h3baa26f9),
	.w6(32'h3c1e3ad2),
	.w7(32'h3b0a5463),
	.w8(32'h3b6fc7a2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4df061),
	.w1(32'hba32d955),
	.w2(32'hbbce4c7c),
	.w3(32'hba628421),
	.w4(32'hbb8343d5),
	.w5(32'hbc4589a9),
	.w6(32'hba8d3953),
	.w7(32'hbba76909),
	.w8(32'hbc0d69c1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bfa3f),
	.w1(32'hbb8923dc),
	.w2(32'h38db176e),
	.w3(32'hbb324876),
	.w4(32'h3bd95cbb),
	.w5(32'hbaffe436),
	.w6(32'hba486bee),
	.w7(32'h3c44e919),
	.w8(32'hbae15a0d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e143d),
	.w1(32'hbaa58f47),
	.w2(32'h3bdccf56),
	.w3(32'hbb7bb991),
	.w4(32'hbb9b2e7c),
	.w5(32'hbb7d9fd5),
	.w6(32'hbb9c292e),
	.w7(32'hbbcd762d),
	.w8(32'hbab2e775),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95f203),
	.w1(32'hbb916c26),
	.w2(32'h3b889df3),
	.w3(32'hbc122cd7),
	.w4(32'hbbf769d7),
	.w5(32'h3b0936cc),
	.w6(32'hbb2ac107),
	.w7(32'h3b8e9b63),
	.w8(32'hba9be769),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389b25d2),
	.w1(32'hbad0bf41),
	.w2(32'hbb0874ec),
	.w3(32'hbb8b84a4),
	.w4(32'hbbddee72),
	.w5(32'hbb1b955e),
	.w6(32'hbafe9786),
	.w7(32'hbc073058),
	.w8(32'hbb557126),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0124fc),
	.w1(32'h3bbacab6),
	.w2(32'h3c4b4e89),
	.w3(32'hb9c1e634),
	.w4(32'h3a8a71ea),
	.w5(32'h3c1b830a),
	.w6(32'hbc18c94d),
	.w7(32'hbb7af77f),
	.w8(32'h3c55f20b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0b753),
	.w1(32'hbc1e1191),
	.w2(32'hbbb68d17),
	.w3(32'hbb5a1417),
	.w4(32'hbc5a1f4d),
	.w5(32'hbb58d222),
	.w6(32'h3b99ab8f),
	.w7(32'hbba68f72),
	.w8(32'hbb167507),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b265934),
	.w1(32'hbbb7d63d),
	.w2(32'h3b535459),
	.w3(32'h3ae18cfd),
	.w4(32'hbb96d3d6),
	.w5(32'h3c2b48ea),
	.w6(32'hba2d9957),
	.w7(32'h3a9d5689),
	.w8(32'h3b6ab707),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07ad7a),
	.w1(32'h3bf76b0d),
	.w2(32'hbaba893d),
	.w3(32'h3c006ce6),
	.w4(32'h3bd4e433),
	.w5(32'h3c010d5c),
	.w6(32'h395d81f0),
	.w7(32'h3ad14891),
	.w8(32'h3bf489f8),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa37605),
	.w1(32'h3b0528f5),
	.w2(32'hbbdcdb2a),
	.w3(32'h3b6cc3a1),
	.w4(32'hba8e5f23),
	.w5(32'hbbaac40c),
	.w6(32'h3bfd641f),
	.w7(32'h3c019a20),
	.w8(32'hbb89cb47),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81646a),
	.w1(32'h3a2b5269),
	.w2(32'hbc020c19),
	.w3(32'hbb925c17),
	.w4(32'h39ca4381),
	.w5(32'hbc052227),
	.w6(32'hbb61d72a),
	.w7(32'h3a80b4ec),
	.w8(32'hbbf26ff8),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab39df7),
	.w1(32'h3b1a9db4),
	.w2(32'h3c178234),
	.w3(32'hbc3e006e),
	.w4(32'hbb584961),
	.w5(32'h3bf4bb87),
	.w6(32'hbc141db1),
	.w7(32'hbb9885cb),
	.w8(32'h3aa8dc89),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4583bb),
	.w1(32'hba99e26d),
	.w2(32'h3c071407),
	.w3(32'hbb2ecfdb),
	.w4(32'hb9a9fb39),
	.w5(32'h3c09dabb),
	.w6(32'hbbc2ab37),
	.w7(32'hbae28472),
	.w8(32'hba13ac77),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9b20e),
	.w1(32'h3b4436af),
	.w2(32'hba9f9613),
	.w3(32'h3c4598f5),
	.w4(32'h3c3e5e38),
	.w5(32'hbb988050),
	.w6(32'h3b8d459d),
	.w7(32'h3b9a8c55),
	.w8(32'hbb8d35af),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01f63a),
	.w1(32'h3b8ecb1a),
	.w2(32'hb94a0401),
	.w3(32'h3befde10),
	.w4(32'h3bf3bf92),
	.w5(32'h3adb74d4),
	.w6(32'hbb1dad0b),
	.w7(32'h3bb1b970),
	.w8(32'hb9de3888),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62d817),
	.w1(32'h3b3d86d3),
	.w2(32'hba5ddeff),
	.w3(32'h3b924b7c),
	.w4(32'h3b21d428),
	.w5(32'hbc053742),
	.w6(32'h3b591741),
	.w7(32'h3b06e023),
	.w8(32'h3ac02e38),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10bb66),
	.w1(32'hbc0b7f8e),
	.w2(32'hbb7831f5),
	.w3(32'h3b475b73),
	.w4(32'h389858b2),
	.w5(32'h39b7a419),
	.w6(32'hba03638f),
	.w7(32'h3ba8ddd6),
	.w8(32'h3b8f522c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbed427),
	.w1(32'h3b74687d),
	.w2(32'h3c6bf1e1),
	.w3(32'h3b148a41),
	.w4(32'h3b87f96b),
	.w5(32'h3c8b80e0),
	.w6(32'hbb8abe86),
	.w7(32'h39e66fc9),
	.w8(32'h3b91c99c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98639d),
	.w1(32'hb9eaa472),
	.w2(32'hbc028083),
	.w3(32'h3c986a90),
	.w4(32'hbba4d993),
	.w5(32'hbbe98a25),
	.w6(32'h3b955ea6),
	.w7(32'hbc3a6529),
	.w8(32'hbb7fa47b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab16361),
	.w1(32'hbbbf1c69),
	.w2(32'h3b89ebaa),
	.w3(32'h39bbf217),
	.w4(32'h3ab1e514),
	.w5(32'hba6927a4),
	.w6(32'hbbf592c4),
	.w7(32'hbc142f01),
	.w8(32'hbbdb85fa),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc161c6),
	.w1(32'h3b31f8c6),
	.w2(32'h3bc2252f),
	.w3(32'h3b96f873),
	.w4(32'hbbd4af02),
	.w5(32'hbba1bff2),
	.w6(32'hbc0ace04),
	.w7(32'hbc3aa1c8),
	.w8(32'hbc26db28),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3707bb),
	.w1(32'h3c477a36),
	.w2(32'hbb60332d),
	.w3(32'hbc23a5fa),
	.w4(32'hb89ec78d),
	.w5(32'hbc1271c7),
	.w6(32'hbbbe3ea1),
	.w7(32'hbb96254c),
	.w8(32'hbb53b760),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d5b7a),
	.w1(32'hbb225676),
	.w2(32'hbb3483a1),
	.w3(32'hbb8c35ef),
	.w4(32'hbb9418e5),
	.w5(32'h3c18ea69),
	.w6(32'h3b29da9f),
	.w7(32'h3bb98097),
	.w8(32'h3b9883bd),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb4d24),
	.w1(32'hbc2ebf82),
	.w2(32'h3b17b259),
	.w3(32'h3b7df186),
	.w4(32'hbbdae085),
	.w5(32'h3bbed00b),
	.w6(32'h3bfe35fa),
	.w7(32'hbb64d591),
	.w8(32'h3a6b7173),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f4f7b),
	.w1(32'hbb3b5970),
	.w2(32'h3a588338),
	.w3(32'hb944ecc7),
	.w4(32'hbbd290f6),
	.w5(32'h3b1880ca),
	.w6(32'hbbeb2a7e),
	.w7(32'hbc18e5b9),
	.w8(32'hbba118a2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e1b3f7),
	.w1(32'hbc0df33f),
	.w2(32'h3b21d19a),
	.w3(32'hb89a87a7),
	.w4(32'hbc1ee75c),
	.w5(32'hbad167b0),
	.w6(32'hbba441d7),
	.w7(32'hbc7c602f),
	.w8(32'hbb4a6de3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a13b7),
	.w1(32'h3b8c82b4),
	.w2(32'hbb520cdc),
	.w3(32'hb995681e),
	.w4(32'hbbcb850d),
	.w5(32'hbbb6b7be),
	.w6(32'hbc741e1e),
	.w7(32'hbc5df13f),
	.w8(32'hb89155e5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77b551),
	.w1(32'h3889fac7),
	.w2(32'h3ba75905),
	.w3(32'h3ac774db),
	.w4(32'h3bc957c5),
	.w5(32'h3c381e7c),
	.w6(32'h3a18e52f),
	.w7(32'h3bed4246),
	.w8(32'h3bfd785e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcc16e),
	.w1(32'h3bb57424),
	.w2(32'h3bd5cd56),
	.w3(32'h3b99ad77),
	.w4(32'h3c223cda),
	.w5(32'h3ab0cb20),
	.w6(32'h3b966f29),
	.w7(32'h3b0f6ce5),
	.w8(32'hbbcbc2ff),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed50c4),
	.w1(32'hbae828f0),
	.w2(32'hb9423a56),
	.w3(32'hbb12f655),
	.w4(32'h38bdb657),
	.w5(32'h3b9d58d2),
	.w6(32'h3b5e03c3),
	.w7(32'hb87fd90c),
	.w8(32'hb9957e42),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac8102),
	.w1(32'h3b15e9a1),
	.w2(32'hbb0aef8d),
	.w3(32'h3b604748),
	.w4(32'hb8a75a35),
	.w5(32'hbbcee98d),
	.w6(32'hba81869d),
	.w7(32'hbb0670e4),
	.w8(32'hba5dadc9),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44fb4a),
	.w1(32'hbb503a90),
	.w2(32'h3a48a2b8),
	.w3(32'hbc38949f),
	.w4(32'hbb94f181),
	.w5(32'hbb0f1d1b),
	.w6(32'hba9450c9),
	.w7(32'h3b11f8b6),
	.w8(32'hbb436cb5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca90a7),
	.w1(32'hba80854f),
	.w2(32'hbb19ba05),
	.w3(32'hbae9de06),
	.w4(32'hba8a2c20),
	.w5(32'hbb1d80f3),
	.w6(32'hbb838c3a),
	.w7(32'hbb19fa2a),
	.w8(32'h399671bd),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d6f6f),
	.w1(32'h3af56cee),
	.w2(32'h3b69db3d),
	.w3(32'hbba911f5),
	.w4(32'h3b400f97),
	.w5(32'h3b5f8a80),
	.w6(32'h3a05a3c9),
	.w7(32'h3bb5e1e4),
	.w8(32'h3ba41855),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b367978),
	.w1(32'h3ae08d05),
	.w2(32'hba55a191),
	.w3(32'h3bdc59bd),
	.w4(32'h3bb76dac),
	.w5(32'hbb0518bb),
	.w6(32'h3a396ed5),
	.w7(32'hbb997204),
	.w8(32'h3b199473),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dd865),
	.w1(32'h39b26e58),
	.w2(32'hbb264dbd),
	.w3(32'hbbc6c375),
	.w4(32'h38ec2077),
	.w5(32'hba85407d),
	.w6(32'h3b0b8fbe),
	.w7(32'h39be92f3),
	.w8(32'hb8cc1367),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12c97b),
	.w1(32'hb9888031),
	.w2(32'hbc1a859e),
	.w3(32'h3a9956ff),
	.w4(32'h3b1662e8),
	.w5(32'hbc97903d),
	.w6(32'h3aeb1451),
	.w7(32'h3b88a637),
	.w8(32'hbc8c53ed),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd36f1c),
	.w1(32'hbb9bf745),
	.w2(32'h3bb76ead),
	.w3(32'hbc233055),
	.w4(32'hbbc7d1cc),
	.w5(32'h3b9dc493),
	.w6(32'hbc75346a),
	.w7(32'hbbacadfb),
	.w8(32'h38db7fb2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e67d6b),
	.w1(32'hbb0967e2),
	.w2(32'h3bb370ce),
	.w3(32'h3b803a74),
	.w4(32'hbb3981a3),
	.w5(32'h3b140cb1),
	.w6(32'hb7723975),
	.w7(32'hbb193cf5),
	.w8(32'hba28376d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfee1f),
	.w1(32'h3b937f5c),
	.w2(32'hbb844a2f),
	.w3(32'h3c1c67e2),
	.w4(32'h3bf5c9b9),
	.w5(32'h39784847),
	.w6(32'h3bb43f62),
	.w7(32'h3b867006),
	.w8(32'h3ad76139),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfca696),
	.w1(32'hbb28fb35),
	.w2(32'hba8440e7),
	.w3(32'hbb7f4c15),
	.w4(32'hbb8f93ed),
	.w5(32'hba53041d),
	.w6(32'hbb9d6159),
	.w7(32'hbb26ebf2),
	.w8(32'hbaa93a09),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2111e),
	.w1(32'hba8d7b6c),
	.w2(32'hbc27ffea),
	.w3(32'h3a682187),
	.w4(32'hbb00261b),
	.w5(32'hbb9700f2),
	.w6(32'hb9a111e8),
	.w7(32'hbb6f87de),
	.w8(32'hbba16b11),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc095ffe),
	.w1(32'hbc57db50),
	.w2(32'hbbd7b6b6),
	.w3(32'hbbcf16d1),
	.w4(32'hbc2dd7af),
	.w5(32'hbc165657),
	.w6(32'hbc0a3e9f),
	.w7(32'hbc29f7a1),
	.w8(32'hbad8c9ec),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ce2f1),
	.w1(32'hbb8bbee2),
	.w2(32'hbab64b1c),
	.w3(32'hbb7d7cb7),
	.w4(32'h3b78b646),
	.w5(32'h3ba00078),
	.w6(32'h3aab8ac3),
	.w7(32'h3be53ebb),
	.w8(32'h3b9358e4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5eccde),
	.w1(32'hbb08ec1e),
	.w2(32'h3a640634),
	.w3(32'h3c34adc3),
	.w4(32'h3c15cae6),
	.w5(32'h3b9a58b8),
	.w6(32'h3b515ca4),
	.w7(32'h3c35a739),
	.w8(32'hbb975c7e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfeef38),
	.w1(32'h3ab2ecd9),
	.w2(32'h3b02328a),
	.w3(32'h3c4a563b),
	.w4(32'h3bd4ca7f),
	.w5(32'h3b92aed5),
	.w6(32'h39bbb339),
	.w7(32'h3aa7867b),
	.w8(32'h3af63e9f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5961a1),
	.w1(32'h3af25693),
	.w2(32'hbb557704),
	.w3(32'h3be810d4),
	.w4(32'h3bb6d35d),
	.w5(32'hbbc54aed),
	.w6(32'h3b56c7dc),
	.w7(32'h3b3fa077),
	.w8(32'hb60fbaa8),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b700f9a),
	.w1(32'h3b10f231),
	.w2(32'h3ac90500),
	.w3(32'h3b9b941b),
	.w4(32'h3aa12523),
	.w5(32'h3a08a13d),
	.w6(32'h3a699341),
	.w7(32'hbb0362cb),
	.w8(32'h3b63e004),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7ee08),
	.w1(32'h3a0ca918),
	.w2(32'hbb39b5f5),
	.w3(32'hbaefdeea),
	.w4(32'h39f45f18),
	.w5(32'hbbf25051),
	.w6(32'h3ac0eee3),
	.w7(32'h3b35e9f8),
	.w8(32'hbb34ebb3),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb944649),
	.w1(32'hbc29755a),
	.w2(32'h3ba350b7),
	.w3(32'hbc13cf7a),
	.w4(32'hbc1e5d44),
	.w5(32'h3c0a0c92),
	.w6(32'hbbae069d),
	.w7(32'hbab6255e),
	.w8(32'hba9b37d8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c171af5),
	.w1(32'h3c207171),
	.w2(32'h3ba2099b),
	.w3(32'h3ab78b2e),
	.w4(32'h3b2de04b),
	.w5(32'h3bacd409),
	.w6(32'h3af1c468),
	.w7(32'h3b2ec48a),
	.w8(32'hbb8e453a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f6114),
	.w1(32'h3a482067),
	.w2(32'h3aa60318),
	.w3(32'h3c59089c),
	.w4(32'h3b551147),
	.w5(32'h3b8e2eab),
	.w6(32'hba433e7a),
	.w7(32'hba0b6db5),
	.w8(32'hbafdea60),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bdcf8),
	.w1(32'h3ab8e92d),
	.w2(32'hbbaa2d5f),
	.w3(32'h3bb296c3),
	.w4(32'h3ad1ce89),
	.w5(32'hbc29c451),
	.w6(32'hb900a484),
	.w7(32'hbb8e201e),
	.w8(32'hbbfae19e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86a87e),
	.w1(32'hbb7ff3bd),
	.w2(32'hbbb7b5c4),
	.w3(32'hbbc679c3),
	.w4(32'hbb89dbfc),
	.w5(32'hbb793da6),
	.w6(32'hbbe97bcf),
	.w7(32'hbb902e4b),
	.w8(32'hbb6a9ddb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc628e),
	.w1(32'hbb888bb8),
	.w2(32'hbb1dabb8),
	.w3(32'hbbd90054),
	.w4(32'hbb8a67d3),
	.w5(32'h3ac629b2),
	.w6(32'hbbc0c1ce),
	.w7(32'hbb5663ac),
	.w8(32'h3c027e37),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21ab7f),
	.w1(32'h3b850b0d),
	.w2(32'h3c09963b),
	.w3(32'h3c2133b7),
	.w4(32'h3b9e7704),
	.w5(32'h3ba1831e),
	.w6(32'h3ba51708),
	.w7(32'hb9390e12),
	.w8(32'h3b6c9a1a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc7dd4),
	.w1(32'h3ba3a7e5),
	.w2(32'h3bf72a06),
	.w3(32'h3c8fb0a4),
	.w4(32'h3b94b0e1),
	.w5(32'h383f5648),
	.w6(32'h3c346015),
	.w7(32'h3ba3e017),
	.w8(32'hbb8b7445),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf2e2a),
	.w1(32'h3b06a18d),
	.w2(32'h3b899c6b),
	.w3(32'hbb8e4fe7),
	.w4(32'hbc032d20),
	.w5(32'hbbd0e635),
	.w6(32'hbc2f3c16),
	.w7(32'hbbe6dd42),
	.w8(32'hbb1c7af5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe649d7),
	.w1(32'hbade395b),
	.w2(32'hbbce0cd7),
	.w3(32'hbc5bb79f),
	.w4(32'hbbf6dd57),
	.w5(32'hbb6ca3a1),
	.w6(32'hbb9e4d44),
	.w7(32'h3b82026e),
	.w8(32'hbbd3214b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3574aa),
	.w1(32'hbb9d6b61),
	.w2(32'hbb90c393),
	.w3(32'h3aa3a753),
	.w4(32'hba98550a),
	.w5(32'hbbda986a),
	.w6(32'hbb131e07),
	.w7(32'hbb4cd702),
	.w8(32'hbb397755),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaee009),
	.w1(32'hbabc18ef),
	.w2(32'h386f9601),
	.w3(32'hbbdca95e),
	.w4(32'hb9e9af73),
	.w5(32'hbb497c8a),
	.w6(32'hbb93176d),
	.w7(32'h3b16934a),
	.w8(32'hbaf12294),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17131a),
	.w1(32'hb9145b83),
	.w2(32'h394a2a09),
	.w3(32'hbb521730),
	.w4(32'h3aee62f4),
	.w5(32'h39b1e407),
	.w6(32'hbb8baf4e),
	.w7(32'hbb3ddee2),
	.w8(32'h3b1a426e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe6384),
	.w1(32'hba1a3a81),
	.w2(32'hbbd3c02e),
	.w3(32'hbb6e9d7a),
	.w4(32'hbbece6d6),
	.w5(32'hba1daff4),
	.w6(32'hbb78eec6),
	.w7(32'h3b711a14),
	.w8(32'hbae8d1af),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8234ec),
	.w1(32'hbc4b5542),
	.w2(32'h3b419f79),
	.w3(32'h3adf2e71),
	.w4(32'hbc221fd6),
	.w5(32'h3c1531b8),
	.w6(32'hbb901357),
	.w7(32'hbbd476a1),
	.w8(32'h3b7ac11a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef862d),
	.w1(32'h3b695472),
	.w2(32'hbae26432),
	.w3(32'h3bc10bc7),
	.w4(32'h3b0a7fe2),
	.w5(32'h3c2156e9),
	.w6(32'h3bf57e6c),
	.w7(32'h3b9c8562),
	.w8(32'h3be9fa79),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fdd51),
	.w1(32'h3acc9823),
	.w2(32'hbbb1924b),
	.w3(32'h3cbc56b0),
	.w4(32'h3c38257f),
	.w5(32'hbb92b056),
	.w6(32'h3ba98d3e),
	.w7(32'h3c13052c),
	.w8(32'hb93df8e2),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16f7c9),
	.w1(32'hbb3ae57d),
	.w2(32'h3767d5d1),
	.w3(32'hbca05cf2),
	.w4(32'hbc72d90b),
	.w5(32'h3bc97549),
	.w6(32'hbc4a826f),
	.w7(32'hbc1df89f),
	.w8(32'hba1d1319),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7875601),
	.w1(32'h3a94ecef),
	.w2(32'hbab5d112),
	.w3(32'h3b960503),
	.w4(32'h3b38ae43),
	.w5(32'h3b7795ce),
	.w6(32'h3b19fbf0),
	.w7(32'h3bac4856),
	.w8(32'h3bc144be),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e917d),
	.w1(32'hbb43b5f6),
	.w2(32'hbb10d861),
	.w3(32'h3c00c609),
	.w4(32'h3c28b712),
	.w5(32'hbb63ad28),
	.w6(32'h3b981e8a),
	.w7(32'h3bf6f47c),
	.w8(32'hbb4e94ab),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8846903),
	.w1(32'hbadf96aa),
	.w2(32'hbaa5a14e),
	.w3(32'h3b09e0ab),
	.w4(32'hbb1d773d),
	.w5(32'h39d1dec0),
	.w6(32'hbabb37e4),
	.w7(32'hbba571f3),
	.w8(32'hbc0ba6a2),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b000b68),
	.w1(32'h3aeb3f23),
	.w2(32'h3b0db71e),
	.w3(32'h39b3092f),
	.w4(32'hbbc6b100),
	.w5(32'h3c385119),
	.w6(32'hbc2a988a),
	.w7(32'hbc38b597),
	.w8(32'h3b2baa4e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf02a0f),
	.w1(32'h3b225932),
	.w2(32'h3af8dd6c),
	.w3(32'h3c662897),
	.w4(32'h3be21dfd),
	.w5(32'h3ba7996c),
	.w6(32'h3c2fc798),
	.w7(32'h3b770f7e),
	.w8(32'h3b575e82),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5685c3),
	.w1(32'hba5108d3),
	.w2(32'h3b7e85df),
	.w3(32'h3c191c83),
	.w4(32'hb7de7dfb),
	.w5(32'h3a39daff),
	.w6(32'h3b34b3da),
	.w7(32'hbb241a9e),
	.w8(32'hbaa507f3),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac080e),
	.w1(32'hbb91f0f5),
	.w2(32'h3ab19746),
	.w3(32'h3ba3ebaa),
	.w4(32'hbb6f7919),
	.w5(32'hbbbefa62),
	.w6(32'hb9b78c37),
	.w7(32'hbbb85f43),
	.w8(32'hbb3a17f1),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fcd02),
	.w1(32'hb938d720),
	.w2(32'h3c0eac3f),
	.w3(32'hbbda90d4),
	.w4(32'hbc07f507),
	.w5(32'h3beaa638),
	.w6(32'hbc290346),
	.w7(32'hbc2686ef),
	.w8(32'h3aed7d47),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc40943),
	.w1(32'hbb36ea7a),
	.w2(32'hbb1aebdb),
	.w3(32'h3b90e392),
	.w4(32'h3aa7d82f),
	.w5(32'h3b3975bd),
	.w6(32'h3afe9715),
	.w7(32'h3b24cb9f),
	.w8(32'h3b92d9ed),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34fea0),
	.w1(32'h3acc9bb4),
	.w2(32'h3b260e7e),
	.w3(32'h3be0c3e5),
	.w4(32'h3b897bd4),
	.w5(32'h3c243d49),
	.w6(32'h3c0142cc),
	.w7(32'h3c649925),
	.w8(32'h3bc1b335),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca2b83),
	.w1(32'hbb80b1a6),
	.w2(32'h39b2c9b0),
	.w3(32'h3b5daa2e),
	.w4(32'h3bd6c8a9),
	.w5(32'h3bb72df9),
	.w6(32'h3bd44682),
	.w7(32'h39b29410),
	.w8(32'h3be7f13d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d1f5f),
	.w1(32'hbbfac85b),
	.w2(32'h3a11383c),
	.w3(32'h3c552bfc),
	.w4(32'h3b7389c0),
	.w5(32'hbb284089),
	.w6(32'h3c01fb17),
	.w7(32'hbb875191),
	.w8(32'h3bed7184),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d9004),
	.w1(32'hba974534),
	.w2(32'h39f74b5b),
	.w3(32'h3c31a7f2),
	.w4(32'h3bb219a8),
	.w5(32'h3c1fdcb7),
	.w6(32'h3b50d366),
	.w7(32'h3b710df2),
	.w8(32'h3c1f620c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1881c1),
	.w1(32'hbb69ac2b),
	.w2(32'hb9a6f88c),
	.w3(32'h3c1e3f54),
	.w4(32'h3c0f8f65),
	.w5(32'hbb46a7b5),
	.w6(32'h3b40ec41),
	.w7(32'h3b5708b9),
	.w8(32'h3b8eca73),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb514dc4),
	.w1(32'h3a70b58a),
	.w2(32'hbb770fff),
	.w3(32'hbb5291d4),
	.w4(32'h3ba27bc9),
	.w5(32'hbbc9667e),
	.w6(32'h3bf88874),
	.w7(32'h3bf87266),
	.w8(32'hbbd6c473),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba56796),
	.w1(32'hbb4129ce),
	.w2(32'h3ae30341),
	.w3(32'hbbe27c86),
	.w4(32'hbbaeac3b),
	.w5(32'hbbe77b73),
	.w6(32'hbc1c2588),
	.w7(32'hbc1cb094),
	.w8(32'hbb65f311),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf5811),
	.w1(32'hbbec374a),
	.w2(32'hbab99f9a),
	.w3(32'hbbede9fb),
	.w4(32'hbc1c1497),
	.w5(32'h3a108c28),
	.w6(32'hbba0feb9),
	.w7(32'hbad8bef8),
	.w8(32'hbbd383bf),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89083b),
	.w1(32'h3b07404e),
	.w2(32'h3bbeee9d),
	.w3(32'h3a77e5b6),
	.w4(32'hb96ea60e),
	.w5(32'h3bf0005e),
	.w6(32'hbbdeeab6),
	.w7(32'hbbb08be8),
	.w8(32'h3c1c661a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d1627),
	.w1(32'h3b3cfff1),
	.w2(32'hbb03a1a8),
	.w3(32'h3c8bbc54),
	.w4(32'h3c8e5dd9),
	.w5(32'h3aabd786),
	.w6(32'h3c413c79),
	.w7(32'h3be93ebe),
	.w8(32'h3a6950f2),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafde49c),
	.w1(32'hb7c21ec9),
	.w2(32'h3a695261),
	.w3(32'hbb052948),
	.w4(32'h3ac3c230),
	.w5(32'hba139e36),
	.w6(32'hbb582b58),
	.w7(32'hba217140),
	.w8(32'hbb02d0ff),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb248625),
	.w1(32'hb99948c3),
	.w2(32'h3a9c2be9),
	.w3(32'hbaaaf83e),
	.w4(32'hbbce68df),
	.w5(32'h39cf3057),
	.w6(32'hbadbfbc0),
	.w7(32'hbaa3bb3f),
	.w8(32'hb97b8908),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1eccc0),
	.w1(32'hbb1ee692),
	.w2(32'h3b0c00fb),
	.w3(32'hbb3bfb1c),
	.w4(32'hbb9a0ca5),
	.w5(32'h3a85ea72),
	.w6(32'hbb21d9e1),
	.w7(32'hbbd8f7cc),
	.w8(32'h3a47eb3e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae50de5),
	.w1(32'hb830d03b),
	.w2(32'hb9d25ff7),
	.w3(32'h3ad7c83e),
	.w4(32'hb95665c0),
	.w5(32'h3b2e9750),
	.w6(32'hbafd108f),
	.w7(32'hbaf7cc62),
	.w8(32'h3b5f0f1e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c426c18),
	.w1(32'h3b824498),
	.w2(32'hba017d13),
	.w3(32'h3cb2ec6f),
	.w4(32'h3c160564),
	.w5(32'hbaedeb5b),
	.w6(32'h3c32a219),
	.w7(32'hbb267e90),
	.w8(32'hbb2693bc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f3a45),
	.w1(32'hbba18f8c),
	.w2(32'h3b0b457d),
	.w3(32'hbb99efea),
	.w4(32'hbb4e5ad9),
	.w5(32'h3c2c7e11),
	.w6(32'hbba0773b),
	.w7(32'hb8ded1d6),
	.w8(32'h3bcfc777),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66204d),
	.w1(32'h3bec7208),
	.w2(32'h3b872d53),
	.w3(32'h3cb629b1),
	.w4(32'h3c639708),
	.w5(32'h3bf6e67b),
	.w6(32'h3bb393ee),
	.w7(32'h3b8f9bbe),
	.w8(32'h3b5ee4b1),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b851321),
	.w1(32'h3c509a11),
	.w2(32'h390dd7b2),
	.w3(32'h3c93fccf),
	.w4(32'h3c613e2e),
	.w5(32'h3b787aac),
	.w6(32'h3bc3fb12),
	.w7(32'h3bd336a2),
	.w8(32'h3bbac63e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93c2ab),
	.w1(32'h3a266136),
	.w2(32'h3c1a0ba6),
	.w3(32'h3baa25c4),
	.w4(32'hbb3ce74d),
	.w5(32'h3c28fcf4),
	.w6(32'hba98e8bf),
	.w7(32'hbb967c88),
	.w8(32'h3b59ddbd),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule