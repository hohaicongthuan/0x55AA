module layer_10_featuremap_133(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba191d38),
	.w1(32'h3ad1582c),
	.w2(32'hba9ebf8c),
	.w3(32'hb993d1fb),
	.w4(32'h3922fe1f),
	.w5(32'h38da2744),
	.w6(32'h3a240658),
	.w7(32'hba42c9b1),
	.w8(32'hba622dcb),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fdfc1),
	.w1(32'hba480543),
	.w2(32'hba952b77),
	.w3(32'hba858faa),
	.w4(32'h3b03066d),
	.w5(32'h3a9976b2),
	.w6(32'hba4955d3),
	.w7(32'h39a056d2),
	.w8(32'hba56e694),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35f05f),
	.w1(32'hb9eb1427),
	.w2(32'hb91b2a1f),
	.w3(32'h3a3114f1),
	.w4(32'h3973a3c9),
	.w5(32'h39dfc1dc),
	.w6(32'hba0097b4),
	.w7(32'hba0d2243),
	.w8(32'h391ea83d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4e5c2),
	.w1(32'hb85db8c6),
	.w2(32'hba8dcebe),
	.w3(32'h3819062c),
	.w4(32'h39d980a2),
	.w5(32'hb9e7c280),
	.w6(32'h3a83db55),
	.w7(32'h3a09f0ed),
	.w8(32'hb9582b42),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fffd4),
	.w1(32'h39cf416e),
	.w2(32'hbad8a8d9),
	.w3(32'h3965585d),
	.w4(32'h39d37a14),
	.w5(32'hba062694),
	.w6(32'h3a4c687e),
	.w7(32'hb76305e3),
	.w8(32'h39228167),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38378d71),
	.w1(32'h3a3f1ea4),
	.w2(32'h3a1c6cdc),
	.w3(32'h39cfd9be),
	.w4(32'h3a9b01fa),
	.w5(32'h39d5ac06),
	.w6(32'h3a1d8e36),
	.w7(32'h39db8a7a),
	.w8(32'h3a380221),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2334e9),
	.w1(32'hbab03a6b),
	.w2(32'hbb5a9655),
	.w3(32'h3b2bbc45),
	.w4(32'hbab8c3a9),
	.w5(32'hbb50a3bc),
	.w6(32'hbadd2029),
	.w7(32'h39d71c38),
	.w8(32'hbb2fb600),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e921e),
	.w1(32'hbc1d0b0c),
	.w2(32'hbbaa185d),
	.w3(32'hbb8dc4b5),
	.w4(32'hbc003335),
	.w5(32'hbc018050),
	.w6(32'hbbc1f264),
	.w7(32'hbb420ba8),
	.w8(32'hba1debb6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389d7bf5),
	.w1(32'h394b6e65),
	.w2(32'hb9aae28a),
	.w3(32'hba107fb5),
	.w4(32'h378ef685),
	.w5(32'hb9541a5b),
	.w6(32'h39abeaba),
	.w7(32'h38a10e7d),
	.w8(32'hb94e1f8d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b400d42),
	.w1(32'h3b957cf0),
	.w2(32'hba279584),
	.w3(32'h3b5d7bf2),
	.w4(32'h3b63d3a5),
	.w5(32'h3a73bbe4),
	.w6(32'hbb59dbdd),
	.w7(32'hbb757b40),
	.w8(32'hbbfcf00b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae04777),
	.w1(32'hba84f894),
	.w2(32'hba704a73),
	.w3(32'h3aaa0401),
	.w4(32'h3a2758d1),
	.w5(32'h39f110be),
	.w6(32'hb9215549),
	.w7(32'h3a04e833),
	.w8(32'h3a6cfb70),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac49c3b),
	.w1(32'h3b331552),
	.w2(32'hbb1d9d9c),
	.w3(32'h3b235143),
	.w4(32'hb8f6396a),
	.w5(32'hbb82da38),
	.w6(32'hbb1a1e74),
	.w7(32'h3ae1b120),
	.w8(32'hbb7c8f8e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2eb91),
	.w1(32'h3b2b08e8),
	.w2(32'hbb2fce8c),
	.w3(32'h3bb01851),
	.w4(32'h3b03779f),
	.w5(32'hbb194c93),
	.w6(32'hbb879dda),
	.w7(32'hbbd32520),
	.w8(32'hbc210e4a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4257a),
	.w1(32'hbb9a948e),
	.w2(32'hbbd51e0d),
	.w3(32'h39def7b8),
	.w4(32'hbaafd07c),
	.w5(32'hbb8dcf98),
	.w6(32'hba0a295a),
	.w7(32'hbb0aa01a),
	.w8(32'hbb0c2e7c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dedcd),
	.w1(32'hbb184142),
	.w2(32'hbb86dd1a),
	.w3(32'hbac4dad5),
	.w4(32'h3b05d8c8),
	.w5(32'hb9732dc8),
	.w6(32'hbb03ec54),
	.w7(32'hba26c27a),
	.w8(32'hbb1799bb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbda2bf),
	.w1(32'hbb6b9f20),
	.w2(32'hbbbb8813),
	.w3(32'h39ec8a8c),
	.w4(32'h3aa0593d),
	.w5(32'hba2fbb33),
	.w6(32'hbb20fe18),
	.w7(32'hbb718f1a),
	.w8(32'hbbf2beea),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e702e),
	.w1(32'hba0be5e8),
	.w2(32'hba9edd78),
	.w3(32'hb8ce14da),
	.w4(32'hb9e4c8be),
	.w5(32'hba6ded10),
	.w6(32'h3a1c6b2c),
	.w7(32'hba8aae06),
	.w8(32'hba6ebfeb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab89f28),
	.w1(32'h3b75570a),
	.w2(32'hbad139af),
	.w3(32'hbb1c94fa),
	.w4(32'hbacb72c5),
	.w5(32'hbb5953ed),
	.w6(32'hbbbed57b),
	.w7(32'hbaa862e2),
	.w8(32'hbbea4342),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6faf72),
	.w1(32'h3b2ed603),
	.w2(32'h3a25826c),
	.w3(32'h3b0c2bf3),
	.w4(32'h3a06dfc9),
	.w5(32'hba3e8aa6),
	.w6(32'hbb4cd122),
	.w7(32'hbb357d7f),
	.w8(32'hbba77ea1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f1902),
	.w1(32'hb998c3fd),
	.w2(32'hb925d599),
	.w3(32'h3817e2d2),
	.w4(32'hb842fc75),
	.w5(32'hb94c31fd),
	.w6(32'h38d652e1),
	.w7(32'hb8fa4c4e),
	.w8(32'hb9cbd056),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba181506),
	.w1(32'hba2ba8d0),
	.w2(32'hbb08c086),
	.w3(32'hba26c1f2),
	.w4(32'h398135bf),
	.w5(32'hbaa3cec1),
	.w6(32'h3869b736),
	.w7(32'hba81c471),
	.w8(32'hb9ba52f4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78fd7c6),
	.w1(32'h3ac302a8),
	.w2(32'h3aca064a),
	.w3(32'h39d65c4a),
	.w4(32'h3b52e425),
	.w5(32'h3ae75a69),
	.w6(32'h39a951a8),
	.w7(32'h3a5680bb),
	.w8(32'hba50e0f3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7dbd7),
	.w1(32'h3ad8c72d),
	.w2(32'hbb8db2ac),
	.w3(32'h3b2348b4),
	.w4(32'h3bbc21c8),
	.w5(32'hba0c0259),
	.w6(32'hbc6c0a40),
	.w7(32'hbc0372ca),
	.w8(32'hbc7ff165),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaeed3b),
	.w1(32'h3af23815),
	.w2(32'hbb4b2094),
	.w3(32'h38e12e81),
	.w4(32'h3acaf6ba),
	.w5(32'hbb19b534),
	.w6(32'hbbdbe0af),
	.w7(32'hbbe37aa7),
	.w8(32'hbc17dbe3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e75a9),
	.w1(32'h3b60230d),
	.w2(32'hba727284),
	.w3(32'hbae3d136),
	.w4(32'h3b39d763),
	.w5(32'h3b0543ce),
	.w6(32'hbb59374e),
	.w7(32'hbbc00630),
	.w8(32'hbc154050),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c0115),
	.w1(32'hba1052e4),
	.w2(32'h39d5eb1a),
	.w3(32'h37a02441),
	.w4(32'hb9f36001),
	.w5(32'hba3664f1),
	.w6(32'h39c7643f),
	.w7(32'hba30411c),
	.w8(32'hba47e5cc),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a295447),
	.w1(32'hba843d34),
	.w2(32'hba6812af),
	.w3(32'hba50dc56),
	.w4(32'hba26f0f7),
	.w5(32'hba5083b3),
	.w6(32'hb9b9cf74),
	.w7(32'hba2efead),
	.w8(32'hba2d2aa9),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e2cac),
	.w1(32'h3a55ff7c),
	.w2(32'h3a3bd476),
	.w3(32'h3c57fa9a),
	.w4(32'hbb9980bc),
	.w5(32'hbb3553f1),
	.w6(32'h3c9f1d4a),
	.w7(32'hbb7233b4),
	.w8(32'hbb4285c8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8055dbd),
	.w1(32'h3a5e1720),
	.w2(32'hbac84742),
	.w3(32'hba0e60f6),
	.w4(32'h3ac6d66b),
	.w5(32'hba3d4f33),
	.w6(32'hb855056a),
	.w7(32'h39d33e81),
	.w8(32'h38f779e5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c581400),
	.w1(32'h3ae88a2d),
	.w2(32'hba577ccb),
	.w3(32'h3c05b96a),
	.w4(32'hba2d4b5b),
	.w5(32'hbb275f48),
	.w6(32'h3c378e1b),
	.w7(32'hbaf00d86),
	.w8(32'hbb9d1ec6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91bc6ae),
	.w1(32'hb9b0152c),
	.w2(32'hba8d0eb1),
	.w3(32'hb96d7f82),
	.w4(32'h379f682c),
	.w5(32'hba39c444),
	.w6(32'h36daaa9e),
	.w7(32'hba0768ff),
	.w8(32'hb9d4de83),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba853c38),
	.w1(32'hba559b54),
	.w2(32'hbaa3289c),
	.w3(32'hba15f228),
	.w4(32'hba113415),
	.w5(32'hbaa20fc4),
	.w6(32'hba1dab5a),
	.w7(32'hba56f67b),
	.w8(32'hb9fc6664),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b4297),
	.w1(32'h3b1042e5),
	.w2(32'h3a7ce8d2),
	.w3(32'h38ccbbd3),
	.w4(32'h3aa6efba),
	.w5(32'h3a5c6b8a),
	.w6(32'hbae7138e),
	.w7(32'hba836225),
	.w8(32'hbb9e8cfb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba524ee2),
	.w1(32'hbb2914db),
	.w2(32'hbb485168),
	.w3(32'hba91ec36),
	.w4(32'hbb0a8884),
	.w5(32'hbb3e2393),
	.w6(32'hbad85e53),
	.w7(32'hbb3edb58),
	.w8(32'hbb45ec4d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba984ab6),
	.w1(32'h3a4a4ac1),
	.w2(32'h3aa05ab2),
	.w3(32'hb99c6795),
	.w4(32'h3a575bc8),
	.w5(32'h39f804dd),
	.w6(32'h3af6cb33),
	.w7(32'h3ac70e84),
	.w8(32'h3a3c4053),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e4352),
	.w1(32'h3aaac3bd),
	.w2(32'hbaf3a849),
	.w3(32'h3b07ed0e),
	.w4(32'h39dcd4ba),
	.w5(32'hbaf2c5c2),
	.w6(32'hbb355cd7),
	.w7(32'hba33a1aa),
	.w8(32'hb964755c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20a147),
	.w1(32'hbb9b54fa),
	.w2(32'hbc742a19),
	.w3(32'h3b11b2d3),
	.w4(32'h3b6ad095),
	.w5(32'hb94dd4ec),
	.w6(32'hbc183bfb),
	.w7(32'h3b85242e),
	.w8(32'hbb85c198),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1dfcf),
	.w1(32'h3be0531b),
	.w2(32'hba5892c4),
	.w3(32'h3b606a59),
	.w4(32'h3bdc07b0),
	.w5(32'h3a9cb951),
	.w6(32'hbaa446dd),
	.w7(32'hbba7e3a5),
	.w8(32'hbc269bdd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f9b0b),
	.w1(32'h3b242d57),
	.w2(32'hbbf7f1c8),
	.w3(32'h3c21a516),
	.w4(32'h3a8fd311),
	.w5(32'hbc05ea0d),
	.w6(32'h3c1c688c),
	.w7(32'hbb375b11),
	.w8(32'hbc2eb2e2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe7bad),
	.w1(32'h3a1b7dd2),
	.w2(32'h39b203c3),
	.w3(32'hba5544e8),
	.w4(32'h3a886081),
	.w5(32'h3a6195aa),
	.w6(32'hbad27939),
	.w7(32'hba5fd980),
	.w8(32'hb9b02bb9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e7b218),
	.w1(32'hb98c5745),
	.w2(32'hba90b1a5),
	.w3(32'h38e1605f),
	.w4(32'hb9496a3b),
	.w5(32'hba669a82),
	.w6(32'hb9d62c9c),
	.w7(32'hba4c9cf9),
	.w8(32'hb88ed09a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a0f4e),
	.w1(32'hbaa10cf1),
	.w2(32'hba8a4413),
	.w3(32'hb9d81ef3),
	.w4(32'hba48be75),
	.w5(32'h38b1ff56),
	.w6(32'hba685ff0),
	.w7(32'hba40888a),
	.w8(32'hb9c2b94b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba927482),
	.w1(32'h3951773c),
	.w2(32'hba95b9a0),
	.w3(32'h399407f0),
	.w4(32'h38b60802),
	.w5(32'hba943f5b),
	.w6(32'h380f57ea),
	.w7(32'h3a5c20f7),
	.w8(32'hb9ba25cd),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a82d6),
	.w1(32'h3b9715dc),
	.w2(32'h3a9d988a),
	.w3(32'h3afdb063),
	.w4(32'h3b51a9f1),
	.w5(32'hba19576c),
	.w6(32'hbb0a7c5a),
	.w7(32'hbb8fc495),
	.w8(32'hbc30412b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9f6b2),
	.w1(32'h3aa99622),
	.w2(32'hbb0f57fc),
	.w3(32'h3b045642),
	.w4(32'h3a3ceef9),
	.w5(32'hba61a1ac),
	.w6(32'hbb88fa63),
	.w7(32'hbbe3bb25),
	.w8(32'hbc1baac8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b4ced),
	.w1(32'h3b943063),
	.w2(32'h3abc4deb),
	.w3(32'hb7eac2a2),
	.w4(32'h3b122a5b),
	.w5(32'hba117976),
	.w6(32'hbc36faca),
	.w7(32'hbc229731),
	.w8(32'hbc3d961d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb736b),
	.w1(32'h3ae186ee),
	.w2(32'hb892d58d),
	.w3(32'h37c2385c),
	.w4(32'h3b328e9f),
	.w5(32'hb8176789),
	.w6(32'hbb028354),
	.w7(32'hbb0329c8),
	.w8(32'hbbb4ad09),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbff90),
	.w1(32'h3bb1c052),
	.w2(32'hbaca495d),
	.w3(32'h3c06c136),
	.w4(32'h3ab0c3f5),
	.w5(32'hbb6e2e48),
	.w6(32'hbbccca6e),
	.w7(32'hbb65f532),
	.w8(32'hbc21d44b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ae3b1),
	.w1(32'hba753d81),
	.w2(32'hba4cd96a),
	.w3(32'h39861cf9),
	.w4(32'hba3e49f0),
	.w5(32'hba682f8a),
	.w6(32'hba46a14f),
	.w7(32'hba9f5c65),
	.w8(32'hba7f3a5a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab714e7),
	.w1(32'hbab65d17),
	.w2(32'hbadd002e),
	.w3(32'hbadc594d),
	.w4(32'hbaa4473a),
	.w5(32'hbab0f3c8),
	.w6(32'hba963180),
	.w7(32'hbabddd1c),
	.w8(32'hba48122a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a27a2),
	.w1(32'hb8427690),
	.w2(32'h39cc9da3),
	.w3(32'hba6aee7c),
	.w4(32'h3a17e444),
	.w5(32'h3a5629e6),
	.w6(32'h39c17d71),
	.w7(32'h39e6c461),
	.w8(32'h3a883788),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3df881),
	.w1(32'h39ca620b),
	.w2(32'hba99736e),
	.w3(32'hb9850bf1),
	.w4(32'hba85eb1d),
	.w5(32'hba5d2413),
	.w6(32'hb99b3623),
	.w7(32'hbb393b73),
	.w8(32'hbbf3fa8f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8562bf),
	.w1(32'h3a6e42a4),
	.w2(32'h39d92e5a),
	.w3(32'h39f9b284),
	.w4(32'h3aa395de),
	.w5(32'hb9d540bf),
	.w6(32'h3693fab2),
	.w7(32'hb785f3c0),
	.w8(32'hba0c3b36),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affd1a9),
	.w1(32'h3ae19fa5),
	.w2(32'hbaa4f5dd),
	.w3(32'h3b2bb2e3),
	.w4(32'hba530b10),
	.w5(32'hbb4ed750),
	.w6(32'hbbb3fdb2),
	.w7(32'hbb91b7d9),
	.w8(32'hbc17db89),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e6ab8),
	.w1(32'h399af8ae),
	.w2(32'hb9ac999f),
	.w3(32'hba0a0b3c),
	.w4(32'hba144072),
	.w5(32'hbac2739f),
	.w6(32'hb82c9a5e),
	.w7(32'hbabcb437),
	.w8(32'hbb20d672),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d56527),
	.w1(32'h3a8169e4),
	.w2(32'hb915402d),
	.w3(32'h38de37e7),
	.w4(32'h3a6aac7d),
	.w5(32'hb98169db),
	.w6(32'h3a8f4cbd),
	.w7(32'h398dd86b),
	.w8(32'h3a8d6905),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3955ea07),
	.w1(32'hb887e89b),
	.w2(32'hb9c4278d),
	.w3(32'h3a13036c),
	.w4(32'hb873cc88),
	.w5(32'h38e4e0cd),
	.w6(32'h395ac6d6),
	.w7(32'hba15359d),
	.w8(32'h38834789),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cb754),
	.w1(32'hb79a0898),
	.w2(32'hbb253729),
	.w3(32'h393ac5ac),
	.w4(32'hb9f138b5),
	.w5(32'hbb34913d),
	.w6(32'hb8f7706e),
	.w7(32'hbb06f5ff),
	.w8(32'hbacea196),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f6436),
	.w1(32'hb92d5424),
	.w2(32'hba4bf8d2),
	.w3(32'hba60c418),
	.w4(32'h38c6a67f),
	.w5(32'hb87ee21c),
	.w6(32'hba287ebb),
	.w7(32'hb9a33399),
	.w8(32'hb8a2cd8b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87c0c3),
	.w1(32'hba28602a),
	.w2(32'hba6d869d),
	.w3(32'h3acb9e58),
	.w4(32'hba47b2d4),
	.w5(32'hbaaafbdc),
	.w6(32'hb9a6957d),
	.w7(32'hba4412ed),
	.w8(32'hba315e45),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39924f88),
	.w1(32'hba5897cd),
	.w2(32'hbb3fb3f7),
	.w3(32'h397ec48b),
	.w4(32'hbad17af7),
	.w5(32'hbb4be24f),
	.w6(32'hbb92d038),
	.w7(32'hbb6209e4),
	.w8(32'hbbc70b2e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab6fc3),
	.w1(32'hbadf3605),
	.w2(32'hbb10ce63),
	.w3(32'h3a45ca34),
	.w4(32'hbab95af6),
	.w5(32'hba61b512),
	.w6(32'h3b8d2567),
	.w7(32'h3b046dd8),
	.w8(32'hbacbe940),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae09ee7),
	.w1(32'h3b012d75),
	.w2(32'h39ea3bb8),
	.w3(32'hb9d78f78),
	.w4(32'hb928b4c0),
	.w5(32'h3ac29424),
	.w6(32'h3ac62b0d),
	.w7(32'h3a5876fc),
	.w8(32'h39c92c6a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3445f7),
	.w1(32'h3a6b8d04),
	.w2(32'h3aa55436),
	.w3(32'h3a94d305),
	.w4(32'h3a46f081),
	.w5(32'h3ab1d539),
	.w6(32'h3aa39174),
	.w7(32'h3a969f79),
	.w8(32'h3abbd53a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addcdf4),
	.w1(32'hba10bdcb),
	.w2(32'hb99a86ff),
	.w3(32'h3ac11099),
	.w4(32'h38bfd8ce),
	.w5(32'h38861428),
	.w6(32'hba33b5ac),
	.w7(32'hb99a67c8),
	.w8(32'hba064a28),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff8dc7),
	.w1(32'hba787c67),
	.w2(32'hbb16fd4a),
	.w3(32'hb89078c6),
	.w4(32'hba9c4a7b),
	.w5(32'hbb365f6a),
	.w6(32'hba92c863),
	.w7(32'hbb24ae00),
	.w8(32'hbb15f978),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc535f6a),
	.w1(32'hbba1a050),
	.w2(32'hbb08b484),
	.w3(32'h3b94b051),
	.w4(32'h3ba92ede),
	.w5(32'h3b89d927),
	.w6(32'h3accd5ba),
	.w7(32'hba702dfc),
	.w8(32'hbb80872a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1577f),
	.w1(32'h3b4fa7b4),
	.w2(32'hba5cd383),
	.w3(32'hbad4263b),
	.w4(32'hba8e3b16),
	.w5(32'hbbd14dce),
	.w6(32'hbc882531),
	.w7(32'hbc44c1ab),
	.w8(32'hbc751804),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90ca08),
	.w1(32'h3b1fc8bb),
	.w2(32'hbb229b5d),
	.w3(32'hbb3db496),
	.w4(32'h3932c4c7),
	.w5(32'hbbd8d94b),
	.w6(32'hbc004d01),
	.w7(32'hbbba5710),
	.w8(32'hbc49509d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16a544),
	.w1(32'h3ba759ca),
	.w2(32'hbb47a516),
	.w3(32'h39d35be7),
	.w4(32'h3acab631),
	.w5(32'hbb5d174e),
	.w6(32'hbc00f310),
	.w7(32'hbc7074a4),
	.w8(32'hbc9c61c4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb000af2),
	.w1(32'hb960765b),
	.w2(32'hb8c6d0c4),
	.w3(32'hbaf23d97),
	.w4(32'hb9bb836f),
	.w5(32'hb8b1e9b4),
	.w6(32'h37970d99),
	.w7(32'hb939d7d0),
	.w8(32'h392285c1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907fe37),
	.w1(32'hba6277b9),
	.w2(32'hba98c3aa),
	.w3(32'h3a037c8f),
	.w4(32'hb9e6c95a),
	.w5(32'hba6bbdd6),
	.w6(32'hba400123),
	.w7(32'hba951e95),
	.w8(32'hb9dadd13),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f87b0),
	.w1(32'hba1ab11a),
	.w2(32'hba5b3fc0),
	.w3(32'hb9a9b247),
	.w4(32'hb9caabbe),
	.w5(32'hba27d9d5),
	.w6(32'hb9d0f1de),
	.w7(32'hba28f901),
	.w8(32'hb8d1b09e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ab3e3),
	.w1(32'hb9b012b2),
	.w2(32'hbac6d175),
	.w3(32'h3a8b7539),
	.w4(32'h3a127e44),
	.w5(32'hbac8951f),
	.w6(32'hbac02e66),
	.w7(32'hbab9d9c2),
	.w8(32'hbaf147a2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad15f0a),
	.w1(32'hbad5a088),
	.w2(32'hba935c26),
	.w3(32'hbab7aeb1),
	.w4(32'hbaae9289),
	.w5(32'hb9971dfb),
	.w6(32'hbab24cb2),
	.w7(32'hba8d7421),
	.w8(32'hba080a93),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97bbf6),
	.w1(32'hbb2461ce),
	.w2(32'h3a86b2fd),
	.w3(32'h39a92de3),
	.w4(32'hbb0dbb1e),
	.w5(32'hbaaa2859),
	.w6(32'hbb5ad724),
	.w7(32'hbb653505),
	.w8(32'hbb8ef2da),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb188bc2),
	.w1(32'hba7c991a),
	.w2(32'hbb1d3db2),
	.w3(32'h3982dd4f),
	.w4(32'hba637cfa),
	.w5(32'hbb7d7cde),
	.w6(32'hbc0e062a),
	.w7(32'hbb723b38),
	.w8(32'hbb44e1ad),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a2965),
	.w1(32'h3b0edbcc),
	.w2(32'hb9defcdc),
	.w3(32'h3ad13d85),
	.w4(32'h3ac4f85e),
	.w5(32'h3a9836be),
	.w6(32'hb9fd290a),
	.w7(32'hbb8fb2ae),
	.w8(32'hbba1a110),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a2638),
	.w1(32'hba4bac43),
	.w2(32'hbace412c),
	.w3(32'h3a13d098),
	.w4(32'hba07ad11),
	.w5(32'hbb03679f),
	.w6(32'hbb50db94),
	.w7(32'hbb3857e1),
	.w8(32'hbb9d921e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e74bf),
	.w1(32'hbb3df8c5),
	.w2(32'hbb90e11e),
	.w3(32'h3afe043f),
	.w4(32'h3a2e2976),
	.w5(32'h39d904cd),
	.w6(32'h3a524356),
	.w7(32'hba15aed5),
	.w8(32'hbace51da),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37584d),
	.w1(32'hb88d8dfa),
	.w2(32'hbad843ec),
	.w3(32'hba7b68f6),
	.w4(32'hb8e78f38),
	.w5(32'hbaac7bf1),
	.w6(32'hba0c61a4),
	.w7(32'hbb28eee8),
	.w8(32'hbb8b1104),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1fdde),
	.w1(32'h3a67ee39),
	.w2(32'hba9a0bff),
	.w3(32'h3b083c45),
	.w4(32'h393e82ec),
	.w5(32'hba56ce56),
	.w6(32'hbb3b1505),
	.w7(32'hbb33fba7),
	.w8(32'hbb872eb7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39976138),
	.w1(32'h3a70a624),
	.w2(32'h39d6d21a),
	.w3(32'h399f683d),
	.w4(32'h3a699951),
	.w5(32'h3a261dc4),
	.w6(32'h3a876118),
	.w7(32'h3a0be712),
	.w8(32'h3a355598),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3935b659),
	.w1(32'hba6f51f8),
	.w2(32'hb9bfb006),
	.w3(32'h39c0856e),
	.w4(32'hb9dc4fc6),
	.w5(32'h3a063d25),
	.w6(32'hba9cec3c),
	.w7(32'hba7bac80),
	.w8(32'hb9bf7c9b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e01280),
	.w1(32'hb9314203),
	.w2(32'h39f65ef8),
	.w3(32'h3a380cbf),
	.w4(32'h391dff46),
	.w5(32'h3a252a47),
	.w6(32'hbac4847c),
	.w7(32'hb983204f),
	.w8(32'hba93a6d1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c205f),
	.w1(32'h3a7be90e),
	.w2(32'h3aa07b8a),
	.w3(32'h3a313202),
	.w4(32'h39b13019),
	.w5(32'h3a1c36b9),
	.w6(32'h3a97d4ea),
	.w7(32'h3a12a052),
	.w8(32'h3a5e192e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e2ef7),
	.w1(32'h3b12715a),
	.w2(32'hba5eeba9),
	.w3(32'hbb02aedf),
	.w4(32'h3aac7eb6),
	.w5(32'hba2a4b6a),
	.w6(32'hbbaabb20),
	.w7(32'hbb626e74),
	.w8(32'hbb9588ed),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925b1ed),
	.w1(32'h3a62a479),
	.w2(32'hba91f370),
	.w3(32'h3901965c),
	.w4(32'h3aa90946),
	.w5(32'hba208f4e),
	.w6(32'h393ed805),
	.w7(32'h39d0c790),
	.w8(32'hb9292695),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d27ad6),
	.w1(32'h3aa1218d),
	.w2(32'h3b2754e3),
	.w3(32'hbb684305),
	.w4(32'hba09492c),
	.w5(32'hb9d28eae),
	.w6(32'hbb8d97d7),
	.w7(32'hbb8c1357),
	.w8(32'hbb5d4a04),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb72b12),
	.w1(32'hbb1ac51c),
	.w2(32'hbb944a56),
	.w3(32'hbb1e6875),
	.w4(32'hbb8031eb),
	.w5(32'hbb9e3bd4),
	.w6(32'hbc39845a),
	.w7(32'hbbb18950),
	.w8(32'hbc0fe573),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd4afb),
	.w1(32'h3af817e4),
	.w2(32'hbb095668),
	.w3(32'h3b8155c2),
	.w4(32'h3a537713),
	.w5(32'hbb318a6b),
	.w6(32'h3bc12a83),
	.w7(32'hba03ede6),
	.w8(32'hbb66626e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbebb08),
	.w1(32'hbb726756),
	.w2(32'hbbad8e62),
	.w3(32'h3b725e8c),
	.w4(32'h3b60a377),
	.w5(32'h3b85d9d3),
	.w6(32'hbbd5bfb8),
	.w7(32'hba6b7ed9),
	.w8(32'hbb977cf6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be455b4),
	.w1(32'h3bcfc91e),
	.w2(32'h3b0fbf98),
	.w3(32'h3b0f46f0),
	.w4(32'h3ab0e85c),
	.w5(32'hba8b7a29),
	.w6(32'hbb2742bd),
	.w7(32'hbb76b1b7),
	.w8(32'hbba23f42),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae4863),
	.w1(32'hbba329f9),
	.w2(32'hbba3dada),
	.w3(32'hbb85df62),
	.w4(32'hbada7dec),
	.w5(32'hbb180b24),
	.w6(32'hbc228999),
	.w7(32'hbbc5526b),
	.w8(32'hbbeea3a8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb749a63),
	.w1(32'hbb819c7c),
	.w2(32'hbb1e41a5),
	.w3(32'h3a565737),
	.w4(32'hba8c7e78),
	.w5(32'hba047271),
	.w6(32'hbab22bdd),
	.w7(32'hbaef5027),
	.w8(32'hbb8caf7b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b174bc2),
	.w1(32'h3a65ae15),
	.w2(32'h3a6f88f8),
	.w3(32'h3b52eca2),
	.w4(32'h3b42147e),
	.w5(32'hb992fc0a),
	.w6(32'h3b8e27db),
	.w7(32'hb9fde4fd),
	.w8(32'hbb86b1ce),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09f77b),
	.w1(32'h3a5501ec),
	.w2(32'h388a2436),
	.w3(32'hb9f56566),
	.w4(32'hb9c00820),
	.w5(32'hb8f3f9cb),
	.w6(32'h3a893777),
	.w7(32'h3aa1fb90),
	.w8(32'hba9d521b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1e687),
	.w1(32'h3b9541c9),
	.w2(32'hba70330e),
	.w3(32'hba2f95eb),
	.w4(32'h398e4fe1),
	.w5(32'hbb0479b6),
	.w6(32'hbb8362f4),
	.w7(32'hbbb625dc),
	.w8(32'hbc18eb6b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949a496),
	.w1(32'hba909299),
	.w2(32'hbb822991),
	.w3(32'h3b9e46b7),
	.w4(32'hbb604595),
	.w5(32'hbb93c3b6),
	.w6(32'hbb8825b5),
	.w7(32'hbc06d14a),
	.w8(32'hbc12b8f5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaba10f),
	.w1(32'h3bd7c15b),
	.w2(32'hbbf3d9cf),
	.w3(32'h3acc8e4d),
	.w4(32'h3b9facd3),
	.w5(32'hbad33b9f),
	.w6(32'hbc512d8d),
	.w7(32'h3a737854),
	.w8(32'hbb72e096),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d8e1f),
	.w1(32'h3bca3c53),
	.w2(32'hbb543c99),
	.w3(32'h3a03666f),
	.w4(32'h3bd7c68b),
	.w5(32'hb93c3b40),
	.w6(32'hbab36bf9),
	.w7(32'hbaac6a8a),
	.w8(32'hbb16afbc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87a503),
	.w1(32'h3b934a57),
	.w2(32'h3af548be),
	.w3(32'hb9b8445e),
	.w4(32'h3a9487e7),
	.w5(32'hbb1077b2),
	.w6(32'hbb444c04),
	.w7(32'hbbc24241),
	.w8(32'hbc0c578b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8241b),
	.w1(32'hbb6b5350),
	.w2(32'hbc1ea936),
	.w3(32'hba977bcc),
	.w4(32'hb8d0bab3),
	.w5(32'hbaf48342),
	.w6(32'hbc12d4e8),
	.w7(32'hba1ac226),
	.w8(32'hbb74dfc9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3ec55),
	.w1(32'hba7cf462),
	.w2(32'hbab99dfe),
	.w3(32'hbab815b0),
	.w4(32'hb9a886d6),
	.w5(32'hba8ab2ed),
	.w6(32'hba1cee9f),
	.w7(32'hba6eab24),
	.w8(32'hb9639e37),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe224ff),
	.w1(32'hbbae8b7d),
	.w2(32'hbc60ce46),
	.w3(32'hba2a1e16),
	.w4(32'h3b7a0a66),
	.w5(32'hbc27104f),
	.w6(32'hbc051a55),
	.w7(32'h3a0dd916),
	.w8(32'hbb4731de),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64c9dc),
	.w1(32'h3b99f52e),
	.w2(32'hbb861c87),
	.w3(32'h3b050b90),
	.w4(32'h39c5dffc),
	.w5(32'hbbbbe22a),
	.w6(32'hbaaec669),
	.w7(32'hbb22534c),
	.w8(32'hbbbb0a19),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b5457),
	.w1(32'hba4e6599),
	.w2(32'hba096675),
	.w3(32'hba5a17f3),
	.w4(32'hb95f4c06),
	.w5(32'hb8b3df31),
	.w6(32'hb956f8c6),
	.w7(32'hb977e6c4),
	.w8(32'hb79c5093),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0d411),
	.w1(32'hba162151),
	.w2(32'hba5d0783),
	.w3(32'hbaca283a),
	.w4(32'hba29a5c7),
	.w5(32'hba6602c8),
	.w6(32'hbb00040e),
	.w7(32'hbad88269),
	.w8(32'hbb373e3c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b841e5e),
	.w1(32'h3b5fb958),
	.w2(32'hba37debe),
	.w3(32'h3b9610e7),
	.w4(32'h3b740bb3),
	.w5(32'hbabcff6e),
	.w6(32'hbb07c907),
	.w7(32'hbb3b8451),
	.w8(32'hbbd484ab),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b713d7e),
	.w1(32'h3b0ada9c),
	.w2(32'hba1549d3),
	.w3(32'h3a4ed2d2),
	.w4(32'h3abbb177),
	.w5(32'h3ab2bb7c),
	.w6(32'hb8ba2c75),
	.w7(32'hbb596141),
	.w8(32'hbb8c5811),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea45c3),
	.w1(32'h39963758),
	.w2(32'h38959902),
	.w3(32'h3b9dfcb6),
	.w4(32'h3abf402d),
	.w5(32'hba5d0ea2),
	.w6(32'h3b83330f),
	.w7(32'hbaec16d6),
	.w8(32'hbb930f36),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bae80),
	.w1(32'h3b00a058),
	.w2(32'hbacfc37d),
	.w3(32'h3b2c348b),
	.w4(32'h3aa0d10e),
	.w5(32'hba9cb2f8),
	.w6(32'h3b00fa65),
	.w7(32'hbb626142),
	.w8(32'hbbb1d59c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97fc1f),
	.w1(32'h3bffb8b0),
	.w2(32'h3b7b2a01),
	.w3(32'hbb8b239b),
	.w4(32'hb9ab793b),
	.w5(32'hbaebe638),
	.w6(32'hbbdd9c1b),
	.w7(32'hbb7211cf),
	.w8(32'hbb60ef1b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea2388),
	.w1(32'hbc083b47),
	.w2(32'hbc06f8da),
	.w3(32'hb9cecc6d),
	.w4(32'hbad15d05),
	.w5(32'hbaf0cea7),
	.w6(32'hbb113174),
	.w7(32'hbade740b),
	.w8(32'hbb878195),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e265d),
	.w1(32'hba6f3fca),
	.w2(32'hbb285afb),
	.w3(32'h388eecc6),
	.w4(32'hbb05016a),
	.w5(32'hbb51eb58),
	.w6(32'hbb7ef002),
	.w7(32'hbb9cce28),
	.w8(32'hbbc28907),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c5c80),
	.w1(32'hba8d72ce),
	.w2(32'hbad75eda),
	.w3(32'hbb3b0903),
	.w4(32'hb9ad5dfb),
	.w5(32'hbaa61b48),
	.w6(32'hba1303fb),
	.w7(32'hba884e6d),
	.w8(32'hb97cdecf),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04eba4),
	.w1(32'hbad1adb5),
	.w2(32'hba9e0797),
	.w3(32'hba98246e),
	.w4(32'h39404f9f),
	.w5(32'hba0fd753),
	.w6(32'hba10f3b5),
	.w7(32'hba34ca66),
	.w8(32'hb97866cf),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4aac29),
	.w1(32'hb9b63ac8),
	.w2(32'hba6a8270),
	.w3(32'hb9f73da4),
	.w4(32'hb90eec33),
	.w5(32'hba54a4bf),
	.w6(32'hb9501acc),
	.w7(32'hba2534ed),
	.w8(32'hb9b000c8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba418c11),
	.w1(32'hbaaadcf8),
	.w2(32'hbacd6514),
	.w3(32'hb9dc92dd),
	.w4(32'h38ce76d3),
	.w5(32'hb9912819),
	.w6(32'hba6626c3),
	.w7(32'hbaba9024),
	.w8(32'hbb0aa8ca),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20f4f3),
	.w1(32'h3aec2d40),
	.w2(32'h390f33bb),
	.w3(32'hba02ef1a),
	.w4(32'h3a7a902a),
	.w5(32'hba173cbd),
	.w6(32'hbb7cfc22),
	.w7(32'hbb959cfa),
	.w8(32'hbbb600b1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0067e2),
	.w1(32'hba096b9e),
	.w2(32'hba8edba7),
	.w3(32'hba812a5b),
	.w4(32'h375a153a),
	.w5(32'hba66e514),
	.w6(32'hb944de49),
	.w7(32'hba49a632),
	.w8(32'hba66b531),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd8f95),
	.w1(32'h3a6d9412),
	.w2(32'hba31a720),
	.w3(32'h39f92898),
	.w4(32'h39f13367),
	.w5(32'h39874b98),
	.w6(32'hbabdf26c),
	.w7(32'hbb0eb13d),
	.w8(32'hbb369da3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf5105),
	.w1(32'h3a336213),
	.w2(32'hbba827d0),
	.w3(32'h3b905990),
	.w4(32'h3b17cc78),
	.w5(32'hbb536eff),
	.w6(32'h3b99cf0f),
	.w7(32'hbb2ddf00),
	.w8(32'hbc11c728),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78294d),
	.w1(32'hb93b1c42),
	.w2(32'h3ae39617),
	.w3(32'hb9b5a518),
	.w4(32'h3a41992e),
	.w5(32'h3a515a83),
	.w6(32'hba37e4ac),
	.w7(32'h3a619eff),
	.w8(32'hba858a7b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8ac99),
	.w1(32'h3b262640),
	.w2(32'h3b24d930),
	.w3(32'hb9d227b8),
	.w4(32'h3b2aa3aa),
	.w5(32'h3ae9707f),
	.w6(32'h3b06c92a),
	.w7(32'h3acacf6c),
	.w8(32'h3ad1f4ba),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08e246),
	.w1(32'hba334225),
	.w2(32'hbac14130),
	.w3(32'h3aa6d903),
	.w4(32'h3820dfb9),
	.w5(32'hba6e2e25),
	.w6(32'hb7ef5693),
	.w7(32'hba435cf7),
	.w8(32'hba04f380),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba133edb),
	.w1(32'h39a3c621),
	.w2(32'hb8eff103),
	.w3(32'hb9e15ac3),
	.w4(32'hb98cbf10),
	.w5(32'hba50ecd5),
	.w6(32'hb9a6055d),
	.w7(32'hba49f85d),
	.w8(32'hba2a9fa7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47247f),
	.w1(32'h3b7c1a6d),
	.w2(32'h39491859),
	.w3(32'hbb032fcd),
	.w4(32'hbbb477a0),
	.w5(32'hbb67b70c),
	.w6(32'hbbe98981),
	.w7(32'hbb613211),
	.w8(32'hbbc61a28),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59f655),
	.w1(32'h3b160dbe),
	.w2(32'hb9101338),
	.w3(32'h3b554e93),
	.w4(32'h3a10dafe),
	.w5(32'hbac61da2),
	.w6(32'hbaad1bec),
	.w7(32'hbb03b10c),
	.w8(32'hbbcdc5f7),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba471c37),
	.w1(32'h3910efac),
	.w2(32'hb98a61c6),
	.w3(32'h3a3a6807),
	.w4(32'h3a84a3dd),
	.w5(32'h39e62605),
	.w6(32'h370c5741),
	.w7(32'h383e87bf),
	.w8(32'hb9a6a388),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff62ad),
	.w1(32'hb9d7d5a9),
	.w2(32'hba48d185),
	.w3(32'h3a4d149e),
	.w4(32'h3a379429),
	.w5(32'hbad0f5a7),
	.w6(32'hbb23cd9b),
	.w7(32'hba90adfa),
	.w8(32'hbab95471),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06beb5),
	.w1(32'hb7e91973),
	.w2(32'hb7562b1b),
	.w3(32'hb887c61e),
	.w4(32'h39f1b9be),
	.w5(32'hb53eafd5),
	.w6(32'h39467b7e),
	.w7(32'hba2c299f),
	.w8(32'hba92d600),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369325ef),
	.w1(32'hb63556ea),
	.w2(32'h388c6074),
	.w3(32'h3a4fe093),
	.w4(32'h3a9ec147),
	.w5(32'h3a94eaeb),
	.w6(32'hbaa7c890),
	.w7(32'hb9a55dc6),
	.w8(32'hba8e7aa7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86750e),
	.w1(32'hbb847d62),
	.w2(32'hbb56219a),
	.w3(32'h38365c05),
	.w4(32'h3903af5c),
	.w5(32'hb9ce1c97),
	.w6(32'h3a5b89c1),
	.w7(32'hb8247403),
	.w8(32'hbb6e65be),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad18603),
	.w1(32'h3ad4ed7f),
	.w2(32'hbb69b74d),
	.w3(32'h3b5d2efb),
	.w4(32'hb9a0f0b8),
	.w5(32'hbad9ebdd),
	.w6(32'hbb4706c1),
	.w7(32'hbb9e5ce9),
	.w8(32'hbc09b732),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93594b),
	.w1(32'h3a904c96),
	.w2(32'hba029cda),
	.w3(32'h3a67e9d7),
	.w4(32'h3a910caf),
	.w5(32'hb59d5b1a),
	.w6(32'h3987b8cb),
	.w7(32'hbb0c0237),
	.w8(32'hbb532d10),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33e81f),
	.w1(32'h39886734),
	.w2(32'hba8f1db2),
	.w3(32'h3a9bcaa7),
	.w4(32'h3a81f4fb),
	.w5(32'h3a0d7af1),
	.w6(32'hbb9290cd),
	.w7(32'hbb151dc5),
	.w8(32'hbb9fd5bf),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaea0e4),
	.w1(32'hbac8b333),
	.w2(32'hbb030f58),
	.w3(32'h39f44e30),
	.w4(32'hba5f17af),
	.w5(32'hba8cc951),
	.w6(32'hbb9ede61),
	.w7(32'hbb4625ab),
	.w8(32'hbb9e36fb),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd411f),
	.w1(32'h3b4e61df),
	.w2(32'h3b257d8d),
	.w3(32'hbad6d7d6),
	.w4(32'h3a88cd2d),
	.w5(32'h3ab6ec10),
	.w6(32'hbbc4926c),
	.w7(32'hbb4d4f2d),
	.w8(32'hbb4dc3b4),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e68c5),
	.w1(32'h39ae785d),
	.w2(32'hba74553c),
	.w3(32'h3b28c944),
	.w4(32'h3a869b3b),
	.w5(32'hba65897d),
	.w6(32'hbaf54f49),
	.w7(32'hbac550c5),
	.w8(32'hbb51df5a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c6cb5),
	.w1(32'h3a4328fc),
	.w2(32'hb99c397a),
	.w3(32'h3a11b862),
	.w4(32'h398b686e),
	.w5(32'hba2c1257),
	.w6(32'hba78dcd7),
	.w7(32'hbaa5d9ee),
	.w8(32'hbaf47575),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b16da),
	.w1(32'hb95ecb3d),
	.w2(32'hb8e4f056),
	.w3(32'h3c23e535),
	.w4(32'hb9ecb07e),
	.w5(32'hbb569b0d),
	.w6(32'h3c47710a),
	.w7(32'hbb1480d4),
	.w8(32'hbbc62541),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cceb51),
	.w1(32'hb95b1f4e),
	.w2(32'hb9bc1e30),
	.w3(32'hba86df9b),
	.w4(32'hba8f0583),
	.w5(32'hba6b23e0),
	.w6(32'hbb1bc9c4),
	.w7(32'hbadbc10f),
	.w8(32'hbb36fb8c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b81bc),
	.w1(32'h39614f14),
	.w2(32'h394d6c80),
	.w3(32'hb99c0177),
	.w4(32'h39264dee),
	.w5(32'h391c7f63),
	.w6(32'h3911cf7c),
	.w7(32'hb7b5ab53),
	.w8(32'hb79c4d9f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3977fdcd),
	.w1(32'hb9ee720f),
	.w2(32'hb877eb0b),
	.w3(32'h3903ccc9),
	.w4(32'hb911365a),
	.w5(32'hb80076b4),
	.w6(32'hba054384),
	.w7(32'hb836ecb8),
	.w8(32'hb92317c7),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac87998),
	.w1(32'h3aa19354),
	.w2(32'hb9a06ee2),
	.w3(32'h3a2623cd),
	.w4(32'h3a8f882a),
	.w5(32'hba153b08),
	.w6(32'hba972a4d),
	.w7(32'hba7614de),
	.w8(32'hbad9f946),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39296135),
	.w1(32'h3a36861e),
	.w2(32'hb9baf168),
	.w3(32'hbab707b2),
	.w4(32'h3a595822),
	.w5(32'hb83e10c4),
	.w6(32'hbb7bfe02),
	.w7(32'hbba99366),
	.w8(32'hbb99558f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf6ff0),
	.w1(32'h3b9dca5e),
	.w2(32'h39b410b3),
	.w3(32'h3b965b90),
	.w4(32'h3b3fcae0),
	.w5(32'hba9fccf0),
	.w6(32'hbb22f815),
	.w7(32'hbb8866a6),
	.w8(32'hbbec1064),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8600e60),
	.w1(32'hba06a2dc),
	.w2(32'hba51f478),
	.w3(32'hb887ac33),
	.w4(32'hba045d89),
	.w5(32'hba1dae93),
	.w6(32'hb9b12bb8),
	.w7(32'hba0d76c7),
	.w8(32'hb92b052a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03102c),
	.w1(32'h3ada9119),
	.w2(32'hba49489e),
	.w3(32'h3b44b73f),
	.w4(32'h3b05f2cd),
	.w5(32'hbaaab5ba),
	.w6(32'hbb0c7088),
	.w7(32'hbb3f8440),
	.w8(32'hbbbb7d37),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03d0bf),
	.w1(32'h3b03a254),
	.w2(32'h397b72b9),
	.w3(32'h3a9bf85b),
	.w4(32'h3a4bb625),
	.w5(32'hb9a78b17),
	.w6(32'hbb1aeb84),
	.w7(32'hbb48d69a),
	.w8(32'hbb8335a1),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb969507),
	.w1(32'hbb865b4b),
	.w2(32'hbb60ed9b),
	.w3(32'hbaa73aeb),
	.w4(32'hb8555871),
	.w5(32'h3b1d09ea),
	.w6(32'hbbb14e90),
	.w7(32'hbb5683ef),
	.w8(32'hbb6a7b67),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c296230),
	.w1(32'h39c1d084),
	.w2(32'h3a804484),
	.w3(32'h3c19b91d),
	.w4(32'h3a1fdf5a),
	.w5(32'hbb12b9d8),
	.w6(32'h3bf80456),
	.w7(32'hbbe4e60b),
	.w8(32'hbc4682ed),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba516c0f),
	.w1(32'hba15d3f8),
	.w2(32'hbae2c0a9),
	.w3(32'hba8e1b9a),
	.w4(32'h3a4ae5f2),
	.w5(32'hb7f6aa6a),
	.w6(32'hba772802),
	.w7(32'h3a0305a2),
	.w8(32'hb850b378),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73b7549),
	.w1(32'h39d44cfe),
	.w2(32'h39b8d04b),
	.w3(32'h38c4135f),
	.w4(32'h398e2e44),
	.w5(32'h399581da),
	.w6(32'h395f3a77),
	.w7(32'h3989a655),
	.w8(32'h399eddca),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e645c),
	.w1(32'h3b327146),
	.w2(32'h3ad8b309),
	.w3(32'h39993801),
	.w4(32'h399ea30b),
	.w5(32'hb81ee6e1),
	.w6(32'hba668b5b),
	.w7(32'hbb18e897),
	.w8(32'hbb454bda),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f83b6),
	.w1(32'h3a7e151a),
	.w2(32'hb9cdceb3),
	.w3(32'hbb1d3659),
	.w4(32'h39e81226),
	.w5(32'hba153fa2),
	.w6(32'hbb4eb67a),
	.w7(32'hba8aaa49),
	.w8(32'hbb36c72e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bc1f9),
	.w1(32'h3ac6cc51),
	.w2(32'hba8ec29e),
	.w3(32'hb9b020c2),
	.w4(32'h3ac3458e),
	.w5(32'hb9a78d3b),
	.w6(32'h385a6458),
	.w7(32'hb9902d61),
	.w8(32'hbb00105f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab4e2e),
	.w1(32'hba00d319),
	.w2(32'hbabbba09),
	.w3(32'h3a32330a),
	.w4(32'h3a55cfa9),
	.w5(32'h39afc4ab),
	.w6(32'hbb00690a),
	.w7(32'hbabddb44),
	.w8(32'hbad9e390),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0937b),
	.w1(32'hb9cc3af0),
	.w2(32'hb9d5cdca),
	.w3(32'hb9cceff4),
	.w4(32'hb995d510),
	.w5(32'hb92c578b),
	.w6(32'hb9cbd4bc),
	.w7(32'hba0af064),
	.w8(32'hb9af3c4e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9173d24),
	.w1(32'h3905d358),
	.w2(32'hb7aa3326),
	.w3(32'h3b1603c5),
	.w4(32'h3a1ae78b),
	.w5(32'hba3edc2f),
	.w6(32'hbb532024),
	.w7(32'hbad7b203),
	.w8(32'hbb702325),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3878f569),
	.w1(32'h36f40358),
	.w2(32'hba906371),
	.w3(32'h3a1e85a8),
	.w4(32'hb9ab408a),
	.w5(32'hb9e155ce),
	.w6(32'h3881e408),
	.w7(32'hba2fabe2),
	.w8(32'hba8642bf),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64dc2b),
	.w1(32'h399fc95a),
	.w2(32'h39b4ed7e),
	.w3(32'h39063a04),
	.w4(32'hbac9fd56),
	.w5(32'hbaecc84f),
	.w6(32'h3a4884c8),
	.w7(32'hbb35ab32),
	.w8(32'hbb85ae61),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bf523e),
	.w1(32'h39313dfc),
	.w2(32'h37a3c672),
	.w3(32'h396c525a),
	.w4(32'h38cae0c6),
	.w5(32'hb8ce54ea),
	.w6(32'h38001d76),
	.w7(32'h38443d91),
	.w8(32'h38227a86),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac81f9),
	.w1(32'h3b9e0237),
	.w2(32'hbb03bf44),
	.w3(32'h3b45445b),
	.w4(32'h3aa5cbb9),
	.w5(32'hbb8b28c2),
	.w6(32'h3ae235a9),
	.w7(32'h3aa3b3b3),
	.w8(32'hbb8cc261),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e75337),
	.w1(32'h39ec8433),
	.w2(32'h3970aea1),
	.w3(32'hb7b2da54),
	.w4(32'h3a01c207),
	.w5(32'h39d55409),
	.w6(32'h39efde83),
	.w7(32'h39a932fb),
	.w8(32'h39ed2bb9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980cd4b),
	.w1(32'hb887c72f),
	.w2(32'h3645703b),
	.w3(32'h39c76c9a),
	.w4(32'hb8f459c3),
	.w5(32'hb94dd3a0),
	.w6(32'hb894c0f0),
	.w7(32'hb8cbdb39),
	.w8(32'hb8b671f9),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a007eb6),
	.w1(32'h3a8343df),
	.w2(32'h3a0c706f),
	.w3(32'hb93b04bf),
	.w4(32'h3ab5563a),
	.w5(32'h3a3145cd),
	.w6(32'hb9dca1bf),
	.w7(32'hba0bcbda),
	.w8(32'hbaca6a6f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83a5e5),
	.w1(32'h3bc7e302),
	.w2(32'h39837154),
	.w3(32'h39051e79),
	.w4(32'h3b48e048),
	.w5(32'hbb7ed0a8),
	.w6(32'hbc3dca2b),
	.w7(32'hbb871cbf),
	.w8(32'hbc00ab7c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38433e97),
	.w1(32'h3a933508),
	.w2(32'hba8f7dd3),
	.w3(32'hb8f1d574),
	.w4(32'h3a5a79ab),
	.w5(32'hbab178a8),
	.w6(32'h38ce47ae),
	.w7(32'h3a319a86),
	.w8(32'hba36457b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48f335),
	.w1(32'h3a81d0f7),
	.w2(32'hba099c3a),
	.w3(32'h3ac5f48c),
	.w4(32'h3a92a871),
	.w5(32'hba5f1d01),
	.w6(32'h3a919fc0),
	.w7(32'hbafd6201),
	.w8(32'hbb91e133),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6c37f),
	.w1(32'h3ad0715e),
	.w2(32'h3a8ffd84),
	.w3(32'h3afb2f1c),
	.w4(32'h3a15045c),
	.w5(32'hba2e3d14),
	.w6(32'h3bab6d83),
	.w7(32'h3af4549e),
	.w8(32'h3a3cda77),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0b809),
	.w1(32'h3b2defc9),
	.w2(32'h3825f0ea),
	.w3(32'hba078010),
	.w4(32'hba24ea6c),
	.w5(32'hbad322ed),
	.w6(32'hbbdfd06e),
	.w7(32'hbbee622f),
	.w8(32'hbc3002e1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb093ca6),
	.w1(32'hba903c85),
	.w2(32'hbba1f2af),
	.w3(32'h3a149c56),
	.w4(32'h3a878ae3),
	.w5(32'hbabf8b0e),
	.w6(32'hbb473342),
	.w7(32'hbb3fee2f),
	.w8(32'hbbba318a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b3d8d),
	.w1(32'h3ab27848),
	.w2(32'hba642bff),
	.w3(32'h3a07beb7),
	.w4(32'hb7f56143),
	.w5(32'hbaaa0d00),
	.w6(32'hbb9e7dcf),
	.w7(32'hbb8207f1),
	.w8(32'hbbed54ce),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386fad17),
	.w1(32'hb993e690),
	.w2(32'hb997f41c),
	.w3(32'h39dd4d15),
	.w4(32'hb7b1c21c),
	.w5(32'h3707c480),
	.w6(32'hb9720f1b),
	.w7(32'h37a55602),
	.w8(32'hb9c808c1),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb885d7e),
	.w1(32'hbb665095),
	.w2(32'hba8238c5),
	.w3(32'hba5a8185),
	.w4(32'hbaaffed1),
	.w5(32'hb9897cdd),
	.w6(32'hba492c41),
	.w7(32'hbadef77d),
	.w8(32'hbb1bbdcb),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb936421d),
	.w1(32'hb9b2e767),
	.w2(32'hb9b9c221),
	.w3(32'hb9603436),
	.w4(32'hb9c6e93a),
	.w5(32'hb9ce0e84),
	.w6(32'hb95bd11a),
	.w7(32'hb99c67b1),
	.w8(32'hb9317c73),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b96f18),
	.w1(32'h39f0e898),
	.w2(32'h374fb38a),
	.w3(32'h39baa9e9),
	.w4(32'h39d9cc86),
	.w5(32'h38860eaf),
	.w6(32'hba39acc4),
	.w7(32'hbaa4f033),
	.w8(32'hbae3aec0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e8da4),
	.w1(32'h3656c070),
	.w2(32'h398e090f),
	.w3(32'hb9c877b8),
	.w4(32'h374c5b73),
	.w5(32'h38a1c181),
	.w6(32'hb8819f3a),
	.w7(32'hba2a0a13),
	.w8(32'hba0f47ca),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb062ae4),
	.w1(32'h386ddb92),
	.w2(32'hbb0c4bbe),
	.w3(32'h399c5339),
	.w4(32'h3ae57122),
	.w5(32'h38ea198f),
	.w6(32'hba57609d),
	.w7(32'hba19fd3e),
	.w8(32'hbb8a14d4),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d611e2),
	.w1(32'h39521e7e),
	.w2(32'h3a339264),
	.w3(32'h393b99fd),
	.w4(32'h39bb51b3),
	.w5(32'h3a560fbe),
	.w6(32'h39758e1e),
	.w7(32'h3a5e74bb),
	.w8(32'h39f70e83),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d074b7),
	.w1(32'hb9b2b704),
	.w2(32'hb96b83ec),
	.w3(32'h39a21aeb),
	.w4(32'hb98b959f),
	.w5(32'hb95be61f),
	.w6(32'hb9793c87),
	.w7(32'h36d8c282),
	.w8(32'hb91512cb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09ab24),
	.w1(32'h39eb9aa2),
	.w2(32'h3a25ddb7),
	.w3(32'h3a3e3443),
	.w4(32'hb9275bae),
	.w5(32'hb9b43ef1),
	.w6(32'h3a19cde5),
	.w7(32'hbab95e1a),
	.w8(32'hbb0f5b0f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a8a66),
	.w1(32'hb9023fb8),
	.w2(32'hbafedea4),
	.w3(32'hba80205e),
	.w4(32'h39f08780),
	.w5(32'hbb399983),
	.w6(32'hbb14034e),
	.w7(32'hbb2249ca),
	.w8(32'hbbbbcacd),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20706c),
	.w1(32'hbb411b33),
	.w2(32'hbbd2c0d5),
	.w3(32'h3a9f47c3),
	.w4(32'hbaab3021),
	.w5(32'hbab534d7),
	.w6(32'hbb4686aa),
	.w7(32'h3a81ae1b),
	.w8(32'hba3ce1fa),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90927e8),
	.w1(32'h3a17570b),
	.w2(32'h39cf0299),
	.w3(32'hb861c5bd),
	.w4(32'h3a32ccc7),
	.w5(32'h39f398dc),
	.w6(32'hba109638),
	.w7(32'hb9455bba),
	.w8(32'h37a17953),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9f8f6),
	.w1(32'hb9558e60),
	.w2(32'hbba8c77c),
	.w3(32'h39b16b77),
	.w4(32'hbb0c8f6e),
	.w5(32'hbbe43040),
	.w6(32'hbc318f82),
	.w7(32'hbc0dddc0),
	.w8(32'hbc6663d9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0ac83),
	.w1(32'hbb1d4550),
	.w2(32'h3a5cf86c),
	.w3(32'h3bde2b93),
	.w4(32'h3afea8d5),
	.w5(32'h3a2f358e),
	.w6(32'h3bded384),
	.w7(32'hbaf0b59d),
	.w8(32'hbbd8ac2c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5b00d),
	.w1(32'hbab8115d),
	.w2(32'hbad1544b),
	.w3(32'h3a846207),
	.w4(32'hb9b4a635),
	.w5(32'hbb02309f),
	.w6(32'hba6ad9f0),
	.w7(32'hba97976f),
	.w8(32'hba897ee1),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f656e6),
	.w1(32'hba07cfdf),
	.w2(32'h3968786b),
	.w3(32'hb9933f65),
	.w4(32'hb99df726),
	.w5(32'hb8f613bf),
	.w6(32'hb9cc2945),
	.w7(32'hb8ee58af),
	.w8(32'hb8fb5c8d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d0b44),
	.w1(32'h3a040e3e),
	.w2(32'h39920127),
	.w3(32'h38dade9b),
	.w4(32'h39fa9bd6),
	.w5(32'h39ea2aaa),
	.w6(32'h3a2411a7),
	.w7(32'h39fd885e),
	.w8(32'h3a2ab4ee),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea3173),
	.w1(32'hb9bc8052),
	.w2(32'hb8be1a5b),
	.w3(32'h39ff963e),
	.w4(32'hb9ca60e3),
	.w5(32'hb8d131f2),
	.w6(32'hb98f3027),
	.w7(32'hb9159280),
	.w8(32'hb8b8e165),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc34fd),
	.w1(32'h3af77bb6),
	.w2(32'hba9ed290),
	.w3(32'h3ae1c39b),
	.w4(32'h3a258d8b),
	.w5(32'hbacf0efd),
	.w6(32'hba4aed21),
	.w7(32'h3a78776e),
	.w8(32'hb9a3f508),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914abff),
	.w1(32'h3a900285),
	.w2(32'h3a2ae188),
	.w3(32'hb9ada3cc),
	.w4(32'h3a6ba660),
	.w5(32'hbaa0b2c2),
	.w6(32'hbba79a17),
	.w7(32'hbb53726e),
	.w8(32'hbb7e4b04),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa375a),
	.w1(32'h3b004394),
	.w2(32'hbb1a07c5),
	.w3(32'h39a021c9),
	.w4(32'h3b2ecde9),
	.w5(32'hb7680dfe),
	.w6(32'hbac2e4cc),
	.w7(32'hbb64a89c),
	.w8(32'hbba8778b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80f8ec),
	.w1(32'h3ac111f9),
	.w2(32'h3a9a0dc2),
	.w3(32'hba01fd39),
	.w4(32'h38fa7490),
	.w5(32'hb8f728d8),
	.w6(32'hb9fc7e35),
	.w7(32'hb9dedb22),
	.w8(32'hba7346e2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a1cf2),
	.w1(32'h3b624c8c),
	.w2(32'hba17ea4e),
	.w3(32'h3b84fe6b),
	.w4(32'h3b2700b5),
	.w5(32'hbaab0ba8),
	.w6(32'hbbace2a4),
	.w7(32'hbb9a4cc6),
	.w8(32'hbbed15ba),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0238e7),
	.w1(32'h3af2f966),
	.w2(32'hba809db4),
	.w3(32'h3aa9b169),
	.w4(32'h39afcc88),
	.w5(32'hbb0b2392),
	.w6(32'hbb042ce4),
	.w7(32'hbac74457),
	.w8(32'hbae92c1a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998ad0e),
	.w1(32'hb894c00a),
	.w2(32'hb89a62ad),
	.w3(32'h3993a6cc),
	.w4(32'hb8d0b5c8),
	.w5(32'hb8ce86f1),
	.w6(32'h381d33e1),
	.w7(32'hb807a35f),
	.w8(32'h38b70112),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e56dc),
	.w1(32'hbb3dc8d0),
	.w2(32'hbb31e459),
	.w3(32'h3a1f60a7),
	.w4(32'hb9dc3976),
	.w5(32'hbb1120bd),
	.w6(32'h3a198a08),
	.w7(32'h3acd1310),
	.w8(32'h3ac51d5c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3810a091),
	.w1(32'hb980c07d),
	.w2(32'hb92d5ec7),
	.w3(32'h36d044b2),
	.w4(32'hb95ba112),
	.w5(32'hb918e5c8),
	.w6(32'h3810f381),
	.w7(32'hb92bd364),
	.w8(32'h38619f56),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf46b76),
	.w1(32'h3bb5c9d7),
	.w2(32'hbac6e73a),
	.w3(32'h3bd0fdfe),
	.w4(32'h3b866a0a),
	.w5(32'hbb54b887),
	.w6(32'hba137f1c),
	.w7(32'hbacb80e1),
	.w8(32'hbbdcf6e6),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b193f3),
	.w1(32'h3b545693),
	.w2(32'hb9721b21),
	.w3(32'hbb14d363),
	.w4(32'h3b23b900),
	.w5(32'hba9facde),
	.w6(32'hbb9191c6),
	.w7(32'hbb1c9fac),
	.w8(32'hbbcbbc38),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e5d33),
	.w1(32'h3ae1235d),
	.w2(32'hba51fb3c),
	.w3(32'hb8add038),
	.w4(32'h3a329510),
	.w5(32'hbab9d9ec),
	.w6(32'hbb58fafc),
	.w7(32'hbb76af02),
	.w8(32'hbbc0bb87),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917a859),
	.w1(32'h3a3dfd19),
	.w2(32'hba4cf2bd),
	.w3(32'hb86d76de),
	.w4(32'h39f3a1ca),
	.w5(32'hba8f89f2),
	.w6(32'hb9cad3e5),
	.w7(32'h38b450c9),
	.w8(32'hba821cde),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b264a83),
	.w1(32'h38ba1903),
	.w2(32'hb9a2bf74),
	.w3(32'h3b345c2f),
	.w4(32'h3b061acd),
	.w5(32'hb9dfffb8),
	.w6(32'h3a984c7a),
	.w7(32'hbb07514d),
	.w8(32'hbbc8cf6a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f35150),
	.w1(32'hb81d2607),
	.w2(32'hbb09f5a0),
	.w3(32'h390a1329),
	.w4(32'h39233e36),
	.w5(32'hba4580b6),
	.w6(32'hbb33ddae),
	.w7(32'hbb2c0895),
	.w8(32'hbb1e4bd1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babf568),
	.w1(32'h3b6d1158),
	.w2(32'hbae7c0a0),
	.w3(32'h3b35202c),
	.w4(32'h3ae8e0d1),
	.w5(32'hbae7fe91),
	.w6(32'hbbac57c7),
	.w7(32'hbbe2dec7),
	.w8(32'hbc18d2d3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa5a0f),
	.w1(32'h393ee315),
	.w2(32'hb8f4ae00),
	.w3(32'hb995a4e4),
	.w4(32'h390ea699),
	.w5(32'h390ca5f1),
	.w6(32'h39581ab8),
	.w7(32'hb8321431),
	.w8(32'h388b6431),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bc7598),
	.w1(32'h37f2ac25),
	.w2(32'hb90a89f9),
	.w3(32'h3919167f),
	.w4(32'hb9a34a30),
	.w5(32'hba225b66),
	.w6(32'h38fbcb31),
	.w7(32'hb80397b0),
	.w8(32'hb9822990),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb25a9e),
	.w1(32'h3bc65d1b),
	.w2(32'h3ab4dce0),
	.w3(32'h3a6c97a3),
	.w4(32'h3b610b0c),
	.w5(32'hbab7d8a5),
	.w6(32'hbc3bfadb),
	.w7(32'hbc03ac6a),
	.w8(32'hbc03a4b7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71c75e),
	.w1(32'h3b1ece4f),
	.w2(32'hbafc168f),
	.w3(32'h3a615217),
	.w4(32'h3a5bc6b6),
	.w5(32'hbb9e5108),
	.w6(32'hbc26b293),
	.w7(32'hbbec5842),
	.w8(32'hbc322768),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1b356),
	.w1(32'h3b063a3c),
	.w2(32'h3a0b4aa3),
	.w3(32'hba4b2ba5),
	.w4(32'h3b113ac3),
	.w5(32'hb9844dea),
	.w6(32'hbba2c646),
	.w7(32'hbb9c4161),
	.w8(32'hbbce00f9),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54c21b),
	.w1(32'hbb0e8989),
	.w2(32'hbabf1efc),
	.w3(32'h3bb50d3a),
	.w4(32'hba99e555),
	.w5(32'h3b070edc),
	.w6(32'h3b56e8f8),
	.w7(32'h3a31d5ee),
	.w8(32'hba461e00),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ea7a0f),
	.w1(32'hba0a7ee2),
	.w2(32'hba517867),
	.w3(32'h397efd07),
	.w4(32'hb9072a1d),
	.w5(32'hb9f95718),
	.w6(32'hba70e3eb),
	.w7(32'hba01d0f6),
	.w8(32'hb9550eba),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba262561),
	.w1(32'hba9c67c9),
	.w2(32'hbaa9e83c),
	.w3(32'h3987f362),
	.w4(32'h39ac4471),
	.w5(32'hb98711a5),
	.w6(32'hb988fca4),
	.w7(32'h39aaa3b6),
	.w8(32'h388ecd0a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25fbed),
	.w1(32'h3b89bede),
	.w2(32'hbbd3c275),
	.w3(32'hba92672f),
	.w4(32'h3a848d1e),
	.w5(32'hbb8e1057),
	.w6(32'hbc202c6e),
	.w7(32'h3a5691bc),
	.w8(32'hbb2b77b8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b77a4),
	.w1(32'h3b1346e0),
	.w2(32'hbac9c1be),
	.w3(32'h3a1ebac8),
	.w4(32'hbaa282f0),
	.w5(32'hbb4e936b),
	.w6(32'hbbe152d5),
	.w7(32'hbba9273d),
	.w8(32'hbc03bcd3),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ada80),
	.w1(32'h39ff936b),
	.w2(32'hbab228bc),
	.w3(32'h3ac298df),
	.w4(32'h3b5d5792),
	.w5(32'h371ec6b4),
	.w6(32'hbbfd3741),
	.w7(32'h3a063193),
	.w8(32'hbb28fd5c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba727eb),
	.w1(32'h3b54a482),
	.w2(32'h3837e3d4),
	.w3(32'h3a8fe56d),
	.w4(32'h3a5faa0f),
	.w5(32'hb9e973fc),
	.w6(32'hba1b29bf),
	.w7(32'hbb39377c),
	.w8(32'hbb8608db),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba686ca6),
	.w1(32'hbb28b036),
	.w2(32'hbb9adbf0),
	.w3(32'hbad72745),
	.w4(32'hba096c38),
	.w5(32'hbb277e4d),
	.w6(32'hbae4adad),
	.w7(32'hbb9f4f42),
	.w8(32'hbbf68e80),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a306b),
	.w1(32'hb8b445c9),
	.w2(32'hb989cb7a),
	.w3(32'hb9a22004),
	.w4(32'hb9063327),
	.w5(32'hb97f959b),
	.w6(32'hb96de02d),
	.w7(32'hb9a2a84f),
	.w8(32'hb930fb2d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946786c),
	.w1(32'h38dc702d),
	.w2(32'h397e83a4),
	.w3(32'hb9655c50),
	.w4(32'h398861ec),
	.w5(32'h397e5307),
	.w6(32'h39fa19ba),
	.w7(32'h3a728935),
	.w8(32'h3a1fa1db),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93fd31),
	.w1(32'h3ac3fa2f),
	.w2(32'h3a7e12bd),
	.w3(32'h3a1ee612),
	.w4(32'hba259170),
	.w5(32'hbaa95cd3),
	.w6(32'h3a8379a6),
	.w7(32'h39bd0299),
	.w8(32'hba0c1017),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcb009),
	.w1(32'hb8ad25ed),
	.w2(32'hb9c9a5b4),
	.w3(32'hb9f6f15e),
	.w4(32'h3927ee31),
	.w5(32'hb95b651f),
	.w6(32'h3815d60c),
	.w7(32'hb961541b),
	.w8(32'hb848aa9d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b819f),
	.w1(32'h3a54b31a),
	.w2(32'hbb084677),
	.w3(32'h3adeebc0),
	.w4(32'h3a618bff),
	.w5(32'hbaa39baf),
	.w6(32'hb88ec4b4),
	.w7(32'hba16ac94),
	.w8(32'hba1b797d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb031fb0),
	.w1(32'hbacce037),
	.w2(32'hbb0e55f2),
	.w3(32'hbace6adc),
	.w4(32'hbaa00618),
	.w5(32'hbb38ef26),
	.w6(32'hbc01bd95),
	.w7(32'hbbb506dc),
	.w8(32'hbbd33910),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e9e12),
	.w1(32'h3b1cfd21),
	.w2(32'h3a9b2147),
	.w3(32'h3a262da9),
	.w4(32'h3a60f847),
	.w5(32'hba20b520),
	.w6(32'hbb28c902),
	.w7(32'hbb0bf625),
	.w8(32'hbb7f916b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d74a7),
	.w1(32'h3a27822d),
	.w2(32'h3a3520cb),
	.w3(32'h397912cf),
	.w4(32'h3a47bab8),
	.w5(32'h3a40f1f6),
	.w6(32'h399cbef5),
	.w7(32'h3a42a604),
	.w8(32'h3ab45485),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39957467),
	.w1(32'h39d0d21b),
	.w2(32'hbb739f32),
	.w3(32'h3a866c52),
	.w4(32'h3a84606b),
	.w5(32'hbb0298d8),
	.w6(32'hbc1fa794),
	.w7(32'hbacf438b),
	.w8(32'hbb55c823),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b0ce5),
	.w1(32'h3a98e728),
	.w2(32'hba02adce),
	.w3(32'h3a904d51),
	.w4(32'h39a37ab2),
	.w5(32'hba30aba4),
	.w6(32'hbb20a8e5),
	.w7(32'hba86554f),
	.w8(32'hbb1fa8b1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2f361),
	.w1(32'hba00d343),
	.w2(32'hb97d87f8),
	.w3(32'hb91c188f),
	.w4(32'hba139439),
	.w5(32'hb99592f0),
	.w6(32'hb9750469),
	.w7(32'hb9447ae4),
	.w8(32'h37c39fd8),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4da4f3),
	.w1(32'h3a8ca98d),
	.w2(32'hb93fe4ba),
	.w3(32'h3af0265a),
	.w4(32'h3a1cba22),
	.w5(32'h390b30ba),
	.w6(32'hbb1dbbef),
	.w7(32'hbb001690),
	.w8(32'hbb2e797f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8649141),
	.w1(32'hb92045d9),
	.w2(32'hb996663b),
	.w3(32'hb8eab111),
	.w4(32'hb962e150),
	.w5(32'hb95bc212),
	.w6(32'hb943b70f),
	.w7(32'hb9caea24),
	.w8(32'hb985f056),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e15ea5),
	.w1(32'hb99fb06d),
	.w2(32'hb9ef590c),
	.w3(32'hb8e320fd),
	.w4(32'hb9648dc0),
	.w5(32'hb9c9409e),
	.w6(32'hba4d150e),
	.w7(32'hba57155a),
	.w8(32'hba16e812),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9916a52),
	.w1(32'hb9744613),
	.w2(32'hb97aa6fb),
	.w3(32'hb956b235),
	.w4(32'hb989f39c),
	.w5(32'hb99537f5),
	.w6(32'hb9527e30),
	.w7(32'hb9658b09),
	.w8(32'hb840e6ab),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb852bdef),
	.w1(32'h37b716b8),
	.w2(32'h399cf11f),
	.w3(32'hb8a83417),
	.w4(32'hb66ea8e6),
	.w5(32'h3986df26),
	.w6(32'h37fa061c),
	.w7(32'h39090d81),
	.w8(32'h38e1e881),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8df211),
	.w1(32'h3a357480),
	.w2(32'hb9a96688),
	.w3(32'hba78d0ed),
	.w4(32'hba6952f4),
	.w5(32'hba73a11d),
	.w6(32'hbaae78f8),
	.w7(32'hbb126603),
	.w8(32'hbb18f21e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89a1fc),
	.w1(32'hbb626ab7),
	.w2(32'hbb665be5),
	.w3(32'h3aa26065),
	.w4(32'hba56ccde),
	.w5(32'hba1b5676),
	.w6(32'hbb4ba06d),
	.w7(32'hbb97a2d8),
	.w8(32'hbc06c15e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a9dc91),
	.w1(32'h39a02fdb),
	.w2(32'hbadcebf2),
	.w3(32'h3a605b81),
	.w4(32'hba3078a0),
	.w5(32'hba93ac7e),
	.w6(32'hbb376216),
	.w7(32'hbb334c2e),
	.w8(32'hbb8430f8),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5cfb2),
	.w1(32'hb965805a),
	.w2(32'hbabf3765),
	.w3(32'h3b117797),
	.w4(32'hba143c82),
	.w5(32'h39ee3868),
	.w6(32'hbb2b4b76),
	.w7(32'hbb911604),
	.w8(32'hbbb1414d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f90b5),
	.w1(32'hba0c467b),
	.w2(32'hb99af8a8),
	.w3(32'hb964dd87),
	.w4(32'hb9feb4bd),
	.w5(32'hb9c7b9ef),
	.w6(32'hba1d4231),
	.w7(32'hb94f09d9),
	.w8(32'hb96b63ae),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e72ebd),
	.w1(32'hba046d0a),
	.w2(32'hb9cdd8db),
	.w3(32'hb9459d08),
	.w4(32'hba0549f3),
	.w5(32'hba0127fe),
	.w6(32'hb8d0fab2),
	.w7(32'h3954c5f8),
	.w8(32'h38e283f7),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9411e),
	.w1(32'hb921a0e5),
	.w2(32'hb935d253),
	.w3(32'hb8fd8fc6),
	.w4(32'hb93b66d8),
	.w5(32'hb980b9c6),
	.w6(32'hb895c18c),
	.w7(32'hb8c97605),
	.w8(32'hb5bc5c5d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3611ef19),
	.w1(32'hb91039f4),
	.w2(32'hb918e5cf),
	.w3(32'hb8820fc7),
	.w4(32'hb9319a36),
	.w5(32'hb9645e8a),
	.w6(32'hb7d0cf4c),
	.w7(32'hb895b252),
	.w8(32'h380f401c),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb425150),
	.w1(32'hbb2493b1),
	.w2(32'hbaa73bfa),
	.w3(32'h3a154360),
	.w4(32'h39e03207),
	.w5(32'hbac77b47),
	.w6(32'hbb5fb031),
	.w7(32'hbb0f385a),
	.w8(32'hbb9f9573),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8843b1d),
	.w1(32'hb95f2f8e),
	.w2(32'hb8ad1821),
	.w3(32'h392120b1),
	.w4(32'hb94a0ed4),
	.w5(32'h38627dab),
	.w6(32'hb99a50db),
	.w7(32'hb826a047),
	.w8(32'hb86be8e0),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c61e04),
	.w1(32'h3a8a2c60),
	.w2(32'hba275e6f),
	.w3(32'hb9f53f7a),
	.w4(32'h39e7a775),
	.w5(32'hba81052d),
	.w6(32'hb984785c),
	.w7(32'h39fd09fd),
	.w8(32'hba5e407f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f68c9e),
	.w1(32'hba311e3b),
	.w2(32'hba7aa4ce),
	.w3(32'hb982a367),
	.w4(32'hb8cbd544),
	.w5(32'hbacaf6ef),
	.w6(32'h3a9e51bc),
	.w7(32'h39128072),
	.w8(32'hba39a947),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76ae1e5),
	.w1(32'hb98100d9),
	.w2(32'hb9815ce1),
	.w3(32'hb828aa78),
	.w4(32'hb990d16f),
	.w5(32'hb9b146b8),
	.w6(32'hb9321e8e),
	.w7(32'hb987edb8),
	.w8(32'hb9292114),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeba5f6),
	.w1(32'h3aa2a12f),
	.w2(32'h39119fbd),
	.w3(32'h3ace943a),
	.w4(32'h3aa8e651),
	.w5(32'hb90821fa),
	.w6(32'hba74c8cf),
	.w7(32'hba8fe0e2),
	.w8(32'hbadfbfdb),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8236f16),
	.w1(32'hb9363f2d),
	.w2(32'hb98d8fdb),
	.w3(32'h39d328f6),
	.w4(32'h39e61944),
	.w5(32'h38809099),
	.w6(32'h39be6001),
	.w7(32'h3a098903),
	.w8(32'h39b30c2e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb70688),
	.w1(32'hbb8f7e4e),
	.w2(32'hbb02206b),
	.w3(32'h3b223c59),
	.w4(32'h3b5113af),
	.w5(32'h3af08cd4),
	.w6(32'h3a46e008),
	.w7(32'h3a794b8a),
	.w8(32'hbb981843),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9506aec),
	.w1(32'h38e2b4e8),
	.w2(32'hb8557e9c),
	.w3(32'hb919ad44),
	.w4(32'h38f10f99),
	.w5(32'hb95fb88d),
	.w6(32'h399db05d),
	.w7(32'h3869ce39),
	.w8(32'h36e13f29),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83a070),
	.w1(32'h3bd01e0c),
	.w2(32'h3b8d6a4e),
	.w3(32'hbb5d8965),
	.w4(32'hba63137c),
	.w5(32'hbb20fa5a),
	.w6(32'hbc027379),
	.w7(32'hbbbbef1e),
	.w8(32'hbba6774a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule