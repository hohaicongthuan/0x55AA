module layer_10_featuremap_284(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d483b),
	.w1(32'hbb29c3ce),
	.w2(32'hba61d298),
	.w3(32'hbb10df8e),
	.w4(32'hbb4e2f93),
	.w5(32'h3ac7fb3a),
	.w6(32'hbb1cf33c),
	.w7(32'h390a4497),
	.w8(32'h3ab47b32),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b4ee2),
	.w1(32'h3b8c2374),
	.w2(32'h3b95b85b),
	.w3(32'h3a5fc2f2),
	.w4(32'h3ba7efc2),
	.w5(32'hb9c50273),
	.w6(32'h3b64b60d),
	.w7(32'h3bb4bdc7),
	.w8(32'hba2878cd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55b1b9),
	.w1(32'hbb62b407),
	.w2(32'hbb8c386f),
	.w3(32'hbb01a32b),
	.w4(32'hbb639c68),
	.w5(32'h3aaa9118),
	.w6(32'hbbd88f7c),
	.w7(32'hbbc09485),
	.w8(32'h3a0b7f33),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac91db1),
	.w1(32'h3aef5f27),
	.w2(32'h3ab53b68),
	.w3(32'h3ac057b5),
	.w4(32'h3a2eb499),
	.w5(32'hb89f8fe5),
	.w6(32'h3afc6934),
	.w7(32'h39034cfb),
	.w8(32'h3bb64f5d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2f4b5),
	.w1(32'h399db91e),
	.w2(32'hbb01fe90),
	.w3(32'h39b36940),
	.w4(32'hbb5dbc10),
	.w5(32'hbb402288),
	.w6(32'h3ad37948),
	.w7(32'h3b6648ba),
	.w8(32'hbb1936de),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53f277),
	.w1(32'hbabb7ae7),
	.w2(32'hb9fbc2bb),
	.w3(32'hbaefbd66),
	.w4(32'hbb01600b),
	.w5(32'hbae53484),
	.w6(32'hb9f50301),
	.w7(32'hba21225e),
	.w8(32'hbb36f0ba),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab33234),
	.w1(32'h3a8436d2),
	.w2(32'hba278056),
	.w3(32'h3ac9f397),
	.w4(32'h3a8fb254),
	.w5(32'hbac93521),
	.w6(32'h3aeb655c),
	.w7(32'h39eae564),
	.w8(32'hba7f547a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998475e),
	.w1(32'hbaeb6fab),
	.w2(32'h3749cd4d),
	.w3(32'hbb0e1770),
	.w4(32'hbaea17d3),
	.w5(32'hbb04a3b7),
	.w6(32'hb9d4851a),
	.w7(32'h394d216d),
	.w8(32'hba8f0deb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe5fed),
	.w1(32'h3934e0c4),
	.w2(32'h38f7b57b),
	.w3(32'hb91759d9),
	.w4(32'h3a3e1b93),
	.w5(32'hbb63b9ed),
	.w6(32'h3b0fc9a6),
	.w7(32'h3b068949),
	.w8(32'hbb59bbc8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67d801),
	.w1(32'hbaee19dd),
	.w2(32'hba962cf9),
	.w3(32'hbb4aac2a),
	.w4(32'hbb512c53),
	.w5(32'hbacdba8c),
	.w6(32'hbaee603f),
	.w7(32'hbb143ea1),
	.w8(32'hbab10c12),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb038309),
	.w1(32'hb9764de6),
	.w2(32'hba84063a),
	.w3(32'hb9d050dd),
	.w4(32'hbb33516a),
	.w5(32'hbb80afc7),
	.w6(32'hb9d7a7fa),
	.w7(32'hbb29c4d7),
	.w8(32'hbbfa7b93),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fb73b),
	.w1(32'hba52835c),
	.w2(32'hbb8b4588),
	.w3(32'hbac13765),
	.w4(32'hb9aeef87),
	.w5(32'h3bcc3220),
	.w6(32'hbbb18e8a),
	.w7(32'hbb935ebe),
	.w8(32'h3c3f4bdd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b0ba6),
	.w1(32'h3c016c85),
	.w2(32'h3bf5ce91),
	.w3(32'h3be2879b),
	.w4(32'h3ba5387d),
	.w5(32'h3b098402),
	.w6(32'h3c0438ee),
	.w7(32'h3c1d07de),
	.w8(32'hbb66bbe0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88947a1),
	.w1(32'h38e39675),
	.w2(32'h3bb6e5d2),
	.w3(32'h3b8bd4f3),
	.w4(32'h3bc88e13),
	.w5(32'h3a8190be),
	.w6(32'hbb414f52),
	.w7(32'h3c1cbb55),
	.w8(32'hbaf8f25d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd8c6),
	.w1(32'hbafbbccb),
	.w2(32'h3a7a4577),
	.w3(32'h3ab04d53),
	.w4(32'hb9a7f6f4),
	.w5(32'h3a191b82),
	.w6(32'h3b153745),
	.w7(32'h39f223c0),
	.w8(32'h39272c2e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae87204),
	.w1(32'hb9ed163d),
	.w2(32'hbb1450c9),
	.w3(32'hbaa9e5d9),
	.w4(32'hbb8ef777),
	.w5(32'hba20c464),
	.w6(32'h3b181e47),
	.w7(32'hbb29ea8a),
	.w8(32'hba8e761c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf8542),
	.w1(32'h397ba009),
	.w2(32'h3adf0ec2),
	.w3(32'hba88dee7),
	.w4(32'hba49f122),
	.w5(32'hb9640504),
	.w6(32'h3a845ccd),
	.w7(32'h3b687df3),
	.w8(32'h3a9c8b8b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f7897),
	.w1(32'hba84a1de),
	.w2(32'hbaf3f896),
	.w3(32'h3ad4acdc),
	.w4(32'h3ad9b9af),
	.w5(32'hb9521e02),
	.w6(32'hba8d2884),
	.w7(32'hbac902b8),
	.w8(32'hba2878d9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c7ffd),
	.w1(32'h3a36f21d),
	.w2(32'h3a3144a9),
	.w3(32'hb8fa26dc),
	.w4(32'hbb67e241),
	.w5(32'hba124010),
	.w6(32'h3b6ab790),
	.w7(32'hba89a479),
	.w8(32'hbbab229a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3f489),
	.w1(32'hbbf586e8),
	.w2(32'hbb11341e),
	.w3(32'h3aa5ad8b),
	.w4(32'h3bb062ce),
	.w5(32'h3b0bb407),
	.w6(32'hbc01182c),
	.w7(32'h38c71863),
	.w8(32'h3ba7d930),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fc86c),
	.w1(32'h3b19bd82),
	.w2(32'hbb6a08d1),
	.w3(32'hba19d5ed),
	.w4(32'hbbb81c9c),
	.w5(32'hbb296ec1),
	.w6(32'h3b97cd5f),
	.w7(32'hbb8dc14e),
	.w8(32'hbb631c0b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad83c9d),
	.w1(32'hbb801635),
	.w2(32'hbb133434),
	.w3(32'hbb817dc0),
	.w4(32'hbb2ca362),
	.w5(32'h3c0167c0),
	.w6(32'hbb990e93),
	.w7(32'hbb7db39c),
	.w8(32'h3b8cd887),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91d290),
	.w1(32'hba342b90),
	.w2(32'hba2d49d6),
	.w3(32'h3b7eb03b),
	.w4(32'hbac320a1),
	.w5(32'h3ba4708b),
	.w6(32'hbad44894),
	.w7(32'hbb477f48),
	.w8(32'h3b8924be),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8ee42),
	.w1(32'h3a82d776),
	.w2(32'hb9b9f30c),
	.w3(32'h3b82a290),
	.w4(32'hbb56ef52),
	.w5(32'hbb15858e),
	.w6(32'h3badcfc4),
	.w7(32'hbb2231ae),
	.w8(32'hbbc7c315),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb695f70),
	.w1(32'hbb88d616),
	.w2(32'hbb0bc1d9),
	.w3(32'hbae34dbc),
	.w4(32'hbb1157ea),
	.w5(32'h38a88a14),
	.w6(32'hbbdb4c54),
	.w7(32'hbbb97b12),
	.w8(32'hbafd9c3c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b19d3),
	.w1(32'hbb273807),
	.w2(32'h39bacf94),
	.w3(32'hba506588),
	.w4(32'hbadeb2a6),
	.w5(32'hb9afaa42),
	.w6(32'hba22d9a4),
	.w7(32'hba085d36),
	.w8(32'hba5d1e8e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c75b9),
	.w1(32'h39eff7bf),
	.w2(32'hb9937db0),
	.w3(32'hba94df0f),
	.w4(32'hbacd2478),
	.w5(32'hbb0bbb9c),
	.w6(32'hb983ad37),
	.w7(32'hba7aaea1),
	.w8(32'h39214118),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c3005),
	.w1(32'hba94fdac),
	.w2(32'h39faed92),
	.w3(32'hbaa38d3d),
	.w4(32'hba4e3d1d),
	.w5(32'h3a12b614),
	.w6(32'h39b10dbd),
	.w7(32'h3b412471),
	.w8(32'hbb8ff445),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e967f),
	.w1(32'hbb8c207c),
	.w2(32'h3abedde0),
	.w3(32'h3b025a4c),
	.w4(32'h3b4930b1),
	.w5(32'h3a2b2b58),
	.w6(32'hbb9a2bd8),
	.w7(32'h3b6dbf89),
	.w8(32'hba8fcfdd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51d70b),
	.w1(32'hba7e6919),
	.w2(32'h3b9e364e),
	.w3(32'h3ac26d86),
	.w4(32'h3b73bcea),
	.w5(32'h38e00ac9),
	.w6(32'hbb8dbf48),
	.w7(32'h3b279f28),
	.w8(32'h3ac5e568),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef6f8e),
	.w1(32'h3b8413f5),
	.w2(32'h3b3f5c8b),
	.w3(32'h3b48e9eb),
	.w4(32'h3b24a877),
	.w5(32'h3acc4485),
	.w6(32'h3bef2c43),
	.w7(32'h3bc6655a),
	.w8(32'h3970e318),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae38ed),
	.w1(32'h3b7ca644),
	.w2(32'h3a129538),
	.w3(32'h3b3f6050),
	.w4(32'h3b9e9da7),
	.w5(32'hbb7930eb),
	.w6(32'hbb22dfcd),
	.w7(32'h3aecea41),
	.w8(32'hbb80d15c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc4691),
	.w1(32'h3aba815f),
	.w2(32'h3a9746aa),
	.w3(32'hbb25b682),
	.w4(32'h3a3d5587),
	.w5(32'h3ad3c7a1),
	.w6(32'hba9569d1),
	.w7(32'hb951ea40),
	.w8(32'h3b8a4af0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391bd1d6),
	.w1(32'h390b128f),
	.w2(32'hb9f36e83),
	.w3(32'h3a9e0745),
	.w4(32'h3affc766),
	.w5(32'h3b25f8b4),
	.w6(32'h3ad27c4c),
	.w7(32'h3a401f59),
	.w8(32'h3bca4128),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42a755),
	.w1(32'h3c117dc1),
	.w2(32'h3b98df05),
	.w3(32'hbab25d50),
	.w4(32'h39b581c0),
	.w5(32'h3b3ea005),
	.w6(32'hbb1f501d),
	.w7(32'hbb650107),
	.w8(32'h3b8b8576),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cdc61),
	.w1(32'hbb52f206),
	.w2(32'hbb87dd11),
	.w3(32'h3b424da0),
	.w4(32'h3a59562b),
	.w5(32'hbb229605),
	.w6(32'h3b918669),
	.w7(32'hbac7dbcb),
	.w8(32'hbb2e6f01),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba155fc5),
	.w1(32'h3b13acfd),
	.w2(32'hba5923bc),
	.w3(32'hbb0c883e),
	.w4(32'hba00e139),
	.w5(32'hba2a0e49),
	.w6(32'h3b14f49a),
	.w7(32'h3a93878d),
	.w8(32'h3a1c24f6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f8f2e),
	.w1(32'h3a6c5112),
	.w2(32'h3b4a26d8),
	.w3(32'h38dc1b4d),
	.w4(32'h3a886739),
	.w5(32'hbb42d2be),
	.w6(32'h3b3dfb79),
	.w7(32'h3b10f1ac),
	.w8(32'hbb0859f5),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16fbfc),
	.w1(32'hbb6303a5),
	.w2(32'hbb563f2f),
	.w3(32'hbab19fc3),
	.w4(32'hbafb0810),
	.w5(32'hbb9a6a13),
	.w6(32'hbb09add9),
	.w7(32'hbaa24887),
	.w8(32'hbbbb74b2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad80566),
	.w1(32'hbb4c3b5e),
	.w2(32'hbaeb866b),
	.w3(32'hbb02fd1f),
	.w4(32'hba820ca0),
	.w5(32'hbbe7e5e4),
	.w6(32'hba152c42),
	.w7(32'hbb8a1e49),
	.w8(32'hbc1ca8b6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2d78e),
	.w1(32'hbbcbc842),
	.w2(32'hbb80bf9f),
	.w3(32'hbc06b7b1),
	.w4(32'hbb9fd865),
	.w5(32'hba9ec86b),
	.w6(32'hbc3a1c29),
	.w7(32'hbbd8b6b2),
	.w8(32'hbb14aae8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95eab3),
	.w1(32'hba179505),
	.w2(32'h3975ccb7),
	.w3(32'hbad5b92b),
	.w4(32'hba812c8a),
	.w5(32'h3b26a4ac),
	.w6(32'hbabaad22),
	.w7(32'hbb1bcf38),
	.w8(32'hba5480f6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b0ef6),
	.w1(32'h3b43722e),
	.w2(32'h3aa25516),
	.w3(32'h3bcf6754),
	.w4(32'h3afb43e5),
	.w5(32'h3b1f50ed),
	.w6(32'h3b8c7d87),
	.w7(32'hba9e9e58),
	.w8(32'h3bc0ddfe),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1c960),
	.w1(32'h3c0d9980),
	.w2(32'h3ac90483),
	.w3(32'h3be36f5f),
	.w4(32'h3b59d753),
	.w5(32'hba24639d),
	.w6(32'h3c17487e),
	.w7(32'h3bba4bbc),
	.w8(32'h3908e5c1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2082c),
	.w1(32'h3b20ac05),
	.w2(32'hb9a41939),
	.w3(32'h3a594ce3),
	.w4(32'hba0bf591),
	.w5(32'h3aeeeb51),
	.w6(32'h3b4d0095),
	.w7(32'hbad52bf7),
	.w8(32'h3b09ff94),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a951f70),
	.w1(32'hba8b4c9e),
	.w2(32'hbadd0e2a),
	.w3(32'hbad34d2b),
	.w4(32'hb9ae81e7),
	.w5(32'hb90bfe14),
	.w6(32'h3ac34511),
	.w7(32'h3a5e506d),
	.w8(32'hb737bc69),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8035c),
	.w1(32'h3b49d21b),
	.w2(32'h3a105a7a),
	.w3(32'hba9f9a6b),
	.w4(32'hba63e59c),
	.w5(32'hbb30baed),
	.w6(32'h3b29e478),
	.w7(32'h39e6f835),
	.w8(32'hbafb5476),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8eb50f),
	.w1(32'hba78ab6b),
	.w2(32'hba38e18d),
	.w3(32'hbb0d3a9c),
	.w4(32'hbb35d92b),
	.w5(32'h3b2ff18d),
	.w6(32'hba11cc96),
	.w7(32'hbac4c966),
	.w8(32'h3c01d76b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7d6cc),
	.w1(32'h3bced324),
	.w2(32'h3b9a01ba),
	.w3(32'h3b9c9aeb),
	.w4(32'h3b8760ad),
	.w5(32'hbb817c51),
	.w6(32'h3bf6f988),
	.w7(32'h3bc79aa3),
	.w8(32'hbba46aaa),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67b23c),
	.w1(32'hbb933121),
	.w2(32'hbb5d8902),
	.w3(32'hbb98c3ac),
	.w4(32'hbb863e9d),
	.w5(32'hbc2d5648),
	.w6(32'hbbc0b723),
	.w7(32'hbba1abad),
	.w8(32'hbc112513),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc32c6d),
	.w1(32'hbb05c2aa),
	.w2(32'h3bf2b6be),
	.w3(32'hbbcb430c),
	.w4(32'h3bdc8760),
	.w5(32'hbab82a48),
	.w6(32'hbbd7c941),
	.w7(32'h3bc1375f),
	.w8(32'hba2f8a21),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c72ca0),
	.w1(32'h398a22a6),
	.w2(32'hbad507c1),
	.w3(32'h39a3927a),
	.w4(32'h3b2cc4d5),
	.w5(32'h39d08864),
	.w6(32'h3838c698),
	.w7(32'hb9104ac5),
	.w8(32'hbb9006c1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32132b),
	.w1(32'h3a05c338),
	.w2(32'h3ba75460),
	.w3(32'h3964e4a8),
	.w4(32'h3ac8ce46),
	.w5(32'h3a7943f2),
	.w6(32'hbc108ae3),
	.w7(32'hba9b5137),
	.w8(32'hbadccfa7),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe02c4),
	.w1(32'hbafb9a7e),
	.w2(32'h3b92b672),
	.w3(32'h3a8d1a36),
	.w4(32'h3b5d0442),
	.w5(32'hbbd7a793),
	.w6(32'hbb939534),
	.w7(32'h3b721df6),
	.w8(32'hbc115d33),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cd0ce),
	.w1(32'hbc0ac33e),
	.w2(32'hbbe217dd),
	.w3(32'hbbe1c225),
	.w4(32'hbb8ca5aa),
	.w5(32'hb88eef94),
	.w6(32'hbc33950b),
	.w7(32'hbc024d91),
	.w8(32'h3a2efeb6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b552856),
	.w1(32'h3b3c05ee),
	.w2(32'h36b82b34),
	.w3(32'hbb23c1c6),
	.w4(32'h3b047079),
	.w5(32'hbb0e5e67),
	.w6(32'hbbbe303c),
	.w7(32'hbb751726),
	.w8(32'hbb50541c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafbfe3),
	.w1(32'hba4eaa39),
	.w2(32'hbab86272),
	.w3(32'hbad09f54),
	.w4(32'h38f4f3a4),
	.w5(32'h3b11d0c1),
	.w6(32'hbaf681cf),
	.w7(32'hbb0e7342),
	.w8(32'h3a046958),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47036a),
	.w1(32'hbaf78bfe),
	.w2(32'h3ac7ccde),
	.w3(32'hb8dcaf59),
	.w4(32'hba8a824b),
	.w5(32'hbb4d8759),
	.w6(32'hbb30438b),
	.w7(32'h3af79c13),
	.w8(32'hbbab0fef),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34a087),
	.w1(32'hbb47d572),
	.w2(32'hbb143f43),
	.w3(32'hbb4f2b5f),
	.w4(32'hbb359af1),
	.w5(32'hbb038bc1),
	.w6(32'hbba33b07),
	.w7(32'hbb86ce1e),
	.w8(32'h39bde10b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dc7dbf),
	.w1(32'hba9bcf42),
	.w2(32'hba679f56),
	.w3(32'h394d2592),
	.w4(32'hba994949),
	.w5(32'h3a450782),
	.w6(32'h3a86e711),
	.w7(32'hba6c7cbb),
	.w8(32'hb859db6f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fbb38),
	.w1(32'hbabf8417),
	.w2(32'h391671f7),
	.w3(32'hba2fd0e0),
	.w4(32'hbab1a952),
	.w5(32'h3a8e46e7),
	.w6(32'hba9115a4),
	.w7(32'hb994342d),
	.w8(32'h3b05650b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc1409),
	.w1(32'hba3ca05f),
	.w2(32'hba281ad8),
	.w3(32'hba9d925a),
	.w4(32'hbacd20a4),
	.w5(32'hba0b8665),
	.w6(32'h3abd3a85),
	.w7(32'hb9930a1c),
	.w8(32'h3b8bef25),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f8775),
	.w1(32'h3c37ec45),
	.w2(32'h3bf0aee5),
	.w3(32'hbb0e2d82),
	.w4(32'hb9cebf9f),
	.w5(32'hbb746530),
	.w6(32'hbb4712a2),
	.w7(32'h398d5c3c),
	.w8(32'hbb4704af),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb081b6e),
	.w1(32'hbb2cc630),
	.w2(32'hbb4a788f),
	.w3(32'hbbe60cf9),
	.w4(32'hbae06581),
	.w5(32'h3b83414e),
	.w6(32'hbbf59c82),
	.w7(32'hbb4733f4),
	.w8(32'h3bef8bad),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d3d45),
	.w1(32'h3ba38d35),
	.w2(32'h3bcab15f),
	.w3(32'hba4afa34),
	.w4(32'h3bb2fe4a),
	.w5(32'hbbac0bf4),
	.w6(32'hbba5da00),
	.w7(32'h386be87f),
	.w8(32'hbc07764f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c5dde),
	.w1(32'hba84c267),
	.w2(32'hba9321ff),
	.w3(32'hbb95cb00),
	.w4(32'hbb480a33),
	.w5(32'hb993abb1),
	.w6(32'hbc274115),
	.w7(32'hbbc517c1),
	.w8(32'hbab7245c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bc4d0),
	.w1(32'hbb437dc2),
	.w2(32'hbb2c0739),
	.w3(32'hb9de33fb),
	.w4(32'hbae9501e),
	.w5(32'hbb1575a2),
	.w6(32'hbb03a5bf),
	.w7(32'hbad88224),
	.w8(32'h39bced50),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eeecb4),
	.w1(32'h3ad5ee84),
	.w2(32'hbb2d75ad),
	.w3(32'h39b52dbd),
	.w4(32'hbaad25ad),
	.w5(32'hbba1b715),
	.w6(32'h3bcca40e),
	.w7(32'h3b1e6d98),
	.w8(32'hbbb9b3c4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe1d7c),
	.w1(32'hbbce3d52),
	.w2(32'hbb488cab),
	.w3(32'hbbee5a62),
	.w4(32'hbabf1c1f),
	.w5(32'h3bf6c6df),
	.w6(32'hbc0f8148),
	.w7(32'hbbb4beed),
	.w8(32'h3c0c638b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c10ba),
	.w1(32'h3c1400ba),
	.w2(32'h3bbc404e),
	.w3(32'h3bda9e3f),
	.w4(32'h3bc7eeb3),
	.w5(32'h3b0727b2),
	.w6(32'h3c736be5),
	.w7(32'h3c0d0952),
	.w8(32'hb9a657ad),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f930f0),
	.w1(32'h3a28c0f1),
	.w2(32'hba34f59e),
	.w3(32'h3a81ded9),
	.w4(32'hbb35d93a),
	.w5(32'hba06c956),
	.w6(32'h3b95b54b),
	.w7(32'hba935fac),
	.w8(32'h3aad756b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3aa226),
	.w1(32'h3ad5846d),
	.w2(32'hbb44462a),
	.w3(32'hba511742),
	.w4(32'hb9e4a721),
	.w5(32'hba924bd3),
	.w6(32'h3b26073f),
	.w7(32'h39ee7672),
	.w8(32'h3a5d7994),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7da67),
	.w1(32'hbae821a8),
	.w2(32'hb9c2594e),
	.w3(32'hb8e1dde6),
	.w4(32'h3a99f42b),
	.w5(32'h3a32b065),
	.w6(32'h3b176a71),
	.w7(32'h3b1788c0),
	.w8(32'h3b20c9f0),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcffc6),
	.w1(32'h3aaafac5),
	.w2(32'h3b5497d1),
	.w3(32'h3a7d74cf),
	.w4(32'h3b9408a3),
	.w5(32'hba81420c),
	.w6(32'h39fa4640),
	.w7(32'h3b86d343),
	.w8(32'hbaf67646),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33c9c2),
	.w1(32'hba65be1c),
	.w2(32'hbb0d4e9e),
	.w3(32'hbb02e5db),
	.w4(32'hbbc88a8b),
	.w5(32'h3b94bf99),
	.w6(32'hba218da9),
	.w7(32'hbb5a2d95),
	.w8(32'h3beada1c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2caf0b),
	.w1(32'h3b2569ca),
	.w2(32'h3b05fb33),
	.w3(32'h3b927648),
	.w4(32'h3ba25977),
	.w5(32'hbb1d2371),
	.w6(32'h3b938f65),
	.w7(32'h3b77ce74),
	.w8(32'hbbba5f92),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb987ef7),
	.w1(32'hbb6957f9),
	.w2(32'hbaf6c6e2),
	.w3(32'hbb741adf),
	.w4(32'hbbb75520),
	.w5(32'hbb31dd82),
	.w6(32'hbc035aa2),
	.w7(32'hbbc9c3c7),
	.w8(32'hbb8054a5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9372ce),
	.w1(32'hbb5fc521),
	.w2(32'hbb7b6b6b),
	.w3(32'hba9dd28a),
	.w4(32'hba69879e),
	.w5(32'h3ae3910e),
	.w6(32'hba879216),
	.w7(32'hbb0e8e9b),
	.w8(32'h3a3465b2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2438d2),
	.w1(32'h3b1ea524),
	.w2(32'h3b855742),
	.w3(32'h3ad335fa),
	.w4(32'h3b3af0a9),
	.w5(32'h3a0df535),
	.w6(32'h3b9dd8d4),
	.w7(32'h3b79c588),
	.w8(32'h3afb257d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5148a3),
	.w1(32'h3a119b49),
	.w2(32'h3a0613fa),
	.w3(32'hb9b53756),
	.w4(32'h39d592ed),
	.w5(32'h3b428441),
	.w6(32'h3b83482d),
	.w7(32'h3b8b6c59),
	.w8(32'h39bf0621),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04441a),
	.w1(32'h3b454b75),
	.w2(32'h3b414839),
	.w3(32'h3afaab8c),
	.w4(32'h3b0b5053),
	.w5(32'h39a515f7),
	.w6(32'h3a89e496),
	.w7(32'hb8879e27),
	.w8(32'h3b13c555),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ed091),
	.w1(32'h3a60a6ad),
	.w2(32'h3a45fc28),
	.w3(32'h3b2aacdd),
	.w4(32'h3b42aa42),
	.w5(32'h3b9f122b),
	.w6(32'h3b3cf782),
	.w7(32'h3b132348),
	.w8(32'h3b9a621d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39faaf25),
	.w1(32'hbaa9e6ad),
	.w2(32'h3b3688d9),
	.w3(32'h3a25eab3),
	.w4(32'h3ac5dc95),
	.w5(32'h3be11f2b),
	.w6(32'hbbdcd449),
	.w7(32'h3a315569),
	.w8(32'h3bcf7bbb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c045bb1),
	.w1(32'h3b56ef71),
	.w2(32'h3b87a332),
	.w3(32'h3b8f5122),
	.w4(32'h3a858958),
	.w5(32'h3c129d7b),
	.w6(32'h3ba1f70b),
	.w7(32'hba02cd13),
	.w8(32'h3becb989),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a623c),
	.w1(32'hbb4aab00),
	.w2(32'h3a8fcce6),
	.w3(32'h3b857e73),
	.w4(32'h3abde1ef),
	.w5(32'h3a029842),
	.w6(32'hbb28c874),
	.w7(32'h3a00f9d0),
	.w8(32'h3b3314de),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b5943),
	.w1(32'h39447269),
	.w2(32'hba9dbaba),
	.w3(32'hba885efc),
	.w4(32'hbb3177a6),
	.w5(32'hbb205437),
	.w6(32'h38817997),
	.w7(32'hb92c6b35),
	.w8(32'hbba17d48),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ba834),
	.w1(32'hbbb1334d),
	.w2(32'h3ae46b04),
	.w3(32'hbab1d6a4),
	.w4(32'h3ae6f8cd),
	.w5(32'h37b178a1),
	.w6(32'hbbab6e27),
	.w7(32'h3b171aa8),
	.w8(32'hbaf043f5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca1af1),
	.w1(32'hbb1fe656),
	.w2(32'hb8eb6626),
	.w3(32'h3ad1fdb4),
	.w4(32'h3af1a963),
	.w5(32'h3a22535f),
	.w6(32'hbb3242d5),
	.w7(32'h3b5a8d47),
	.w8(32'h3a0b084c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f13063),
	.w1(32'h3afe1563),
	.w2(32'h3b1fb43b),
	.w3(32'h3af2434c),
	.w4(32'h3ae686bf),
	.w5(32'hbb31f4d7),
	.w6(32'h3b860640),
	.w7(32'h3b3fa925),
	.w8(32'hbbc9112c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b4c03),
	.w1(32'hbb6efef8),
	.w2(32'hba920bee),
	.w3(32'hbb3a9723),
	.w4(32'hbb2be7ff),
	.w5(32'h3acebe8f),
	.w6(32'hbb86ca9c),
	.w7(32'h39038039),
	.w8(32'h3b55a4f3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ba74c),
	.w1(32'h3ae29c4e),
	.w2(32'h3b20ef91),
	.w3(32'h3b1fd152),
	.w4(32'h3b3eb596),
	.w5(32'h3b8c50a6),
	.w6(32'h3ba5d433),
	.w7(32'h3b75881a),
	.w8(32'h3be11237),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b8371),
	.w1(32'h3a88e022),
	.w2(32'h39f9a4a2),
	.w3(32'h3b7ca0a7),
	.w4(32'h3b3ed89d),
	.w5(32'h3b613c1b),
	.w6(32'hba98ed45),
	.w7(32'hb915ec5b),
	.w8(32'h3b8e1093),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa127e0),
	.w1(32'h3bc0b54c),
	.w2(32'hba004b8b),
	.w3(32'h3bc3fedd),
	.w4(32'h3ba642a7),
	.w5(32'hba550e32),
	.w6(32'hbaadda49),
	.w7(32'hb8e4a79c),
	.w8(32'h3a0ab873),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d994a),
	.w1(32'hbb424dc0),
	.w2(32'hbb511925),
	.w3(32'hbb70e059),
	.w4(32'hbb845268),
	.w5(32'hba8a0aac),
	.w6(32'hbad93855),
	.w7(32'hbae7e2ef),
	.w8(32'hbaf0bacc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02a4f3),
	.w1(32'hbac5cfbe),
	.w2(32'hb939f741),
	.w3(32'hbab85282),
	.w4(32'hbb0e2bb1),
	.w5(32'h3b02f4f3),
	.w6(32'hb99f4b0e),
	.w7(32'hba93bfb8),
	.w8(32'h3b195691),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba9039),
	.w1(32'h3bb39c56),
	.w2(32'h3b2f328c),
	.w3(32'h3b7520a7),
	.w4(32'h3aa782a2),
	.w5(32'hba8e0c4a),
	.w6(32'h3b886483),
	.w7(32'h3afd21a0),
	.w8(32'hba8a02ad),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b084ed7),
	.w1(32'h3a45a8c7),
	.w2(32'h3b33a88c),
	.w3(32'h38a1ba6d),
	.w4(32'h3bb99a35),
	.w5(32'hbb7aaf7d),
	.w6(32'h3b1e5032),
	.w7(32'h3b28db9c),
	.w8(32'hbb6bd0b5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e0f82),
	.w1(32'h3b11d1b1),
	.w2(32'h3a7e4bfd),
	.w3(32'hba1903fd),
	.w4(32'hba31599f),
	.w5(32'h3ad8857b),
	.w6(32'hbb6f69d5),
	.w7(32'hba9957f8),
	.w8(32'h3a9d4200),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b24ce5),
	.w1(32'hb9ce39bf),
	.w2(32'h3aaac668),
	.w3(32'h3b0c99aa),
	.w4(32'h3b5a5115),
	.w5(32'hbba83e0b),
	.w6(32'h3a73d82e),
	.w7(32'h3b67a0d6),
	.w8(32'hbbab71cb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a949e61),
	.w1(32'h3a5fe47c),
	.w2(32'h3ac041f7),
	.w3(32'hbbe87818),
	.w4(32'hbb11ed97),
	.w5(32'hbb5c338b),
	.w6(32'h38ec3b02),
	.w7(32'hbab5d713),
	.w8(32'h3a275ce4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f4c03),
	.w1(32'h3bcda409),
	.w2(32'h3b97a9be),
	.w3(32'hbb9258e4),
	.w4(32'hbb7230fc),
	.w5(32'hbb020ba1),
	.w6(32'hbb55e4e3),
	.w7(32'h3a9cd2f2),
	.w8(32'h3c408b18),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb0143),
	.w1(32'h3acebd20),
	.w2(32'h383a79f3),
	.w3(32'h3bd289c2),
	.w4(32'h3c0af10b),
	.w5(32'hba85883c),
	.w6(32'h3c319b07),
	.w7(32'h3c7531e4),
	.w8(32'hbb8669fe),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d1f28),
	.w1(32'hbb890477),
	.w2(32'hbac094d8),
	.w3(32'hbba82545),
	.w4(32'hba0d435d),
	.w5(32'hbb82540f),
	.w6(32'hbae0d06a),
	.w7(32'hb823675f),
	.w8(32'hba8e5fbd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ee4a2),
	.w1(32'h3b6122b9),
	.w2(32'h3ab99de5),
	.w3(32'hbbacdd85),
	.w4(32'hbb90047a),
	.w5(32'h3a0663d4),
	.w6(32'hbb049505),
	.w7(32'hbb77283a),
	.w8(32'hbadbc920),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e92754),
	.w1(32'hbab34ecd),
	.w2(32'hba187259),
	.w3(32'h3a2f0bae),
	.w4(32'h3b234ac4),
	.w5(32'hba7a42a4),
	.w6(32'h3b9b12ef),
	.w7(32'hbb4377b1),
	.w8(32'hbaf70a36),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6858e2),
	.w1(32'h3b3350de),
	.w2(32'h3ab959da),
	.w3(32'hbaed1cac),
	.w4(32'hbadb7f81),
	.w5(32'hbb3c496d),
	.w6(32'hbaf39609),
	.w7(32'h395d0f0a),
	.w8(32'h3aa90e7c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b130364),
	.w1(32'hbab19a27),
	.w2(32'hbb43a6a6),
	.w3(32'hbb9eeddb),
	.w4(32'h3ba0ae66),
	.w5(32'hbac6e968),
	.w6(32'h3c15fb09),
	.w7(32'h3c10cecb),
	.w8(32'hb9937d71),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988a263),
	.w1(32'h3b667c8f),
	.w2(32'h3b51a5b0),
	.w3(32'hba5dd7c0),
	.w4(32'h3b60e354),
	.w5(32'h3b393efb),
	.w6(32'hbaaeaba1),
	.w7(32'h3b07e64e),
	.w8(32'h3aee6e4a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98f2d6),
	.w1(32'hba777245),
	.w2(32'h3b14db63),
	.w3(32'h3b231ee5),
	.w4(32'h3b0d322d),
	.w5(32'hba248d65),
	.w6(32'h3747969e),
	.w7(32'h3b8b9ffb),
	.w8(32'hbb2830cd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb924682),
	.w1(32'hbb902199),
	.w2(32'hbbd19df9),
	.w3(32'hbaa66d6b),
	.w4(32'hba8a78c3),
	.w5(32'hbb57a38c),
	.w6(32'hbaf9743a),
	.w7(32'hbb2870b0),
	.w8(32'hba84607a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b002d81),
	.w1(32'hba5470a9),
	.w2(32'h3b0e92b5),
	.w3(32'hbbd9cb3c),
	.w4(32'hb8832353),
	.w5(32'hbb327a83),
	.w6(32'h385bb1c8),
	.w7(32'h3b5a3bdb),
	.w8(32'hbc25b011),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4999ae),
	.w1(32'h3b313770),
	.w2(32'hbb4d1471),
	.w3(32'h3b5f11ad),
	.w4(32'h3bd9e0a5),
	.w5(32'hbae1d4a1),
	.w6(32'h3b9d6209),
	.w7(32'hbb49812d),
	.w8(32'hb9aafaf7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a133549),
	.w1(32'h39135ab2),
	.w2(32'h3ab2b4c6),
	.w3(32'hbb3e5035),
	.w4(32'h3b05b5f3),
	.w5(32'h3b173549),
	.w6(32'h399ef9e5),
	.w7(32'h3b912c45),
	.w8(32'h3a8605bf),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f8fb1),
	.w1(32'hba8e85ee),
	.w2(32'h3b4489c8),
	.w3(32'h3b69d649),
	.w4(32'hba470c4a),
	.w5(32'h3b652457),
	.w6(32'h3b0b4491),
	.w7(32'h3b3e342c),
	.w8(32'h3a7c082a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b4360),
	.w1(32'hba39d17d),
	.w2(32'hbb0c0c4a),
	.w3(32'h3ac31af8),
	.w4(32'hbb0e34fa),
	.w5(32'hbb08941c),
	.w6(32'hbb906ef9),
	.w7(32'hbb33f79d),
	.w8(32'hbafc99ec),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca1fe5),
	.w1(32'h3b4d19f9),
	.w2(32'hba20c134),
	.w3(32'h3bbeb43e),
	.w4(32'h3c5b709b),
	.w5(32'hbb244bb9),
	.w6(32'h3bf546dc),
	.w7(32'h3c0ecc8d),
	.w8(32'hba0a01a4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6cae8),
	.w1(32'h3adb698f),
	.w2(32'h3b8f9935),
	.w3(32'hbb6b9024),
	.w4(32'hbb8a76fe),
	.w5(32'hbb063bb7),
	.w6(32'hbad129e6),
	.w7(32'hbb083cd7),
	.w8(32'hba8b24df),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f3301),
	.w1(32'hbaa9a756),
	.w2(32'h3abc28ff),
	.w3(32'hbba05a8a),
	.w4(32'hbb4f55ad),
	.w5(32'h3ae1b9eb),
	.w6(32'hbac7c050),
	.w7(32'hbbd3403d),
	.w8(32'hbb8caf28),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84a3710),
	.w1(32'hbad7963b),
	.w2(32'h37c53db1),
	.w3(32'hba97c9ce),
	.w4(32'h3b51afa7),
	.w5(32'hbb18546a),
	.w6(32'hbb6fddb1),
	.w7(32'hbac4ddf4),
	.w8(32'h3b90d8fc),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b2e3d),
	.w1(32'h3b1e24ed),
	.w2(32'h3b91dfd1),
	.w3(32'hbb96736f),
	.w4(32'hbb4caee9),
	.w5(32'hbad1c6f4),
	.w6(32'hbaf95982),
	.w7(32'h3b11bea6),
	.w8(32'hbb768bf2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eaf2c),
	.w1(32'h3bd7986a),
	.w2(32'h3bc6e711),
	.w3(32'hbac31058),
	.w4(32'h3816779d),
	.w5(32'hbac743a9),
	.w6(32'h38850931),
	.w7(32'h3b1c04f6),
	.w8(32'h3aa25dc6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3967c9c9),
	.w1(32'hb9bd3036),
	.w2(32'hbad14ddf),
	.w3(32'hb9dbf162),
	.w4(32'hbb0bab1c),
	.w5(32'hbb45ee45),
	.w6(32'hb92d1c9a),
	.w7(32'hba89a2b7),
	.w8(32'hbbd0c2de),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb963d73),
	.w1(32'hbaf168aa),
	.w2(32'hbb9c0d5e),
	.w3(32'hbb6e4fed),
	.w4(32'hbbf019d9),
	.w5(32'h3b0dd11b),
	.w6(32'hbbccab7d),
	.w7(32'hbc1c1bdf),
	.w8(32'h3b7d0392),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a061999),
	.w1(32'hbabe2d13),
	.w2(32'hba060b41),
	.w3(32'h3b5c5908),
	.w4(32'h3945b9b8),
	.w5(32'h3a701409),
	.w6(32'h3a7462be),
	.w7(32'h3af670b2),
	.w8(32'hbb51c359),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba639ab),
	.w1(32'hbb9e2f40),
	.w2(32'hbb5a02e9),
	.w3(32'h3a823306),
	.w4(32'hbb55f2c2),
	.w5(32'hbb5df3ba),
	.w6(32'hbb75ff49),
	.w7(32'hbbfa6560),
	.w8(32'h3b590121),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb006b9),
	.w1(32'hbb115b7b),
	.w2(32'hbb658a4b),
	.w3(32'hbbe5ecc4),
	.w4(32'hbc2cb638),
	.w5(32'h3a4b8cf6),
	.w6(32'hb92df14b),
	.w7(32'hbb97ca00),
	.w8(32'h3b80015c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17cbe9),
	.w1(32'h397ed241),
	.w2(32'h39c2c794),
	.w3(32'h3a50fc9c),
	.w4(32'hb960a5e3),
	.w5(32'h3b77ee55),
	.w6(32'h3b86545a),
	.w7(32'h3b852667),
	.w8(32'hbaa5f61e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07ac7b),
	.w1(32'h39c77973),
	.w2(32'hb9c54df3),
	.w3(32'h3b8a5add),
	.w4(32'hb93dde5b),
	.w5(32'h3b395b2e),
	.w6(32'hba18a2d8),
	.w7(32'hb9b1c118),
	.w8(32'h398ecd97),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9c567),
	.w1(32'hbb85eb30),
	.w2(32'hbb49858a),
	.w3(32'h3b873f35),
	.w4(32'h3bbb29e9),
	.w5(32'hba4d2125),
	.w6(32'hbac39fe3),
	.w7(32'hba22fdbc),
	.w8(32'hba08a8c0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d6ac0),
	.w1(32'hb8e42e65),
	.w2(32'hbadc3755),
	.w3(32'h3afea634),
	.w4(32'hb91d6a83),
	.w5(32'hbb530fec),
	.w6(32'hb9662065),
	.w7(32'hbb13dbaa),
	.w8(32'h3b9e7c64),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bdab2),
	.w1(32'h3c9106b0),
	.w2(32'h3bdf16e6),
	.w3(32'hba7a09af),
	.w4(32'h3c14e3a7),
	.w5(32'hb97c63da),
	.w6(32'h3c47df27),
	.w7(32'h3c8d1ee8),
	.w8(32'hba44297a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c76ad),
	.w1(32'h3afb89a7),
	.w2(32'h3ade2c40),
	.w3(32'h395aca3b),
	.w4(32'h3a63b393),
	.w5(32'h3b9bfe59),
	.w6(32'h3afeca37),
	.w7(32'h3aa49b88),
	.w8(32'h3c7bbfae),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78eeba7),
	.w1(32'hbaecd140),
	.w2(32'hbb0f815c),
	.w3(32'h3a0e63cf),
	.w4(32'h3b11bb5e),
	.w5(32'h3907bcc3),
	.w6(32'h3c37aa7c),
	.w7(32'h3c202364),
	.w8(32'hba843cbf),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb544082),
	.w1(32'hbb226279),
	.w2(32'hbb220734),
	.w3(32'hb98282fa),
	.w4(32'h39b3b00d),
	.w5(32'hbb51df3d),
	.w6(32'h3a5aa56b),
	.w7(32'h396bc8c9),
	.w8(32'h3aad018a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac86e3d),
	.w1(32'hba651617),
	.w2(32'hba8a9d31),
	.w3(32'hba527ff7),
	.w4(32'h36c538ba),
	.w5(32'hba19676a),
	.w6(32'h3a64f1ee),
	.w7(32'h3a83d091),
	.w8(32'hbb276137),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc0180),
	.w1(32'h3ab10ae9),
	.w2(32'h3af8e387),
	.w3(32'h3aa74d73),
	.w4(32'h3b32171c),
	.w5(32'hbaa06d59),
	.w6(32'hba479d75),
	.w7(32'hb97cc4ce),
	.w8(32'h3996444a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1813e),
	.w1(32'hb9709bd7),
	.w2(32'h3a873644),
	.w3(32'hbb3f719d),
	.w4(32'hba9a3537),
	.w5(32'h3af3e70e),
	.w6(32'hb9f48bd6),
	.w7(32'h3ab17a75),
	.w8(32'h3898354a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb615ba7),
	.w1(32'hbb1768d7),
	.w2(32'hbb460cf9),
	.w3(32'h3ae6580c),
	.w4(32'h3b2e52b9),
	.w5(32'h3aca57a1),
	.w6(32'h3afb8efc),
	.w7(32'h3a82e124),
	.w8(32'hba032cad),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f03cdb),
	.w1(32'h3b2a5f5e),
	.w2(32'h3b33a1bd),
	.w3(32'h3b71117f),
	.w4(32'h3ba6e992),
	.w5(32'h3a997427),
	.w6(32'h3b5059ab),
	.w7(32'h3aafce30),
	.w8(32'hbb38cf9b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cecfed),
	.w1(32'h3b3336bf),
	.w2(32'h3a7334f9),
	.w3(32'h3af44281),
	.w4(32'hb8fd2c17),
	.w5(32'hba82a1dd),
	.w6(32'hbbc8df2f),
	.w7(32'h3b346f02),
	.w8(32'hbb8b9d63),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a209164),
	.w1(32'h3a924b01),
	.w2(32'hba31e1b2),
	.w3(32'h3b83aab2),
	.w4(32'h3abf692a),
	.w5(32'hbb89dcd8),
	.w6(32'hb94d2cc0),
	.w7(32'hbb87c390),
	.w8(32'hbb4157f6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39500547),
	.w1(32'hbba22c79),
	.w2(32'hbaff8241),
	.w3(32'hbbceff5c),
	.w4(32'hb9daa5a0),
	.w5(32'hbb5cf161),
	.w6(32'hbb345479),
	.w7(32'hbabd9323),
	.w8(32'hbb38372b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04f0d0),
	.w1(32'hbaf27c2c),
	.w2(32'h394064d3),
	.w3(32'hbb9c4e1a),
	.w4(32'hba43ad7e),
	.w5(32'hbb37b7c7),
	.w6(32'h39ed7f2a),
	.w7(32'h3b7a7137),
	.w8(32'hbbcaf760),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ee2f9),
	.w1(32'hbb29d45a),
	.w2(32'hb609601d),
	.w3(32'hba78c0ba),
	.w4(32'h38d02efd),
	.w5(32'hbb026854),
	.w6(32'hbabfc190),
	.w7(32'hb90dd0db),
	.w8(32'h3a90bb40),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ba09b),
	.w1(32'h3b444711),
	.w2(32'h3b0e140c),
	.w3(32'hbaf1758b),
	.w4(32'hbab3cd82),
	.w5(32'hba9ea574),
	.w6(32'h3b6ca555),
	.w7(32'h3b867daa),
	.w8(32'h3ac6e9fe),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba065534),
	.w1(32'h3ae1b003),
	.w2(32'h3ad7f16d),
	.w3(32'h3afaf3b6),
	.w4(32'h3a0732ae),
	.w5(32'hbb801d90),
	.w6(32'h3b2e1829),
	.w7(32'h39f5c6e9),
	.w8(32'hb910ab6d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9617f2e),
	.w1(32'hba05080d),
	.w2(32'h3b17e9c9),
	.w3(32'hbb8f31ba),
	.w4(32'hbb4c2ca5),
	.w5(32'h39e1e110),
	.w6(32'hbb313550),
	.w7(32'hbaed34aa),
	.w8(32'h3a5ab73b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997b53e),
	.w1(32'h3ac4f383),
	.w2(32'hbb445044),
	.w3(32'hbaa76f3d),
	.w4(32'hbb5f5b2b),
	.w5(32'hbb5878e5),
	.w6(32'hbaac739b),
	.w7(32'hbbd4905b),
	.w8(32'hb9c6668b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dbbb0),
	.w1(32'h3a9713cf),
	.w2(32'h3910dcf8),
	.w3(32'hbb69c286),
	.w4(32'hbb390833),
	.w5(32'hbb4008f3),
	.w6(32'hba11be0b),
	.w7(32'h3a463100),
	.w8(32'hbae6e799),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef046c),
	.w1(32'h3abb923b),
	.w2(32'h3b7c9047),
	.w3(32'hbb9c0d05),
	.w4(32'hbb8d6eac),
	.w5(32'hba8dd67e),
	.w6(32'hbb197571),
	.w7(32'hbb0dd9c6),
	.w8(32'hbb33a09c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb660fd8),
	.w1(32'hbbcc6caa),
	.w2(32'hbbcb6baf),
	.w3(32'hbb387788),
	.w4(32'h38eb205c),
	.w5(32'h392a8cde),
	.w6(32'h3a9ef29d),
	.w7(32'h3ab618fa),
	.w8(32'h3b65b8f2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ace75),
	.w1(32'h3b0cd7ce),
	.w2(32'h3a8a607a),
	.w3(32'h3bbff249),
	.w4(32'h3b9b5e66),
	.w5(32'h38d08570),
	.w6(32'h3bddcbbd),
	.w7(32'h3a92494e),
	.w8(32'h3c54609c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af97040),
	.w1(32'hbb0f607a),
	.w2(32'h3a4e29d8),
	.w3(32'hbb76cb8f),
	.w4(32'hbb8a2b9b),
	.w5(32'hbb2b3126),
	.w6(32'hbbb0e4ba),
	.w7(32'h3c2fe6d1),
	.w8(32'hba6855c3),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba183f77),
	.w1(32'h3a825712),
	.w2(32'h3afb5c8c),
	.w3(32'hbbc65af5),
	.w4(32'hbb52c180),
	.w5(32'hbaa385fa),
	.w6(32'hb8b5cc6d),
	.w7(32'h3b51dbad),
	.w8(32'h3ad46283),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17071f),
	.w1(32'h390def0c),
	.w2(32'hba077784),
	.w3(32'hbb53fc4d),
	.w4(32'hbb0cb691),
	.w5(32'hba40b73d),
	.w6(32'hbad9c440),
	.w7(32'h3b38bcbf),
	.w8(32'hba968265),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67a14f),
	.w1(32'hbbba9aa8),
	.w2(32'hbbb86a4b),
	.w3(32'hbb20cdf4),
	.w4(32'hbaf185cd),
	.w5(32'h3c02e0c8),
	.w6(32'hbb5a46a0),
	.w7(32'hbadefa23),
	.w8(32'h3c6a1512),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94ea21),
	.w1(32'h3b224436),
	.w2(32'h3b81b63d),
	.w3(32'h3bcf7a8e),
	.w4(32'h39ed7cea),
	.w5(32'hba9d1fcc),
	.w6(32'h3bb98777),
	.w7(32'hbb06215e),
	.w8(32'h3ab14053),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09fd0a),
	.w1(32'hba1b0e1a),
	.w2(32'hbb2fbf34),
	.w3(32'h3a1b584d),
	.w4(32'h39e317ca),
	.w5(32'hba27b6f4),
	.w6(32'hb9e612db),
	.w7(32'hb9e92d8f),
	.w8(32'h3afd80b7),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff3379),
	.w1(32'h3b98a1fb),
	.w2(32'h3c24be96),
	.w3(32'h3b8b0af8),
	.w4(32'hbbbc48a4),
	.w5(32'h3a9f5876),
	.w6(32'h3afd9191),
	.w7(32'h39381a52),
	.w8(32'h3b999cbb),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2433f),
	.w1(32'h3c11dc79),
	.w2(32'h3bac3b25),
	.w3(32'hbbbb8fe3),
	.w4(32'hbc11fb51),
	.w5(32'hbb84c607),
	.w6(32'h3b11886b),
	.w7(32'hba5948b6),
	.w8(32'hbacdabda),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14c888),
	.w1(32'hbb8c816d),
	.w2(32'hbb4c0899),
	.w3(32'h3b66f783),
	.w4(32'hba954f52),
	.w5(32'hbb847d4a),
	.w6(32'hbb3f5bed),
	.w7(32'hbbdb62a2),
	.w8(32'hba8fe1bd),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc84aa),
	.w1(32'hba494b4c),
	.w2(32'h39daa129),
	.w3(32'h39f77deb),
	.w4(32'h39c91604),
	.w5(32'h3a55bbae),
	.w6(32'h3a87b7f4),
	.w7(32'hb98a0d1c),
	.w8(32'h3b9a2ed3),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae59308),
	.w1(32'h3b5b3ea1),
	.w2(32'h3a1f66dd),
	.w3(32'hbb1d1ab9),
	.w4(32'hbc13e0f8),
	.w5(32'hba9fcdbb),
	.w6(32'h3b398f41),
	.w7(32'hbb3a3a43),
	.w8(32'h3b31c640),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad98c6),
	.w1(32'h3ad36092),
	.w2(32'h3b7fd16a),
	.w3(32'h3aa20e12),
	.w4(32'h3c288684),
	.w5(32'hb9a2a512),
	.w6(32'h3c093387),
	.w7(32'h3c17c0b1),
	.w8(32'hbb4cc195),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7372f4),
	.w1(32'hba581248),
	.w2(32'hbac88ef6),
	.w3(32'h3b22331e),
	.w4(32'hb956f450),
	.w5(32'h3b3f73ed),
	.w6(32'hbbba876f),
	.w7(32'hbbc2152b),
	.w8(32'hba910271),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0dfd2),
	.w1(32'h39b89d6b),
	.w2(32'h3b0e025d),
	.w3(32'h3b0654d0),
	.w4(32'h3b424ae2),
	.w5(32'h3bd68c7e),
	.w6(32'h3a0848e7),
	.w7(32'h3b930c62),
	.w8(32'hb97ede4b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e4eee),
	.w1(32'hbb40de23),
	.w2(32'hbb086b36),
	.w3(32'h3bb8cae9),
	.w4(32'h3c083985),
	.w5(32'h3a8d61a0),
	.w6(32'h3a2d2ab4),
	.w7(32'h3a91ec80),
	.w8(32'h39f628df),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b396d24),
	.w1(32'h3a5c1ab2),
	.w2(32'h3b7ae2d7),
	.w3(32'hbaa3b68e),
	.w4(32'h39c7374f),
	.w5(32'h3acd3ed3),
	.w6(32'hb816a5e9),
	.w7(32'hbb0d1d15),
	.w8(32'hb790bf7f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b676f09),
	.w1(32'h3b138cf9),
	.w2(32'hbb3c5436),
	.w3(32'h3ae40ca3),
	.w4(32'h3a974e3d),
	.w5(32'hbb11571c),
	.w6(32'hbb7f333a),
	.w7(32'hba9f0990),
	.w8(32'h3a07e29e),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3114a),
	.w1(32'h3b78adad),
	.w2(32'h3b284feb),
	.w3(32'hbafb365b),
	.w4(32'h391ec735),
	.w5(32'h3b3922a3),
	.w6(32'h3b1e0f08),
	.w7(32'h3bc34477),
	.w8(32'h3b46a53c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abee888),
	.w1(32'h3b4e97fb),
	.w2(32'h3bb593c2),
	.w3(32'hba49cbd0),
	.w4(32'hbb6ead7a),
	.w5(32'hb8f5523c),
	.w6(32'hbb233d5d),
	.w7(32'h3936ea32),
	.w8(32'h3b58f96f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7f013),
	.w1(32'h3a4d37ec),
	.w2(32'h39ed7f30),
	.w3(32'h3a35613b),
	.w4(32'hbb9e2887),
	.w5(32'hbb45aa32),
	.w6(32'h3bdf9b18),
	.w7(32'h3b195a60),
	.w8(32'h3b1214ed),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3734bc),
	.w1(32'h3b904c4e),
	.w2(32'h3b7fcf91),
	.w3(32'hbb7831a1),
	.w4(32'hbaad2790),
	.w5(32'hbb9f4af2),
	.w6(32'hba2d059f),
	.w7(32'hba9350a8),
	.w8(32'hbbb8cc76),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5b855),
	.w1(32'hba312ce9),
	.w2(32'hbac010dd),
	.w3(32'hbb85cd47),
	.w4(32'hbaf190c0),
	.w5(32'hbb55bb30),
	.w6(32'hbbb37746),
	.w7(32'hbb87fa89),
	.w8(32'hbb226a46),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9211ab),
	.w1(32'h3b210d46),
	.w2(32'hb9199caa),
	.w3(32'hbb3ab593),
	.w4(32'hb8732b14),
	.w5(32'hba70ee1c),
	.w6(32'hbb82b247),
	.w7(32'hbaaed62d),
	.w8(32'h3aa8b723),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba55ccd),
	.w1(32'h3ae46325),
	.w2(32'h3b87a6db),
	.w3(32'hbb5ed3f2),
	.w4(32'hbb89d437),
	.w5(32'h3b76f8e5),
	.w6(32'h38c4dc63),
	.w7(32'h3aa77345),
	.w8(32'h3b4308c4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a85fd),
	.w1(32'h3a1df033),
	.w2(32'hba9399fe),
	.w3(32'h3bf3748d),
	.w4(32'h3b96543e),
	.w5(32'hbb7940c4),
	.w6(32'h3b1927c3),
	.w7(32'h3a5267b3),
	.w8(32'hbb0b7a93),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdbc5e),
	.w1(32'h3aa98da1),
	.w2(32'h3b710f43),
	.w3(32'hbbcd3d4c),
	.w4(32'hbbae34e6),
	.w5(32'h3b43e910),
	.w6(32'hbb807eea),
	.w7(32'hba62f071),
	.w8(32'h3c13f0ad),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea8bf7),
	.w1(32'hbbfef7da),
	.w2(32'hbb8ac649),
	.w3(32'hbb2d2627),
	.w4(32'hb9c8d97c),
	.w5(32'h3a07bda3),
	.w6(32'h3b13c912),
	.w7(32'h3b7edeb9),
	.w8(32'h3b22ac0d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d8579),
	.w1(32'h3b16cfe6),
	.w2(32'h3b342058),
	.w3(32'h36dcc0c0),
	.w4(32'hb9dd3023),
	.w5(32'h3b61d664),
	.w6(32'hb9841462),
	.w7(32'hbb4ece1f),
	.w8(32'hbb83f5b9),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13a345),
	.w1(32'hbafe8ab6),
	.w2(32'h3bd72311),
	.w3(32'hba334968),
	.w4(32'hb69ca81b),
	.w5(32'hbbccc8ba),
	.w6(32'hbba2a51e),
	.w7(32'h3adc601e),
	.w8(32'h3a450c30),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12231c),
	.w1(32'hbb4dba96),
	.w2(32'hbba0d9b5),
	.w3(32'hbb98bd33),
	.w4(32'h39f6e551),
	.w5(32'h3b139c3c),
	.w6(32'hbb97eb2a),
	.w7(32'hba9db6c0),
	.w8(32'hbb8fda6c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9365498),
	.w1(32'h39cfa541),
	.w2(32'h37b4ef60),
	.w3(32'h3b9af33d),
	.w4(32'h3b2db8d1),
	.w5(32'h3ba95bf8),
	.w6(32'hbbba6197),
	.w7(32'hbbe31f54),
	.w8(32'h3c822f14),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92962e),
	.w1(32'h3c289020),
	.w2(32'h3bdcf033),
	.w3(32'h3ab29d58),
	.w4(32'hbbcc726d),
	.w5(32'h3ac1e981),
	.w6(32'h3c518a69),
	.w7(32'h3b989563),
	.w8(32'h3baa56bc),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cc9eb),
	.w1(32'h3b137e9d),
	.w2(32'h3ad31979),
	.w3(32'h3a309b09),
	.w4(32'hbb4a02b4),
	.w5(32'hbadb4724),
	.w6(32'h3b127ef7),
	.w7(32'hbb165c6e),
	.w8(32'hba9c0a73),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9b93c),
	.w1(32'h3ad45906),
	.w2(32'h39081eb8),
	.w3(32'hba962321),
	.w4(32'h3c2b7cb6),
	.w5(32'hbb522383),
	.w6(32'h3bfd5f0f),
	.w7(32'h3bc97642),
	.w8(32'hb99f77c3),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68c876),
	.w1(32'h3aa2c68b),
	.w2(32'h3b50eda0),
	.w3(32'hbbb58867),
	.w4(32'hbbcc9684),
	.w5(32'h3b5317c7),
	.w6(32'hbb4b5fdf),
	.w7(32'h3aadb959),
	.w8(32'h3b92e699),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0a18b),
	.w1(32'h3b70f08b),
	.w2(32'h3c1a9aa0),
	.w3(32'hba86c7a7),
	.w4(32'hbadbf54a),
	.w5(32'h3b41cf67),
	.w6(32'h3b0843a3),
	.w7(32'h3bde116c),
	.w8(32'h3970fe45),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f05a3),
	.w1(32'hbb143ad7),
	.w2(32'h39940cfd),
	.w3(32'h3abf0746),
	.w4(32'h3b9ce2ec),
	.w5(32'hbb5c5e12),
	.w6(32'hb987f45f),
	.w7(32'h39b19dd0),
	.w8(32'h39fceb19),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a62996),
	.w1(32'hb905bd43),
	.w2(32'h3a87501a),
	.w3(32'hbb9e5036),
	.w4(32'hbaba573f),
	.w5(32'hbb87224f),
	.w6(32'h3abb924f),
	.w7(32'h3b85a67b),
	.w8(32'h3c159e62),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f0e09),
	.w1(32'h3b6d3678),
	.w2(32'hba2dd6e5),
	.w3(32'hbbfb246d),
	.w4(32'hbc22e717),
	.w5(32'h3b16d868),
	.w6(32'h3bca5047),
	.w7(32'h3af2bef8),
	.w8(32'h3b38c324),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8d98e),
	.w1(32'hba384d83),
	.w2(32'hbbabbdc0),
	.w3(32'h3b3f82da),
	.w4(32'h3a608fea),
	.w5(32'hbb2b6eca),
	.w6(32'hba313b13),
	.w7(32'hbba3ec54),
	.w8(32'hba86ff49),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a9020),
	.w1(32'hbb2f1f7e),
	.w2(32'hbbe72a7e),
	.w3(32'hbb208cb1),
	.w4(32'hb9dbdb67),
	.w5(32'h3bef92f1),
	.w6(32'hbb664e2c),
	.w7(32'hbc10052d),
	.w8(32'hbc547a7b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af47c09),
	.w1(32'hba8779f9),
	.w2(32'h3b4097e2),
	.w3(32'h3c056bd7),
	.w4(32'h3b3681d5),
	.w5(32'hbad4f859),
	.w6(32'hbc417ce3),
	.w7(32'hbc33c1b5),
	.w8(32'hbaa5f6e8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9b38c),
	.w1(32'h3a7444b0),
	.w2(32'hb9afdcef),
	.w3(32'hbad0d2d9),
	.w4(32'h3b0ea69c),
	.w5(32'hb981033f),
	.w6(32'h3b2ed67e),
	.w7(32'h3b732395),
	.w8(32'hbb611ea2),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4c1b7),
	.w1(32'hbb11cc59),
	.w2(32'hbb5a9121),
	.w3(32'hb96119b6),
	.w4(32'h3aad3865),
	.w5(32'h3b2df133),
	.w6(32'h3b213cb7),
	.w7(32'h38937028),
	.w8(32'hb99a1fe4),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4315f),
	.w1(32'hbc1a99b9),
	.w2(32'hbbae4b9f),
	.w3(32'h3c402e38),
	.w4(32'h3c2d3380),
	.w5(32'hba16b20d),
	.w6(32'h3aacc60a),
	.w7(32'hbb34d205),
	.w8(32'hbae57a52),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b4fe1),
	.w1(32'h39e6a867),
	.w2(32'hba5702f0),
	.w3(32'hbae8a4d8),
	.w4(32'hbb8361f5),
	.w5(32'hbb0e248d),
	.w6(32'hbbc8b1fa),
	.w7(32'hba7a198b),
	.w8(32'h3a58b037),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c0041),
	.w1(32'h3b253db3),
	.w2(32'h3b4e77ff),
	.w3(32'hbb695046),
	.w4(32'hbb834755),
	.w5(32'hbb321f4e),
	.w6(32'hbac25e3a),
	.w7(32'h3a36ccbb),
	.w8(32'hba704226),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a7d39),
	.w1(32'h3b783c6d),
	.w2(32'hb8b94581),
	.w3(32'hbb751516),
	.w4(32'h39ece30b),
	.w5(32'h3b092bc3),
	.w6(32'h3ba03676),
	.w7(32'h3b217a14),
	.w8(32'h3c03ca87),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb163f1b),
	.w1(32'hbb0c9225),
	.w2(32'hbb55b3e4),
	.w3(32'h3a8c5843),
	.w4(32'h39ccc2bd),
	.w5(32'h3b030662),
	.w6(32'h3c1d30c1),
	.w7(32'h3bdd0e3a),
	.w8(32'h39f9fed2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1259e),
	.w1(32'h3a3f1deb),
	.w2(32'hbb03d5c8),
	.w3(32'hba93eb55),
	.w4(32'hb8f46242),
	.w5(32'hb88fe88e),
	.w6(32'hb9972432),
	.w7(32'hbba6b64f),
	.w8(32'hbb1a64d1),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1a52d),
	.w1(32'hbaa9bfd1),
	.w2(32'hba673c14),
	.w3(32'hba1ade0a),
	.w4(32'h3aab94d0),
	.w5(32'hbaa1ac22),
	.w6(32'hba16011e),
	.w7(32'h3aaed63f),
	.w8(32'h3ab32ec9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add2159),
	.w1(32'h3a4daa3b),
	.w2(32'hb910eeba),
	.w3(32'hba11c417),
	.w4(32'hbb2a0d6a),
	.w5(32'h3b7677e9),
	.w6(32'h3ab28e98),
	.w7(32'hbb3f63d3),
	.w8(32'hbbef8aaa),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea2f09),
	.w1(32'hbb492093),
	.w2(32'h3b2f5992),
	.w3(32'h39368aa4),
	.w4(32'hba9931ff),
	.w5(32'hbb414fa1),
	.w6(32'hbbf69748),
	.w7(32'hbab07c9d),
	.w8(32'h38ef6edf),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b6b44),
	.w1(32'h3a8fe97b),
	.w2(32'h3b425170),
	.w3(32'h3a390912),
	.w4(32'hb9c8b44f),
	.w5(32'hbb1d74e1),
	.w6(32'h3b115d86),
	.w7(32'h39d9ece4),
	.w8(32'hbb570322),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa499be),
	.w1(32'h38ee0594),
	.w2(32'hbade6b5b),
	.w3(32'hbb1bf351),
	.w4(32'h390445c4),
	.w5(32'hbad3b112),
	.w6(32'h3a02885e),
	.w7(32'hbabf6e37),
	.w8(32'h3aa51f7f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bd45b),
	.w1(32'hbb07f0d8),
	.w2(32'hbb0a3d4e),
	.w3(32'hbb13686c),
	.w4(32'h3990777d),
	.w5(32'hba040207),
	.w6(32'h3ba2da0f),
	.w7(32'h3b50a0eb),
	.w8(32'hb941f18a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba10e18),
	.w1(32'h3b1d1c06),
	.w2(32'h3a998959),
	.w3(32'hbae5ff13),
	.w4(32'hbb544e72),
	.w5(32'h3a677336),
	.w6(32'hba5d904d),
	.w7(32'hbb5d4481),
	.w8(32'hb7fd1141),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e7522),
	.w1(32'h3947a63b),
	.w2(32'hba47df28),
	.w3(32'h3a3170c6),
	.w4(32'hb98a644c),
	.w5(32'hbb82f9f9),
	.w6(32'hba98956a),
	.w7(32'hba912641),
	.w8(32'hbb37bc5d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989a657),
	.w1(32'h3b226589),
	.w2(32'hba85dbde),
	.w3(32'h3ba50b6b),
	.w4(32'h3c14dd3e),
	.w5(32'hbb00d2ca),
	.w6(32'h3c2fddcd),
	.w7(32'h3a3e6361),
	.w8(32'hbbc1728d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed5bcf),
	.w1(32'hbb1f38cf),
	.w2(32'hbbbeac31),
	.w3(32'hbac3f906),
	.w4(32'hbb5869b0),
	.w5(32'hbb884813),
	.w6(32'hbbc8eccd),
	.w7(32'hbbf09fe9),
	.w8(32'hbacb881a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b3b03),
	.w1(32'h3b03e122),
	.w2(32'hbb4e3263),
	.w3(32'hbae14e42),
	.w4(32'hb9d32c80),
	.w5(32'h3b618a34),
	.w6(32'h3b935a5c),
	.w7(32'h3a237d30),
	.w8(32'hba79126a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf04697),
	.w1(32'hbb164f4a),
	.w2(32'h3ad0c34d),
	.w3(32'h3b5dc76e),
	.w4(32'h3afff093),
	.w5(32'hbbc0b52e),
	.w6(32'h38fac56d),
	.w7(32'hb9775958),
	.w8(32'h3ad35428),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee911c),
	.w1(32'h3c4612aa),
	.w2(32'h39961ce5),
	.w3(32'hbb5b57c2),
	.w4(32'h3c005030),
	.w5(32'hbaa0a29b),
	.w6(32'h3c32f96a),
	.w7(32'h3c1af95f),
	.w8(32'hbb46f16a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba679137),
	.w1(32'hbaa857d4),
	.w2(32'h3a917e20),
	.w3(32'hba837761),
	.w4(32'hbb52dd9d),
	.w5(32'hbb82d3f0),
	.w6(32'hbac9d2cf),
	.w7(32'hbc19d8f9),
	.w8(32'hbaa9b861),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e73f5),
	.w1(32'h3a485bd8),
	.w2(32'h3aadb77a),
	.w3(32'hbb76ea1c),
	.w4(32'hbb09425d),
	.w5(32'h3b6a6fc5),
	.w6(32'h3b05e0d5),
	.w7(32'h3b197e31),
	.w8(32'h3b6c3874),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5868d2),
	.w1(32'h3b8e1d33),
	.w2(32'h3ab5e2b3),
	.w3(32'h39fd7eb2),
	.w4(32'h3a58466e),
	.w5(32'hba8dc3ba),
	.w6(32'hba8cf028),
	.w7(32'h3b42fc81),
	.w8(32'h3b4021f7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba130c55),
	.w1(32'h3b0921a7),
	.w2(32'hbaa08139),
	.w3(32'hbab93f4e),
	.w4(32'hba7d85bb),
	.w5(32'hbac5fbdc),
	.w6(32'hbb0275aa),
	.w7(32'hbb92de67),
	.w8(32'h3af4b800),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa422a8),
	.w1(32'h38de32e1),
	.w2(32'hba9ae9e8),
	.w3(32'hbbae521d),
	.w4(32'hba1de579),
	.w5(32'hbb01ba81),
	.w6(32'h3a10487e),
	.w7(32'h39c7a476),
	.w8(32'h3c1c400e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d6964),
	.w1(32'h3ab168a5),
	.w2(32'hbbd31d84),
	.w3(32'hbacf1bb0),
	.w4(32'hbba38df1),
	.w5(32'hbb2c89dd),
	.w6(32'h3b3ee753),
	.w7(32'h391ca56e),
	.w8(32'h3b90d7ba),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba621dcf),
	.w1(32'hbbe12842),
	.w2(32'hbb614d8f),
	.w3(32'hbb93e7a5),
	.w4(32'h3a2dc538),
	.w5(32'h3a677bbe),
	.w6(32'h3c21b374),
	.w7(32'h3bf342c0),
	.w8(32'hbaeb10c3),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a4d7e),
	.w1(32'hbb268876),
	.w2(32'hbb9aa31d),
	.w3(32'h3b926675),
	.w4(32'h3b3eaf55),
	.w5(32'h3b06f509),
	.w6(32'h3a786d09),
	.w7(32'h3b04a511),
	.w8(32'h3a0de644),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81a056),
	.w1(32'h3a8005b2),
	.w2(32'h3ae4d293),
	.w3(32'h3a0c1fcb),
	.w4(32'hba8b17fb),
	.w5(32'h3a0fd13c),
	.w6(32'h3ae14735),
	.w7(32'h3bd4a3bc),
	.w8(32'hbb77f705),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e902c),
	.w1(32'h39d21bbe),
	.w2(32'h3ac25071),
	.w3(32'hb9824bdc),
	.w4(32'hbb413c19),
	.w5(32'hbaf06fac),
	.w6(32'hbb4dbee3),
	.w7(32'hbb75ed05),
	.w8(32'h3aba36a8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be57624),
	.w1(32'h3b9c537b),
	.w2(32'h3c0c66d5),
	.w3(32'hbb212090),
	.w4(32'hbb553682),
	.w5(32'h358019fb),
	.w6(32'hba84d15e),
	.w7(32'h3b4f9319),
	.w8(32'h391833b5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3f765),
	.w1(32'h39f0bd77),
	.w2(32'h3a019928),
	.w3(32'hb92415d7),
	.w4(32'h3af4da23),
	.w5(32'hbb99d51f),
	.w6(32'hba30bb31),
	.w7(32'h3a7fec53),
	.w8(32'hbacd62f3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39787a01),
	.w1(32'hbb7294ce),
	.w2(32'h37525e80),
	.w3(32'hbaaefcee),
	.w4(32'hb97a76c0),
	.w5(32'hb9787b03),
	.w6(32'hb935c5b1),
	.w7(32'hba6aeec6),
	.w8(32'hbb98e88a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a479839),
	.w1(32'h3b702d18),
	.w2(32'hba7e33ef),
	.w3(32'h3b65b352),
	.w4(32'h3afa7316),
	.w5(32'hbc057108),
	.w6(32'hbb8a20e2),
	.w7(32'hb8c7a7ef),
	.w8(32'hb9d704a0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd468e2),
	.w1(32'hbb0d0c4d),
	.w2(32'hb6f3779b),
	.w3(32'hbb0a05d8),
	.w4(32'h3b8b925b),
	.w5(32'hbadb6110),
	.w6(32'h3c172010),
	.w7(32'h3bfee7ec),
	.w8(32'hbb15c387),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea9eef),
	.w1(32'hb9dbc047),
	.w2(32'h3c07a786),
	.w3(32'hb9f0b65f),
	.w4(32'h39a94ccd),
	.w5(32'hbba7b603),
	.w6(32'hbb87225e),
	.w7(32'h3adca346),
	.w8(32'hbb18fd74),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ec230b),
	.w1(32'h3b64bf9e),
	.w2(32'hb9e6c581),
	.w3(32'hbbcb011b),
	.w4(32'h3af9dafd),
	.w5(32'h3bbb6298),
	.w6(32'hb957cac9),
	.w7(32'hbb4b35be),
	.w8(32'hbbb82619),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba0646),
	.w1(32'hbbc758bd),
	.w2(32'h3af4963a),
	.w3(32'h3b201602),
	.w4(32'h3b7e6e12),
	.w5(32'h3bddc904),
	.w6(32'h3a0a1fcd),
	.w7(32'h3b186627),
	.w8(32'h3b4f43ab),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a714e97),
	.w1(32'hba980839),
	.w2(32'hbb2184c8),
	.w3(32'h3bd79f55),
	.w4(32'h3bcdf04a),
	.w5(32'hbb8408b0),
	.w6(32'h3c03376f),
	.w7(32'h3b328c6c),
	.w8(32'hbb9e3cfa),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b799225),
	.w1(32'hbb82b3ec),
	.w2(32'hba1cc842),
	.w3(32'hbb58f2a2),
	.w4(32'hb9bda925),
	.w5(32'hbb03acbf),
	.w6(32'hba8f7767),
	.w7(32'hb9fa9b22),
	.w8(32'hbb62665e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9962db3),
	.w1(32'hbbb7a598),
	.w2(32'h3ae2650b),
	.w3(32'hbb2828d6),
	.w4(32'hba814b27),
	.w5(32'hbb5c4a9a),
	.w6(32'hb91c5fac),
	.w7(32'hbb5af47f),
	.w8(32'hbaf58032),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba424979),
	.w1(32'hba79d8ab),
	.w2(32'hbb0eef5a),
	.w3(32'hbb9ced3d),
	.w4(32'hb9d77ce4),
	.w5(32'h3c3331f3),
	.w6(32'hbb8e8016),
	.w7(32'hbb4e56c6),
	.w8(32'h3ba9264e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad6f1c),
	.w1(32'hbb081a79),
	.w2(32'hba0be6eb),
	.w3(32'h3c12fe44),
	.w4(32'h3bb8918b),
	.w5(32'hbb58e760),
	.w6(32'h3c17fe28),
	.w7(32'h3b8b89d8),
	.w8(32'hba447c65),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba03ef8),
	.w1(32'hbb4fd4ef),
	.w2(32'h3b367399),
	.w3(32'hbb2514eb),
	.w4(32'h388d8490),
	.w5(32'hbbbafeb4),
	.w6(32'hbb6e01f4),
	.w7(32'hbb8fdd77),
	.w8(32'hbbb44ec4),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7c968),
	.w1(32'hbb21b24c),
	.w2(32'h3b347e53),
	.w3(32'hbac49115),
	.w4(32'h3aafb73e),
	.w5(32'h3bb1878a),
	.w6(32'hbb5d4641),
	.w7(32'h3989dde5),
	.w8(32'h3aab7b39),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4a903),
	.w1(32'hbb24f924),
	.w2(32'hbab5dcbc),
	.w3(32'h3b62a49d),
	.w4(32'h3b0cdf74),
	.w5(32'h3b3ca9a6),
	.w6(32'h3bc1fa33),
	.w7(32'h3b483ecf),
	.w8(32'hb80460cb),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e61ab),
	.w1(32'hbad4b16f),
	.w2(32'h3ab56bbe),
	.w3(32'h3ae56ae4),
	.w4(32'h3ad729ed),
	.w5(32'h3aeba56f),
	.w6(32'hbad98ace),
	.w7(32'hbb0b900a),
	.w8(32'h3b7cb652),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03c214),
	.w1(32'hbabfe0b0),
	.w2(32'hbb06f715),
	.w3(32'hbb9c09ca),
	.w4(32'h3abfe189),
	.w5(32'hbc09c402),
	.w6(32'hbab896af),
	.w7(32'h386e22bb),
	.w8(32'hbb318e66),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf55e97),
	.w1(32'hbb8c4cd4),
	.w2(32'h3af08cd7),
	.w3(32'hbb4d5775),
	.w4(32'h3ad3b224),
	.w5(32'h3b338ef4),
	.w6(32'hba7348c1),
	.w7(32'h3a918356),
	.w8(32'hba91bfd8),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a2cb5),
	.w1(32'h3b7d68b4),
	.w2(32'h3bd456c0),
	.w3(32'hbb5e17dd),
	.w4(32'h3b6d9a2d),
	.w5(32'h3bb7f809),
	.w6(32'hbb4fb9ab),
	.w7(32'h3b09e48f),
	.w8(32'h3b30e371),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab2a20),
	.w1(32'h3a0b0466),
	.w2(32'hba5087b5),
	.w3(32'h3b977692),
	.w4(32'h3a74608c),
	.w5(32'h3b949ab1),
	.w6(32'h3c0bd509),
	.w7(32'h3adab022),
	.w8(32'h3adae387),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c60ac),
	.w1(32'hbb25a9ab),
	.w2(32'hbaec1d04),
	.w3(32'h3b2a9c78),
	.w4(32'h3b9e0e17),
	.w5(32'hbbbc40b7),
	.w6(32'hbb04cf17),
	.w7(32'hb9ed46b4),
	.w8(32'hbc066ff4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba16dea),
	.w1(32'hbb803c41),
	.w2(32'hbba300be),
	.w3(32'hbb7f0eda),
	.w4(32'hbb47b36e),
	.w5(32'hba9b0a60),
	.w6(32'hbbfdf510),
	.w7(32'hbc04d53b),
	.w8(32'h3b25f1e0),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d70cb),
	.w1(32'h3b2be759),
	.w2(32'h3ac85304),
	.w3(32'hb8c4bae1),
	.w4(32'h3a6fc04a),
	.w5(32'hbba94f43),
	.w6(32'h3b6f45f3),
	.w7(32'hbaa9e739),
	.w8(32'hbbefd3b5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66c68e),
	.w1(32'h3a9474b3),
	.w2(32'h3bc4d87c),
	.w3(32'h3bfce14b),
	.w4(32'hba572b15),
	.w5(32'h3a6e37a3),
	.w6(32'h3b8e7492),
	.w7(32'h396bb63e),
	.w8(32'h3c3bbf64),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b511cbe),
	.w1(32'h3c33b500),
	.w2(32'hbc60742e),
	.w3(32'h3c8f1ed4),
	.w4(32'h3a761d48),
	.w5(32'hba623989),
	.w6(32'hbb59ace4),
	.w7(32'hb9230a7b),
	.w8(32'hbc1014be),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f18be),
	.w1(32'hbbbbf444),
	.w2(32'h3a1f2493),
	.w3(32'hbb3d9b47),
	.w4(32'hba99253c),
	.w5(32'h37e9b44f),
	.w6(32'h3c96f7a7),
	.w7(32'hbbc7d177),
	.w8(32'h3b6fd585),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8652c),
	.w1(32'h3b0e770f),
	.w2(32'hbbd31abf),
	.w3(32'h3c838573),
	.w4(32'hbaf8c5bd),
	.w5(32'hba8ad1a5),
	.w6(32'hbb74cb89),
	.w7(32'h3b908b81),
	.w8(32'hbbb3bb00),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dbdeb4),
	.w1(32'hbb323c72),
	.w2(32'hbb142567),
	.w3(32'h3a98279c),
	.w4(32'hb903ec65),
	.w5(32'h396c067d),
	.w6(32'h3b28c490),
	.w7(32'h39a0ca53),
	.w8(32'hbbea7416),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c95f0),
	.w1(32'hbc077475),
	.w2(32'hbb86a5fa),
	.w3(32'h3b4eeb14),
	.w4(32'h3b4e146b),
	.w5(32'hb98b15aa),
	.w6(32'hbb6eb561),
	.w7(32'hb77d80e6),
	.w8(32'hbb276d45),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc36d0),
	.w1(32'hbad6da68),
	.w2(32'h3adcd300),
	.w3(32'hb88a8338),
	.w4(32'hbb1e7532),
	.w5(32'hba6ed2cc),
	.w6(32'hba5b2233),
	.w7(32'hb951ac4a),
	.w8(32'h3b0ff445),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule