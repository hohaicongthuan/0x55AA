module layer_10_featuremap_234(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba72c09),
	.w1(32'h3bee7463),
	.w2(32'h3c998f17),
	.w3(32'h3c1eb6b5),
	.w4(32'hbabdebc1),
	.w5(32'h3a36a390),
	.w6(32'hbb96a838),
	.w7(32'h3bf60c67),
	.w8(32'h3afb7ceb),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b180a),
	.w1(32'h3bbe3e6b),
	.w2(32'h3bc8f745),
	.w3(32'h3a33f76f),
	.w4(32'hbbf4d08d),
	.w5(32'hbb781885),
	.w6(32'hbbf2a1a0),
	.w7(32'hbb3a8ba3),
	.w8(32'h3c4f6f2f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6438),
	.w1(32'h3b1045a2),
	.w2(32'hbbc9605f),
	.w3(32'h3be57296),
	.w4(32'hbc86ec6d),
	.w5(32'hbc294026),
	.w6(32'h3c30a636),
	.w7(32'hbba1360d),
	.w8(32'h3bf4773a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d9a16),
	.w1(32'hbc3fb0f4),
	.w2(32'hbb656f42),
	.w3(32'h3c9d51d9),
	.w4(32'hb8b50a9c),
	.w5(32'hbbe7795d),
	.w6(32'hbbae37f9),
	.w7(32'hbb14f3a3),
	.w8(32'hbbbd5847),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a499bf),
	.w1(32'hbc87d073),
	.w2(32'hbbb46bd3),
	.w3(32'h3b1eb93b),
	.w4(32'h3a2b45dc),
	.w5(32'hba247246),
	.w6(32'h3b849082),
	.w7(32'hbb05ef23),
	.w8(32'h3b4083da),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0b54d),
	.w1(32'h3cb111c0),
	.w2(32'hbb9e22c3),
	.w3(32'hbc0ab2f9),
	.w4(32'hbb6f25b2),
	.w5(32'h3b877ca3),
	.w6(32'h3bf8fd2d),
	.w7(32'h3bfe16af),
	.w8(32'hbc1aebd1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9d403),
	.w1(32'hbc607018),
	.w2(32'hbb136030),
	.w3(32'h3b1e3060),
	.w4(32'h3c63a4be),
	.w5(32'h3ad05354),
	.w6(32'hbc600814),
	.w7(32'h3c0bbe26),
	.w8(32'h3b6c3d50),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cda6e6a),
	.w1(32'hba1863d1),
	.w2(32'h3ba0214e),
	.w3(32'hbb45d379),
	.w4(32'hbb853d7e),
	.w5(32'h3b512b38),
	.w6(32'h3b3dd33a),
	.w7(32'hbb9ac862),
	.w8(32'h3c236381),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c2c7c),
	.w1(32'h3ba8a1ce),
	.w2(32'h3a9d18e3),
	.w3(32'hbb3d1498),
	.w4(32'hbc180a49),
	.w5(32'h3befcb58),
	.w6(32'hbc50f10f),
	.w7(32'h3b52fa58),
	.w8(32'hbadc508b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba513fe),
	.w1(32'hb84cf397),
	.w2(32'h3b873662),
	.w3(32'hba8bf698),
	.w4(32'hbb113c59),
	.w5(32'h3b0848f7),
	.w6(32'hbad50799),
	.w7(32'hbb3eab42),
	.w8(32'h3c84a3da),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f2763),
	.w1(32'h3aed857b),
	.w2(32'hbba4a558),
	.w3(32'hbc8777ee),
	.w4(32'h3c0819ad),
	.w5(32'h3bad8af1),
	.w6(32'hbbdc4aaa),
	.w7(32'h3b6c04cb),
	.w8(32'hbb30818e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce78dd),
	.w1(32'h3b22034d),
	.w2(32'h3c10b9f6),
	.w3(32'hbabd5a44),
	.w4(32'h3c2f3a64),
	.w5(32'hb9a0dad4),
	.w6(32'hbb2090a3),
	.w7(32'hb96ab051),
	.w8(32'h3c066e0d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5204d),
	.w1(32'hba383f61),
	.w2(32'hbc636c1e),
	.w3(32'hbb96c4a4),
	.w4(32'h3aaae1f6),
	.w5(32'h3ca0af7b),
	.w6(32'h3b7d9c7e),
	.w7(32'h3b12594d),
	.w8(32'h3c22d1a1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b9a13),
	.w1(32'h3bafbd63),
	.w2(32'hbbee3afd),
	.w3(32'h3c1665a5),
	.w4(32'h3a24cbf3),
	.w5(32'h3c20eedb),
	.w6(32'h3bf9f0f2),
	.w7(32'hbba04ae5),
	.w8(32'h3b6e0dcb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4a784),
	.w1(32'h38cf502d),
	.w2(32'hbbf7cb7b),
	.w3(32'h3933ee9f),
	.w4(32'h3ad1357e),
	.w5(32'hbb390ee4),
	.w6(32'hbba92a7d),
	.w7(32'hbbf0a644),
	.w8(32'h3ab1100a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cb52a),
	.w1(32'h3b3f70c4),
	.w2(32'h3ca76503),
	.w3(32'hbbdfa489),
	.w4(32'h3b623e2e),
	.w5(32'hbb43add3),
	.w6(32'hba2d7bdd),
	.w7(32'h3a647ca2),
	.w8(32'h3aa52784),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad601ec),
	.w1(32'hbc26ca49),
	.w2(32'h3cf4fd1e),
	.w3(32'h39ef1ff2),
	.w4(32'h36179572),
	.w5(32'hbae6dc88),
	.w6(32'hbaae9b54),
	.w7(32'h3b10c4fd),
	.w8(32'h3b443332),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace3da6),
	.w1(32'hbbd5b907),
	.w2(32'hbc118061),
	.w3(32'hbbe97a0a),
	.w4(32'h3ba165eb),
	.w5(32'hb94907b0),
	.w6(32'h3c157b73),
	.w7(32'hbbbfa08a),
	.w8(32'h3b5ba39b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2f6a3),
	.w1(32'hbbb41fa0),
	.w2(32'hbb153810),
	.w3(32'hb9924489),
	.w4(32'h3b7b9520),
	.w5(32'h3c4f7b11),
	.w6(32'hbc53e7b7),
	.w7(32'hbc41afb5),
	.w8(32'h3a5129d7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8d773),
	.w1(32'h3bfcabea),
	.w2(32'h3bf472a7),
	.w3(32'hbc17d4ab),
	.w4(32'hbba103cf),
	.w5(32'hbc04eb20),
	.w6(32'h3c2b6eba),
	.w7(32'h3c6b8ea0),
	.w8(32'hba012997),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05e132),
	.w1(32'hba62b707),
	.w2(32'h3c436592),
	.w3(32'hbba41c67),
	.w4(32'hbb3be9e8),
	.w5(32'hbabc6b17),
	.w6(32'hbb9a5cb5),
	.w7(32'h3c312f60),
	.w8(32'h3c1bad93),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc319d16),
	.w1(32'h3aac3ddd),
	.w2(32'hbc8095da),
	.w3(32'hbac80962),
	.w4(32'h3b7a4f84),
	.w5(32'hb9d59109),
	.w6(32'h3bc8ba2b),
	.w7(32'h38de86f0),
	.w8(32'h3b3fcda7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5db552),
	.w1(32'hba0267c6),
	.w2(32'h3bb8c022),
	.w3(32'h3bc17430),
	.w4(32'hba1d596f),
	.w5(32'hbbbc6b48),
	.w6(32'h3afa128a),
	.w7(32'h3c8cce1a),
	.w8(32'h3c7ab1a2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7632f5),
	.w1(32'h3c57bce7),
	.w2(32'h3bb7bf34),
	.w3(32'h3cc52ce9),
	.w4(32'hbb1cbfd4),
	.w5(32'hbc987f40),
	.w6(32'h3aa33de9),
	.w7(32'h3cb50cb0),
	.w8(32'hba3286af),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a62a5),
	.w1(32'hbbebfffc),
	.w2(32'h3b9c8399),
	.w3(32'h3d0a7d2b),
	.w4(32'h3bfc5748),
	.w5(32'h3c4b5845),
	.w6(32'h3b9da2a4),
	.w7(32'hbc34a864),
	.w8(32'h3c4153f6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc211ffc),
	.w1(32'hbaf3ff4a),
	.w2(32'hbc3a0c07),
	.w3(32'h3c7ac3f9),
	.w4(32'h3c5eb8f5),
	.w5(32'h3c261fcd),
	.w6(32'h3c0ac9d4),
	.w7(32'h3c564c9f),
	.w8(32'hbb29c847),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59656e),
	.w1(32'h3c072683),
	.w2(32'h3bef0834),
	.w3(32'hbbdce2aa),
	.w4(32'h3a102833),
	.w5(32'h3a3502a7),
	.w6(32'h3ba99bb7),
	.w7(32'hb96c52c6),
	.w8(32'h3a5f9b34),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0085f4),
	.w1(32'hb9ff6eb9),
	.w2(32'h3bf5ffd6),
	.w3(32'h3ad7eb4d),
	.w4(32'hba531bec),
	.w5(32'hbb22cc2e),
	.w6(32'h3bffaba7),
	.w7(32'hbc5eb8ba),
	.w8(32'hbb500315),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b284489),
	.w1(32'h3c365e44),
	.w2(32'hbbb38300),
	.w3(32'h3c0bf472),
	.w4(32'hbb117b5a),
	.w5(32'h3b88e2a5),
	.w6(32'h3cbd8ecf),
	.w7(32'h3c059723),
	.w8(32'h3b02f0e5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0f2dc),
	.w1(32'h3b99eac4),
	.w2(32'hbc4f37f3),
	.w3(32'hbbf7079c),
	.w4(32'h3aacdcdd),
	.w5(32'hbc2b8f26),
	.w6(32'h3c34cd8e),
	.w7(32'h3bb4170d),
	.w8(32'hba96d20f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3c853),
	.w1(32'h3c09c1ec),
	.w2(32'h3b539bc5),
	.w3(32'hbb5ab0a1),
	.w4(32'hbb0624c6),
	.w5(32'h3c8fa664),
	.w6(32'h3a96a249),
	.w7(32'h3b9af721),
	.w8(32'h3ac90ef4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1399f),
	.w1(32'h3c528fb4),
	.w2(32'hbbe99892),
	.w3(32'hbc7e7dc9),
	.w4(32'h3b404849),
	.w5(32'h3ba16585),
	.w6(32'h3c067e38),
	.w7(32'h3b6e306a),
	.w8(32'h3b2de93e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c087ac8),
	.w1(32'h3a2c3652),
	.w2(32'h3bafd8a4),
	.w3(32'hbb9182ce),
	.w4(32'hbb8a3cfb),
	.w5(32'h3c9b1171),
	.w6(32'hbc5c03f4),
	.w7(32'hb9e9cd3d),
	.w8(32'hbb21f922),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80aa26),
	.w1(32'hbca1c193),
	.w2(32'h3c36a7b5),
	.w3(32'hb9037aad),
	.w4(32'hbb67f4ef),
	.w5(32'hbbce149d),
	.w6(32'h3acc8848),
	.w7(32'h3bdbc69a),
	.w8(32'h3a27015a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd57d7),
	.w1(32'h3bd6f9ea),
	.w2(32'h3c27f339),
	.w3(32'h3c95cda1),
	.w4(32'h3a8cbb70),
	.w5(32'hbb873769),
	.w6(32'hbbd15cce),
	.w7(32'h3c2e70b5),
	.w8(32'h3c8aab82),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cffeb),
	.w1(32'hbb2d53e9),
	.w2(32'hbc5785cf),
	.w3(32'h3ca3c4db),
	.w4(32'h3b6d6b35),
	.w5(32'h3c8bed2e),
	.w6(32'hbc1967d6),
	.w7(32'h3baf62ee),
	.w8(32'hbabb857c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf20271),
	.w1(32'h3a90f892),
	.w2(32'h3ab94456),
	.w3(32'hbbf2f3f3),
	.w4(32'hbc1ce323),
	.w5(32'hbbcdf0a1),
	.w6(32'hba8bd87b),
	.w7(32'h3bb75971),
	.w8(32'h39e084bd),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfaa60d),
	.w1(32'hba8bfca0),
	.w2(32'h3b21b488),
	.w3(32'h3c660551),
	.w4(32'hbbcf3915),
	.w5(32'h3909e04a),
	.w6(32'hbba123fc),
	.w7(32'hbb854088),
	.w8(32'h3b9b30d7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47f1e9),
	.w1(32'h3c5c2fb7),
	.w2(32'hbbd53e03),
	.w3(32'hbc9b41ec),
	.w4(32'hbc36dd95),
	.w5(32'h38c4d371),
	.w6(32'h3ba227ae),
	.w7(32'h3c1608cf),
	.w8(32'hbc050488),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac507d1),
	.w1(32'h3a94f949),
	.w2(32'h3aa4b150),
	.w3(32'h3bae6ec2),
	.w4(32'h3b5b113c),
	.w5(32'h3a49e9fb),
	.w6(32'hbc1c3cf0),
	.w7(32'hb89cb97b),
	.w8(32'h3bd76f6f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36795290),
	.w1(32'hbbb9eb3c),
	.w2(32'h3b7533f7),
	.w3(32'hbc4dda8e),
	.w4(32'h3bf8dbb1),
	.w5(32'hbbad5ca8),
	.w6(32'hbb5e8ce0),
	.w7(32'hbb2a76eb),
	.w8(32'hbb42fb2b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07e82f),
	.w1(32'hbb0616a9),
	.w2(32'h3c051d2c),
	.w3(32'hbaca7148),
	.w4(32'h3b206029),
	.w5(32'hbb15bbc6),
	.w6(32'hbc3494a8),
	.w7(32'hbb2f4a2b),
	.w8(32'h3c329d9a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53939c),
	.w1(32'h3c593977),
	.w2(32'hba956138),
	.w3(32'h3c5f43e9),
	.w4(32'hbaf244aa),
	.w5(32'hbbb284db),
	.w6(32'h3c26b528),
	.w7(32'h3c478bc8),
	.w8(32'hbb50305d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34d0d6),
	.w1(32'h3bc75653),
	.w2(32'h3c987c33),
	.w3(32'hbb963bf7),
	.w4(32'hbb42a213),
	.w5(32'hbb2ae4a0),
	.w6(32'hbc118941),
	.w7(32'h3c01f5c9),
	.w8(32'h3a83846f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb855f),
	.w1(32'hba69bda9),
	.w2(32'h3c48f2cd),
	.w3(32'hbbcebc47),
	.w4(32'h3c5c9879),
	.w5(32'h3b93b633),
	.w6(32'h3943ed7c),
	.w7(32'hba7506a6),
	.w8(32'hb8c7e324),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb936f),
	.w1(32'hbbf76697),
	.w2(32'hbcd1397f),
	.w3(32'h3b98309e),
	.w4(32'hbc217db4),
	.w5(32'h3c2ca39d),
	.w6(32'hbbd099a2),
	.w7(32'h3b0a1ee3),
	.w8(32'h3b3d10a6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca02b5b),
	.w1(32'h3bb49617),
	.w2(32'h3bc26ff8),
	.w3(32'h3b249c12),
	.w4(32'h3c046189),
	.w5(32'hb935e9ad),
	.w6(32'hba3d7bb1),
	.w7(32'hba5933ad),
	.w8(32'h3a1b043f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb601400),
	.w1(32'h3c0edfde),
	.w2(32'hbc48b08e),
	.w3(32'h3ccd933d),
	.w4(32'hbabf1ef6),
	.w5(32'h3be3cab9),
	.w6(32'h3bd729dd),
	.w7(32'hbbe6e6b7),
	.w8(32'h3d0ffb9c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8423fb),
	.w1(32'h3bf6e359),
	.w2(32'h3c12a901),
	.w3(32'hbbbb7d78),
	.w4(32'h3b55ea0c),
	.w5(32'h3bc99421),
	.w6(32'hbabf1e7f),
	.w7(32'hbba4b697),
	.w8(32'hbba749f1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc84b00),
	.w1(32'hbb90a255),
	.w2(32'hbc46cbca),
	.w3(32'hbbf1d5d8),
	.w4(32'h3b9d7dc9),
	.w5(32'h3b2cd9f0),
	.w6(32'hbc469409),
	.w7(32'h3a0968b9),
	.w8(32'h3c043784),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7df1c6f),
	.w1(32'hbb5a6c20),
	.w2(32'h3b3feb72),
	.w3(32'hba3b51da),
	.w4(32'h3b0d7809),
	.w5(32'hba839b6f),
	.w6(32'h39830beb),
	.w7(32'h3ada256c),
	.w8(32'hbadf2d40),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29ff19),
	.w1(32'hbc27c819),
	.w2(32'h3ab5d674),
	.w3(32'hbc78bfbb),
	.w4(32'hbbb1687d),
	.w5(32'hbb2de2f1),
	.w6(32'h3c950083),
	.w7(32'h3c3e00de),
	.w8(32'hbb93273e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf866f1),
	.w1(32'h39cf6d30),
	.w2(32'hbc453696),
	.w3(32'hbc520684),
	.w4(32'h3b8481e7),
	.w5(32'h3c988880),
	.w6(32'hbb442ce2),
	.w7(32'h3ca7ec76),
	.w8(32'hbbfbdd92),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08fc86),
	.w1(32'h3b73f5c7),
	.w2(32'h3a6e0c24),
	.w3(32'hbacf181a),
	.w4(32'hbb30c366),
	.w5(32'h3b3e231c),
	.w6(32'hb9151ad1),
	.w7(32'h3aab7bb2),
	.w8(32'h3c00111f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca14ec5),
	.w1(32'h3c1eadca),
	.w2(32'h3bc49969),
	.w3(32'h3c9895b8),
	.w4(32'h3c8e0b70),
	.w5(32'hbc3f3828),
	.w6(32'hbbb90b50),
	.w7(32'hbbc840d9),
	.w8(32'hbb95eb1c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca61495),
	.w1(32'h3b4b2f5b),
	.w2(32'h3b8745b3),
	.w3(32'hbbfcf3f6),
	.w4(32'hbb839e74),
	.w5(32'hbb75ddb8),
	.w6(32'h3a0e9738),
	.w7(32'hbb9b4219),
	.w8(32'h3b743b1f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61c5ab),
	.w1(32'h3a8a7ed1),
	.w2(32'hbaf6524e),
	.w3(32'hbbb74e04),
	.w4(32'hbb29eb64),
	.w5(32'hbbbdd911),
	.w6(32'hb88bc3f3),
	.w7(32'hba912877),
	.w8(32'h3b238a17),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb997d12),
	.w1(32'hbb382057),
	.w2(32'h36b113d6),
	.w3(32'h3c08df7f),
	.w4(32'h3aaa8089),
	.w5(32'hbacc23cd),
	.w6(32'hbc2e6e87),
	.w7(32'hbb696b21),
	.w8(32'hbd0700f4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2c0c3),
	.w1(32'hb9c5d4fe),
	.w2(32'h3b1f6cb2),
	.w3(32'h3b36e82b),
	.w4(32'hbba40221),
	.w5(32'hbabebea3),
	.w6(32'h3b97622f),
	.w7(32'h3866e12f),
	.w8(32'h3b2b1d57),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd9083),
	.w1(32'h3ab047d6),
	.w2(32'h3c0af2f0),
	.w3(32'hbca8bf24),
	.w4(32'hbb94f597),
	.w5(32'hbb11ccae),
	.w6(32'hbb279e40),
	.w7(32'h3a84c6e7),
	.w8(32'hba23dafd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d002432),
	.w1(32'h3bf0ee52),
	.w2(32'h3a9015eb),
	.w3(32'hbb6e19fc),
	.w4(32'h3bbafce7),
	.w5(32'h3b309e78),
	.w6(32'hbbd2484f),
	.w7(32'h3a5cd8cc),
	.w8(32'hbaf553a4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45a767),
	.w1(32'hbaf8784c),
	.w2(32'hba1c31cb),
	.w3(32'h3c104c6f),
	.w4(32'hba4d4457),
	.w5(32'hbc6fb749),
	.w6(32'hbb3b2f25),
	.w7(32'h3a06ad01),
	.w8(32'h3b6cbecf),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19164e),
	.w1(32'hb9651be0),
	.w2(32'h3c09fa43),
	.w3(32'h3c00ba81),
	.w4(32'h3c0f02d1),
	.w5(32'h3bd376e1),
	.w6(32'hbbc9c6b6),
	.w7(32'hbbe0ab9b),
	.w8(32'hbac77b36),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ead0b),
	.w1(32'h3b6f0d7c),
	.w2(32'hbd06303f),
	.w3(32'hbb8164e1),
	.w4(32'hbb9e1d20),
	.w5(32'hbbc2952e),
	.w6(32'hba8acc5d),
	.w7(32'h3b09d82e),
	.w8(32'h3b118e7f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7da52),
	.w1(32'hba5c1bcb),
	.w2(32'h3a9d930a),
	.w3(32'hbc4719c6),
	.w4(32'hbae91805),
	.w5(32'hbc2034ec),
	.w6(32'hbb4443d8),
	.w7(32'hb9b09ad4),
	.w8(32'hbc7c233b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7047b6),
	.w1(32'hba5edc76),
	.w2(32'h3c311251),
	.w3(32'hbad70936),
	.w4(32'hbb16acca),
	.w5(32'h39a7299e),
	.w6(32'hbc7a7743),
	.w7(32'hbb902e1f),
	.w8(32'h3c8008ea),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb5767),
	.w1(32'h3b357144),
	.w2(32'hbb6af2fd),
	.w3(32'hbb725369),
	.w4(32'h39f4063a),
	.w5(32'hbb653c57),
	.w6(32'h38901cff),
	.w7(32'h3b6d8d41),
	.w8(32'h393c1693),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb812b10f),
	.w1(32'h3b846f40),
	.w2(32'h3d74903b),
	.w3(32'h3bcee387),
	.w4(32'hbaeb1fb3),
	.w5(32'hbab559f7),
	.w6(32'hbb0b58d2),
	.w7(32'hbbbc9b3d),
	.w8(32'h3c05d109),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb813009a),
	.w1(32'hbb6f6ca5),
	.w2(32'h3a9f87c2),
	.w3(32'h3bc43501),
	.w4(32'h371682f2),
	.w5(32'h3c1e6c50),
	.w6(32'hbaddcbec),
	.w7(32'h3c930860),
	.w8(32'hbba91598),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ed4d4),
	.w1(32'h3a61c807),
	.w2(32'hbc197160),
	.w3(32'h3b6e0f7e),
	.w4(32'h3a03f588),
	.w5(32'hbcaf9051),
	.w6(32'hbb39eeb2),
	.w7(32'h3a82b7b1),
	.w8(32'h3c20d072),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9afd8b),
	.w1(32'hbcf6d0c4),
	.w2(32'hbc76a2e0),
	.w3(32'hbbf82d5c),
	.w4(32'hbbe5df1e),
	.w5(32'h397ecd5b),
	.w6(32'h3c33cf35),
	.w7(32'hbaa361c1),
	.w8(32'h3d1fa269),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb69de),
	.w1(32'h3ae83209),
	.w2(32'h3b57c9ae),
	.w3(32'hbad2bc7f),
	.w4(32'hbbf75d1a),
	.w5(32'hbb22f457),
	.w6(32'hbb184057),
	.w7(32'h3ade4392),
	.w8(32'h3b6bf86e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefebaa),
	.w1(32'hbb2ad335),
	.w2(32'hbb83525c),
	.w3(32'hbb9ec745),
	.w4(32'hbb47ec14),
	.w5(32'hbcb47e64),
	.w6(32'h3a144dc8),
	.w7(32'hbbf48965),
	.w8(32'hbb20d2e8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86f5092),
	.w1(32'hb7e15811),
	.w2(32'h3be44d83),
	.w3(32'h3aa41d45),
	.w4(32'hbb8d81e9),
	.w5(32'h38df6a5d),
	.w6(32'hbc3222f4),
	.w7(32'hbb809748),
	.w8(32'h3a718ecd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395480ff),
	.w1(32'h3b09d335),
	.w2(32'h390ed07d),
	.w3(32'h3bc5bb4a),
	.w4(32'h3bd40ca7),
	.w5(32'hbb83054d),
	.w6(32'h3c8591b8),
	.w7(32'hba79c5c6),
	.w8(32'h3bd0f66d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada1a4a),
	.w1(32'hbb818a72),
	.w2(32'h3d0526c5),
	.w3(32'hbbcb25b1),
	.w4(32'h3be5ec4a),
	.w5(32'hbb149971),
	.w6(32'hbbe11b73),
	.w7(32'hbb12c111),
	.w8(32'h3c32a4c0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ef76),
	.w1(32'h3c1530ac),
	.w2(32'h3b5254f5),
	.w3(32'h3bf02e2f),
	.w4(32'hbb42efc1),
	.w5(32'hbbf82a61),
	.w6(32'hbc04a42a),
	.w7(32'h3bf93a55),
	.w8(32'h3c174fad),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab40aa4),
	.w1(32'h3b7b8d60),
	.w2(32'h3b8e3c29),
	.w3(32'hbc4590d5),
	.w4(32'hbbcba1fd),
	.w5(32'h3bde018a),
	.w6(32'h3abb4358),
	.w7(32'hbc0c581b),
	.w8(32'hbb83c6f2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b3f5d),
	.w1(32'hbb79e599),
	.w2(32'hba3b60f5),
	.w3(32'hbc0bb6e7),
	.w4(32'h388c7bd5),
	.w5(32'h3c2b97b1),
	.w6(32'h3c674c4c),
	.w7(32'hbb655624),
	.w8(32'hbb05f7b5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5573a),
	.w1(32'h3adb8417),
	.w2(32'h3c31b2ba),
	.w3(32'hbaa3f170),
	.w4(32'hbafcbca3),
	.w5(32'hbbadb21b),
	.w6(32'h39a29bbf),
	.w7(32'hbcd720fb),
	.w8(32'hbc64c02a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb369ed3),
	.w1(32'hbb90c691),
	.w2(32'h3b5fa7c2),
	.w3(32'hbb6d9b66),
	.w4(32'h3c1dd04a),
	.w5(32'hb9fb7f0e),
	.w6(32'h3be9fa79),
	.w7(32'hbb15d9ee),
	.w8(32'h3bb332a6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a51df),
	.w1(32'hbb938108),
	.w2(32'h3b26b2ef),
	.w3(32'h3bc29325),
	.w4(32'h39a367c2),
	.w5(32'hbc422bb9),
	.w6(32'hbbc2730c),
	.w7(32'h3c415159),
	.w8(32'h3c2b4c06),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16bfaf),
	.w1(32'h3b4ed9ce),
	.w2(32'h3ac15c35),
	.w3(32'hbb205e4d),
	.w4(32'hba6991b6),
	.w5(32'hbb0e8b0f),
	.w6(32'hbba8d99c),
	.w7(32'h3ba98df2),
	.w8(32'hbc2fd0da),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd6224),
	.w1(32'h3b44918f),
	.w2(32'hbb40ea18),
	.w3(32'h3ad41534),
	.w4(32'hb9ca9de8),
	.w5(32'hba05f0da),
	.w6(32'hbc20a22b),
	.w7(32'hbbab3f35),
	.w8(32'h3b4ec481),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acce671),
	.w1(32'h3b305f4f),
	.w2(32'hbb8c86c8),
	.w3(32'h3bb9efae),
	.w4(32'hb9c997e1),
	.w5(32'h3a9b5b52),
	.w6(32'h3a08df76),
	.w7(32'hb9ad658f),
	.w8(32'hbab6ebc1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba19491),
	.w1(32'h3b9f0450),
	.w2(32'hbb1deb8b),
	.w3(32'h3b07f22b),
	.w4(32'h3a68fdbb),
	.w5(32'hba662bc7),
	.w6(32'h3b6c9ddd),
	.w7(32'hbb13a6db),
	.w8(32'h3b82015c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae08d68),
	.w1(32'hbbb6f593),
	.w2(32'hbb01808c),
	.w3(32'h3c9339c5),
	.w4(32'hbbcae0ea),
	.w5(32'h3cc39c0a),
	.w6(32'h3c0d1644),
	.w7(32'hbb1e06a8),
	.w8(32'h3994efa8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53975b),
	.w1(32'h3b62b898),
	.w2(32'h3b8bedee),
	.w3(32'h3bbd71a3),
	.w4(32'hb985aa72),
	.w5(32'h3c8d0bf4),
	.w6(32'h3bbeabaf),
	.w7(32'h3be33793),
	.w8(32'hbba56039),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba13c15),
	.w1(32'hbb8e79da),
	.w2(32'h3b9b38fc),
	.w3(32'h3aa9ffa1),
	.w4(32'h3c18e3af),
	.w5(32'hbb13dc69),
	.w6(32'h3b787d3c),
	.w7(32'hbbf41cfd),
	.w8(32'hbb88bece),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4681ee),
	.w1(32'h3aa26f63),
	.w2(32'h3b213333),
	.w3(32'h3aa230a8),
	.w4(32'h39ea98da),
	.w5(32'hbae34a2b),
	.w6(32'h3d24aea7),
	.w7(32'hbaca7258),
	.w8(32'hbbcf1853),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ce0c9),
	.w1(32'hbb4a05d7),
	.w2(32'hbc0ed3f1),
	.w3(32'h3b235185),
	.w4(32'h3c00c82e),
	.w5(32'hb9e4d126),
	.w6(32'hbaed2779),
	.w7(32'h3bbf61cf),
	.w8(32'h3c17c5ed),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9863849),
	.w1(32'h389aaafb),
	.w2(32'hbcec4629),
	.w3(32'h3bcaa056),
	.w4(32'hbc90fb50),
	.w5(32'hb9d9b913),
	.w6(32'hbb3cdc27),
	.w7(32'h3a7029af),
	.w8(32'h3b55ea70),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34600a),
	.w1(32'h3c324714),
	.w2(32'h3c261524),
	.w3(32'h3b7f87e1),
	.w4(32'h3b728fbe),
	.w5(32'h3b872265),
	.w6(32'h3b7bfea1),
	.w7(32'hbb371341),
	.w8(32'hbc8165d8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27705c),
	.w1(32'h3a4468cc),
	.w2(32'hb92792af),
	.w3(32'hbaa6bc9e),
	.w4(32'h37d3b93e),
	.w5(32'hbc254302),
	.w6(32'hba7acee6),
	.w7(32'hbbf3ba4e),
	.w8(32'h3b550f35),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80c906),
	.w1(32'hbb7f6977),
	.w2(32'h38b573c0),
	.w3(32'h3b7e1526),
	.w4(32'h3ae68ef0),
	.w5(32'hbbd313f4),
	.w6(32'hba75438c),
	.w7(32'h3c32391f),
	.w8(32'hb93ff060),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9253e2),
	.w1(32'hba873b53),
	.w2(32'hbb1e6a75),
	.w3(32'hbc07e12d),
	.w4(32'h3c685b38),
	.w5(32'hbaeb6335),
	.w6(32'h3bff7ab1),
	.w7(32'hba0bb54f),
	.w8(32'h3bb5f611),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98c7a7),
	.w1(32'h3beb5d06),
	.w2(32'hbbe74d93),
	.w3(32'hbacb6b90),
	.w4(32'hbb88f989),
	.w5(32'h3a5c4c27),
	.w6(32'hbbf31123),
	.w7(32'h3bd3280a),
	.w8(32'hb4d6f4da),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb861),
	.w1(32'hbc793c7b),
	.w2(32'hba6b1c9b),
	.w3(32'hba84e9ae),
	.w4(32'h3b3d9eec),
	.w5(32'h3a7a2a38),
	.w6(32'hbc30a5d3),
	.w7(32'h3a24b206),
	.w8(32'h3be0b968),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf71a2),
	.w1(32'hbb4fb783),
	.w2(32'h39a23971),
	.w3(32'h3a878c59),
	.w4(32'hbc054fe2),
	.w5(32'h3ab655cb),
	.w6(32'h3bb9a217),
	.w7(32'hbc1342b4),
	.w8(32'h3a721056),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04dc82),
	.w1(32'h3b8ffde6),
	.w2(32'hbc2077a9),
	.w3(32'h3b56e1be),
	.w4(32'hbb9f9723),
	.w5(32'hb85a2106),
	.w6(32'h3a8fdd94),
	.w7(32'h3ae8a5fb),
	.w8(32'h3c63ce96),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23115e),
	.w1(32'hba83384b),
	.w2(32'hbac04d3e),
	.w3(32'h3c319252),
	.w4(32'hbb0cca76),
	.w5(32'h3b4d93a6),
	.w6(32'h3b6213ba),
	.w7(32'h389612b1),
	.w8(32'h3c08a6f8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb276659),
	.w1(32'h375623cd),
	.w2(32'h3b2a1c40),
	.w3(32'hbb91bbc5),
	.w4(32'hbaff4d78),
	.w5(32'h395a94ee),
	.w6(32'hbbe88256),
	.w7(32'h3bdc53bd),
	.w8(32'h3abea4e4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34e18c),
	.w1(32'h3ad2805d),
	.w2(32'hbc0978fb),
	.w3(32'hbb01f03f),
	.w4(32'h3c2eb95c),
	.w5(32'h3b41cee4),
	.w6(32'hbbd5d280),
	.w7(32'hbb4da31c),
	.w8(32'hba9863b3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5bfe1),
	.w1(32'h392e86ce),
	.w2(32'hbb575640),
	.w3(32'hba115530),
	.w4(32'h3bedc5c0),
	.w5(32'hbc099608),
	.w6(32'h3bec48bc),
	.w7(32'h3c3809f5),
	.w8(32'h3b83e296),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fe822),
	.w1(32'hbb86c19b),
	.w2(32'hbba79082),
	.w3(32'h3bbf57d6),
	.w4(32'hbb90e178),
	.w5(32'h3b851b08),
	.w6(32'h3bf999f4),
	.w7(32'hbb1cf5f7),
	.w8(32'hbb15aa20),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76df5c),
	.w1(32'h3c0bbe47),
	.w2(32'h3a5fce01),
	.w3(32'h3b09b26b),
	.w4(32'hbb87930a),
	.w5(32'h3afa9f15),
	.w6(32'hbb318d47),
	.w7(32'hbb3c1aa1),
	.w8(32'hbb1fc446),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc859d4d),
	.w1(32'h3bc181dd),
	.w2(32'hbb1abab5),
	.w3(32'hbc8640aa),
	.w4(32'hba332ed1),
	.w5(32'h3ab3e6c5),
	.w6(32'hbb4661e4),
	.w7(32'hbbaa4950),
	.w8(32'hb92fdbdd),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba786e83),
	.w1(32'hba8f7f35),
	.w2(32'h391a1135),
	.w3(32'h3a796ee5),
	.w4(32'hbb3ca3e4),
	.w5(32'hb9abdd17),
	.w6(32'h3b85d86b),
	.w7(32'hbb3f4513),
	.w8(32'hbbd7dd31),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc133c68),
	.w1(32'h37a49d53),
	.w2(32'h3c8c49eb),
	.w3(32'hbbffd30d),
	.w4(32'h3b8e5421),
	.w5(32'h3a8632fe),
	.w6(32'hbbaa5d7f),
	.w7(32'hbb91383b),
	.w8(32'hba8ed4a8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396358e8),
	.w1(32'h3b0feed7),
	.w2(32'hbb52fae5),
	.w3(32'hb9654f23),
	.w4(32'h3c4e6803),
	.w5(32'h3ba32f28),
	.w6(32'hbadceae3),
	.w7(32'hbb7b7f79),
	.w8(32'h3c46c8c6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77bdfa),
	.w1(32'h3b12c0e9),
	.w2(32'h3c3ff784),
	.w3(32'hbb909096),
	.w4(32'hbbbed69d),
	.w5(32'hb930f435),
	.w6(32'h3bd55ab2),
	.w7(32'h3882402d),
	.w8(32'h3b9422fe),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b13c4),
	.w1(32'h3d30aca9),
	.w2(32'hba9a5877),
	.w3(32'hba1fc3fe),
	.w4(32'h3c00c010),
	.w5(32'hbc01e506),
	.w6(32'h3c270c91),
	.w7(32'h3c6a35dd),
	.w8(32'hbb90d8f2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0197ee),
	.w1(32'h3b1eaf21),
	.w2(32'hbb60d948),
	.w3(32'h3afda922),
	.w4(32'hb9a0d52e),
	.w5(32'h3c7647a4),
	.w6(32'hbb62b731),
	.w7(32'hbba23804),
	.w8(32'hbc3acb51),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cce6a03),
	.w1(32'hbaeb60fb),
	.w2(32'hbc3d2270),
	.w3(32'hbc0376ee),
	.w4(32'h3b8ee530),
	.w5(32'hbab74c5d),
	.w6(32'hbaa6939e),
	.w7(32'hbb273c4c),
	.w8(32'h3a6a600f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc44c80),
	.w1(32'h3bc17b4c),
	.w2(32'hbbad6f96),
	.w3(32'h3c8d2cf6),
	.w4(32'h3a600fec),
	.w5(32'h3a1a51e0),
	.w6(32'h3b840cb5),
	.w7(32'hbbd004c1),
	.w8(32'hbbe3e516),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce70cf2),
	.w1(32'hbbfe3130),
	.w2(32'hbaf11a92),
	.w3(32'hbb677d39),
	.w4(32'hbbd91791),
	.w5(32'hbb90d833),
	.w6(32'h3b0c66bc),
	.w7(32'hba259d94),
	.w8(32'h39b594b6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addda32),
	.w1(32'h3c3ac399),
	.w2(32'h3bd1512e),
	.w3(32'hbc0fa33e),
	.w4(32'hbbd4c7b9),
	.w5(32'hbc283665),
	.w6(32'hbb4eb819),
	.w7(32'h3a5b7233),
	.w8(32'hbc5b8624),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb710fca),
	.w1(32'h3bce7429),
	.w2(32'hbc20faab),
	.w3(32'hbd0a4e05),
	.w4(32'h3bddaacb),
	.w5(32'h3b2a629f),
	.w6(32'h3bf139e6),
	.w7(32'h3b917148),
	.w8(32'hb9271fee),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2e0dd),
	.w1(32'hbc3d4bd2),
	.w2(32'h3c7a8251),
	.w3(32'hb722fa75),
	.w4(32'h3bd27235),
	.w5(32'h3b136157),
	.w6(32'hbb615053),
	.w7(32'hbb0ac2a4),
	.w8(32'hbc4163a4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a9259),
	.w1(32'hbc0c9404),
	.w2(32'hba52df05),
	.w3(32'h3c2089a5),
	.w4(32'hb9763c20),
	.w5(32'hbb8d3967),
	.w6(32'h3b96ff26),
	.w7(32'h3c26b63a),
	.w8(32'h3bbcfdf1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6a1f6),
	.w1(32'h3c3587dc),
	.w2(32'hbc013c05),
	.w3(32'hbb538cc9),
	.w4(32'hbb1f957b),
	.w5(32'h3c8f2ecc),
	.w6(32'hbccda83c),
	.w7(32'hbc0f0c00),
	.w8(32'hbb251a2f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eab0a),
	.w1(32'h3b4530f2),
	.w2(32'hbc2398f4),
	.w3(32'hbc0bbd10),
	.w4(32'hbb8bbecb),
	.w5(32'h3c759b1f),
	.w6(32'h3b212ef2),
	.w7(32'h3a6fbe57),
	.w8(32'h3c588ab9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d101e1d),
	.w1(32'hbb81c383),
	.w2(32'hbb519100),
	.w3(32'hbbb24401),
	.w4(32'hbad55cbd),
	.w5(32'hbc13f04f),
	.w6(32'hbc305abe),
	.w7(32'hbba160d0),
	.w8(32'h3bc2bd28),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad54953),
	.w1(32'hbb93d324),
	.w2(32'hbac21d73),
	.w3(32'h3841d812),
	.w4(32'h3bbd2b06),
	.w5(32'hbbdcfe4a),
	.w6(32'h3b07370d),
	.w7(32'hba2452be),
	.w8(32'h3c7e865e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77ad49),
	.w1(32'hbadfc7c6),
	.w2(32'h3bb222fe),
	.w3(32'h3bda96f4),
	.w4(32'hba745c26),
	.w5(32'h3b6b11c7),
	.w6(32'h3c23baae),
	.w7(32'h3b86c0b1),
	.w8(32'h3c8b3720),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abffd2c),
	.w1(32'hb51e824a),
	.w2(32'h3c4b1e4f),
	.w3(32'h3b936936),
	.w4(32'h3ac42fec),
	.w5(32'hbbee2eed),
	.w6(32'h3c3b738e),
	.w7(32'hb8391834),
	.w8(32'h3b81e4e0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a4d5),
	.w1(32'hbc7e8e95),
	.w2(32'hbbc65422),
	.w3(32'hbb9b7e01),
	.w4(32'hbc4cd5bd),
	.w5(32'hbc2cd5f0),
	.w6(32'hbbe7011a),
	.w7(32'h3c26c1fd),
	.w8(32'hbb997e2b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c9b40),
	.w1(32'hbb01d915),
	.w2(32'h3bddf4f3),
	.w3(32'hba9993d9),
	.w4(32'hbc65610f),
	.w5(32'h3bbb07c5),
	.w6(32'h3b8b07c4),
	.w7(32'hbc2a8388),
	.w8(32'hbb8a89a6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07d0e3),
	.w1(32'hbc0cdce4),
	.w2(32'hba529f40),
	.w3(32'h3b607857),
	.w4(32'hbc03a671),
	.w5(32'hbc9c4808),
	.w6(32'hbbe33145),
	.w7(32'hbb717364),
	.w8(32'hbc820866),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc967af6),
	.w1(32'hbbb8214e),
	.w2(32'h3c23afe1),
	.w3(32'hbbef3f07),
	.w4(32'hbc0c766f),
	.w5(32'hbbdbc5ed),
	.w6(32'hbb689c06),
	.w7(32'hbb361353),
	.w8(32'hbb38d8c7),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc329b49),
	.w1(32'hbb824989),
	.w2(32'h3aef0053),
	.w3(32'h3b39ee38),
	.w4(32'hbc5afc62),
	.w5(32'h3bcaa8ca),
	.w6(32'hb76382ae),
	.w7(32'hbb015c75),
	.w8(32'hbbaaf781),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70afa2),
	.w1(32'h3d0ca8bf),
	.w2(32'hbc31405c),
	.w3(32'h3ba413c3),
	.w4(32'hbca04edc),
	.w5(32'h3a2f7ae2),
	.w6(32'hbbb131db),
	.w7(32'hba3bc35e),
	.w8(32'hbc3db808),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5aec7),
	.w1(32'h3d1fd60c),
	.w2(32'hbbda9579),
	.w3(32'h3c64da4a),
	.w4(32'h3b1c09d1),
	.w5(32'hbb2c850e),
	.w6(32'hbb619d79),
	.w7(32'hbb90cdf7),
	.w8(32'hbb7bc6c2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb28ed),
	.w1(32'hba1f6413),
	.w2(32'h3abcfdf0),
	.w3(32'hbc160245),
	.w4(32'h3b2d31d8),
	.w5(32'h3bccd349),
	.w6(32'hbb42053c),
	.w7(32'h3c05a8d4),
	.w8(32'h3b94053b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc429b04),
	.w1(32'hbc168c44),
	.w2(32'h3c6dce5a),
	.w3(32'hbc02818f),
	.w4(32'hbc2baa56),
	.w5(32'hbb44c66e),
	.w6(32'h3c114df4),
	.w7(32'h3c100975),
	.w8(32'hbb334b93),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac679d),
	.w1(32'hb90173f3),
	.w2(32'h3b9d366c),
	.w3(32'h3c92a03c),
	.w4(32'h3c31864a),
	.w5(32'hbbae13ec),
	.w6(32'hbbbb8852),
	.w7(32'hba45aaf4),
	.w8(32'hb9df736b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b1bff),
	.w1(32'hbae168ae),
	.w2(32'h3916e4a7),
	.w3(32'hba0292bc),
	.w4(32'hba21bcd9),
	.w5(32'hb986adbf),
	.w6(32'hbb6d9d33),
	.w7(32'hba33a647),
	.w8(32'hbb9b53fb),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdfa5d),
	.w1(32'hba2e71d3),
	.w2(32'hb99bef7a),
	.w3(32'h3ac2e54c),
	.w4(32'h3c588040),
	.w5(32'hbbd193c5),
	.w6(32'h3bcda6f1),
	.w7(32'h3a3873f1),
	.w8(32'h3c2e4dd1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13888a),
	.w1(32'hba4f66c3),
	.w2(32'hbcf2d58d),
	.w3(32'hbba07190),
	.w4(32'h3b2c7ae3),
	.w5(32'h39beeb98),
	.w6(32'h3cd0169b),
	.w7(32'h38c6e607),
	.w8(32'hbb6f1f69),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a499d),
	.w1(32'h3902c712),
	.w2(32'hbc81d4bb),
	.w3(32'hbc21b697),
	.w4(32'h3b71115e),
	.w5(32'hbbee53c3),
	.w6(32'h3c06c604),
	.w7(32'h3b8b44f4),
	.w8(32'hbc461ed2),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39914589),
	.w1(32'hbaa8c22a),
	.w2(32'hbc0c0680),
	.w3(32'hbc235fa8),
	.w4(32'h3bddd412),
	.w5(32'h3b62c98c),
	.w6(32'hbb992174),
	.w7(32'hb8c3abc0),
	.w8(32'hbbb4973d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace2655),
	.w1(32'h3c02e0f3),
	.w2(32'hb9932468),
	.w3(32'hbb2b38f1),
	.w4(32'hbbb311cc),
	.w5(32'hbaaf121b),
	.w6(32'hbb1a01bf),
	.w7(32'h3c0e7c3e),
	.w8(32'hbbce7231),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf9d8e),
	.w1(32'hbb235e8d),
	.w2(32'hbb88dbac),
	.w3(32'hbbe165a6),
	.w4(32'hbbb5b3d2),
	.w5(32'hbc78c7df),
	.w6(32'h3b05e568),
	.w7(32'h3c172404),
	.w8(32'hbc038222),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d6bc0),
	.w1(32'hba2b7b62),
	.w2(32'h3b01e7e0),
	.w3(32'hba0b54c8),
	.w4(32'hbc04e207),
	.w5(32'hbba5b0d6),
	.w6(32'hbb8f3327),
	.w7(32'hba20174b),
	.w8(32'hbb0701ff),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b325df8),
	.w1(32'hba9e9f9c),
	.w2(32'hba001392),
	.w3(32'hbbcf29f5),
	.w4(32'h3b71a91c),
	.w5(32'hbb7be2eb),
	.w6(32'h3c984075),
	.w7(32'h3aa9d585),
	.w8(32'hbc273883),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8f7e4),
	.w1(32'hbc2c2e9c),
	.w2(32'hbb86eb98),
	.w3(32'h3bf16d06),
	.w4(32'hbc174694),
	.w5(32'hbb913a3c),
	.w6(32'hbb12a600),
	.w7(32'hbbc7ac30),
	.w8(32'h3ba703c5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e1c88),
	.w1(32'hbb552a48),
	.w2(32'hbaa07500),
	.w3(32'hbc4aaf07),
	.w4(32'hbc31ee82),
	.w5(32'hbb2c981d),
	.w6(32'hbc2e9535),
	.w7(32'h3c672063),
	.w8(32'h3a5ed5e5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fa304),
	.w1(32'h3bb84336),
	.w2(32'h3b727faa),
	.w3(32'hbbf83e58),
	.w4(32'hbb339901),
	.w5(32'hbbd3011a),
	.w6(32'hbc803e60),
	.w7(32'hbaeb231c),
	.w8(32'hb8964f62),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11f6a6),
	.w1(32'hba20dff1),
	.w2(32'hbc3a85f9),
	.w3(32'hbb377583),
	.w4(32'h3b6a686e),
	.w5(32'h3a681606),
	.w6(32'hbb122646),
	.w7(32'hbc7e4653),
	.w8(32'hbbbe59f2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0207ba),
	.w1(32'hbc1d58ac),
	.w2(32'h3cea23df),
	.w3(32'hbb32b108),
	.w4(32'h3be6e1f9),
	.w5(32'h3bc12605),
	.w6(32'h3b8573d6),
	.w7(32'h3abe3225),
	.w8(32'h3c216af6),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5945b1),
	.w1(32'h3bac5de2),
	.w2(32'hbc70055a),
	.w3(32'h3bcf689b),
	.w4(32'h3b4bb7f0),
	.w5(32'hba2f9cd3),
	.w6(32'hbc45df9c),
	.w7(32'h3b70c1fb),
	.w8(32'h3ca41854),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda253e),
	.w1(32'h3b9fcbb0),
	.w2(32'h3d147180),
	.w3(32'h3a5a4984),
	.w4(32'h3bb9f74a),
	.w5(32'h3a709535),
	.w6(32'hbad685fa),
	.w7(32'hb8e6a453),
	.w8(32'hbb845e90),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd90aa),
	.w1(32'hbb615e17),
	.w2(32'hba75143b),
	.w3(32'hbb30ae3f),
	.w4(32'hbb7041aa),
	.w5(32'hbbb580c7),
	.w6(32'h3c466319),
	.w7(32'h3bba9dd6),
	.w8(32'h3c14cc16),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb64b4),
	.w1(32'h3beb0097),
	.w2(32'h3abd85e3),
	.w3(32'h3bd16ce0),
	.w4(32'h3a697a68),
	.w5(32'h3623f640),
	.w6(32'hbb1e2005),
	.w7(32'hbc2b4454),
	.w8(32'h3ab0cced),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9974cc),
	.w1(32'h3b28cd14),
	.w2(32'hbbe121a3),
	.w3(32'h3c48b9bc),
	.w4(32'h3be3cf81),
	.w5(32'hbb23f286),
	.w6(32'hbc325b48),
	.w7(32'h3b2f0488),
	.w8(32'hbba48747),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5cd59),
	.w1(32'hbb6491b7),
	.w2(32'h3b9cf91d),
	.w3(32'h3a823163),
	.w4(32'h3c2a6314),
	.w5(32'h3b94d1bb),
	.w6(32'hbafad0ea),
	.w7(32'h3a0092cb),
	.w8(32'hbbd7f675),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ed22f),
	.w1(32'hbbabe041),
	.w2(32'hbb353968),
	.w3(32'h3b867d6b),
	.w4(32'h3bff8af5),
	.w5(32'hbb815d2c),
	.w6(32'h3b8d7a10),
	.w7(32'hbbab31e7),
	.w8(32'h3ac6e13a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf06057),
	.w1(32'hbb9a33db),
	.w2(32'hbb903d34),
	.w3(32'h39c26846),
	.w4(32'h3c82830a),
	.w5(32'h3c099ea2),
	.w6(32'h3b99342c),
	.w7(32'h3a840e61),
	.w8(32'hbc873376),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab53bc8),
	.w1(32'hbb896087),
	.w2(32'hb83b036f),
	.w3(32'h3b73b124),
	.w4(32'h3b291b68),
	.w5(32'hbc05b929),
	.w6(32'hbbafb739),
	.w7(32'hbc4e184f),
	.w8(32'hbc0a9d45),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e304b),
	.w1(32'hbbf0c062),
	.w2(32'hbc063e8c),
	.w3(32'hbab13e05),
	.w4(32'h3d283088),
	.w5(32'hbb39b9ee),
	.w6(32'h3b8605fb),
	.w7(32'h3a74dc69),
	.w8(32'hbc0f11aa),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12bf6f),
	.w1(32'hbbcc88a0),
	.w2(32'hbc72704f),
	.w3(32'hbb958338),
	.w4(32'hbb88ae9a),
	.w5(32'hbc3cf75a),
	.w6(32'hbb242d8c),
	.w7(32'h3b945a17),
	.w8(32'hbb2a83e3),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf69fb3),
	.w1(32'h3cb05a86),
	.w2(32'h3b77617e),
	.w3(32'h3a33b903),
	.w4(32'hb9cc145e),
	.w5(32'hbbd43c97),
	.w6(32'h3a6833bd),
	.w7(32'hbc308080),
	.w8(32'hbb6222b7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7d88a),
	.w1(32'hbc209191),
	.w2(32'hbc2b6907),
	.w3(32'hbc3b096c),
	.w4(32'hbb747c94),
	.w5(32'hba0db9fa),
	.w6(32'h3c24ffb9),
	.w7(32'h3aa2ea1e),
	.w8(32'hbc96435c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c625583),
	.w1(32'hbb015852),
	.w2(32'hbb57518c),
	.w3(32'h3c1c7982),
	.w4(32'hbc35345a),
	.w5(32'hb97073a4),
	.w6(32'hbbcd9f19),
	.w7(32'hbc4358a6),
	.w8(32'h3bcb1b41),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40cc1c),
	.w1(32'h3ad46130),
	.w2(32'h3a2c9a04),
	.w3(32'h38afc88e),
	.w4(32'h3a82731f),
	.w5(32'hbb4b86c4),
	.w6(32'hbae1bee6),
	.w7(32'h398a299a),
	.w8(32'h3b13f500),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c519370),
	.w1(32'hbc1e4a55),
	.w2(32'h3b52f442),
	.w3(32'hbbae893f),
	.w4(32'h388d6e05),
	.w5(32'hb990624a),
	.w6(32'hb9c0b964),
	.w7(32'h3b9f3b64),
	.w8(32'h3d0a894b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39b30d),
	.w1(32'h3c07615c),
	.w2(32'h39606822),
	.w3(32'h3ba2f6b7),
	.w4(32'h3b82f42b),
	.w5(32'hbb950111),
	.w6(32'hbc5cee9f),
	.w7(32'hbc5665d0),
	.w8(32'h3b8bff56),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f762d),
	.w1(32'hbb30452c),
	.w2(32'hbc0e4f2a),
	.w3(32'hbcbc3784),
	.w4(32'hbb751a51),
	.w5(32'hb9abcd77),
	.w6(32'h3ac8dacc),
	.w7(32'hb9b5b293),
	.w8(32'hbbf7b3f6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cfd21),
	.w1(32'h3b653c7a),
	.w2(32'h3a7acac5),
	.w3(32'h3b1a41f4),
	.w4(32'hbbcc337a),
	.w5(32'h3bb51c59),
	.w6(32'hbb049116),
	.w7(32'hb92a0ce9),
	.w8(32'h3bf3abdd),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e242e),
	.w1(32'h3b1f26f1),
	.w2(32'hbc42e5ca),
	.w3(32'hba3cff3b),
	.w4(32'h3be8c245),
	.w5(32'h3bd2be9a),
	.w6(32'h3a1830d4),
	.w7(32'hbb022a5b),
	.w8(32'h3ccf6646),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81fe5f),
	.w1(32'h3b3e572b),
	.w2(32'hba170ab6),
	.w3(32'h3a8a0723),
	.w4(32'hb986a51e),
	.w5(32'hbbdbef61),
	.w6(32'hbb90fff1),
	.w7(32'hbbd3a915),
	.w8(32'hbbbc81b2),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cfb3a),
	.w1(32'hbb3ce063),
	.w2(32'h3b8391fd),
	.w3(32'hbc13ea3e),
	.w4(32'h3cdf0674),
	.w5(32'h38d64bad),
	.w6(32'hbc9eda7e),
	.w7(32'h3c30536d),
	.w8(32'h3b55a550),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc580a),
	.w1(32'hbc176bee),
	.w2(32'hbb07ad5b),
	.w3(32'h3c0def68),
	.w4(32'hbbc6762c),
	.w5(32'hbb431671),
	.w6(32'h39bb90c4),
	.w7(32'hbbdace79),
	.w8(32'hbb9ee3ec),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb070092),
	.w1(32'hbb91767f),
	.w2(32'h3a754dbb),
	.w3(32'hbc6d1f22),
	.w4(32'h3c0a4f15),
	.w5(32'h3b7d7078),
	.w6(32'h3b3cf197),
	.w7(32'hbbf57af6),
	.w8(32'h3b844bfd),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9e161),
	.w1(32'hbc4febcf),
	.w2(32'hbc129d48),
	.w3(32'h3c02ad8a),
	.w4(32'hba13e65a),
	.w5(32'h3abea8e6),
	.w6(32'hb9f32bd8),
	.w7(32'hbb948ad9),
	.w8(32'hb923771c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcac3b1),
	.w1(32'hbc8480da),
	.w2(32'hbcb21b01),
	.w3(32'h3b41e870),
	.w4(32'h38cb0a94),
	.w5(32'hbc899ef0),
	.w6(32'h3bb22387),
	.w7(32'hbb5e760b),
	.w8(32'hbc2fd290),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71fcfa),
	.w1(32'hbbd3c2e1),
	.w2(32'hbb46f89b),
	.w3(32'hba4e7143),
	.w4(32'h3a83bb0e),
	.w5(32'h3bf2c38d),
	.w6(32'h3b3874d0),
	.w7(32'h3caf267e),
	.w8(32'hbb84b70d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fe65c),
	.w1(32'h3ad92b96),
	.w2(32'hbca336ac),
	.w3(32'hbbe2d40a),
	.w4(32'h39dd50de),
	.w5(32'hbb0839e3),
	.w6(32'hbc3ee869),
	.w7(32'h3bb50885),
	.w8(32'hbc05f5e1),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f372c6),
	.w1(32'hbb0c61b2),
	.w2(32'h3c830c32),
	.w3(32'hbb3068ae),
	.w4(32'hbad14b47),
	.w5(32'h3aa2fc6b),
	.w6(32'h39e854fc),
	.w7(32'hbb8bcf6f),
	.w8(32'h3b8025ad),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba95e9a),
	.w1(32'hbc31442f),
	.w2(32'h3bbe1d39),
	.w3(32'hbbd6da6a),
	.w4(32'hbbdd6d9d),
	.w5(32'hbb4e9e9f),
	.w6(32'hba4c9b7c),
	.w7(32'hb9b7fe33),
	.w8(32'h3aa9b2e3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7f641),
	.w1(32'h3c9a2012),
	.w2(32'hbb4c8718),
	.w3(32'hbba25278),
	.w4(32'h3b7c53ab),
	.w5(32'hbb0156da),
	.w6(32'h3bfda0df),
	.w7(32'h3c9bed45),
	.w8(32'h3bd1a84a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a10fc1),
	.w1(32'hbb3d2a68),
	.w2(32'hbaa3fbd9),
	.w3(32'hbbb5567e),
	.w4(32'h3a0bff19),
	.w5(32'h3c01ab27),
	.w6(32'hbb03d0df),
	.w7(32'h3aae48c3),
	.w8(32'hbbdb01e8),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa44e17),
	.w1(32'hbc12b431),
	.w2(32'hbc01da63),
	.w3(32'h3ba23efb),
	.w4(32'h3ab2ad5e),
	.w5(32'hbb1284f2),
	.w6(32'h35999e5d),
	.w7(32'hbbc01ae0),
	.w8(32'hbad423dc),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2208e),
	.w1(32'h3b1e10e5),
	.w2(32'h3b85cb46),
	.w3(32'h3adaa9f5),
	.w4(32'h3c7eee6c),
	.w5(32'hbb87c3da),
	.w6(32'hbb7b9912),
	.w7(32'hbbd63835),
	.w8(32'h3bc50a28),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15d149),
	.w1(32'h3c4f91d6),
	.w2(32'h3b26bb97),
	.w3(32'h3b6d679a),
	.w4(32'hbbe030a0),
	.w5(32'h39d80a16),
	.w6(32'hbb893755),
	.w7(32'h3b9b5bb3),
	.w8(32'hbc7416bb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad25d19),
	.w1(32'h3a05ec4b),
	.w2(32'h3d25d760),
	.w3(32'h3c86ff5f),
	.w4(32'hbb349e89),
	.w5(32'hbc03ca2e),
	.w6(32'hb8c89eb1),
	.w7(32'hbb9659ce),
	.w8(32'h3a34c666),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab400c8),
	.w1(32'h3b4c8459),
	.w2(32'h3bc2c6d5),
	.w3(32'h3b941368),
	.w4(32'h3c2daeba),
	.w5(32'h3b22d1c7),
	.w6(32'hbbe81320),
	.w7(32'h3c81a95e),
	.w8(32'h3b7a13b0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89c6ad),
	.w1(32'h3a588291),
	.w2(32'hbba9f35d),
	.w3(32'h39010966),
	.w4(32'hbbfec2b8),
	.w5(32'hbc1e5d9e),
	.w6(32'h3b576d3b),
	.w7(32'hbba361af),
	.w8(32'h3bc3462e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4a58f),
	.w1(32'hbbd24dd0),
	.w2(32'hb9a6a9f9),
	.w3(32'h398c3634),
	.w4(32'h394bf1c6),
	.w5(32'hbaec8dc6),
	.w6(32'h3cae0712),
	.w7(32'h3b1026dd),
	.w8(32'h3b493dc9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a98f3e),
	.w1(32'hbb3e2ff2),
	.w2(32'h3a8086a6),
	.w3(32'h3be06324),
	.w4(32'hbbcd64fd),
	.w5(32'h3bbfdf50),
	.w6(32'h3b961e1a),
	.w7(32'h3b61a1e3),
	.w8(32'h3bd34996),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33bb74),
	.w1(32'h3c81cd13),
	.w2(32'hbc09a5f5),
	.w3(32'h3c8737a6),
	.w4(32'hbb85806b),
	.w5(32'hbc2a473b),
	.w6(32'hbb83693c),
	.w7(32'h3b24f36d),
	.w8(32'hbcaac758),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2eb4c),
	.w1(32'h3b100d50),
	.w2(32'h3c09da67),
	.w3(32'hbb60cc66),
	.w4(32'hbcc4d964),
	.w5(32'h3afb6f3a),
	.w6(32'hbb4d0a42),
	.w7(32'h3cbc41d0),
	.w8(32'h3cd82d44),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78847f),
	.w1(32'hbae83e30),
	.w2(32'hba3989f6),
	.w3(32'h3b70fe47),
	.w4(32'hba2b6077),
	.w5(32'hbb80c19b),
	.w6(32'h383701ed),
	.w7(32'h3c7d9604),
	.w8(32'h3b4b9930),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee2992),
	.w1(32'h3c4ac6ff),
	.w2(32'h3cc278c8),
	.w3(32'hbb7df554),
	.w4(32'hbc96d636),
	.w5(32'hbc75e6b7),
	.w6(32'hbb9495dd),
	.w7(32'h39dad733),
	.w8(32'hbc6567c9),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae3ead),
	.w1(32'hbcbf79c3),
	.w2(32'hbab8a725),
	.w3(32'hbba7905a),
	.w4(32'hbc544e02),
	.w5(32'hbab926df),
	.w6(32'hb97b33e5),
	.w7(32'h3b86af1a),
	.w8(32'hbb31780f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad80239),
	.w1(32'h3923187b),
	.w2(32'hbbe80bbd),
	.w3(32'h3cc5b369),
	.w4(32'h3c9a7665),
	.w5(32'h3ab04ae3),
	.w6(32'h3c13407f),
	.w7(32'h3cf18bf9),
	.w8(32'hb9a48282),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6beb0f),
	.w1(32'h3bc33547),
	.w2(32'hbc159412),
	.w3(32'hbc981948),
	.w4(32'h3ac2c96a),
	.w5(32'h3b671e0b),
	.w6(32'hbb779540),
	.w7(32'hbc8228a6),
	.w8(32'h3c2c9279),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17e5b3),
	.w1(32'h3c29dd7b),
	.w2(32'hb997ca2a),
	.w3(32'h3a961760),
	.w4(32'hbb40882f),
	.w5(32'hba9b1666),
	.w6(32'hb9b3755e),
	.w7(32'h3b1523bd),
	.w8(32'hb9248666),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13c515),
	.w1(32'h3c3b9519),
	.w2(32'h3c644a98),
	.w3(32'hbb9422d2),
	.w4(32'h3b2f0bce),
	.w5(32'h3aed2142),
	.w6(32'hbb1e017e),
	.w7(32'hba9c9b4f),
	.w8(32'h3cc863c4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e8d85),
	.w1(32'hbc0e4e7f),
	.w2(32'h3cd57aef),
	.w3(32'h3b459550),
	.w4(32'h3c01d12c),
	.w5(32'hbc14164c),
	.w6(32'h3baaa4e7),
	.w7(32'hbb7f105d),
	.w8(32'h3c4ecab8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa15784),
	.w1(32'h3b8bb360),
	.w2(32'h3ca1acde),
	.w3(32'hbc1e4dff),
	.w4(32'h3aef2414),
	.w5(32'hba13db2b),
	.w6(32'h3c1bc3ba),
	.w7(32'h3c93a40f),
	.w8(32'hbb049b12),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f77c0),
	.w1(32'h3c493f27),
	.w2(32'h3c920401),
	.w3(32'hbc5af9b4),
	.w4(32'h3c015e57),
	.w5(32'hbc91b561),
	.w6(32'h3c43606e),
	.w7(32'h3ccbbbac),
	.w8(32'h3bde548f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23f5e2),
	.w1(32'hbad9629e),
	.w2(32'hbb887693),
	.w3(32'hbc05bd33),
	.w4(32'h3c81d8b6),
	.w5(32'hbc1d6533),
	.w6(32'h3bf2fc77),
	.w7(32'h3c2f9a01),
	.w8(32'h3b89c968),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5435cf),
	.w1(32'hbb2cf54b),
	.w2(32'h3c122c7a),
	.w3(32'hbc8e331e),
	.w4(32'h3bd2f5ce),
	.w5(32'h3b8e4c6d),
	.w6(32'h3a494eeb),
	.w7(32'h3a38278b),
	.w8(32'hbaf881e7),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79e5d3),
	.w1(32'hbb9e0e4b),
	.w2(32'hbb09da57),
	.w3(32'hbbefd804),
	.w4(32'hbbba7f22),
	.w5(32'h3a5287f6),
	.w6(32'h3bfa05f2),
	.w7(32'hbb8aa085),
	.w8(32'h3b039bc1),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe3e88),
	.w1(32'hbc5c8dca),
	.w2(32'hbbac0017),
	.w3(32'h39853520),
	.w4(32'hbca0a2c2),
	.w5(32'h3b4bbff3),
	.w6(32'hbc0bbba2),
	.w7(32'h3b388724),
	.w8(32'hbc179752),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0405ba),
	.w1(32'hbac611e7),
	.w2(32'hbb9ad1a0),
	.w3(32'hbc03cce7),
	.w4(32'h3b581029),
	.w5(32'hbc166261),
	.w6(32'hbc465192),
	.w7(32'hb89da49c),
	.w8(32'hbb275f2e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b805109),
	.w1(32'hbb8e6a2d),
	.w2(32'hbbc2f306),
	.w3(32'h3b5f15ac),
	.w4(32'hbc83461a),
	.w5(32'h3c783be4),
	.w6(32'hbc0791ab),
	.w7(32'hbc1bc174),
	.w8(32'h3ab2758a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46e8fc),
	.w1(32'h3ca2777a),
	.w2(32'h3c363644),
	.w3(32'hbc25fbb8),
	.w4(32'hb8f55312),
	.w5(32'h3bdf3f39),
	.w6(32'hbc101873),
	.w7(32'hbb195d90),
	.w8(32'hba5d0ba8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5448be),
	.w1(32'hbc347452),
	.w2(32'h3beecbb6),
	.w3(32'hbaeb6187),
	.w4(32'h3b2f317c),
	.w5(32'h3c0746da),
	.w6(32'hbbf1cc69),
	.w7(32'h3935a3e0),
	.w8(32'h3b93e0fe),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb06d90),
	.w1(32'hbaae475e),
	.w2(32'h372f4390),
	.w3(32'hbc0e58c2),
	.w4(32'h3bba215a),
	.w5(32'hbbba538c),
	.w6(32'h3b78c0c6),
	.w7(32'h3bbc8805),
	.w8(32'hba0871de),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c809012),
	.w1(32'h3b8503e3),
	.w2(32'hbc0f1ecd),
	.w3(32'hbb3d62fb),
	.w4(32'h3b03eea1),
	.w5(32'h3c936dfc),
	.w6(32'h3b413952),
	.w7(32'h3a328563),
	.w8(32'h3c4540f8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd169cc),
	.w1(32'hba143ba9),
	.w2(32'h3bdfd234),
	.w3(32'hbc0dea60),
	.w4(32'h3b5e23ca),
	.w5(32'hbc3a4a28),
	.w6(32'hbb0ed8c7),
	.w7(32'h3accdb01),
	.w8(32'hbac7279d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b31e0),
	.w1(32'hbc128050),
	.w2(32'h3aab4d0d),
	.w3(32'h3c2ee7ab),
	.w4(32'h3d2a0f75),
	.w5(32'h3aee75a1),
	.w6(32'hba876989),
	.w7(32'h3c066dbe),
	.w8(32'h3c405777),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2aea8),
	.w1(32'h3c3495a1),
	.w2(32'hbb4afa23),
	.w3(32'h3c9fa079),
	.w4(32'h3ab58735),
	.w5(32'h3c828018),
	.w6(32'hbc08d9bb),
	.w7(32'h3bd1f22c),
	.w8(32'hbb660ac5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48013a),
	.w1(32'h3ba9ace4),
	.w2(32'h3b5e3f76),
	.w3(32'h3b831efd),
	.w4(32'h3bde1838),
	.w5(32'h3a588004),
	.w6(32'h3a7a8c7b),
	.w7(32'hb5bf9584),
	.w8(32'hbba3a796),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb651e87),
	.w1(32'h3cc7b0f9),
	.w2(32'hba88f220),
	.w3(32'hbb7501d7),
	.w4(32'h3925433a),
	.w5(32'h3b39b734),
	.w6(32'h3bf0d0fb),
	.w7(32'h3bf1e6bc),
	.w8(32'h3a017722),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26e71b),
	.w1(32'h3c480eac),
	.w2(32'hbaa99689),
	.w3(32'h3b79185a),
	.w4(32'hbc178697),
	.w5(32'h3bf3f7cf),
	.w6(32'h3cc2a051),
	.w7(32'h3ad3ac9b),
	.w8(32'h3caf967a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07057e),
	.w1(32'hbc8084a6),
	.w2(32'hbb83780e),
	.w3(32'hba98337c),
	.w4(32'h3c7251d7),
	.w5(32'h3a8f4b51),
	.w6(32'hbb30df8d),
	.w7(32'h3c01afa4),
	.w8(32'h3bfdf1b5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a58cb),
	.w1(32'hbc41b2dd),
	.w2(32'hbb731e7c),
	.w3(32'hbb8d08d3),
	.w4(32'h3a234857),
	.w5(32'hbc099fcf),
	.w6(32'h3ad52a0a),
	.w7(32'h3b4f06f9),
	.w8(32'hbcc1232c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3427ce),
	.w1(32'hbb2ab15d),
	.w2(32'h36a87e71),
	.w3(32'hbbe840cc),
	.w4(32'hbc28a802),
	.w5(32'h3c170e35),
	.w6(32'h3a16bf31),
	.w7(32'hba90e995),
	.w8(32'h3bde7846),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca63eac),
	.w1(32'h3aff582e),
	.w2(32'hbc4ee01f),
	.w3(32'h3ca3eb47),
	.w4(32'hba8269d5),
	.w5(32'h3c9d20b3),
	.w6(32'h3a2714b3),
	.w7(32'hba8029e9),
	.w8(32'h3c2f4f65),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4c513),
	.w1(32'h3a99d28e),
	.w2(32'h3b96598b),
	.w3(32'h3b175460),
	.w4(32'h3c47aa50),
	.w5(32'h3a4f4d46),
	.w6(32'h3bb0efeb),
	.w7(32'hbb66344b),
	.w8(32'h383c19e1),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a790680),
	.w1(32'hbc3464ec),
	.w2(32'h3c998a38),
	.w3(32'h3b198d50),
	.w4(32'h3a554ce7),
	.w5(32'hbbaa1ca3),
	.w6(32'h3c845ee8),
	.w7(32'h3c0c4622),
	.w8(32'h3cc3439e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd051e9),
	.w1(32'h3bed4e49),
	.w2(32'h3bca2649),
	.w3(32'h3c666ad8),
	.w4(32'h3bc384bb),
	.w5(32'h3ca1b3f5),
	.w6(32'h3c5d9363),
	.w7(32'h3b948641),
	.w8(32'hbb668177),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9dc2b),
	.w1(32'h3cd31b80),
	.w2(32'h3b63f477),
	.w3(32'h3c85dc50),
	.w4(32'hbbfba9ce),
	.w5(32'hbc4b43c6),
	.w6(32'h3c614709),
	.w7(32'hb9a2b87e),
	.w8(32'h3b21559c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b0cf1),
	.w1(32'h3c73cf2b),
	.w2(32'h3c5699ef),
	.w3(32'h3bce251a),
	.w4(32'h3c1d8e73),
	.w5(32'h3c0cb723),
	.w6(32'h3c4a7f95),
	.w7(32'hb9a2ad4e),
	.w8(32'h3c8d9748),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3a604),
	.w1(32'hbc23f022),
	.w2(32'hbb591bd3),
	.w3(32'hbbe36247),
	.w4(32'hb96777ba),
	.w5(32'h3b1f8353),
	.w6(32'h3b8b08fb),
	.w7(32'h3c758e1b),
	.w8(32'h3b49e00c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae37b71),
	.w1(32'hba8bc8ca),
	.w2(32'hbc386b04),
	.w3(32'hbb5554fa),
	.w4(32'h3aae14cb),
	.w5(32'h3b48332d),
	.w6(32'hbc2b13ae),
	.w7(32'h3b8a425b),
	.w8(32'hbbc8ec1e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc019e70),
	.w1(32'h3b802fd5),
	.w2(32'h3c818d24),
	.w3(32'h3c44a536),
	.w4(32'h3ca2bbd7),
	.w5(32'h3cd5868f),
	.w6(32'hbb370493),
	.w7(32'h3b26dbb2),
	.w8(32'hba82a7c6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc2b0f6),
	.w1(32'h3c1a7269),
	.w2(32'hbbf5b0f5),
	.w3(32'hbb6518e9),
	.w4(32'h397f6853),
	.w5(32'hbc37bebc),
	.w6(32'hbca1a53f),
	.w7(32'h3c126c01),
	.w8(32'hbb675d79),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedbb25),
	.w1(32'hbaae258e),
	.w2(32'h3b82ae93),
	.w3(32'h3caa5d4a),
	.w4(32'hba7f507d),
	.w5(32'hbb47d475),
	.w6(32'h3b3e0764),
	.w7(32'h3c0902b1),
	.w8(32'hbc5dcce1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babd5ce),
	.w1(32'h3ab9d332),
	.w2(32'h3a4a138b),
	.w3(32'hb99c420c),
	.w4(32'h3c945acb),
	.w5(32'h3c398637),
	.w6(32'h3a26d5a6),
	.w7(32'hbc112149),
	.w8(32'hbb366817),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66fd34),
	.w1(32'h3cbc9b82),
	.w2(32'hbae280be),
	.w3(32'hbb881248),
	.w4(32'h3d654e12),
	.w5(32'hbbd327b6),
	.w6(32'h3c4041a9),
	.w7(32'h3ae1a0dc),
	.w8(32'h3bfd7fa0),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0ed91b),
	.w1(32'hbc28f2c1),
	.w2(32'h3b8679e1),
	.w3(32'hbac31020),
	.w4(32'h3b7e0e14),
	.w5(32'hbb8d12e1),
	.w6(32'h3bdb3b57),
	.w7(32'h3c199193),
	.w8(32'h3b064dc0),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb751e6f),
	.w1(32'h3b1cdafd),
	.w2(32'h3baca454),
	.w3(32'hbadbfe1f),
	.w4(32'hbc2099d9),
	.w5(32'hbbd5327c),
	.w6(32'h3ca5b52c),
	.w7(32'h3bade0c6),
	.w8(32'hbbfc9710),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b612c28),
	.w1(32'hbbc50ecd),
	.w2(32'h3cc982f1),
	.w3(32'h3cc325ff),
	.w4(32'h39b9f449),
	.w5(32'h3aa4144c),
	.w6(32'h3cbc59c5),
	.w7(32'h3c9b962b),
	.w8(32'hb8147543),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9e8b7),
	.w1(32'h3d2f770d),
	.w2(32'h3c3ba3b0),
	.w3(32'h3a6b6878),
	.w4(32'h3bd6f8e1),
	.w5(32'h3be83b53),
	.w6(32'h3ba13652),
	.w7(32'hbb8c7969),
	.w8(32'hbb2d28e4),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3152c),
	.w1(32'hbba7c166),
	.w2(32'hbc3fac13),
	.w3(32'h3c066771),
	.w4(32'h3a6d9fb4),
	.w5(32'h3b896dba),
	.w6(32'hbb2bbe13),
	.w7(32'hbba7f747),
	.w8(32'hbb0d4d93),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a03b3),
	.w1(32'h39d4193e),
	.w2(32'h3bbebee5),
	.w3(32'h36a8a992),
	.w4(32'h3c102b63),
	.w5(32'hbb4076d5),
	.w6(32'h3a9d37b5),
	.w7(32'hbc8eff82),
	.w8(32'hbba19c80),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9189fd),
	.w1(32'h3bfc1b4f),
	.w2(32'hbba71085),
	.w3(32'h3c1b8147),
	.w4(32'h3b1183f0),
	.w5(32'h3b94954c),
	.w6(32'h3b52df19),
	.w7(32'h3b013850),
	.w8(32'hbb3847fa),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce6741c),
	.w1(32'h3c064ab0),
	.w2(32'hbc090536),
	.w3(32'h3af9e27d),
	.w4(32'h3bdacc49),
	.w5(32'hbb84e276),
	.w6(32'h3c9d2ee6),
	.w7(32'h3bd2b014),
	.w8(32'hbb856dd8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3238d0),
	.w1(32'h3c04f4ed),
	.w2(32'hbb43aadd),
	.w3(32'h3b3369fe),
	.w4(32'hbaedb394),
	.w5(32'h3b364da8),
	.w6(32'h3bfe3e7f),
	.w7(32'h39d68037),
	.w8(32'hb8c24a55),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1f1d9),
	.w1(32'h3bd3800f),
	.w2(32'hbb8f6923),
	.w3(32'h3a3b8ca7),
	.w4(32'h3bc6ebcd),
	.w5(32'h3ae2b8e8),
	.w6(32'hba81834d),
	.w7(32'h3c3d8b8c),
	.w8(32'h3a995506),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3536b3a8),
	.w1(32'h3bfc5aef),
	.w2(32'hba455b32),
	.w3(32'h3afda375),
	.w4(32'h3b9d1e4a),
	.w5(32'hbb36a5bf),
	.w6(32'hbb7e81ac),
	.w7(32'hbc4ec291),
	.w8(32'h3b7cd8f8),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c1a84),
	.w1(32'hba0bddd9),
	.w2(32'hbc5af4be),
	.w3(32'h3c41e825),
	.w4(32'hbb8ca1e0),
	.w5(32'hbc905faa),
	.w6(32'h3bc7f840),
	.w7(32'hbbbd891f),
	.w8(32'hbba859ab),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca66f66),
	.w1(32'hbb362a60),
	.w2(32'hba6fe27c),
	.w3(32'h3c34a2d7),
	.w4(32'h3834f470),
	.w5(32'h3bdcdcbd),
	.w6(32'h3ba73539),
	.w7(32'h3b9b3a9b),
	.w8(32'hb9bb17f3),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ea3e9),
	.w1(32'h3c90695f),
	.w2(32'hbb476d84),
	.w3(32'hbc552457),
	.w4(32'hbbb42bd8),
	.w5(32'hbbb709cd),
	.w6(32'h3b41e841),
	.w7(32'h3b812e6d),
	.w8(32'h3c04bcf6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39fd00),
	.w1(32'hbb99ccea),
	.w2(32'hbaf00e93),
	.w3(32'h3a8054ec),
	.w4(32'hbbb1eda8),
	.w5(32'h3af4fa0d),
	.w6(32'h3d0fcf9e),
	.w7(32'hbb51bb71),
	.w8(32'h3c255422),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec697c),
	.w1(32'hbb471124),
	.w2(32'hbaf81fa6),
	.w3(32'h3932323f),
	.w4(32'hb8e842e1),
	.w5(32'h39299222),
	.w6(32'hbb7843f5),
	.w7(32'hbad1aa7f),
	.w8(32'hb9c80e36),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b667262),
	.w1(32'h3bb07527),
	.w2(32'hbc7218fe),
	.w3(32'h3b52c843),
	.w4(32'hbb7e003e),
	.w5(32'hbc65fb9d),
	.w6(32'h3c3e1e61),
	.w7(32'h3bd8398c),
	.w8(32'h3c86f889),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc521b9a),
	.w1(32'h3afa2a66),
	.w2(32'h3abaaa30),
	.w3(32'h3bdd1117),
	.w4(32'h3c856a6c),
	.w5(32'hbbf34fc7),
	.w6(32'hbc2e26b7),
	.w7(32'hbc4d930d),
	.w8(32'hbc26b01d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be19ba9),
	.w1(32'hbb9285a3),
	.w2(32'hbb173aa2),
	.w3(32'h3c8f653b),
	.w4(32'hbbd0de16),
	.w5(32'hbb655ec2),
	.w6(32'h3cf77534),
	.w7(32'hbc2fddd1),
	.w8(32'hbc28a37d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba113db),
	.w1(32'h3c14d75d),
	.w2(32'hbaf3513f),
	.w3(32'hbb33b011),
	.w4(32'hbba9db83),
	.w5(32'hb7f0f346),
	.w6(32'h3bde879c),
	.w7(32'h395212fe),
	.w8(32'h3bace824),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3945e8),
	.w1(32'hbabbfaa3),
	.w2(32'h3a7a5254),
	.w3(32'hbc1910f1),
	.w4(32'h3b73df64),
	.w5(32'hbb9d7797),
	.w6(32'hbbf805ce),
	.w7(32'h3c1a57b1),
	.w8(32'h3b6e0bf3),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03d258),
	.w1(32'h3ad8119d),
	.w2(32'h3c6a35b6),
	.w3(32'hbbbbbaab),
	.w4(32'h3b8a4660),
	.w5(32'h3a0f35fd),
	.w6(32'h3c9a500d),
	.w7(32'hb9fbb7bf),
	.w8(32'hbbeb8740),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule