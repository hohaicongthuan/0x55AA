module layer_8_featuremap_161(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba55d6b),
	.w1(32'h3c37a70f),
	.w2(32'h3c3e7945),
	.w3(32'h3c0e39d9),
	.w4(32'h3bed3c78),
	.w5(32'h3c13dc61),
	.w6(32'h3c039d41),
	.w7(32'h39e14817),
	.w8(32'hbb8f6783),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2e088),
	.w1(32'hbbae4777),
	.w2(32'hbbf54f72),
	.w3(32'h3c6d0511),
	.w4(32'h39c80bad),
	.w5(32'hb890af81),
	.w6(32'h3ac95768),
	.w7(32'hbae5338f),
	.w8(32'h39e67fbc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc030263),
	.w1(32'hbc1ca4dc),
	.w2(32'hbc0204f7),
	.w3(32'hb9fa221b),
	.w4(32'h3a3d28df),
	.w5(32'h3c554619),
	.w6(32'h3a5e5a12),
	.w7(32'hbc497463),
	.w8(32'h3b8a4d96),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07786),
	.w1(32'hbb025247),
	.w2(32'hbc7c7c7a),
	.w3(32'h3c99ad8f),
	.w4(32'h3ba1d925),
	.w5(32'h39c7345c),
	.w6(32'h3c365ec8),
	.w7(32'hbac6ffc9),
	.w8(32'hbb7a7ef7),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42dbe4),
	.w1(32'hbba21460),
	.w2(32'hbbf84fbd),
	.w3(32'h3bac529f),
	.w4(32'h3af7b593),
	.w5(32'hba0ca8c4),
	.w6(32'h3b8d15a1),
	.w7(32'h3b67140f),
	.w8(32'h3a614e7f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2331f5),
	.w1(32'h3c4b45f3),
	.w2(32'h3c22dc95),
	.w3(32'hbb629b5d),
	.w4(32'h3b00fa70),
	.w5(32'h3c25278d),
	.w6(32'h3bbeab6c),
	.w7(32'h3c7bfcd6),
	.w8(32'h3c306ed2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a7b5b),
	.w1(32'h3b44e84b),
	.w2(32'hbbb1bc3e),
	.w3(32'h3c771b12),
	.w4(32'hbba6d377),
	.w5(32'hbc37581a),
	.w6(32'h3b3bce5c),
	.w7(32'h3b01c533),
	.w8(32'h3ab25ee8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb175034),
	.w1(32'hbb617487),
	.w2(32'hbc8cb1f7),
	.w3(32'hbc00c834),
	.w4(32'h3b817b3d),
	.w5(32'hbc67e275),
	.w6(32'hbc242b69),
	.w7(32'hbb1fac7d),
	.w8(32'h3b216c91),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca77419),
	.w1(32'h3b3c03a8),
	.w2(32'hbbb614a6),
	.w3(32'hbc761d13),
	.w4(32'h3a77c670),
	.w5(32'hbbb8147e),
	.w6(32'h3c74ba23),
	.w7(32'h3c321f6a),
	.w8(32'h3beb91ab),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e5d89),
	.w1(32'hbba89a3e),
	.w2(32'h3c2822f8),
	.w3(32'hbbc61d9d),
	.w4(32'hba95b3e3),
	.w5(32'h3c7d4e2d),
	.w6(32'hba5a747d),
	.w7(32'hbbbe5334),
	.w8(32'h3704d6ea),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9421e),
	.w1(32'h3919f11e),
	.w2(32'hbc0b966a),
	.w3(32'h3c137ad1),
	.w4(32'h3a9d538e),
	.w5(32'hbc818218),
	.w6(32'h3c72e934),
	.w7(32'h3c2f79f1),
	.w8(32'hbbac2308),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f7707),
	.w1(32'hbc152ebe),
	.w2(32'hbc0d6063),
	.w3(32'hbc51f573),
	.w4(32'hbc169c63),
	.w5(32'hbc472a6e),
	.w6(32'hbc29368e),
	.w7(32'hbbdcf08a),
	.w8(32'h3b283354),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4801c1),
	.w1(32'hbbde6c77),
	.w2(32'hba1382de),
	.w3(32'hbc184330),
	.w4(32'hbb58f3de),
	.w5(32'h398e7177),
	.w6(32'hbbf3d8be),
	.w7(32'hbad78246),
	.w8(32'hb8b95394),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5cce2),
	.w1(32'hba25b923),
	.w2(32'h3abc8c5a),
	.w3(32'hb9d66b9f),
	.w4(32'h3babb70f),
	.w5(32'h3c51b5d8),
	.w6(32'hbafb2375),
	.w7(32'hbb24ad59),
	.w8(32'h3c157744),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89de2b),
	.w1(32'h3b6110ba),
	.w2(32'hb9d0e607),
	.w3(32'h3ba6fcc3),
	.w4(32'h3823f137),
	.w5(32'hba920ec3),
	.w6(32'hb7daab2e),
	.w7(32'hbbad2e3b),
	.w8(32'hbbbc8ab1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5477e1),
	.w1(32'h3ab24712),
	.w2(32'hbb5999a2),
	.w3(32'hbadf8ffd),
	.w4(32'hbcc40ab8),
	.w5(32'hbc198a3b),
	.w6(32'h3c738b64),
	.w7(32'h3c56ec72),
	.w8(32'hbaaae865),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5dca4),
	.w1(32'h3c30407f),
	.w2(32'h3c1f988e),
	.w3(32'h3c1a4a7d),
	.w4(32'h3bdb813b),
	.w5(32'h3c8f137c),
	.w6(32'h3cad8e7a),
	.w7(32'h3b1d6e57),
	.w8(32'h3b11c4be),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a600bae),
	.w1(32'hbacf1691),
	.w2(32'hbbfa470c),
	.w3(32'hbb4a0dcc),
	.w4(32'hba78fa47),
	.w5(32'hbc689af2),
	.w6(32'hbb27a428),
	.w7(32'h3b394ed7),
	.w8(32'h3b9c726f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95f1f2),
	.w1(32'hbc771922),
	.w2(32'hbc75e4df),
	.w3(32'hbbcd79cf),
	.w4(32'h3baa9eba),
	.w5(32'h3a1c3e6b),
	.w6(32'h3a8f9b92),
	.w7(32'h3c4e48c1),
	.w8(32'h3c4034b8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9364c0),
	.w1(32'h3b5f17c1),
	.w2(32'h3b11aec7),
	.w3(32'hbc8d572d),
	.w4(32'hbb9fcaf7),
	.w5(32'hbbec5ed1),
	.w6(32'h3a390266),
	.w7(32'h3a6853b0),
	.w8(32'hbad7ce0b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bf764),
	.w1(32'h39a82048),
	.w2(32'hbb51f168),
	.w3(32'hbc368f5b),
	.w4(32'h3bb2fce0),
	.w5(32'h3c37d7ef),
	.w6(32'hbc062a68),
	.w7(32'hbc637075),
	.w8(32'h3b018f82),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ba4e5),
	.w1(32'h3c534e50),
	.w2(32'h3d102877),
	.w3(32'h3b3ea680),
	.w4(32'h3bea95af),
	.w5(32'h3c8da904),
	.w6(32'hbb7d7539),
	.w7(32'h3c41cc99),
	.w8(32'h3c7a76f8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3188a),
	.w1(32'h3c571e68),
	.w2(32'h3ce069c9),
	.w3(32'h3bea8180),
	.w4(32'h3c7691f5),
	.w5(32'h3c98fd3e),
	.w6(32'h3c3f0de4),
	.w7(32'h3c8a885b),
	.w8(32'h3cbc9967),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29bd2c),
	.w1(32'h3b4a0384),
	.w2(32'h3cb5fb39),
	.w3(32'h3bafe057),
	.w4(32'h3ba1501f),
	.w5(32'h3c912f02),
	.w6(32'h3af4c182),
	.w7(32'h3bf93719),
	.w8(32'h3bd8aac6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b7e42),
	.w1(32'hbbf5aaae),
	.w2(32'h3b507a79),
	.w3(32'hbbf6445d),
	.w4(32'hbb8585fa),
	.w5(32'h3b9a1193),
	.w6(32'hbc1de220),
	.w7(32'hbbf7ebbe),
	.w8(32'h3b40ed1b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fc0b3c),
	.w1(32'hbb2c4f03),
	.w2(32'h3bad0d18),
	.w3(32'hbb55e1d7),
	.w4(32'hbbd03bf2),
	.w5(32'hbb234a43),
	.w6(32'hbbe0e64f),
	.w7(32'h3b53b1e3),
	.w8(32'h39f1a2b9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb511ec),
	.w1(32'hbc97f8fb),
	.w2(32'hbd4467a0),
	.w3(32'h3bb6aaf1),
	.w4(32'hbc9cdf06),
	.w5(32'hbcb724dc),
	.w6(32'hba9042c0),
	.w7(32'hbc007702),
	.w8(32'hbb952d5f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd31de98),
	.w1(32'hbc4e34e9),
	.w2(32'hbc43f8dc),
	.w3(32'hbc014f17),
	.w4(32'hbb63bf3c),
	.w5(32'hbc09dab5),
	.w6(32'hbb5f5a77),
	.w7(32'h3c0fef75),
	.w8(32'h3c12ae7f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc12f57),
	.w1(32'h3c2fbefd),
	.w2(32'hb9aecb2c),
	.w3(32'hbbcbff1c),
	.w4(32'h3bdd0f61),
	.w5(32'hbba6b562),
	.w6(32'h3bc8f19c),
	.w7(32'h3b3d3c2c),
	.w8(32'h3b24aa14),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8aa49),
	.w1(32'hbb3b7486),
	.w2(32'hbb14fea5),
	.w3(32'hbb01e6f8),
	.w4(32'hbc8f113b),
	.w5(32'hbc6e0338),
	.w6(32'hbaeed33e),
	.w7(32'hbae55752),
	.w8(32'h39a2984d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393139e0),
	.w1(32'hba99dcd9),
	.w2(32'hbb61a717),
	.w3(32'hbc7e5e66),
	.w4(32'hbbca3f03),
	.w5(32'hbc021194),
	.w6(32'h3a904f52),
	.w7(32'h3b97f609),
	.w8(32'h39bb052a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0292da),
	.w1(32'hbc15182f),
	.w2(32'h3beabdae),
	.w3(32'hbb2744b4),
	.w4(32'hbb2f990d),
	.w5(32'h3b639109),
	.w6(32'hbc77ad93),
	.w7(32'hbb84724e),
	.w8(32'hbb0df676),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f3a64),
	.w1(32'hbba053d3),
	.w2(32'hbac0343d),
	.w3(32'hbba0b6b8),
	.w4(32'hba3ac807),
	.w5(32'hbc6ddd07),
	.w6(32'h3bc8c11f),
	.w7(32'h3bd502de),
	.w8(32'h3b154dac),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1361c),
	.w1(32'h3d041356),
	.w2(32'h3d892da3),
	.w3(32'hbc8d34d7),
	.w4(32'h3c916de4),
	.w5(32'h3cf0f8dc),
	.w6(32'h3d067ef4),
	.w7(32'h3d424979),
	.w8(32'h3c8c1ea3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03e501),
	.w1(32'hbb2cbdbd),
	.w2(32'hbb75f7af),
	.w3(32'h3c8c7029),
	.w4(32'h3c1c606e),
	.w5(32'h3c3736bf),
	.w6(32'h3baf9fcc),
	.w7(32'h3b4cf03c),
	.w8(32'h3c208294),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9455ae),
	.w1(32'hbd607eb5),
	.w2(32'hbdb20ae5),
	.w3(32'h3c23479f),
	.w4(32'hbce44323),
	.w5(32'hbd26b609),
	.w6(32'hbcdc2804),
	.w7(32'hbd178832),
	.w8(32'hbccb2f9c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd55cf52),
	.w1(32'hbb89491d),
	.w2(32'h39f2e914),
	.w3(32'hbca72f28),
	.w4(32'hbbd9a3da),
	.w5(32'hbb6b180a),
	.w6(32'h3ac2e0bb),
	.w7(32'h3b82d3dc),
	.w8(32'h3bab458f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18161e),
	.w1(32'h3ba4061d),
	.w2(32'h3c121d01),
	.w3(32'h3b7dcc58),
	.w4(32'h3bf871d5),
	.w5(32'h3c4f0ea7),
	.w6(32'h3afc4ef5),
	.w7(32'h3b1d75d9),
	.w8(32'hbaf0da68),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8dc9c),
	.w1(32'h3c38f237),
	.w2(32'h3c9a9977),
	.w3(32'h3bc48ba5),
	.w4(32'h3be6829e),
	.w5(32'h3c6f9ca0),
	.w6(32'h3c56e8f2),
	.w7(32'h3c68c8dd),
	.w8(32'h3c27f550),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c773c64),
	.w1(32'h3c021a05),
	.w2(32'h3bc275cf),
	.w3(32'h3c3c24ae),
	.w4(32'h3b2f2482),
	.w5(32'h3bf8e21f),
	.w6(32'h3bbe2849),
	.w7(32'h3b7ef39e),
	.w8(32'h39f3d486),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba7419),
	.w1(32'hbb626e90),
	.w2(32'hbba66d20),
	.w3(32'h3a3b65a9),
	.w4(32'hb95dc062),
	.w5(32'hbb169e1a),
	.w6(32'hbb7d9dc4),
	.w7(32'hbbf26ea1),
	.w8(32'hb9b662a8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb830ee8),
	.w1(32'hbb47515a),
	.w2(32'h3bd64c65),
	.w3(32'hbb0c6088),
	.w4(32'hbabdf20b),
	.w5(32'hbaeed1b6),
	.w6(32'hb9d9ca9a),
	.w7(32'h3c2ade01),
	.w8(32'h3b1fad92),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe9647),
	.w1(32'hbaa7d7a0),
	.w2(32'h3b37de96),
	.w3(32'hbad8cadc),
	.w4(32'hbba8d788),
	.w5(32'hbbf78fa6),
	.w6(32'h3a8a560c),
	.w7(32'h3a0751ea),
	.w8(32'hbb1ab4e6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b0585),
	.w1(32'hbbc579cc),
	.w2(32'hbc4909ad),
	.w3(32'hbb4b2847),
	.w4(32'h3b0082bc),
	.w5(32'hbc67f5d0),
	.w6(32'hbbddd15d),
	.w7(32'hbb03484d),
	.w8(32'h3b60d06a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0a6b),
	.w1(32'hbcba020f),
	.w2(32'hbd242030),
	.w3(32'hbc53547b),
	.w4(32'hbc1b6a7d),
	.w5(32'h3a170c4e),
	.w6(32'hbcb3d878),
	.w7(32'hbcd796f1),
	.w8(32'hbc9b4684),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc01b76),
	.w1(32'h3b895411),
	.w2(32'hbc01750f),
	.w3(32'h3a4633f8),
	.w4(32'h3928cb3e),
	.w5(32'hbbec8a78),
	.w6(32'h3c07e675),
	.w7(32'h3b2f6036),
	.w8(32'h3bc34e6a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d32f0),
	.w1(32'hbb92ce33),
	.w2(32'hbbf08cd7),
	.w3(32'hbba2374d),
	.w4(32'h3bc31741),
	.w5(32'h3a779108),
	.w6(32'h3a81f80c),
	.w7(32'hbc39c90d),
	.w8(32'hbbc7f76c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42c6a8),
	.w1(32'hbcd2f50c),
	.w2(32'hbd2c22bc),
	.w3(32'hbab84a41),
	.w4(32'hbc967ba6),
	.w5(32'hbbe7dee6),
	.w6(32'hbc498197),
	.w7(32'hbceb470f),
	.w8(32'hbccb79fe),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bd84d),
	.w1(32'hbc507090),
	.w2(32'hbca5c1e3),
	.w3(32'h3b7ac9a0),
	.w4(32'hbc62983d),
	.w5(32'hbaa261db),
	.w6(32'hbc0368bf),
	.w7(32'hbce29613),
	.w8(32'hbc77c88b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8894a0),
	.w1(32'h38ca9704),
	.w2(32'hbbe2b861),
	.w3(32'h3c8010bb),
	.w4(32'hbc534c02),
	.w5(32'hbca87e5d),
	.w6(32'h3c1bf990),
	.w7(32'h3b49e6e1),
	.w8(32'h3be7da7d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386e102e),
	.w1(32'hbb94bd22),
	.w2(32'hbbe37a70),
	.w3(32'hbc606396),
	.w4(32'hbb4ab011),
	.w5(32'hbaf8fe07),
	.w6(32'hbc2b7064),
	.w7(32'hbc0b884b),
	.w8(32'h3a598042),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ce29a),
	.w1(32'hbb2628c8),
	.w2(32'hbaaaf6ea),
	.w3(32'hbb81e5ae),
	.w4(32'hbb0c7093),
	.w5(32'hbbab4edb),
	.w6(32'hbbe83812),
	.w7(32'h3babd9bc),
	.w8(32'h3bf6bdc4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ec01b),
	.w1(32'hbbb93ace),
	.w2(32'hbc1c362d),
	.w3(32'hbbf7d7f0),
	.w4(32'h3afc7404),
	.w5(32'h3b1c77e3),
	.w6(32'hbaf014e8),
	.w7(32'hbc01b69b),
	.w8(32'hbb85c03f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f3945),
	.w1(32'h38fadbb7),
	.w2(32'h3bb423f5),
	.w3(32'h3b4d4c4f),
	.w4(32'h3c927ce9),
	.w5(32'hbb982be7),
	.w6(32'hbc64ec1b),
	.w7(32'hbb4e51b4),
	.w8(32'h3c80665e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0fe8f),
	.w1(32'h39b6d9eb),
	.w2(32'hbb4b1117),
	.w3(32'hbc909b6b),
	.w4(32'hbb374a21),
	.w5(32'hbc547de7),
	.w6(32'h3c268dd4),
	.w7(32'h3bfd0edd),
	.w8(32'h3bd57ca6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b195e),
	.w1(32'h3b3b9d24),
	.w2(32'h3bc08894),
	.w3(32'hbca15adf),
	.w4(32'h3bc1ab0b),
	.w5(32'h3b9e783b),
	.w6(32'hbb16d0b7),
	.w7(32'h3c291e89),
	.w8(32'h3b65e652),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1bffc),
	.w1(32'hbaa07ab4),
	.w2(32'h3bfe3b33),
	.w3(32'hbc44e8ee),
	.w4(32'hbb877e69),
	.w5(32'h3ba7701b),
	.w6(32'h3c43815b),
	.w7(32'h3c441d73),
	.w8(32'h3c17aebb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84aee7),
	.w1(32'hbbed723f),
	.w2(32'h3b8de573),
	.w3(32'h3bf57bdd),
	.w4(32'hb9f3da72),
	.w5(32'h3b8d11ad),
	.w6(32'hbb7e65d0),
	.w7(32'h3b744122),
	.w8(32'h368055e0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb622c51),
	.w1(32'hba9ed078),
	.w2(32'hbb68d098),
	.w3(32'h3a67eee7),
	.w4(32'h3a6782b4),
	.w5(32'h3b5bae67),
	.w6(32'hbade2b4d),
	.w7(32'hbaf02f5f),
	.w8(32'hbb7e4e74),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04700a),
	.w1(32'h3c8da269),
	.w2(32'h3d152137),
	.w3(32'hbabd7a36),
	.w4(32'h3b2808fd),
	.w5(32'h3c862867),
	.w6(32'h3c1e3141),
	.w7(32'h3ca40d57),
	.w8(32'h3c011d88),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca18ca5),
	.w1(32'hbbe72c81),
	.w2(32'hbc06a2ac),
	.w3(32'h3c19607e),
	.w4(32'hbc12f373),
	.w5(32'h3c606311),
	.w6(32'h3b8a0841),
	.w7(32'h3bd03e5f),
	.w8(32'hba69e6f6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e3341),
	.w1(32'h3bb3b72d),
	.w2(32'h3b94f1a6),
	.w3(32'hbba66816),
	.w4(32'h3bd4b3b2),
	.w5(32'h3af1edf1),
	.w6(32'h3bf14938),
	.w7(32'hbb07ca38),
	.w8(32'h3b6801fb),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7346f8),
	.w1(32'h3c338c1a),
	.w2(32'h3caaae53),
	.w3(32'hbb7d471c),
	.w4(32'h3b8c2b8a),
	.w5(32'h3bbec2c1),
	.w6(32'hbb305848),
	.w7(32'h3c86c4b3),
	.w8(32'h3c709eb0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44a6a1),
	.w1(32'hbbefaf6f),
	.w2(32'hbbcd69be),
	.w3(32'h3c3581b0),
	.w4(32'hbb70d7e3),
	.w5(32'hb9b88ac0),
	.w6(32'hbbd3af16),
	.w7(32'hbb8c2096),
	.w8(32'hbb9aa706),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba10554),
	.w1(32'h3b559183),
	.w2(32'h3b652610),
	.w3(32'hbaab1bfe),
	.w4(32'h3ae54c37),
	.w5(32'h3afe09b0),
	.w6(32'hbaa4d6fe),
	.w7(32'hbb34779b),
	.w8(32'hbb14142d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb271641),
	.w1(32'h3bb2abf1),
	.w2(32'h3bebd30b),
	.w3(32'hba119f72),
	.w4(32'h3bbb4ce1),
	.w5(32'h3c26cd5a),
	.w6(32'h3c12dc2c),
	.w7(32'h3b6afdab),
	.w8(32'h3c20c4e1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bdaf4),
	.w1(32'hbc92dbea),
	.w2(32'hbc1cb6c1),
	.w3(32'hba0ec1f0),
	.w4(32'hbbb291cc),
	.w5(32'h3c7e8121),
	.w6(32'h3a884c51),
	.w7(32'hbbc106e7),
	.w8(32'h3bc6355d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b514341),
	.w1(32'h3bbda203),
	.w2(32'h3bbc0c1d),
	.w3(32'h3c07e6fb),
	.w4(32'h3c6a537b),
	.w5(32'h3c2c571c),
	.w6(32'hbb2bacb7),
	.w7(32'hbb95f96e),
	.w8(32'h3b1e0d8d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9459e0),
	.w1(32'h3c9720f0),
	.w2(32'h3d36fb59),
	.w3(32'hba2a14fe),
	.w4(32'hbb1c49d2),
	.w5(32'h3c2b8726),
	.w6(32'h3cc12c93),
	.w7(32'h3ced2d94),
	.w8(32'h3c39a2e6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd54a77),
	.w1(32'h3c0738f5),
	.w2(32'h3bc8b697),
	.w3(32'hbbf6dfaf),
	.w4(32'h3b97a8f8),
	.w5(32'h3c93014e),
	.w6(32'h3c1b996f),
	.w7(32'h3b58a8b9),
	.w8(32'h3cacd33f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c912abe),
	.w1(32'h3bcce42c),
	.w2(32'h3ab7d6e0),
	.w3(32'h3ccbe4f6),
	.w4(32'h3a976fa1),
	.w5(32'hbb2f0092),
	.w6(32'h3c00d086),
	.w7(32'h3b56bdbe),
	.w8(32'hbb040f37),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a3151),
	.w1(32'hbd1aa11c),
	.w2(32'hbd6e1e12),
	.w3(32'hbc136130),
	.w4(32'hbaca91c0),
	.w5(32'hbc1a6ebb),
	.w6(32'hbd25fc70),
	.w7(32'hbd5d96d9),
	.w8(32'hbc26d5bf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb13ed6),
	.w1(32'hbd301cfe),
	.w2(32'hbd9d7db1),
	.w3(32'h3b9d941d),
	.w4(32'hbc63251d),
	.w5(32'hbcae138b),
	.w6(32'hbcf650c6),
	.w7(32'hbd5458d0),
	.w8(32'hbcccf280),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2be81e),
	.w1(32'h3bf56ac7),
	.w2(32'h3c210313),
	.w3(32'h3baa2405),
	.w4(32'hb98bdead),
	.w5(32'h3b6aca39),
	.w6(32'hbacc9dd9),
	.w7(32'h3bd62f7e),
	.w8(32'hbb8f61f4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1c7f3),
	.w1(32'hbc18b093),
	.w2(32'h39f11fbd),
	.w3(32'hbb4fbe9c),
	.w4(32'h3b6ddf9f),
	.w5(32'h3b7a39b2),
	.w6(32'hbb7fe608),
	.w7(32'hb947f104),
	.w8(32'h3b1e8d4f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd734db),
	.w1(32'h3b80f496),
	.w2(32'h3bf97247),
	.w3(32'hbaa4516d),
	.w4(32'hbb5eadc5),
	.w5(32'hba345cd7),
	.w6(32'h3c038fd0),
	.w7(32'h3c80df18),
	.w8(32'h3cb35cb1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c545b11),
	.w1(32'h3b635904),
	.w2(32'h3ad1d916),
	.w3(32'h3bbe298d),
	.w4(32'h3bd6229d),
	.w5(32'h3a05dd22),
	.w6(32'hbb4fd660),
	.w7(32'h3bc0fe65),
	.w8(32'h39c6be3f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b32b5),
	.w1(32'h3ac36863),
	.w2(32'h3b43cba0),
	.w3(32'hbc003a94),
	.w4(32'h3c28ee4b),
	.w5(32'h3afb5167),
	.w6(32'h3af7ddc9),
	.w7(32'h3c2836c0),
	.w8(32'h3bb92b7d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba978b78),
	.w1(32'hbac305a6),
	.w2(32'hbbeaa472),
	.w3(32'hbb3d135a),
	.w4(32'hbb857188),
	.w5(32'hb9180363),
	.w6(32'h3ba41064),
	.w7(32'h3bc6ac22),
	.w8(32'h3b34eb61),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab4827),
	.w1(32'h3c1be47b),
	.w2(32'h3b99b8e2),
	.w3(32'hbbc6222a),
	.w4(32'hba04b189),
	.w5(32'hbc1e65fa),
	.w6(32'hba84999f),
	.w7(32'h3c652f43),
	.w8(32'h3b27e556),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38eb7d),
	.w1(32'hbba870d3),
	.w2(32'hbc9216d3),
	.w3(32'hbc71d6be),
	.w4(32'hbb442e40),
	.w5(32'h3c00253d),
	.w6(32'hbbb5599f),
	.w7(32'hbc16eddb),
	.w8(32'h3bcc06d9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb934a9e),
	.w1(32'h3c423c95),
	.w2(32'h3d042787),
	.w3(32'h3c011550),
	.w4(32'hbb92306d),
	.w5(32'h3c0a7409),
	.w6(32'h3c90737f),
	.w7(32'h3ca50001),
	.w8(32'h3bd6b240),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde1c9b),
	.w1(32'hbbdfe64f),
	.w2(32'hbc208841),
	.w3(32'hba033e8b),
	.w4(32'h3c4213b2),
	.w5(32'h3a8dcc69),
	.w6(32'hbb79877d),
	.w7(32'hba98ba02),
	.w8(32'h3c634c0b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf47778),
	.w1(32'h3c485bcf),
	.w2(32'h3ccaf326),
	.w3(32'h3bc1d99d),
	.w4(32'h3c261792),
	.w5(32'h3cc3325f),
	.w6(32'h3b9bd557),
	.w7(32'h3c2ee322),
	.w8(32'h3c7b6fa1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b908727),
	.w1(32'hbc07b700),
	.w2(32'hbb770e85),
	.w3(32'h38ee0328),
	.w4(32'h3bb32079),
	.w5(32'h3c650820),
	.w6(32'hbb1f8c15),
	.w7(32'h3bf0aa78),
	.w8(32'h3b391325),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b141249),
	.w1(32'hbb08f9ef),
	.w2(32'hbc879c87),
	.w3(32'h3bc347ea),
	.w4(32'hbbe7c0e5),
	.w5(32'hbbd50f19),
	.w6(32'h3aae76f5),
	.w7(32'h3bccf0ec),
	.w8(32'h3aa364da),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23d5f1),
	.w1(32'h3907733f),
	.w2(32'hbab3259c),
	.w3(32'h3c71184d),
	.w4(32'hbae7f0da),
	.w5(32'hba936e79),
	.w6(32'h3a152db1),
	.w7(32'hba923d4f),
	.w8(32'h3b5f0cd5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5df86f),
	.w1(32'hba8104c9),
	.w2(32'hbb0063f3),
	.w3(32'hbb8fbadd),
	.w4(32'h3b64baf0),
	.w5(32'hbb9a210f),
	.w6(32'h3c00e481),
	.w7(32'h3b57e2a4),
	.w8(32'h3b85fccc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee6843),
	.w1(32'hbb8c2dfe),
	.w2(32'hbb5e944b),
	.w3(32'hbc1e0b79),
	.w4(32'hbbec53a8),
	.w5(32'hbb6930c0),
	.w6(32'h3b101fb7),
	.w7(32'h3a09ad6d),
	.w8(32'h3be11e97),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae75c21),
	.w1(32'h3a7d3a5d),
	.w2(32'hbbb135a7),
	.w3(32'hbaac900f),
	.w4(32'hbbad249c),
	.w5(32'h3c98317f),
	.w6(32'hbb4759ac),
	.w7(32'hbb80cc5d),
	.w8(32'h3baf0abd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf3611),
	.w1(32'hbd2329d0),
	.w2(32'hbdabe7e8),
	.w3(32'h3cb4764e),
	.w4(32'hbc45ca9c),
	.w5(32'hbd00340a),
	.w6(32'hbcf7de37),
	.w7(32'hbd4587cc),
	.w8(32'hbcb7ecfd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd413d92),
	.w1(32'h3cf0e0c6),
	.w2(32'h3d6d5aa9),
	.w3(32'hbc4b59b2),
	.w4(32'h3c4c0072),
	.w5(32'h3d1e2b56),
	.w6(32'h3ceddc00),
	.w7(32'h3d05ab62),
	.w8(32'h3c7a5626),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d205367),
	.w1(32'h3a9aaade),
	.w2(32'h3b71d60c),
	.w3(32'h3d037a9e),
	.w4(32'hba0ec6d3),
	.w5(32'hbabb5d98),
	.w6(32'h39fb8b29),
	.w7(32'h3b1acfc5),
	.w8(32'h3b66db22),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0996f),
	.w1(32'h39764de7),
	.w2(32'h3ad8e832),
	.w3(32'h39830828),
	.w4(32'h3bd83fc0),
	.w5(32'h3bde5031),
	.w6(32'h3b45ec65),
	.w7(32'h3b46c41f),
	.w8(32'h3b97196d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa966fe),
	.w1(32'h3bea0118),
	.w2(32'h3c8011f7),
	.w3(32'h3b1b4ed1),
	.w4(32'h3b239260),
	.w5(32'h3a8537e9),
	.w6(32'h3c03614a),
	.w7(32'h3be1696f),
	.w8(32'h3c639323),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba523ab),
	.w1(32'hbaf86554),
	.w2(32'hbab8e074),
	.w3(32'h3b530bbd),
	.w4(32'h3a96124d),
	.w5(32'h3b30e347),
	.w6(32'hbb8be243),
	.w7(32'hbab75c84),
	.w8(32'h3b62d69f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16624f),
	.w1(32'h3cb32cb6),
	.w2(32'h3ce096d6),
	.w3(32'h3b9fac26),
	.w4(32'h3ca8b0ef),
	.w5(32'h3c6ab790),
	.w6(32'h3c5aa76d),
	.w7(32'h3c9e411a),
	.w8(32'h3c9b54e8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdbae8c),
	.w1(32'h3be60ff2),
	.w2(32'h3bd1c4c8),
	.w3(32'h3c8068c3),
	.w4(32'h3c0707c0),
	.w5(32'h3bd29af8),
	.w6(32'h3c31eace),
	.w7(32'h3c28a46c),
	.w8(32'h3c39fe43),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c555cb9),
	.w1(32'h3bddb702),
	.w2(32'h3be5fe38),
	.w3(32'h3be64284),
	.w4(32'h3bc46af3),
	.w5(32'hbb1f504f),
	.w6(32'h3b2c6b0a),
	.w7(32'h3b832cfc),
	.w8(32'h3c68bf86),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35e8c6),
	.w1(32'hbbc3e4f6),
	.w2(32'hbbb64719),
	.w3(32'h3c35e17e),
	.w4(32'h3b5c7d3c),
	.w5(32'hb88c6d1a),
	.w6(32'h3bbed3a9),
	.w7(32'h3bf4049f),
	.w8(32'hb8f8e559),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95699b),
	.w1(32'hbb9995c1),
	.w2(32'h3b8e9474),
	.w3(32'hbbdc964d),
	.w4(32'h3bcea73c),
	.w5(32'hbb0d175b),
	.w6(32'h3b845eff),
	.w7(32'h3c8122a6),
	.w8(32'h3c778fc5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04846a),
	.w1(32'hbc4496aa),
	.w2(32'hbc8862d2),
	.w3(32'hbc30bc1c),
	.w4(32'hbc82eab7),
	.w5(32'hbc9634fe),
	.w6(32'hbc60e4ca),
	.w7(32'hbc2ec941),
	.w8(32'hbc116462),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7327f0),
	.w1(32'h3bab538e),
	.w2(32'h3bc4282c),
	.w3(32'hbc53a143),
	.w4(32'h3abc5486),
	.w5(32'h3c58f3e5),
	.w6(32'h3b9976e2),
	.w7(32'h39b53388),
	.w8(32'h3c315f1b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b61641),
	.w1(32'hbbc3e53c),
	.w2(32'h3c603e02),
	.w3(32'h3be76f87),
	.w4(32'h3b2a9167),
	.w5(32'h3c8b5871),
	.w6(32'hb9cd1c33),
	.w7(32'hbc2cbf51),
	.w8(32'h3bc77b95),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dc5c0),
	.w1(32'hbbdf63d8),
	.w2(32'hbc845889),
	.w3(32'hba26f91c),
	.w4(32'hbc7a3b0a),
	.w5(32'hbc8a395f),
	.w6(32'h3a9c32dd),
	.w7(32'hbb167f0d),
	.w8(32'h3ae8aede),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc236298),
	.w1(32'h3a93ffcb),
	.w2(32'hbc310c12),
	.w3(32'hbbf78ae0),
	.w4(32'h3b6a82b3),
	.w5(32'hbbd34bd9),
	.w6(32'hba3fc849),
	.w7(32'hbc050469),
	.w8(32'hba038526),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a046511),
	.w1(32'hbbe1c804),
	.w2(32'hbc24ff59),
	.w3(32'h39bbcbeb),
	.w4(32'hbb650e4d),
	.w5(32'h3ba504ab),
	.w6(32'h394832cf),
	.w7(32'hbbbc0292),
	.w8(32'hba8630ae),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d46e0),
	.w1(32'hbbc71515),
	.w2(32'hbb8b89cd),
	.w3(32'h3c333dc5),
	.w4(32'hbb3402a3),
	.w5(32'h3a8575b5),
	.w6(32'hbaa1d799),
	.w7(32'hbbc386b4),
	.w8(32'hbc4804de),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb0e8f),
	.w1(32'hbbf9913b),
	.w2(32'hbc3f66d2),
	.w3(32'h3b55f3f9),
	.w4(32'hbbf0b064),
	.w5(32'hbc16da66),
	.w6(32'hbc28d5da),
	.w7(32'hbc15ce0c),
	.w8(32'hbc52127a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e36ff),
	.w1(32'h39377282),
	.w2(32'h3b6a2741),
	.w3(32'hbc1b2197),
	.w4(32'h3bbbc854),
	.w5(32'h3c135f16),
	.w6(32'h3a98afe7),
	.w7(32'h3aecd72c),
	.w8(32'h3b2264e3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9909f76),
	.w1(32'hbca1fd49),
	.w2(32'hbcad0d9a),
	.w3(32'h3bc09fcf),
	.w4(32'hbb7dee34),
	.w5(32'h3bd0707c),
	.w6(32'hbc2053d4),
	.w7(32'hbc85839f),
	.w8(32'h393f72f1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a03cb),
	.w1(32'hbb437d77),
	.w2(32'hbbc2eef2),
	.w3(32'hbb8330e7),
	.w4(32'hbbf957d1),
	.w5(32'hbc1e9ac0),
	.w6(32'hb8db2d39),
	.w7(32'hbb735925),
	.w8(32'hbb5b12ae),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0de496),
	.w1(32'hbbeca7d4),
	.w2(32'hbc24e012),
	.w3(32'hbc44102a),
	.w4(32'hbbd46a08),
	.w5(32'h3b06c0bd),
	.w6(32'hbb9a5aff),
	.w7(32'h3b753268),
	.w8(32'hbc2fa79b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f8fb9),
	.w1(32'hbb88f383),
	.w2(32'hbb0aa212),
	.w3(32'hbbe762df),
	.w4(32'h3bed173f),
	.w5(32'hb8fb400a),
	.w6(32'hbc9ab3e0),
	.w7(32'hbcbffcc1),
	.w8(32'h3b95acb9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e6ec1),
	.w1(32'hbbc9464d),
	.w2(32'hbbd6f443),
	.w3(32'hb8e90882),
	.w4(32'hbc1585ea),
	.w5(32'hbc19dd65),
	.w6(32'hbb425329),
	.w7(32'hbb3afbbf),
	.w8(32'hbb625b14),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9c0e2),
	.w1(32'h3aac419f),
	.w2(32'h3b7a1fe2),
	.w3(32'hbb7ee337),
	.w4(32'h3b6c55cf),
	.w5(32'h3bb66fec),
	.w6(32'h395061e2),
	.w7(32'h3a841927),
	.w8(32'h3b0fa89a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5caae4),
	.w1(32'h3acc5134),
	.w2(32'h3ba49b6b),
	.w3(32'h3b83cead),
	.w4(32'h3c0a702a),
	.w5(32'h3b4fd1be),
	.w6(32'h3c15f862),
	.w7(32'h3bf67ca9),
	.w8(32'h3c122ed7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92447d),
	.w1(32'hbb8557e0),
	.w2(32'h3b9f4893),
	.w3(32'h3b9e6c51),
	.w4(32'hbc032b9c),
	.w5(32'h3b01a78e),
	.w6(32'hbb90c088),
	.w7(32'h3b84dabc),
	.w8(32'hbb39ebac),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9830c6),
	.w1(32'h3bce7b43),
	.w2(32'h3c9877db),
	.w3(32'hbbb325ac),
	.w4(32'h3b9fef10),
	.w5(32'h3b93be95),
	.w6(32'h3c29c9ba),
	.w7(32'h3bf5de94),
	.w8(32'h3bc359f5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68b74d),
	.w1(32'hbb84f6f5),
	.w2(32'h39ab8c04),
	.w3(32'h3b006fd9),
	.w4(32'h3b8738ff),
	.w5(32'h3bbfa14e),
	.w6(32'hbadc38c5),
	.w7(32'h39e2eff8),
	.w8(32'h3a77d162),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c67eb),
	.w1(32'h3c79478b),
	.w2(32'h3d35b563),
	.w3(32'hb98ea484),
	.w4(32'hbb838fb9),
	.w5(32'h3c038f20),
	.w6(32'h3c3d6e9d),
	.w7(32'h3d035060),
	.w8(32'h3b34c479),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb57ca6),
	.w1(32'hbb132845),
	.w2(32'hbb491401),
	.w3(32'h3ac80b68),
	.w4(32'h3bc35b88),
	.w5(32'h3bb4f2f3),
	.w6(32'h3c13d960),
	.w7(32'hbbbeca4c),
	.w8(32'hbb4710ec),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00fe95),
	.w1(32'hbc10073c),
	.w2(32'hbc3d1730),
	.w3(32'hbab609f0),
	.w4(32'hbb1e23cc),
	.w5(32'hbb6f337b),
	.w6(32'hbb06770d),
	.w7(32'hbb83aa55),
	.w8(32'hba51b16b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12ec2c),
	.w1(32'hbc80af36),
	.w2(32'hbbf956b2),
	.w3(32'hbb04a29b),
	.w4(32'hbc3906e4),
	.w5(32'hbb5622a7),
	.w6(32'hbc38db5b),
	.w7(32'hbba2b8fe),
	.w8(32'hbbb77d27),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce72a9),
	.w1(32'h3bc8c7d8),
	.w2(32'h3ca38497),
	.w3(32'hbbb1b632),
	.w4(32'h3c8361b5),
	.w5(32'h3c94fe18),
	.w6(32'hbbb5d4ae),
	.w7(32'h3b2d7c2d),
	.w8(32'h3c45bd55),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67c8fd),
	.w1(32'hbc7a8ee7),
	.w2(32'hbc9b7115),
	.w3(32'h3b742cfb),
	.w4(32'hbca132ab),
	.w5(32'hbbea0975),
	.w6(32'hbc226c8c),
	.w7(32'hbc74a5bf),
	.w8(32'hbc66ff62),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1445a),
	.w1(32'hbaaae72b),
	.w2(32'hbb3822ae),
	.w3(32'hb9e49953),
	.w4(32'hba31a419),
	.w5(32'hbb115365),
	.w6(32'hbb1460c3),
	.w7(32'hbb4802ca),
	.w8(32'hba26b4da),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eaded),
	.w1(32'h3b3fdc4b),
	.w2(32'h3b502c6c),
	.w3(32'hbad339e9),
	.w4(32'h386780d2),
	.w5(32'hbb06a92f),
	.w6(32'h3a27c625),
	.w7(32'h3b23edbd),
	.w8(32'hbb5abed1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule