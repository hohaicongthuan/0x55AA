module layer_10_featuremap_202(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e4e37),
	.w1(32'hbb0e3462),
	.w2(32'hbb85b566),
	.w3(32'hba1ee514),
	.w4(32'hb9604465),
	.w5(32'hba775b14),
	.w6(32'hbad08bbe),
	.w7(32'hbb03510b),
	.w8(32'hba70bcdd),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb293588),
	.w1(32'h39ac3c8e),
	.w2(32'h3a0b630d),
	.w3(32'hbb030492),
	.w4(32'h3989e96b),
	.w5(32'h39b400b7),
	.w6(32'h397c8e97),
	.w7(32'h39db0006),
	.w8(32'h38dfcabe),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0ad0c),
	.w1(32'hbab3869f),
	.w2(32'hba69af9c),
	.w3(32'h39796c53),
	.w4(32'hb9c55688),
	.w5(32'h3961ed55),
	.w6(32'hbab607e8),
	.w7(32'hba6c98c0),
	.w8(32'hba2a44fa),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9356b82),
	.w1(32'hb973de31),
	.w2(32'h3af5461c),
	.w3(32'h3a16e90d),
	.w4(32'hb9a88cf8),
	.w5(32'hba704a27),
	.w6(32'hbac56a26),
	.w7(32'hbaff2785),
	.w8(32'hbb30f557),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0dd58),
	.w1(32'hba1bc7cc),
	.w2(32'h3a313528),
	.w3(32'hb8c126ac),
	.w4(32'hba2165eb),
	.w5(32'hb97fed9e),
	.w6(32'h3a04a25a),
	.w7(32'h3972c761),
	.w8(32'h38fde8a1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92fc2a9),
	.w1(32'h39193bb7),
	.w2(32'h3ab878bd),
	.w3(32'hba7038de),
	.w4(32'h3a4341df),
	.w5(32'h3a58c73a),
	.w6(32'h39b49c95),
	.w7(32'h3a02887d),
	.w8(32'hba1cc36c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3920b024),
	.w1(32'hb9fbbcff),
	.w2(32'h39356726),
	.w3(32'h39545e04),
	.w4(32'hba009d09),
	.w5(32'hb9552f4b),
	.w6(32'hb98a2086),
	.w7(32'h37d636e2),
	.w8(32'h39d62e23),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38700b4e),
	.w1(32'h39049e7f),
	.w2(32'h3a44c5ef),
	.w3(32'h39ef6891),
	.w4(32'h39bcf410),
	.w5(32'hb7d8611d),
	.w6(32'h38b026e1),
	.w7(32'h39a0e2a6),
	.w8(32'h39daaca3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef91ca),
	.w1(32'hba132a39),
	.w2(32'hba1ed796),
	.w3(32'h38a8d7cd),
	.w4(32'hba6093b7),
	.w5(32'hbaaa05ef),
	.w6(32'hba374097),
	.w7(32'hba24c553),
	.w8(32'hb9a0e15c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b0444),
	.w1(32'hbaaffd80),
	.w2(32'hb9dd5241),
	.w3(32'hba980fcf),
	.w4(32'hba9080b5),
	.w5(32'hba5ce209),
	.w6(32'hbac689ca),
	.w7(32'hbac1b978),
	.w8(32'hb929542a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02527d),
	.w1(32'hbb3741e1),
	.w2(32'hbb045ef6),
	.w3(32'h38b03a85),
	.w4(32'hba4af08c),
	.w5(32'hb9dd3387),
	.w6(32'hbad51091),
	.w7(32'hbb0d411d),
	.w8(32'hbac4fa30),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9efb3df),
	.w1(32'hbb020afe),
	.w2(32'hba05b510),
	.w3(32'h39693d9b),
	.w4(32'hbb0718c8),
	.w5(32'hbadb43d7),
	.w6(32'hba1e390c),
	.w7(32'h39d70ba3),
	.w8(32'hb95545fc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aa0e6e),
	.w1(32'hba7032d6),
	.w2(32'hb9db294e),
	.w3(32'hbab2caa9),
	.w4(32'hba28005f),
	.w5(32'hba11a138),
	.w6(32'hba61c84b),
	.w7(32'hba0173ee),
	.w8(32'hba3d7e56),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dd406),
	.w1(32'h3996a427),
	.w2(32'h3a12a224),
	.w3(32'hba1f178e),
	.w4(32'hb7609fdc),
	.w5(32'hb992bf50),
	.w6(32'hb98d08ac),
	.w7(32'h39a0e132),
	.w8(32'h3a06fa2c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a245ff4),
	.w1(32'hbb514619),
	.w2(32'hba68bf7c),
	.w3(32'hba216497),
	.w4(32'hbb39d659),
	.w5(32'hbb253654),
	.w6(32'hba5dec10),
	.w7(32'hba552704),
	.w8(32'hb7cd2dc5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0543a2),
	.w1(32'hb87dcebb),
	.w2(32'h3967ae15),
	.w3(32'hbb0d25bb),
	.w4(32'hba403189),
	.w5(32'hba105b0f),
	.w6(32'hb933be7d),
	.w7(32'hb95e7906),
	.w8(32'hb8310ab6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9991c2d),
	.w1(32'h3a3e83a0),
	.w2(32'h3a8b4170),
	.w3(32'hba54f327),
	.w4(32'h3b804f52),
	.w5(32'h3b9b4e07),
	.w6(32'h3a817fca),
	.w7(32'h3b028f6f),
	.w8(32'hba8bf4a1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b200e),
	.w1(32'hb9e6535a),
	.w2(32'h3913fea1),
	.w3(32'h3abba0a6),
	.w4(32'hba1bcc55),
	.w5(32'hb94b34aa),
	.w6(32'hba0ebf78),
	.w7(32'hba37448a),
	.w8(32'hb869d42b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99310f9),
	.w1(32'hba3fd67a),
	.w2(32'h39403c8f),
	.w3(32'h39c9f819),
	.w4(32'hba2c1b16),
	.w5(32'hb82a3a35),
	.w6(32'hba28d9d2),
	.w7(32'hb8b62b2e),
	.w8(32'h3a7d4f68),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aae6a8),
	.w1(32'hba602788),
	.w2(32'hb9dd462b),
	.w3(32'h38829392),
	.w4(32'hba8728b0),
	.w5(32'hba71a775),
	.w6(32'hba5298f5),
	.w7(32'hba4e78d2),
	.w8(32'hba9e3659),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a84e9),
	.w1(32'hb9175e62),
	.w2(32'h3ae6f84e),
	.w3(32'hba95c3db),
	.w4(32'hb9f81aba),
	.w5(32'hb87bcd38),
	.w6(32'h39b13499),
	.w7(32'h3a91812c),
	.w8(32'hba28f056),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e848f7),
	.w1(32'hbb9fbaca),
	.w2(32'hbb9cfb2d),
	.w3(32'hba543160),
	.w4(32'hbadfd66f),
	.w5(32'hb8b9e6cf),
	.w6(32'hbb901b91),
	.w7(32'hbb9769a5),
	.w8(32'hbb5429d3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2bff0),
	.w1(32'h3b773bfe),
	.w2(32'h3ba7494d),
	.w3(32'hb7c172e8),
	.w4(32'h3a9de88e),
	.w5(32'h3afcbb7f),
	.w6(32'hba0803de),
	.w7(32'h3987e6e7),
	.w8(32'hbb1edf33),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d94a5),
	.w1(32'h38ef82b4),
	.w2(32'h3a097fa4),
	.w3(32'h39e215a5),
	.w4(32'hb99042c8),
	.w5(32'hb91aabac),
	.w6(32'hb8a01c56),
	.w7(32'h39173cd1),
	.w8(32'h39d7f430),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2a3c8),
	.w1(32'h3a83c834),
	.w2(32'h3a6da6de),
	.w3(32'hb950395c),
	.w4(32'h3a567fa4),
	.w5(32'h38fc1898),
	.w6(32'hb8bfb356),
	.w7(32'hb9c71fbf),
	.w8(32'hba992383),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c79010),
	.w1(32'hb9ef40dc),
	.w2(32'hba54ee6e),
	.w3(32'hba069791),
	.w4(32'h3b1ee6ce),
	.w5(32'h3ad367da),
	.w6(32'hba3b4806),
	.w7(32'hba684797),
	.w8(32'hbac5f5d3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90858c1),
	.w1(32'hba973d7f),
	.w2(32'hba226795),
	.w3(32'h3aef55f0),
	.w4(32'hba977a1c),
	.w5(32'hba7e8d15),
	.w6(32'hba411377),
	.w7(32'hba2b1c74),
	.w8(32'hba9d4899),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bc472),
	.w1(32'hbabef8ce),
	.w2(32'hbaa2a5d7),
	.w3(32'hba6218e4),
	.w4(32'hbad8023e),
	.w5(32'hbae2c68b),
	.w6(32'hba8a0b42),
	.w7(32'hbac5e435),
	.w8(32'hbabd17c8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc65ad),
	.w1(32'h3addbe06),
	.w2(32'h3af54434),
	.w3(32'hba7f6ee8),
	.w4(32'h3b5e3c80),
	.w5(32'h3b363a3c),
	.w6(32'h3a2fc647),
	.w7(32'h3a6994eb),
	.w8(32'hb9ae54a0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a509c86),
	.w1(32'h3b80eb97),
	.w2(32'h3b4f642b),
	.w3(32'h3ae09173),
	.w4(32'h3bbc9b5c),
	.w5(32'h3b9323f6),
	.w6(32'h3b58553c),
	.w7(32'h3b54f861),
	.w8(32'h3a84f90e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b095626),
	.w1(32'hba4f7f1f),
	.w2(32'h393fe112),
	.w3(32'h3b3fa409),
	.w4(32'hba67fb10),
	.w5(32'hba111378),
	.w6(32'hb721c0b8),
	.w7(32'h39d9fdc0),
	.w8(32'hb9d9703b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27ac1e),
	.w1(32'hba86d21d),
	.w2(32'hb905e470),
	.w3(32'hba4dd4e2),
	.w4(32'hba2d4741),
	.w5(32'hb9bb2645),
	.w6(32'hba3788b4),
	.w7(32'hb9ee24a5),
	.w8(32'hbaaa1c85),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba719607),
	.w1(32'hbb328f1d),
	.w2(32'hbb03dde1),
	.w3(32'hba5f7803),
	.w4(32'hbb61b5a5),
	.w5(32'hbb2b6759),
	.w6(32'hbb3e384f),
	.w7(32'hbae85bb3),
	.w8(32'hbadccc85),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b1e2f),
	.w1(32'hba772be6),
	.w2(32'hba97f0d7),
	.w3(32'hbb21f7e2),
	.w4(32'hba8308dc),
	.w5(32'hbadba70d),
	.w6(32'hba6232bc),
	.w7(32'hb9ef8ccd),
	.w8(32'h38a040d6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d97b2a),
	.w1(32'hbb0d579e),
	.w2(32'hbab8ff12),
	.w3(32'hb8ece267),
	.w4(32'hbb04084e),
	.w5(32'hbad1872b),
	.w6(32'hbae3e5e4),
	.w7(32'hbadb6de4),
	.w8(32'hbaa9417a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba895226),
	.w1(32'hba86bc08),
	.w2(32'h390f06f2),
	.w3(32'hbabeb341),
	.w4(32'hba4c5ae0),
	.w5(32'hb9fe1b31),
	.w6(32'hba4e465c),
	.w7(32'hb8db7642),
	.w8(32'hba839753),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba362504),
	.w1(32'hba20b81a),
	.w2(32'h3a6d55d4),
	.w3(32'hbac6b2cd),
	.w4(32'hba106c1e),
	.w5(32'h37f1b6fe),
	.w6(32'h38c7a041),
	.w7(32'h3943b67d),
	.w8(32'h39a7ffe2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9df106),
	.w1(32'h390619c5),
	.w2(32'h351620cd),
	.w3(32'h3a9dcad2),
	.w4(32'h39fd5cb1),
	.w5(32'h3a137d9c),
	.w6(32'h3a46eef8),
	.w7(32'h39dfa676),
	.w8(32'hba135368),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932a6c8),
	.w1(32'hba053b78),
	.w2(32'hb9aa218f),
	.w3(32'h3a0120b7),
	.w4(32'hba03edc5),
	.w5(32'hba5892dc),
	.w6(32'h39fb4112),
	.w7(32'h3975e71e),
	.w8(32'hba02dd4e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb958c597),
	.w1(32'h3982ab74),
	.w2(32'h3a3b2ed8),
	.w3(32'hba13dabf),
	.w4(32'hb8678f55),
	.w5(32'h395e31f2),
	.w6(32'h39c07170),
	.w7(32'h3a24f746),
	.w8(32'h3a40d7ca),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56a689),
	.w1(32'h3b854344),
	.w2(32'h3b9aecc6),
	.w3(32'h3a0b5076),
	.w4(32'h3bc3b51c),
	.w5(32'h3bc7f643),
	.w6(32'h3afbf80a),
	.w7(32'h3b9010ec),
	.w8(32'h3abb00a9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f9f88),
	.w1(32'hba93a5a7),
	.w2(32'hba4d3066),
	.w3(32'h3b737490),
	.w4(32'hbad8df53),
	.w5(32'hbabf87ee),
	.w6(32'hba469c06),
	.w7(32'hb7cc2a68),
	.w8(32'h3a13503e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39587e06),
	.w1(32'hba467572),
	.w2(32'hb9ab433e),
	.w3(32'hb996fc1b),
	.w4(32'hb96f7a9e),
	.w5(32'hb9a40587),
	.w6(32'hba751096),
	.w7(32'hba74dbe7),
	.w8(32'hbae24d10),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9964c0),
	.w1(32'hb9aff714),
	.w2(32'h39a0269d),
	.w3(32'hba8adefd),
	.w4(32'h3805ed8d),
	.w5(32'h395c951e),
	.w6(32'h379272f7),
	.w7(32'hba059884),
	.w8(32'h3ad32103),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22e32e),
	.w1(32'hba953983),
	.w2(32'hbad83813),
	.w3(32'h3ae215d6),
	.w4(32'hbaf22e4d),
	.w5(32'hba945581),
	.w6(32'hbad6fdbc),
	.w7(32'hbb1d2a1b),
	.w8(32'hba786cf3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba751cf6),
	.w1(32'hbadfd071),
	.w2(32'hbac78470),
	.w3(32'hba5307ef),
	.w4(32'hbb24fb62),
	.w5(32'hbb06cbfb),
	.w6(32'hbadcbcfa),
	.w7(32'hbac16197),
	.w8(32'hb99402ee),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa86c6d),
	.w1(32'hba1de8b6),
	.w2(32'h3ab9ad86),
	.w3(32'hbaa14c6a),
	.w4(32'hbacffd2e),
	.w5(32'hbaaa13f5),
	.w6(32'h395dccac),
	.w7(32'h3a754df3),
	.w8(32'h3ad9e85a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ec391),
	.w1(32'h3b013577),
	.w2(32'hb9c6a240),
	.w3(32'h395d97ef),
	.w4(32'h3ba165d3),
	.w5(32'h3b1b504c),
	.w6(32'h398ab83d),
	.w7(32'hbaa0d187),
	.w8(32'hba28f4cd),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a206bec),
	.w1(32'hba889d6f),
	.w2(32'hb90f5d24),
	.w3(32'h3b5e49fa),
	.w4(32'hb9a537c1),
	.w5(32'h38a00480),
	.w6(32'hbaa249b9),
	.w7(32'hba6edc2b),
	.w8(32'hbae97466),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba910293),
	.w1(32'h39d74f70),
	.w2(32'h3a178b0e),
	.w3(32'hba365a82),
	.w4(32'hb8f3b8c2),
	.w5(32'hb888dc52),
	.w6(32'h39d7f9ca),
	.w7(32'h3a53a036),
	.w8(32'h3a81af14),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46f0a0),
	.w1(32'hb9edec58),
	.w2(32'hb917f625),
	.w3(32'h39058659),
	.w4(32'hba2cb19f),
	.w5(32'hba21470c),
	.w6(32'hb91a0946),
	.w7(32'h39a2a9c5),
	.w8(32'h3a924d26),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71fd56),
	.w1(32'hba7e6785),
	.w2(32'hba9ca529),
	.w3(32'hb90aa049),
	.w4(32'hbb4d7661),
	.w5(32'hbb8ecb9e),
	.w6(32'hbb167340),
	.w7(32'hbacf50eb),
	.w8(32'hbaf59d75),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c4562),
	.w1(32'h3a85bb8b),
	.w2(32'h3b025f14),
	.w3(32'hbb4c684e),
	.w4(32'h3aaa970c),
	.w5(32'h3a7eb9bc),
	.w6(32'h3a46ddf4),
	.w7(32'h3a5469b3),
	.w8(32'hb9788e04),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab98074),
	.w1(32'h3977fce9),
	.w2(32'h3aaad037),
	.w3(32'h3a8ea157),
	.w4(32'h394957e0),
	.w5(32'h39220069),
	.w6(32'h39fd75a4),
	.w7(32'h3a3c6cbd),
	.w8(32'hb8fa2c64),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9072e1),
	.w1(32'h3a00f2b5),
	.w2(32'h3ac1154f),
	.w3(32'hba249aa1),
	.w4(32'h3ab86b5e),
	.w5(32'h3aee993b),
	.w6(32'hb971c0b8),
	.w7(32'h39c77e9e),
	.w8(32'hba9b511b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38646416),
	.w1(32'h3b9357a5),
	.w2(32'h3b8e5394),
	.w3(32'h39ae5f1c),
	.w4(32'h3b5855bd),
	.w5(32'h3b175f5c),
	.w6(32'h3b2b825d),
	.w7(32'h3b58aea3),
	.w8(32'h39a479e5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b014a93),
	.w1(32'h3a5a79c9),
	.w2(32'h39d3f14f),
	.w3(32'hba0e90cc),
	.w4(32'h3a91458f),
	.w5(32'h39388a4c),
	.w6(32'hb9e2fab5),
	.w7(32'hba0a0496),
	.w8(32'hbaa00e1b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dade8f),
	.w1(32'hbb0e88bf),
	.w2(32'hbaad803c),
	.w3(32'hb9cfcf60),
	.w4(32'hbb0477c2),
	.w5(32'hbb28f970),
	.w6(32'hba78bad4),
	.w7(32'hba81bc6f),
	.w8(32'hba4d9e3b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e7ab2),
	.w1(32'hb9a49cf6),
	.w2(32'hb9b83b4d),
	.w3(32'hbb165d35),
	.w4(32'hb97b0798),
	.w5(32'hb99108b3),
	.w6(32'hb8e6e34f),
	.w7(32'hb9a8ca70),
	.w8(32'hb9d47849),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9acd441),
	.w1(32'hba3adbb4),
	.w2(32'hb9eb1b98),
	.w3(32'h385633b8),
	.w4(32'hba301d51),
	.w5(32'hba3bf477),
	.w6(32'hb9fd3367),
	.w7(32'hb98ea9b1),
	.w8(32'hb98d290a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba073d44),
	.w1(32'hb7a3b54b),
	.w2(32'h3a21fa7a),
	.w3(32'hba64d934),
	.w4(32'h38ecf840),
	.w5(32'h39ac750c),
	.w6(32'hb91e246b),
	.w7(32'h39b88a5c),
	.w8(32'h3a4f5b61),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09f1d0),
	.w1(32'hba51949c),
	.w2(32'hba0eb682),
	.w3(32'h3a14fa90),
	.w4(32'hba354b59),
	.w5(32'hba0c6a99),
	.w6(32'hb8ce6bb0),
	.w7(32'h37ca7285),
	.w8(32'h3a0c02fe),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea68ad),
	.w1(32'hbb273cd2),
	.w2(32'hbb7cb0ff),
	.w3(32'hb995e701),
	.w4(32'hbb39074b),
	.w5(32'hbb53dcd0),
	.w6(32'hbb7d3ebf),
	.w7(32'hbb603eaf),
	.w8(32'hbb3fb5df),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89b5a0),
	.w1(32'hba210fff),
	.w2(32'hb99cc04e),
	.w3(32'hbb4992d0),
	.w4(32'hb91ab0c7),
	.w5(32'hb96a65e4),
	.w6(32'hb8f69284),
	.w7(32'hb9aa1bbf),
	.w8(32'h3a111168),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9947a9),
	.w1(32'hba9bda00),
	.w2(32'hba208f74),
	.w3(32'h3a83e3ec),
	.w4(32'hba88422a),
	.w5(32'hba884347),
	.w6(32'hba83c5eb),
	.w7(32'hba398ebb),
	.w8(32'hb983ac8e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f88f32),
	.w1(32'hba9ed2e1),
	.w2(32'h38939b87),
	.w3(32'hba20ed23),
	.w4(32'hba34fb67),
	.w5(32'hbaafcfe1),
	.w6(32'hbac7a7e7),
	.w7(32'hba7c8f23),
	.w8(32'hbab20bc8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0790e5),
	.w1(32'h3aac10c1),
	.w2(32'h3b01c6fa),
	.w3(32'hbaacf733),
	.w4(32'h3b1b9f6e),
	.w5(32'h3b0fc7b4),
	.w6(32'h3b21832e),
	.w7(32'h3b3e1029),
	.w8(32'h3ae422fc),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5818f),
	.w1(32'h3bb5eaaa),
	.w2(32'h3bd67b81),
	.w3(32'h393adcee),
	.w4(32'h3bd6ed1b),
	.w5(32'h3bc99bb8),
	.w6(32'h39d64366),
	.w7(32'h3b1edf03),
	.w8(32'hb965a6ee),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd069ec),
	.w1(32'hba10ce54),
	.w2(32'h3a041ca3),
	.w3(32'h3ba1c0dc),
	.w4(32'hba8051b0),
	.w5(32'hb9d19d40),
	.w6(32'hb8e9b49c),
	.w7(32'h394d63c9),
	.w8(32'hb996a2e4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b98f7f),
	.w1(32'hbb274e4a),
	.w2(32'hbacceb48),
	.w3(32'hba1c4bc7),
	.w4(32'hbb15bdca),
	.w5(32'hbb350828),
	.w6(32'hbac1e33e),
	.w7(32'hba745fef),
	.w8(32'h38c89c14),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7952c7),
	.w1(32'hba4237d7),
	.w2(32'hba2a1cf2),
	.w3(32'hbad6e6f1),
	.w4(32'hba47cae8),
	.w5(32'hba325a62),
	.w6(32'hba2e6854),
	.w7(32'hba50a13f),
	.w8(32'hba66bead),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d9d07),
	.w1(32'hba32f21c),
	.w2(32'hb824617e),
	.w3(32'hb9dfd26f),
	.w4(32'hba2f6386),
	.w5(32'hba0121a9),
	.w6(32'hb9be5337),
	.w7(32'hb81ce0f1),
	.w8(32'hb9dc2109),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27fb16),
	.w1(32'hb9ebb8ab),
	.w2(32'hb902d958),
	.w3(32'hba672de5),
	.w4(32'hba192eb1),
	.w5(32'hba232e11),
	.w6(32'hb9cd335a),
	.w7(32'hb979ed03),
	.w8(32'hb98be2ab),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6c334),
	.w1(32'hba8b335f),
	.w2(32'h3899423b),
	.w3(32'hba56265d),
	.w4(32'hba27c04f),
	.w5(32'hb98ef6da),
	.w6(32'hba6cad54),
	.w7(32'hb974dfab),
	.w8(32'hbade0ea0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d79ac),
	.w1(32'h3a051b05),
	.w2(32'h3a2eeb54),
	.w3(32'hba87d0a4),
	.w4(32'hb8d0fd5e),
	.w5(32'h36cada11),
	.w6(32'h3989075b),
	.w7(32'h39867c79),
	.w8(32'h3a32622d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2afa23),
	.w1(32'hba5ad1e5),
	.w2(32'hba5ae681),
	.w3(32'h3a37de0c),
	.w4(32'hbb29a657),
	.w5(32'hbb645535),
	.w6(32'hbb06efb1),
	.w7(32'h393a9ad5),
	.w8(32'hb9dabaa5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad94d08),
	.w1(32'hb87c3775),
	.w2(32'h3a77ac59),
	.w3(32'hbb2a031d),
	.w4(32'hb8d12776),
	.w5(32'h399ef3de),
	.w6(32'h3918e391),
	.w7(32'h39d75cac),
	.w8(32'h3a5f6f57),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d8251),
	.w1(32'hba565789),
	.w2(32'hb9e48d8e),
	.w3(32'h392cae26),
	.w4(32'hba4e591b),
	.w5(32'hba03d1cd),
	.w6(32'hba925849),
	.w7(32'hba2912d8),
	.w8(32'hb8996f00),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cef83e),
	.w1(32'h3a6ae688),
	.w2(32'h3adde33a),
	.w3(32'h39891bfd),
	.w4(32'h3b678d6d),
	.w5(32'h3b7834e8),
	.w6(32'hba239bc3),
	.w7(32'h3a017dc7),
	.w8(32'hbab86275),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4efd7c),
	.w1(32'hba8dbb31),
	.w2(32'h3a2bf152),
	.w3(32'h3aa3553e),
	.w4(32'hbaa92e5d),
	.w5(32'hba5b521a),
	.w6(32'h38538cf7),
	.w7(32'h39ddf4b8),
	.w8(32'hba3a8bef),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73bd03),
	.w1(32'h3b9e9391),
	.w2(32'h3bb985ac),
	.w3(32'hbabff8c5),
	.w4(32'h3b8dba66),
	.w5(32'h3b83ec73),
	.w6(32'h3ad03e4a),
	.w7(32'h3b3e16fc),
	.w8(32'h3ab1f821),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdc246),
	.w1(32'hb9ccf2f6),
	.w2(32'h398b6bd2),
	.w3(32'h3b38e897),
	.w4(32'hb9e80472),
	.w5(32'hb92038de),
	.w6(32'h398fd27b),
	.w7(32'h3a132feb),
	.w8(32'h3a8df3bd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a127014),
	.w1(32'h3a9c8d44),
	.w2(32'h3a0fef69),
	.w3(32'h39827df8),
	.w4(32'h3aa6ed35),
	.w5(32'h3a0b7fe8),
	.w6(32'h38e4bdfa),
	.w7(32'hb9881ff6),
	.w8(32'hba927cbd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbf969),
	.w1(32'h39a18250),
	.w2(32'h39973cf8),
	.w3(32'hb8a69b1e),
	.w4(32'h39e11a12),
	.w5(32'h3a0c8520),
	.w6(32'h399a7b77),
	.w7(32'h3914c070),
	.w8(32'h39a0fe8a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b681cc),
	.w1(32'h39b44b4e),
	.w2(32'hba0135de),
	.w3(32'h3a271417),
	.w4(32'h3b595d88),
	.w5(32'h3b271118),
	.w6(32'hb88c1620),
	.w7(32'hba54c187),
	.w8(32'hbb25b9b3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dabd7),
	.w1(32'h3ae92a74),
	.w2(32'h3b042579),
	.w3(32'h3ae4652d),
	.w4(32'h3ab71973),
	.w5(32'h3ac35865),
	.w6(32'h3b0b41c7),
	.w7(32'h3b18fb59),
	.w8(32'h3ab59486),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f1b9c),
	.w1(32'hba170046),
	.w2(32'hbaf1f59a),
	.w3(32'h39da0777),
	.w4(32'hba871ddf),
	.w5(32'hbb1c184d),
	.w6(32'hbaa68b8d),
	.w7(32'hba9327d9),
	.w8(32'hba83f023),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd0d89),
	.w1(32'hba6fd78a),
	.w2(32'h388ced5b),
	.w3(32'hbaeb367b),
	.w4(32'hba804777),
	.w5(32'hba1d3ca1),
	.w6(32'hb8b7dd07),
	.w7(32'h398bb2e2),
	.w8(32'hba222e83),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969308a),
	.w1(32'h39f92e0b),
	.w2(32'h3ab718ae),
	.w3(32'hba765121),
	.w4(32'h3a91c4b1),
	.w5(32'h3aad2baa),
	.w6(32'hba357a34),
	.w7(32'h377df6b3),
	.w8(32'hbaa18018),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3911ad20),
	.w1(32'hba80e712),
	.w2(32'h3a2fc8da),
	.w3(32'h397ceed6),
	.w4(32'hba98b2ad),
	.w5(32'hba0c3a14),
	.w6(32'h360107e1),
	.w7(32'h39ef40ca),
	.w8(32'hba45189f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01cf4a),
	.w1(32'hba403ac5),
	.w2(32'hb90a0614),
	.w3(32'hba5cc3c1),
	.w4(32'hba4278cd),
	.w5(32'hba071c5e),
	.w6(32'hb99e32aa),
	.w7(32'hb9b87a0a),
	.w8(32'hba8d525c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398aa551),
	.w1(32'h3a61ee46),
	.w2(32'h3a5553b5),
	.w3(32'hb986b9da),
	.w4(32'h391c7f5a),
	.w5(32'h39373cf3),
	.w6(32'h3a4c0d80),
	.w7(32'h3a29d6b6),
	.w8(32'hb9548776),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87f2a3),
	.w1(32'h3a536d5d),
	.w2(32'h3ace1da2),
	.w3(32'h3a9291c1),
	.w4(32'h3a96022f),
	.w5(32'h3ab91734),
	.w6(32'h3a319a37),
	.w7(32'h3a62dd1f),
	.w8(32'hb9c3a2b3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b282e),
	.w1(32'h3bd058b1),
	.w2(32'h3bf10f73),
	.w3(32'h3ade0902),
	.w4(32'h3b9c2308),
	.w5(32'h3b6f474d),
	.w6(32'h3aabb348),
	.w7(32'h3b5d7e60),
	.w8(32'h3a3e0c68),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1edea),
	.w1(32'hba36db13),
	.w2(32'hb9c7a0de),
	.w3(32'h3b00dcac),
	.w4(32'hb9ac5301),
	.w5(32'h39f16e58),
	.w6(32'hba825000),
	.w7(32'hba4a5598),
	.w8(32'h38d9fedd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57422e),
	.w1(32'hb9c62bc0),
	.w2(32'hba50adfe),
	.w3(32'h3a8d4cf3),
	.w4(32'h39b1c620),
	.w5(32'hb835353f),
	.w6(32'hb9899d67),
	.w7(32'hb9ef35dd),
	.w8(32'hba643c70),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec499a),
	.w1(32'h3b4e9eac),
	.w2(32'h3b83ef81),
	.w3(32'hb97a9487),
	.w4(32'h39cf1f73),
	.w5(32'h3b05abf6),
	.w6(32'hba8836b5),
	.w7(32'h3aa38fdc),
	.w8(32'hbad27b22),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cd9c5),
	.w1(32'hbb0122e3),
	.w2(32'hbae69939),
	.w3(32'hb97d72f6),
	.w4(32'hbb0b95e2),
	.w5(32'hbb04dfcb),
	.w6(32'hbb25991a),
	.w7(32'hbb21c55e),
	.w8(32'hba85f615),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef892d),
	.w1(32'h37c34edc),
	.w2(32'h3a5f7c1d),
	.w3(32'hbab09a3c),
	.w4(32'hb91a6f10),
	.w5(32'h388939d0),
	.w6(32'hb994d5fb),
	.w7(32'h3a4e18de),
	.w8(32'h3a8db97b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23d44c),
	.w1(32'h3ad76490),
	.w2(32'h3b07bbf9),
	.w3(32'hb8ec3090),
	.w4(32'h3ab78ebd),
	.w5(32'h3aa28e07),
	.w6(32'h3a91562f),
	.w7(32'h3a21427b),
	.w8(32'hba1f3cae),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4db55a),
	.w1(32'hbb139c35),
	.w2(32'hba463d8d),
	.w3(32'h3aff8015),
	.w4(32'hbb5691a8),
	.w5(32'hbb5ecbe9),
	.w6(32'hbb145e3d),
	.w7(32'hba8bdee8),
	.w8(32'hbb47ea21),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6f22),
	.w1(32'hbb577d49),
	.w2(32'hbaa69d78),
	.w3(32'hbb5f2508),
	.w4(32'hbb5b2947),
	.w5(32'hbaf06151),
	.w6(32'hbb2ff432),
	.w7(32'hba4d28d8),
	.w8(32'hbab979fc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74c056),
	.w1(32'h3a143e55),
	.w2(32'h3afc3983),
	.w3(32'hbae1f192),
	.w4(32'h3998e780),
	.w5(32'h39814c49),
	.w6(32'h39ef95ba),
	.w7(32'h3a7619b6),
	.w8(32'h3aa6be90),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4533e),
	.w1(32'hba57562d),
	.w2(32'h398fc230),
	.w3(32'h39b69e01),
	.w4(32'hba7d1f9f),
	.w5(32'hba631b41),
	.w6(32'hb936c867),
	.w7(32'hb885bdaa),
	.w8(32'hba32fdc2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9938869),
	.w1(32'h3933838d),
	.w2(32'h3a2637d2),
	.w3(32'hbae9dc11),
	.w4(32'hb8bb5009),
	.w5(32'hb954c3e2),
	.w6(32'h38b06256),
	.w7(32'h39b750ba),
	.w8(32'h3993bdb7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21c31e),
	.w1(32'hbab34021),
	.w2(32'hba2859e1),
	.w3(32'hb8b206a0),
	.w4(32'hbac3d53e),
	.w5(32'hbaa23ae7),
	.w6(32'hba9d16ac),
	.w7(32'hba96aa50),
	.w8(32'hbad146cc),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aae22),
	.w1(32'hba0a9d7e),
	.w2(32'hba09fd80),
	.w3(32'hba9cbc5d),
	.w4(32'hb8bd1acb),
	.w5(32'h3732478c),
	.w6(32'hba165372),
	.w7(32'hb9fcf373),
	.w8(32'hb9b28206),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eb4bf0),
	.w1(32'hba19d691),
	.w2(32'h3a5b7155),
	.w3(32'h399816d9),
	.w4(32'hba4884eb),
	.w5(32'hb9168bd2),
	.w6(32'hb9a26252),
	.w7(32'h39e175ed),
	.w8(32'hba4ddc7d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba1e8f),
	.w1(32'h3917f187),
	.w2(32'h3a534e24),
	.w3(32'hba8b01f3),
	.w4(32'hb95f0968),
	.w5(32'hb84969c4),
	.w6(32'h38d454ce),
	.w7(32'h395f9440),
	.w8(32'h3a1f1fbe),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e3285),
	.w1(32'hba96433c),
	.w2(32'hba5f6e47),
	.w3(32'h38a091b8),
	.w4(32'hbaab2c02),
	.w5(32'hba8caeb4),
	.w6(32'hbaf65db2),
	.w7(32'hbae67b42),
	.w8(32'hba1c6f91),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f5629),
	.w1(32'h37713b95),
	.w2(32'h38f44d2f),
	.w3(32'hba6f6383),
	.w4(32'hbab23ead),
	.w5(32'hbad1d7db),
	.w6(32'hba8a4da2),
	.w7(32'hbaa32975),
	.w8(32'hba896c4d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d56d3),
	.w1(32'hbaa2ff95),
	.w2(32'hbb285f25),
	.w3(32'hbaa096d6),
	.w4(32'hba5af3fc),
	.w5(32'hbb2cbbc7),
	.w6(32'hbb00ce5f),
	.w7(32'hbaaa66e3),
	.w8(32'hbac0787a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bd451),
	.w1(32'hb9ca5c9a),
	.w2(32'hb9075e7c),
	.w3(32'hbb66aab9),
	.w4(32'hba5333ae),
	.w5(32'hba8d31b0),
	.w6(32'h370d22ab),
	.w7(32'hb9f1e89d),
	.w8(32'hba2b6255),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d19f4d),
	.w1(32'hba78456c),
	.w2(32'hba121b4d),
	.w3(32'hba8d80d2),
	.w4(32'hbaa46e88),
	.w5(32'hba4ce72f),
	.w6(32'hba79b0ef),
	.w7(32'hba43835f),
	.w8(32'hba1493aa),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e092b4),
	.w1(32'hb91d0c94),
	.w2(32'hba7ba8ba),
	.w3(32'hb9c0a6e2),
	.w4(32'hba4b0e29),
	.w5(32'hbadfa96b),
	.w6(32'hba47e1f0),
	.w7(32'hba8e014d),
	.w8(32'hba8d2f33),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9ce0b),
	.w1(32'h3989d15a),
	.w2(32'h3a88b3b7),
	.w3(32'hbaebf50a),
	.w4(32'h38e3b8e6),
	.w5(32'h38e892e7),
	.w6(32'h3a06961c),
	.w7(32'h3a47b367),
	.w8(32'h3a48fe06),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a969074),
	.w1(32'hb90b721e),
	.w2(32'h3a060271),
	.w3(32'h39659e25),
	.w4(32'hb85ebca8),
	.w5(32'h39737f7e),
	.w6(32'h38928c27),
	.w7(32'h39db1621),
	.w8(32'h39018179),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38138006),
	.w1(32'hb91a18fe),
	.w2(32'h3a15fadd),
	.w3(32'h3794165e),
	.w4(32'hb880f01c),
	.w5(32'h39877611),
	.w6(32'h38b87e26),
	.w7(32'h39d51b2c),
	.w8(32'h392cd048),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ef19ff),
	.w1(32'hbb3f5fab),
	.w2(32'hbb25bb98),
	.w3(32'h37abd3d4),
	.w4(32'hba214dea),
	.w5(32'h392ab53f),
	.w6(32'hbae030eb),
	.w7(32'hbabbc85c),
	.w8(32'hb734441f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacee152),
	.w1(32'hba46ce5d),
	.w2(32'hb833f6c2),
	.w3(32'h3837fa13),
	.w4(32'hbac2f1b1),
	.w5(32'hbab887a1),
	.w6(32'hba633985),
	.w7(32'hb9fe8690),
	.w8(32'h3a8e856a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14cbf1),
	.w1(32'hb9b81166),
	.w2(32'h38c8a02e),
	.w3(32'h38ef8330),
	.w4(32'hba4c11c5),
	.w5(32'hba9d9dfa),
	.w6(32'hb9c1b0fd),
	.w7(32'hba70399a),
	.w8(32'hba9990bb),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d9110),
	.w1(32'hba9c86d1),
	.w2(32'hba501ba5),
	.w3(32'hba7676c8),
	.w4(32'hbacd9455),
	.w5(32'hba832325),
	.w6(32'hbaa6a707),
	.w7(32'hbabdd496),
	.w8(32'hba9cc432),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a35f4),
	.w1(32'hb93f3aa3),
	.w2(32'h391f775a),
	.w3(32'hba25d111),
	.w4(32'hb9976bac),
	.w5(32'hb9c8a592),
	.w6(32'h389dad17),
	.w7(32'h39b7b14d),
	.w8(32'h38396e5c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7049c38),
	.w1(32'hbb4df068),
	.w2(32'hbb5366c6),
	.w3(32'hb9d6d27b),
	.w4(32'hbac5ef51),
	.w5(32'hb9b9e981),
	.w6(32'hbb421657),
	.w7(32'hbafd82f9),
	.w8(32'hba5646fa),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb327333),
	.w1(32'h3a2145b2),
	.w2(32'h3accdbb7),
	.w3(32'hb9e1afd0),
	.w4(32'h3aa985d5),
	.w5(32'h3aa48c47),
	.w6(32'h3a84d722),
	.w7(32'h3a3e0e1b),
	.w8(32'hb9c522d9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac8424),
	.w1(32'hbab13dd0),
	.w2(32'h380bbd94),
	.w3(32'h3a164da3),
	.w4(32'hbac09c53),
	.w5(32'hba94b6cd),
	.w6(32'hb9de1c92),
	.w7(32'h372c4696),
	.w8(32'hba8163c5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba891176),
	.w1(32'hba0cdcae),
	.w2(32'hba4fcf7b),
	.w3(32'hbabc3c18),
	.w4(32'hb90f43c6),
	.w5(32'hb931ddd5),
	.w6(32'hb992d20b),
	.w7(32'h3798ee84),
	.w8(32'h396be22b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eeb083),
	.w1(32'h397d80fe),
	.w2(32'h3a0f4585),
	.w3(32'hb9e1d49a),
	.w4(32'h3a2bf8d0),
	.w5(32'h3a39ede8),
	.w6(32'hb813247a),
	.w7(32'h3952e840),
	.w8(32'h3a095dff),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998ee97),
	.w1(32'h3b135530),
	.w2(32'h3aa48463),
	.w3(32'h3a2fe247),
	.w4(32'h3ab8a42d),
	.w5(32'h3a6301d1),
	.w6(32'h3a66b779),
	.w7(32'hbaa0e441),
	.w8(32'h3a4aeaa2),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06f1c0),
	.w1(32'h38eeedff),
	.w2(32'hb915dcd0),
	.w3(32'h3a96fa60),
	.w4(32'h3a186352),
	.w5(32'h39d983e8),
	.w6(32'h39b46ba9),
	.w7(32'h392dbc85),
	.w8(32'h39b9c23b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fda0d4),
	.w1(32'hb9f44f45),
	.w2(32'hb9ddcce3),
	.w3(32'h39fd172d),
	.w4(32'h39eaa067),
	.w5(32'h39b398a9),
	.w6(32'h399bcd5b),
	.w7(32'hb8668e20),
	.w8(32'hb8664de6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff5f7d),
	.w1(32'hb95e8689),
	.w2(32'h39275f6a),
	.w3(32'h389f857c),
	.w4(32'h3a5b638d),
	.w5(32'h39ed01a0),
	.w6(32'h39e49862),
	.w7(32'hb88264c6),
	.w8(32'h39e223bf),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d6975),
	.w1(32'hb98be6d6),
	.w2(32'hbac52094),
	.w3(32'h39dbdccb),
	.w4(32'h396be871),
	.w5(32'h39b06d3f),
	.w6(32'hba14fad4),
	.w7(32'hb801066b),
	.w8(32'h3a062f2e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18b402),
	.w1(32'h393372a4),
	.w2(32'h38ad2eea),
	.w3(32'h3a45618e),
	.w4(32'h3a5366eb),
	.w5(32'h3aa70bb8),
	.w6(32'h398deb8d),
	.w7(32'h3a7fc50f),
	.w8(32'h3ab406b4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09526b),
	.w1(32'h3867ca4d),
	.w2(32'hb73a392b),
	.w3(32'h3a39f66f),
	.w4(32'h39f04307),
	.w5(32'h3a2b51c8),
	.w6(32'h398c5d92),
	.w7(32'h397184e6),
	.w8(32'h39984379),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fd786),
	.w1(32'h3986678e),
	.w2(32'h3954f64a),
	.w3(32'h3a0828d3),
	.w4(32'h394d0750),
	.w5(32'h399e010a),
	.w6(32'h38b3fb6b),
	.w7(32'h38bcc6aa),
	.w8(32'h3842f029),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38962b89),
	.w1(32'h38177bf1),
	.w2(32'h382f1083),
	.w3(32'h397e4a82),
	.w4(32'h39b63cb6),
	.w5(32'h3a2d8a82),
	.w6(32'h39b08592),
	.w7(32'h39ead3be),
	.w8(32'h39a5122e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30182a),
	.w1(32'h393c1258),
	.w2(32'h38be4801),
	.w3(32'h3a1346d0),
	.w4(32'h39e493f0),
	.w5(32'h39f9c469),
	.w6(32'h3985a632),
	.w7(32'h39a08ded),
	.w8(32'h3a45f8e7),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e47d97),
	.w1(32'h382623e9),
	.w2(32'h3a0cdf2f),
	.w3(32'h3a2e80bb),
	.w4(32'h3a2726db),
	.w5(32'h38772f33),
	.w6(32'h3a2d744b),
	.w7(32'h3a20c4de),
	.w8(32'h3a993798),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379029ec),
	.w1(32'hb9b5ad0a),
	.w2(32'h3a8fc267),
	.w3(32'h383efb8b),
	.w4(32'hb71c8a67),
	.w5(32'h3a118de8),
	.w6(32'h38d79ef0),
	.w7(32'h3a251be5),
	.w8(32'h3a15c23b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7aec1),
	.w1(32'hb95ad3dd),
	.w2(32'hb863781f),
	.w3(32'h39a5f31d),
	.w4(32'hb92154fd),
	.w5(32'hb99765a2),
	.w6(32'hb9a7f304),
	.w7(32'hb99fecda),
	.w8(32'h38ad7a80),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aaf9d6),
	.w1(32'h39870fd3),
	.w2(32'h39718701),
	.w3(32'hb98fac21),
	.w4(32'h3953fc74),
	.w5(32'h3881182c),
	.w6(32'h3a027e8d),
	.w7(32'h3a32a952),
	.w8(32'h39a1eb75),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ce2f8),
	.w1(32'hba5a2178),
	.w2(32'h3a1f9884),
	.w3(32'hb907a4bb),
	.w4(32'h397e837f),
	.w5(32'h3a5a0c90),
	.w6(32'hb924ff24),
	.w7(32'h3987557f),
	.w8(32'h3a893a6f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b4bfc),
	.w1(32'h39f942e3),
	.w2(32'h39e2a2bb),
	.w3(32'h3a960fa4),
	.w4(32'h3a5beccc),
	.w5(32'h3a75964b),
	.w6(32'h3a5e4a20),
	.w7(32'h3a4effcf),
	.w8(32'h3a1f86d9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15e8ac),
	.w1(32'h38cb2b1d),
	.w2(32'h399efe47),
	.w3(32'h3a4375c9),
	.w4(32'h395d74e9),
	.w5(32'hb95d47e2),
	.w6(32'hb89c0eba),
	.w7(32'hb82c2355),
	.w8(32'hb9bf9e01),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1efcc8),
	.w1(32'hb93c6044),
	.w2(32'hb9c4e266),
	.w3(32'hb9c07f04),
	.w4(32'h39da3632),
	.w5(32'h3a01f673),
	.w6(32'h394f802b),
	.w7(32'h395e93dc),
	.w8(32'h39d22a20),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39afd1e6),
	.w1(32'h39ca077e),
	.w2(32'h3962ee4b),
	.w3(32'h39fa1dd0),
	.w4(32'h398f402a),
	.w5(32'h38b3903e),
	.w6(32'h395ddccb),
	.w7(32'hb88b7dcb),
	.w8(32'hb939f9cf),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a052316),
	.w1(32'h39c3af1c),
	.w2(32'hb7d7b5de),
	.w3(32'h3a117f18),
	.w4(32'h3a565530),
	.w5(32'h39d215cb),
	.w6(32'h39ed6baf),
	.w7(32'h3a591393),
	.w8(32'h39872932),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394544d3),
	.w1(32'hb94fb7ef),
	.w2(32'hb9b5a733),
	.w3(32'h390bf859),
	.w4(32'h39759ac8),
	.w5(32'h397c0fb4),
	.w6(32'h38ec340f),
	.w7(32'h38f0a245),
	.w8(32'hb9b0593e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea874c),
	.w1(32'hb5a78139),
	.w2(32'h3a9d402e),
	.w3(32'hb9ab81e6),
	.w4(32'hba006a47),
	.w5(32'hb926c31d),
	.w6(32'hb9deafef),
	.w7(32'h39cc921c),
	.w8(32'h3a778904),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13d621),
	.w1(32'hb9f4777d),
	.w2(32'hb9aa9de6),
	.w3(32'hba2023f8),
	.w4(32'hbab57f6f),
	.w5(32'hba8ed4a1),
	.w6(32'hba20965b),
	.w7(32'hb9e418d6),
	.w8(32'hba6b4711),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a04c1),
	.w1(32'hb8e0f0ff),
	.w2(32'hb88a8112),
	.w3(32'hbab82f4c),
	.w4(32'h387651a0),
	.w5(32'h38d46244),
	.w6(32'hb8f5f7b0),
	.w7(32'h3992c357),
	.w8(32'hb87e6a3d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38738e67),
	.w1(32'h3975be38),
	.w2(32'h38ad8b01),
	.w3(32'h39b62667),
	.w4(32'h3a20f383),
	.w5(32'h39b7332a),
	.w6(32'h3a60b455),
	.w7(32'h3995e29a),
	.w8(32'h39b88ce3),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d69763),
	.w1(32'hb8e3c453),
	.w2(32'h3890be86),
	.w3(32'h3a21dc45),
	.w4(32'h39fe3d6a),
	.w5(32'h39abb4a9),
	.w6(32'h39e85493),
	.w7(32'h3a2b4f6b),
	.w8(32'h39360829),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2065f),
	.w1(32'hb9223fad),
	.w2(32'hb908fc4b),
	.w3(32'h39163efa),
	.w4(32'h396f06f9),
	.w5(32'h3963e906),
	.w6(32'h388d4123),
	.w7(32'h388d0dd2),
	.w8(32'hb950672f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb909fbb0),
	.w1(32'hba1e60ed),
	.w2(32'hb9dae06b),
	.w3(32'hb8ea0d41),
	.w4(32'hb85cd560),
	.w5(32'h391bbd41),
	.w6(32'hba17be31),
	.w7(32'hba44dab2),
	.w8(32'hb98f346b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9086720),
	.w1(32'hb98248dd),
	.w2(32'h39b10941),
	.w3(32'hba02d126),
	.w4(32'hb9a5c560),
	.w5(32'h399a5b2f),
	.w6(32'hba873683),
	.w7(32'h3a9fa243),
	.w8(32'h3999b03f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba344d97),
	.w1(32'hb9491b1d),
	.w2(32'hba82c4fd),
	.w3(32'hb8abc2a2),
	.w4(32'h38319aee),
	.w5(32'hba8aa1db),
	.w6(32'hb9299580),
	.w7(32'hba673033),
	.w8(32'hba40d8f2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990b6e8),
	.w1(32'hb8ee000d),
	.w2(32'hb9099c09),
	.w3(32'hb9e1c22d),
	.w4(32'h39381f43),
	.w5(32'h393a2f94),
	.w6(32'hb7a97d29),
	.w7(32'h38d9881d),
	.w8(32'hb87cd5c0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953abdb),
	.w1(32'hb9379b08),
	.w2(32'hb884695e),
	.w3(32'hb8288be8),
	.w4(32'h391c2e88),
	.w5(32'h39184501),
	.w6(32'hb93136b3),
	.w7(32'hb85ab5ad),
	.w8(32'hb8a49296),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb850006b),
	.w1(32'h3a13a15f),
	.w2(32'hba91b244),
	.w3(32'hb756e8fb),
	.w4(32'h3931967a),
	.w5(32'hba2cac06),
	.w6(32'hb8a5dc16),
	.w7(32'hba4ca401),
	.w8(32'h3a0762e7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a491e66),
	.w1(32'h399f526e),
	.w2(32'hba2c9477),
	.w3(32'h3a0e3381),
	.w4(32'h3a077d04),
	.w5(32'h394cde42),
	.w6(32'hb92cb95e),
	.w7(32'hb9fa8377),
	.w8(32'h39b22ed0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949807c),
	.w1(32'hb9dba641),
	.w2(32'hb9e3d02e),
	.w3(32'h3995ca04),
	.w4(32'h3a20e02b),
	.w5(32'h3a341257),
	.w6(32'h399e7526),
	.w7(32'h3951f17c),
	.w8(32'h3a0b30ed),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390573c0),
	.w1(32'hb999db34),
	.w2(32'hb916fe78),
	.w3(32'h39f4eb21),
	.w4(32'h39391620),
	.w5(32'h38fd5a6c),
	.w6(32'hb805cdc3),
	.w7(32'h372d2f54),
	.w8(32'hb94d581c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ce6032),
	.w1(32'hb9dc33a1),
	.w2(32'hba300608),
	.w3(32'h3918496f),
	.w4(32'h39f2dda4),
	.w5(32'h39568267),
	.w6(32'h39d70c31),
	.w7(32'h3930d2cc),
	.w8(32'h38a8c14f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84c00bb),
	.w1(32'h3930a9ca),
	.w2(32'hb9ba86cd),
	.w3(32'h39467eb9),
	.w4(32'h3a3b49c6),
	.w5(32'h3a02853f),
	.w6(32'h3a058ef4),
	.w7(32'h39d8dc72),
	.w8(32'h39dbffa6),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c2da4),
	.w1(32'h399d248e),
	.w2(32'h39b4132f),
	.w3(32'h3a1dda62),
	.w4(32'h3a2bfb3f),
	.w5(32'h39dbf179),
	.w6(32'h39f6cda7),
	.w7(32'h3a21193d),
	.w8(32'h39b35427),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d5c2a),
	.w1(32'h39ddd354),
	.w2(32'h39cb0eda),
	.w3(32'h39e8f2ae),
	.w4(32'h398bc108),
	.w5(32'h395148d4),
	.w6(32'h3909bcf1),
	.w7(32'hb93b8661),
	.w8(32'hb906d47a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a23b03),
	.w1(32'h391fe6f9),
	.w2(32'hba29d6ac),
	.w3(32'hb8ff455b),
	.w4(32'hb9b65bb8),
	.w5(32'hb9f69518),
	.w6(32'hba18cd91),
	.w7(32'hba916537),
	.w8(32'h3803c9ec),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34659a),
	.w1(32'h394e3a32),
	.w2(32'h39dda6de),
	.w3(32'hb9af78a0),
	.w4(32'h3a3a8857),
	.w5(32'h3a130f26),
	.w6(32'h39c16215),
	.w7(32'h38898c7c),
	.w8(32'h39a1bb1b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb894e92a),
	.w1(32'hb96cbce2),
	.w2(32'hb7c6e3ab),
	.w3(32'hb9f4a613),
	.w4(32'hba276b70),
	.w5(32'hb9b557ad),
	.w6(32'hba853baf),
	.w7(32'hba3b9607),
	.w8(32'hba26bf67),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb974e4eb),
	.w1(32'h3924200a),
	.w2(32'h3926b547),
	.w3(32'hb8b646e1),
	.w4(32'h393b20ec),
	.w5(32'h3a029f9e),
	.w6(32'h3a45959e),
	.w7(32'h3a6edfa7),
	.w8(32'h3aacc8d9),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32c334),
	.w1(32'h39f4e25f),
	.w2(32'hb950857d),
	.w3(32'h3a749171),
	.w4(32'h39a3e1b1),
	.w5(32'h39e8bf7a),
	.w6(32'h3a7c4f85),
	.w7(32'h3a59a2be),
	.w8(32'h3ab68cf2),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a193a4a),
	.w1(32'h38431094),
	.w2(32'h37df14f1),
	.w3(32'h3aa88fd6),
	.w4(32'h396eb1dd),
	.w5(32'h39f5d734),
	.w6(32'h3a0e21c2),
	.w7(32'h3a819154),
	.w8(32'h3a0a6984),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26501d),
	.w1(32'hba5c59ad),
	.w2(32'h3b07c1bd),
	.w3(32'hb8e1f5ff),
	.w4(32'hba4eeed2),
	.w5(32'h3885ff10),
	.w6(32'hb9916f01),
	.w7(32'hb94c9959),
	.w8(32'h3a70b255),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a636a2b),
	.w1(32'hba068ebe),
	.w2(32'hba2349b3),
	.w3(32'h39e75fd1),
	.w4(32'hb9b02366),
	.w5(32'hb815d3a6),
	.w6(32'hb9973a1b),
	.w7(32'hb9e043d5),
	.w8(32'hb9ca9112),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0498b5),
	.w1(32'h386ea149),
	.w2(32'h392deb3a),
	.w3(32'hb815352e),
	.w4(32'hb99ed9cc),
	.w5(32'hb8ebd494),
	.w6(32'hba187e5c),
	.w7(32'hb9b0d8bd),
	.w8(32'hb91e1a4f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb931a667),
	.w1(32'hb89f7f3f),
	.w2(32'hb8087eb8),
	.w3(32'hb8ff4c93),
	.w4(32'h3752104d),
	.w5(32'h38f83b55),
	.w6(32'hb8277d68),
	.w7(32'h3901ef56),
	.w8(32'h36bb0b1e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f7d172),
	.w1(32'h39924b2e),
	.w2(32'h3a3edbfe),
	.w3(32'h3893f37d),
	.w4(32'h394eb845),
	.w5(32'h39211a82),
	.w6(32'h39d371fa),
	.w7(32'h3a1d7cfd),
	.w8(32'h39070908),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4933e),
	.w1(32'h3b01b4df),
	.w2(32'h38c9b839),
	.w3(32'hb9785ee2),
	.w4(32'h3ad1cf53),
	.w5(32'h3911c680),
	.w6(32'h3afcce31),
	.w7(32'h3a5969f6),
	.w8(32'h3aa48cff),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c9cec),
	.w1(32'h3ace0236),
	.w2(32'h3a94b14e),
	.w3(32'h3a0c45a6),
	.w4(32'h3abdbe1a),
	.w5(32'h3aafd6da),
	.w6(32'h3abf46ff),
	.w7(32'h3aa2a5f5),
	.w8(32'h3a8066d7),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab30c29),
	.w1(32'hb887991a),
	.w2(32'hba8674f7),
	.w3(32'h3a9ee84a),
	.w4(32'h38b664ed),
	.w5(32'h39a56a07),
	.w6(32'hb9a690f7),
	.w7(32'h3a249ecf),
	.w8(32'h39e97317),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ecc5b),
	.w1(32'h39a63ef6),
	.w2(32'hb9abcc1c),
	.w3(32'h3a85e16f),
	.w4(32'h3985676e),
	.w5(32'h3897ae3c),
	.w6(32'h3943f430),
	.w7(32'h37fa7a02),
	.w8(32'h394299f0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921495e),
	.w1(32'hba2dfe4b),
	.w2(32'hb94d091d),
	.w3(32'h39c27fd6),
	.w4(32'h3899b693),
	.w5(32'hb9b57c7d),
	.w6(32'hb9c21347),
	.w7(32'hb9c52418),
	.w8(32'hb9a36f08),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb49fd464),
	.w1(32'hb97ab260),
	.w2(32'hb8c48b80),
	.w3(32'hba094f29),
	.w4(32'h38edb846),
	.w5(32'h392f4712),
	.w6(32'h38a5d4e0),
	.w7(32'h3990a797),
	.w8(32'hb98a738e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba114e60),
	.w1(32'h37c31dcb),
	.w2(32'hba43d94a),
	.w3(32'hb9dd2f58),
	.w4(32'h392daec8),
	.w5(32'hb7f70bc6),
	.w6(32'hb9b4b6a8),
	.w7(32'h39829af1),
	.w8(32'h399ef379),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d1059),
	.w1(32'h3a2724fa),
	.w2(32'hb86b31d2),
	.w3(32'h3a563d22),
	.w4(32'h3a85903c),
	.w5(32'h3a0bfa65),
	.w6(32'h3a3605da),
	.w7(32'h39ab1d5b),
	.w8(32'h3a1e8b48),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93085e4),
	.w1(32'h38d7d235),
	.w2(32'h3a022fa6),
	.w3(32'h3899ca83),
	.w4(32'h393a5f04),
	.w5(32'h3a053609),
	.w6(32'hb90009f9),
	.w7(32'h39824817),
	.w8(32'h3a29626d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6cede),
	.w1(32'h38866cf6),
	.w2(32'h39f9247d),
	.w3(32'h3907df98),
	.w4(32'h3a3047f9),
	.w5(32'h3a4372ca),
	.w6(32'hb8416890),
	.w7(32'hb9bc03ff),
	.w8(32'h39603ec7),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398cb838),
	.w1(32'hb9364d4a),
	.w2(32'hb9529299),
	.w3(32'h39d901ff),
	.w4(32'h372218e3),
	.w5(32'hb81a011f),
	.w6(32'hb7027af5),
	.w7(32'h39248425),
	.w8(32'h395ede3b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5f94d),
	.w1(32'h3aac099f),
	.w2(32'hbaef0f00),
	.w3(32'hb92074c5),
	.w4(32'h3a53cc78),
	.w5(32'hb9baf827),
	.w6(32'hb706541b),
	.w7(32'hba750408),
	.w8(32'h3a8ab2e2),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a392def),
	.w1(32'h37acce39),
	.w2(32'h3873278c),
	.w3(32'h3a7a3dd9),
	.w4(32'h39021343),
	.w5(32'h39a32537),
	.w6(32'h39ef71f6),
	.w7(32'h3a13510b),
	.w8(32'h3a6ae1e0),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9c4b6),
	.w1(32'hba0088f7),
	.w2(32'hba08f707),
	.w3(32'h3a131ca6),
	.w4(32'hb832c672),
	.w5(32'hb957554d),
	.w6(32'hb99b8302),
	.w7(32'hb994b221),
	.w8(32'h38df26f8),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394888b7),
	.w1(32'h39f6b719),
	.w2(32'hb99b746c),
	.w3(32'h39316ab5),
	.w4(32'hb98628f6),
	.w5(32'hb9c58aff),
	.w6(32'hb9a9117e),
	.w7(32'h39834ee3),
	.w8(32'h383ebf03),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384e4508),
	.w1(32'h3a3d7a35),
	.w2(32'hb919d1c4),
	.w3(32'hb87f7b12),
	.w4(32'h3a0bf3e0),
	.w5(32'hb8dea199),
	.w6(32'h38d7d325),
	.w7(32'h380a903a),
	.w8(32'h39bca20d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb881853e),
	.w1(32'hb92c69c3),
	.w2(32'hba61446d),
	.w3(32'hb9b23e62),
	.w4(32'hba0ee21b),
	.w5(32'hba405664),
	.w6(32'hb9c46c67),
	.w7(32'hba135677),
	.w8(32'hb9fa07ed),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4796e),
	.w1(32'h3a828ceb),
	.w2(32'h3a39a962),
	.w3(32'hba14ce13),
	.w4(32'h3a5aa024),
	.w5(32'h3a185a2c),
	.w6(32'h3a64b0c2),
	.w7(32'h3a87070f),
	.w8(32'h3a3e8eca),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e2b5c),
	.w1(32'hb9da7c49),
	.w2(32'h391f8c79),
	.w3(32'h39e0a2cf),
	.w4(32'hb9e86b2a),
	.w5(32'h3948baa7),
	.w6(32'hba04c756),
	.w7(32'h37e19410),
	.w8(32'h391eb23f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3880e46f),
	.w1(32'hb96be716),
	.w2(32'hb9b10e74),
	.w3(32'hb94eb6f4),
	.w4(32'h39be1a25),
	.w5(32'h39b6cf0e),
	.w6(32'h395f7c6c),
	.w7(32'h3962be69),
	.w8(32'h396dd7f5),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc4371),
	.w1(32'h38fd2315),
	.w2(32'h390e46e4),
	.w3(32'h397bb5cf),
	.w4(32'h399cb1de),
	.w5(32'h3987fcdc),
	.w6(32'hb89fe144),
	.w7(32'h38c2314f),
	.w8(32'h3953775e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394fd390),
	.w1(32'h3916818e),
	.w2(32'h393e6697),
	.w3(32'h395ff7b7),
	.w4(32'h39ea7d9d),
	.w5(32'h39d57c54),
	.w6(32'h39ad1e32),
	.w7(32'h396cbfd6),
	.w8(32'h3646fddf),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392286a9),
	.w1(32'hb9684bcd),
	.w2(32'hb8c6f5ef),
	.w3(32'h398c2035),
	.w4(32'h398678bd),
	.w5(32'h3998b998),
	.w6(32'hb8f255f4),
	.w7(32'h37a0eda2),
	.w8(32'hb99a12a2),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7588121),
	.w1(32'h399ce0f6),
	.w2(32'h38a29310),
	.w3(32'h38c71971),
	.w4(32'h3a37c841),
	.w5(32'h39e01c05),
	.w6(32'h39a453bc),
	.w7(32'h37cd2097),
	.w8(32'h39c882fa),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c62c6),
	.w1(32'h3a61b695),
	.w2(32'h3b0705b0),
	.w3(32'h38d1c98c),
	.w4(32'hb8a043ff),
	.w5(32'hba8a66ee),
	.w6(32'h3a2348ea),
	.w7(32'hb99e832a),
	.w8(32'h3924289d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd3e33),
	.w1(32'h384b0a0b),
	.w2(32'h3960ba3c),
	.w3(32'hb9161af2),
	.w4(32'hb89c0160),
	.w5(32'h38f08758),
	.w6(32'hb916a2df),
	.w7(32'h38f930e4),
	.w8(32'h3990fb65),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8655e58),
	.w1(32'h3a6bb39a),
	.w2(32'hb98a4517),
	.w3(32'h39402a47),
	.w4(32'h3a94ebeb),
	.w5(32'h3a025863),
	.w6(32'h3a3a973f),
	.w7(32'h38e4ea44),
	.w8(32'h3a27f395),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af6bd9),
	.w1(32'h3991efa4),
	.w2(32'h38ab74bb),
	.w3(32'h3a1270af),
	.w4(32'h39488aee),
	.w5(32'hb9441f2d),
	.w6(32'hb7a102a5),
	.w7(32'h38f5154b),
	.w8(32'hb8f0275c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a8d07f),
	.w1(32'hba0e54f4),
	.w2(32'hb9a20797),
	.w3(32'hb9a75e77),
	.w4(32'hb8e094e5),
	.w5(32'h3894e1dc),
	.w6(32'hb982b730),
	.w7(32'hb8ab104d),
	.w8(32'hb84c1f3f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03f9a0),
	.w1(32'hb9913e13),
	.w2(32'hba19244c),
	.w3(32'hb8316285),
	.w4(32'hb9a86904),
	.w5(32'hb90f442b),
	.w6(32'hba074d4b),
	.w7(32'hb99e2457),
	.w8(32'hb91b245d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba022ec4),
	.w1(32'h3a5c1c4a),
	.w2(32'h39bb98be),
	.w3(32'hb9eb2d46),
	.w4(32'h3a8f6ab6),
	.w5(32'h3a55ed46),
	.w6(32'h3a1d6204),
	.w7(32'h3a0b8054),
	.w8(32'h39f29914),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0dc08),
	.w1(32'h3936f9b2),
	.w2(32'h379eff41),
	.w3(32'h3a0b6924),
	.w4(32'h3840c79c),
	.w5(32'h38dc7881),
	.w6(32'hb8534974),
	.w7(32'hb91aaa19),
	.w8(32'hb8895b18),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394105e3),
	.w1(32'h3a1c018b),
	.w2(32'h39f059d9),
	.w3(32'hb8acbe18),
	.w4(32'h3a635a4d),
	.w5(32'h3a2329b8),
	.w6(32'h3a1f116e),
	.w7(32'h3988d5e1),
	.w8(32'h39fd298b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992a0ba),
	.w1(32'hb9b9fe46),
	.w2(32'hb9d64a62),
	.w3(32'h3764c8ba),
	.w4(32'hba3ae4bb),
	.w5(32'hba0cae65),
	.w6(32'hb785e69b),
	.w7(32'hba1e9d86),
	.w8(32'h3a067395),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b0649),
	.w1(32'h3a493fb8),
	.w2(32'h39db7169),
	.w3(32'hb8f86115),
	.w4(32'h3a092c47),
	.w5(32'h39c22c48),
	.w6(32'h39d95bee),
	.w7(32'h39e3b1ff),
	.w8(32'h3a003f07),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e64a4),
	.w1(32'hb9806065),
	.w2(32'hb9f24578),
	.w3(32'h39387faa),
	.w4(32'hb9e9a7df),
	.w5(32'hb9fc0278),
	.w6(32'hb9a7296d),
	.w7(32'hba2613c2),
	.w8(32'hb903b933),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8216bdb),
	.w1(32'hb84c706a),
	.w2(32'hb9219fc8),
	.w3(32'hb9ed7d55),
	.w4(32'h3985b47e),
	.w5(32'h398211c6),
	.w6(32'h38e3e986),
	.w7(32'h391421f8),
	.w8(32'hb92ce0ed),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982924d),
	.w1(32'h39b6d584),
	.w2(32'hb97b496d),
	.w3(32'h387a2a66),
	.w4(32'h39d5d9e3),
	.w5(32'h39a9161c),
	.w6(32'h39aa9c99),
	.w7(32'h388fe1ca),
	.w8(32'h398bc3b2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38efd56f),
	.w1(32'hb9e036fe),
	.w2(32'hb9708b8d),
	.w3(32'h399d1d06),
	.w4(32'h396b1e9e),
	.w5(32'h39905cee),
	.w6(32'h38b80734),
	.w7(32'hb61356a1),
	.w8(32'hb972b624),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b81644),
	.w1(32'h398852e8),
	.w2(32'h3a1b1a46),
	.w3(32'hb92da485),
	.w4(32'h3a118ef3),
	.w5(32'h39b70240),
	.w6(32'h375af45c),
	.w7(32'h3969c45c),
	.w8(32'h38a822e6),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb908ba7f),
	.w1(32'h3950d1ac),
	.w2(32'hb8fd8edc),
	.w3(32'hb94370e7),
	.w4(32'h3956197f),
	.w5(32'h39a353f2),
	.w6(32'h39d1c1ed),
	.w7(32'h3a165fe5),
	.w8(32'h3a2db558),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a14012),
	.w1(32'h3967eff1),
	.w2(32'hb962906e),
	.w3(32'h3a2c6d98),
	.w4(32'h3a081e61),
	.w5(32'h39760349),
	.w6(32'h39661d8e),
	.w7(32'hb7de4a0f),
	.w8(32'h39a6c9d1),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f776c3),
	.w1(32'hba01eb17),
	.w2(32'hb9a6de35),
	.w3(32'h3a1f4a61),
	.w4(32'hba1ade5b),
	.w5(32'hb9910c4a),
	.w6(32'hb9bfe743),
	.w7(32'hb96aa258),
	.w8(32'hb9f7eadd),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eccd1d),
	.w1(32'hba0573a9),
	.w2(32'hb9b79053),
	.w3(32'hb9da7c17),
	.w4(32'h3933b187),
	.w5(32'h392a4ca4),
	.w6(32'h3860f32d),
	.w7(32'hb85161d8),
	.w8(32'h375a24bd),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfb05e),
	.w1(32'h3a79aacf),
	.w2(32'h3ace51f7),
	.w3(32'hb96e5123),
	.w4(32'hb86d0b35),
	.w5(32'h39b3850f),
	.w6(32'h3984f460),
	.w7(32'h3a15dd45),
	.w8(32'h3a0c32d2),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa82d02),
	.w1(32'h391b1320),
	.w2(32'hba1926a1),
	.w3(32'h3a6ef035),
	.w4(32'hb9dcc339),
	.w5(32'hb9817fee),
	.w6(32'hb90bc650),
	.w7(32'hb81b408c),
	.w8(32'hbaa7b41a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba710e2b),
	.w1(32'h38b082c1),
	.w2(32'hba71cd1e),
	.w3(32'hbaa8a6c4),
	.w4(32'h3a078f57),
	.w5(32'hb90f9149),
	.w6(32'h38611e9c),
	.w7(32'hba16dbae),
	.w8(32'h39515068),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c0107),
	.w1(32'h39ddd72d),
	.w2(32'h396ccf5a),
	.w3(32'h39d96833),
	.w4(32'h3a2e0f30),
	.w5(32'h3a36e73d),
	.w6(32'h397242ae),
	.w7(32'h39a4dd35),
	.w8(32'h39e67d8a),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a4560),
	.w1(32'h3995271f),
	.w2(32'h38b2c4f0),
	.w3(32'h398b9298),
	.w4(32'h39b90a14),
	.w5(32'h39ece6d7),
	.w6(32'h39daae7d),
	.w7(32'hb780c067),
	.w8(32'h391d3827),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39655433),
	.w1(32'hb99d5f9a),
	.w2(32'hba98aa17),
	.w3(32'h3994822c),
	.w4(32'hb9e4fa75),
	.w5(32'hba158715),
	.w6(32'hbaa5ae7f),
	.w7(32'hb903c3bc),
	.w8(32'h397a43d1),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393295e6),
	.w1(32'h3a986c7f),
	.w2(32'h3a902299),
	.w3(32'h399e06b2),
	.w4(32'h395cc9a0),
	.w5(32'hb9ccc51b),
	.w6(32'hba420b4f),
	.w7(32'h3aadcf1c),
	.w8(32'h39fe6fce),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfc021),
	.w1(32'hb9d0a93b),
	.w2(32'h394a75cc),
	.w3(32'h371a103a),
	.w4(32'hb98fbe48),
	.w5(32'h3957c73b),
	.w6(32'hb9a7213a),
	.w7(32'h3971499f),
	.w8(32'h3a0cba44),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991fa8e),
	.w1(32'hb8df5680),
	.w2(32'h38a35d53),
	.w3(32'h38a69c2a),
	.w4(32'h39b220b9),
	.w5(32'h39db8a4c),
	.w6(32'hb99dc723),
	.w7(32'h37c4ee37),
	.w8(32'h39a0a8ea),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d7739b),
	.w1(32'hb984d525),
	.w2(32'hb96396fb),
	.w3(32'h39a19140),
	.w4(32'hb9647f9c),
	.w5(32'hb8d50e54),
	.w6(32'hb95846c6),
	.w7(32'hb79c7451),
	.w8(32'h388f3e1a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76aa854),
	.w1(32'hb92d7e8b),
	.w2(32'hb8cb4f8a),
	.w3(32'h38f9fedc),
	.w4(32'h392db847),
	.w5(32'h39aa63a4),
	.w6(32'h386b9d8c),
	.w7(32'h385ba890),
	.w8(32'hb91f01ab),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e2bce2),
	.w1(32'hb98f99d3),
	.w2(32'hb9fe54dc),
	.w3(32'hb613e290),
	.w4(32'h39e746e5),
	.w5(32'h39f985f7),
	.w6(32'h3924a2e8),
	.w7(32'h38a93de9),
	.w8(32'h3919d165),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e6648),
	.w1(32'h39118a14),
	.w2(32'hb8d47634),
	.w3(32'h3951ceee),
	.w4(32'h39944bc7),
	.w5(32'h391752c2),
	.w6(32'h3937d078),
	.w7(32'hb87d7d56),
	.w8(32'hb9ff0241),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e61c4),
	.w1(32'hb92f7641),
	.w2(32'hb81be74a),
	.w3(32'hb9284e50),
	.w4(32'hb8a4e5cb),
	.w5(32'h38861dbe),
	.w6(32'hb8baf908),
	.w7(32'h394490d8),
	.w8(32'h398cf74d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85827b5),
	.w1(32'h3a66c780),
	.w2(32'h39acd72d),
	.w3(32'h3907883f),
	.w4(32'h3a405512),
	.w5(32'h3a36b853),
	.w6(32'h3a241ab5),
	.w7(32'h39fd1494),
	.w8(32'h3a5fffbc),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f8038),
	.w1(32'h3a050086),
	.w2(32'h39988664),
	.w3(32'h3aa78b6b),
	.w4(32'h3aa89830),
	.w5(32'h3a557e02),
	.w6(32'h3ab0efac),
	.w7(32'h3a8038a5),
	.w8(32'h39e2ff6e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb813eae8),
	.w1(32'h3a9d6549),
	.w2(32'hbaf630c6),
	.w3(32'hb7a4d632),
	.w4(32'h397e9cc2),
	.w5(32'hba4ec524),
	.w6(32'h3962b203),
	.w7(32'hbaa18ee7),
	.w8(32'h3a30d359),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a069e19),
	.w1(32'h3a748e4c),
	.w2(32'h3a3d7860),
	.w3(32'h3a1b3a24),
	.w4(32'h3a9d87dd),
	.w5(32'h3a6900b5),
	.w6(32'h3a744785),
	.w7(32'h3a61c1cf),
	.w8(32'h3a667f5e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a602b),
	.w1(32'hba00f7ff),
	.w2(32'hb8fb046e),
	.w3(32'h3a07e02b),
	.w4(32'h38f3854b),
	.w5(32'h39100870),
	.w6(32'hb9178ac6),
	.w7(32'hb9891b1f),
	.w8(32'h39aeb46f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3786004b),
	.w1(32'hba6f66fa),
	.w2(32'hba7df2b4),
	.w3(32'hb91b5f80),
	.w4(32'hba2ca7f4),
	.w5(32'hba600f6d),
	.w6(32'hba210da9),
	.w7(32'hb9fed1f1),
	.w8(32'hba12567d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fccbf),
	.w1(32'hb970f64b),
	.w2(32'hb6d67eee),
	.w3(32'hba4e1a83),
	.w4(32'hb8c86991),
	.w5(32'h38ed2672),
	.w6(32'hb916942a),
	.w7(32'h3969d645),
	.w8(32'h39954e69),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8741def),
	.w1(32'h389ff754),
	.w2(32'h3908ad27),
	.w3(32'h393e0cad),
	.w4(32'h397fbef0),
	.w5(32'h396952f7),
	.w6(32'h3838ba2b),
	.w7(32'h396555d3),
	.w8(32'h3996fbd0),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39500306),
	.w1(32'h37ea9bcd),
	.w2(32'h38dc27a9),
	.w3(32'h39a218ad),
	.w4(32'h39925be3),
	.w5(32'h399dc399),
	.w6(32'hb483e4b2),
	.w7(32'h3936a301),
	.w8(32'h3985f485),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38868a55),
	.w1(32'hb9bb04f3),
	.w2(32'h398e707e),
	.w3(32'h389829f6),
	.w4(32'hb9a280b1),
	.w5(32'hb8bb4984),
	.w6(32'hb9cea16e),
	.w7(32'hb85d49e1),
	.w8(32'h39e88965),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4423d6),
	.w1(32'hb998507a),
	.w2(32'hba2172c8),
	.w3(32'h38217c88),
	.w4(32'hb8f6226a),
	.w5(32'hb9b6c287),
	.w6(32'hb912722b),
	.w7(32'hb83aa567),
	.w8(32'hba0b9bd7),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8991c08),
	.w1(32'hb8f5aa4d),
	.w2(32'h398e934c),
	.w3(32'hb9c32333),
	.w4(32'h39f1a522),
	.w5(32'h3a38cecb),
	.w6(32'h3995f498),
	.w7(32'h39d3671d),
	.w8(32'h39ebb36f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be92e0),
	.w1(32'h3a00f576),
	.w2(32'h39d44900),
	.w3(32'h3a029c5e),
	.w4(32'h3a02e415),
	.w5(32'h3a2fe93a),
	.w6(32'h39c84268),
	.w7(32'h38fe95b2),
	.w8(32'hb870e9a3),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ffcb54),
	.w1(32'h381f1bfa),
	.w2(32'h39090cdc),
	.w3(32'h39e7b92a),
	.w4(32'h398eaee5),
	.w5(32'h398888cd),
	.w6(32'h3904063a),
	.w7(32'h395757e1),
	.w8(32'h388c93af),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d2024e),
	.w1(32'h39b5d551),
	.w2(32'h3aa60e95),
	.w3(32'h38c2db29),
	.w4(32'hb9913086),
	.w5(32'h390bd86f),
	.w6(32'hb99db2cd),
	.w7(32'h3a642727),
	.w8(32'h3a25ab01),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3976794b),
	.w1(32'h3ad3c367),
	.w2(32'h3ac3dba6),
	.w3(32'h3a73eb44),
	.w4(32'h3ac21c47),
	.w5(32'h3ac6f523),
	.w6(32'h3a852562),
	.w7(32'h3ab2d75b),
	.w8(32'h3a9a200b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02d2ce),
	.w1(32'h39d76234),
	.w2(32'h39884d3c),
	.w3(32'h3ad7bbae),
	.w4(32'h3992c382),
	.w5(32'h39dd9d6e),
	.w6(32'hb7df5319),
	.w7(32'h39418823),
	.w8(32'hb99108be),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d4a0b),
	.w1(32'hbb80d0ed),
	.w2(32'hbba01ccc),
	.w3(32'h37c154ca),
	.w4(32'h3bff7aae),
	.w5(32'hbaa7b678),
	.w6(32'h3b9f2411),
	.w7(32'h3ae4e367),
	.w8(32'hbba77c05),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c9db8),
	.w1(32'hbca78308),
	.w2(32'h3adb9e1a),
	.w3(32'hbb8752b9),
	.w4(32'hbbfbf41f),
	.w5(32'hbc17d375),
	.w6(32'hbba74ee8),
	.w7(32'h3c30775f),
	.w8(32'h3c564a7c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule