module layer_10_featuremap_330(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53280c),
	.w1(32'h3aaa52d9),
	.w2(32'hbb5c04a3),
	.w3(32'hbaea8746),
	.w4(32'hbb7a9087),
	.w5(32'hbacd5005),
	.w6(32'h3c019458),
	.w7(32'hbb8a4999),
	.w8(32'hbb2c9bc3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba207e9),
	.w1(32'hbb8f75b3),
	.w2(32'hb9222b64),
	.w3(32'hbc0621e2),
	.w4(32'hbc1216a3),
	.w5(32'h3b1f7a87),
	.w6(32'h3b517130),
	.w7(32'hbba383e6),
	.w8(32'h3b9c27b4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2badd1),
	.w1(32'h3b51fc9d),
	.w2(32'h3b0200b9),
	.w3(32'hba8e0200),
	.w4(32'h3bca7e4e),
	.w5(32'h3bb3316f),
	.w6(32'hbaf2668c),
	.w7(32'h3c21760d),
	.w8(32'h3bf1e803),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3263a6),
	.w1(32'h3b8a0b18),
	.w2(32'h3ba10196),
	.w3(32'h3a37868e),
	.w4(32'h3b778f9b),
	.w5(32'h3a788b10),
	.w6(32'h3b18e6e5),
	.w7(32'h3b2be10d),
	.w8(32'h3b848950),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91dbc9),
	.w1(32'hbc2ba075),
	.w2(32'hb9bff1fd),
	.w3(32'hbbc7e7ad),
	.w4(32'hbab2ba5b),
	.w5(32'h3b41ac8b),
	.w6(32'hbb197a7c),
	.w7(32'h3b12af11),
	.w8(32'h3b8c8aa3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30d8be),
	.w1(32'h3bbd462c),
	.w2(32'hba7b9e8a),
	.w3(32'h3b9c3caa),
	.w4(32'h3b188696),
	.w5(32'hba9158c4),
	.w6(32'h3bcffa14),
	.w7(32'h3b38057d),
	.w8(32'h3a8e1666),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6815c),
	.w1(32'hbb11ea17),
	.w2(32'hbb99195e),
	.w3(32'hbb976e85),
	.w4(32'h3ad03e84),
	.w5(32'hba09cadb),
	.w6(32'hbb497554),
	.w7(32'hbb35b9e1),
	.w8(32'h3b2899e4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bb09f),
	.w1(32'hbb4d5edc),
	.w2(32'h3acbb5b5),
	.w3(32'hb9788a3b),
	.w4(32'h3c119847),
	.w5(32'h3ba30430),
	.w6(32'hbc3ae594),
	.w7(32'hbb877df7),
	.w8(32'h3b12f127),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84b53c),
	.w1(32'h3b8de2a7),
	.w2(32'h39a45b80),
	.w3(32'h3b87cba5),
	.w4(32'h3b94ef03),
	.w5(32'h3b309301),
	.w6(32'h3bbc758a),
	.w7(32'h3a1918bb),
	.w8(32'h3b21ba66),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8911ff),
	.w1(32'h3bde8232),
	.w2(32'h3b33de1c),
	.w3(32'h3c117aa1),
	.w4(32'h3b7863b5),
	.w5(32'h3c15e88a),
	.w6(32'h3c1a7b0d),
	.w7(32'h3aef6e94),
	.w8(32'h3c2c09d3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6659c4),
	.w1(32'h3b785121),
	.w2(32'h391454ed),
	.w3(32'h3b892e85),
	.w4(32'h3b910bac),
	.w5(32'h3a2dd0da),
	.w6(32'h3930c058),
	.w7(32'hba53560d),
	.w8(32'h3b86fccd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc016e4b),
	.w1(32'hb9e457f0),
	.w2(32'hbaad8d38),
	.w3(32'hbbbd1d0c),
	.w4(32'hbbb2a00a),
	.w5(32'hbbf40a73),
	.w6(32'hbc27d4bb),
	.w7(32'h3a32e982),
	.w8(32'hbbc3fa9d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf5ab2),
	.w1(32'h3b9cf505),
	.w2(32'h3a88310f),
	.w3(32'hbb3f0177),
	.w4(32'hbb9bafc2),
	.w5(32'hbb54da47),
	.w6(32'h3c40b963),
	.w7(32'hbadc5f25),
	.w8(32'h3a9507a0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadc953),
	.w1(32'h38fdbf5c),
	.w2(32'h3ba85a61),
	.w3(32'hba8dd844),
	.w4(32'h3aa1e9fb),
	.w5(32'h3acac436),
	.w6(32'h3be1354c),
	.w7(32'hb979838e),
	.w8(32'h3b1aa25a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69b5bd),
	.w1(32'h3b9fd0c9),
	.w2(32'h3b52df09),
	.w3(32'h3bcebd34),
	.w4(32'h3be97198),
	.w5(32'hbbcea018),
	.w6(32'h39c55321),
	.w7(32'h3b3476f1),
	.w8(32'hbb37c517),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe2f8f),
	.w1(32'h3c3d7c75),
	.w2(32'h3af2bdb2),
	.w3(32'hb7c867ee),
	.w4(32'h3a449d8c),
	.w5(32'h3b17b907),
	.w6(32'h3c96da33),
	.w7(32'hbba0afdf),
	.w8(32'h3b577bf4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a0c4c),
	.w1(32'h3c145620),
	.w2(32'hbabe9e72),
	.w3(32'hbb9b2190),
	.w4(32'hbb419e9c),
	.w5(32'h3aa04ee0),
	.w6(32'h3b974298),
	.w7(32'hb9f29c65),
	.w8(32'h3b015ecd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad775c5),
	.w1(32'h3b6e8846),
	.w2(32'hbaca546c),
	.w3(32'h3aeaae2b),
	.w4(32'h3a9db737),
	.w5(32'h3abb0d7a),
	.w6(32'h3bad425b),
	.w7(32'hbb05d596),
	.w8(32'h3b00ad07),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d0e0),
	.w1(32'hba2a4ae5),
	.w2(32'h3b423ca8),
	.w3(32'hbade8ff9),
	.w4(32'h3b0c97f5),
	.w5(32'h3ab9f541),
	.w6(32'hbb053df2),
	.w7(32'h3a004cca),
	.w8(32'h3b473a12),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a383bb2),
	.w1(32'hb96f3f4a),
	.w2(32'hba9a22f8),
	.w3(32'hbaa2b503),
	.w4(32'h3b64a37a),
	.w5(32'hbbd41886),
	.w6(32'h3b1d46e0),
	.w7(32'h3a978065),
	.w8(32'hbbb0936d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8ca1b),
	.w1(32'h3c2d4eeb),
	.w2(32'hbb48dcd7),
	.w3(32'hbad07355),
	.w4(32'hbc06d4bc),
	.w5(32'h3b6b3771),
	.w6(32'h3cda6587),
	.w7(32'hbb9c83ce),
	.w8(32'h3b380970),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a9905),
	.w1(32'hbb65efc7),
	.w2(32'h3afb14e5),
	.w3(32'hbb03d47a),
	.w4(32'h38fb90b4),
	.w5(32'hba9edcf4),
	.w6(32'hbbdbf466),
	.w7(32'hb9751cb2),
	.w8(32'h3ba33285),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd000f1),
	.w1(32'h3a9986ec),
	.w2(32'h3baa055b),
	.w3(32'h3b4f99a2),
	.w4(32'h3a8e5552),
	.w5(32'hbac76084),
	.w6(32'hbb130f1c),
	.w7(32'h3aa4c822),
	.w8(32'h3bc66803),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ce196),
	.w1(32'h3a0a77d7),
	.w2(32'hbb2a9a5b),
	.w3(32'h3c005cf1),
	.w4(32'h3b8da3f2),
	.w5(32'h3b9dede4),
	.w6(32'h3c8d7bea),
	.w7(32'hbbf3cb74),
	.w8(32'h3a12c767),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb777dc),
	.w1(32'hbab50bad),
	.w2(32'h3b31e3a1),
	.w3(32'h3b02c087),
	.w4(32'hbb617bef),
	.w5(32'hbbb2d0a2),
	.w6(32'hb8c72ae5),
	.w7(32'h3b83d824),
	.w8(32'hbb97684b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4420ba),
	.w1(32'h3b5c4c2b),
	.w2(32'hbb385bda),
	.w3(32'h3b3b183a),
	.w4(32'hbb0d564b),
	.w5(32'hbab8fcc5),
	.w6(32'h3b7de5fa),
	.w7(32'hbb66a5ed),
	.w8(32'hbb2645ff),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab32010),
	.w1(32'hbad98ac6),
	.w2(32'hbada7e01),
	.w3(32'hbadbd1c9),
	.w4(32'h3ad29e05),
	.w5(32'hb95c9cad),
	.w6(32'hbb87e75e),
	.w7(32'h393f7adb),
	.w8(32'hbb61defe),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb971cfc),
	.w1(32'h3b84e56f),
	.w2(32'h3b1128cb),
	.w3(32'h3bea3074),
	.w4(32'hba889ae8),
	.w5(32'h39be672b),
	.w6(32'h3c9ebbe1),
	.w7(32'h3b94c098),
	.w8(32'h3ae9d134),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb448463),
	.w1(32'hbb88f186),
	.w2(32'hbb1ba122),
	.w3(32'hbb94ec68),
	.w4(32'hbbb69470),
	.w5(32'hbb2a9eef),
	.w6(32'h39683dfe),
	.w7(32'hbb26eb35),
	.w8(32'hbb84d7d8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ac76c),
	.w1(32'h39ad9690),
	.w2(32'h3b23cac2),
	.w3(32'h3b866045),
	.w4(32'hbbd362b7),
	.w5(32'h3a71016e),
	.w6(32'h3c634ccb),
	.w7(32'hbaf03dfe),
	.w8(32'hbbb81ed1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa53a45),
	.w1(32'hbc386ec1),
	.w2(32'h3a8a9ff9),
	.w3(32'h3c464643),
	.w4(32'hbadae9e5),
	.w5(32'hbaee13bb),
	.w6(32'hbbdb5d88),
	.w7(32'hba55fea8),
	.w8(32'h3baa0822),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7c1fc),
	.w1(32'h3b1dcb49),
	.w2(32'hbba03671),
	.w3(32'hbb8e62cb),
	.w4(32'hbab60439),
	.w5(32'hbbd1c704),
	.w6(32'hbc14bcc4),
	.w7(32'h3ab13dc9),
	.w8(32'hbac41230),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbe594),
	.w1(32'hbb370cf8),
	.w2(32'h3a3b1fe2),
	.w3(32'hbbad9ece),
	.w4(32'hbb43bc80),
	.w5(32'hbb05d0da),
	.w6(32'hbba1510d),
	.w7(32'hbb9cd03b),
	.w8(32'hbb2b9b45),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3975e3ba),
	.w1(32'hba8a0af7),
	.w2(32'hbb8d8725),
	.w3(32'hb973fc52),
	.w4(32'hbbf5766f),
	.w5(32'h3b2b4ac4),
	.w6(32'h3bbbff43),
	.w7(32'hbbb5ec8f),
	.w8(32'hb9845f1d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee292c),
	.w1(32'hbbb9e9b1),
	.w2(32'hba8d5067),
	.w3(32'hbb5454fc),
	.w4(32'hbb3d53fa),
	.w5(32'hbb8ae512),
	.w6(32'hbbd2ffae),
	.w7(32'h3a9d3aa8),
	.w8(32'hba405c24),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85c5c7),
	.w1(32'hbbc53507),
	.w2(32'hbbd7bb30),
	.w3(32'hbbefe0f1),
	.w4(32'hba3662aa),
	.w5(32'hbba36d7f),
	.w6(32'h3bf72723),
	.w7(32'hbb92c7a5),
	.w8(32'hbb474cf9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f0f4e),
	.w1(32'hbafd2f7a),
	.w2(32'h3b8af3f9),
	.w3(32'hba656661),
	.w4(32'hbbe8f63b),
	.w5(32'h3b814a6e),
	.w6(32'hbb6df9f7),
	.w7(32'h3b1b8d42),
	.w8(32'hbb89954c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84f3a0),
	.w1(32'hba8b23df),
	.w2(32'h3add742a),
	.w3(32'hbafd10f9),
	.w4(32'h3b85dde0),
	.w5(32'hbb94b140),
	.w6(32'hbaa05841),
	.w7(32'hbb1aa083),
	.w8(32'hbba0049e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab896a),
	.w1(32'hbc371e13),
	.w2(32'hbbb98fb6),
	.w3(32'h3a404329),
	.w4(32'hbbb99e07),
	.w5(32'hbaba6bf8),
	.w6(32'hbbed5893),
	.w7(32'hbb8f0b60),
	.w8(32'h3a5dfcfa),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7d5f9),
	.w1(32'h3a96f76a),
	.w2(32'h3ad848b7),
	.w3(32'h3b544a3d),
	.w4(32'h3a1f3641),
	.w5(32'h38a1e5d4),
	.w6(32'h3b0159fa),
	.w7(32'hba5d314f),
	.w8(32'h3b992516),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb261b26),
	.w1(32'hbb0df498),
	.w2(32'h3bceecde),
	.w3(32'hbae2b808),
	.w4(32'hbb242216),
	.w5(32'hbaf996d1),
	.w6(32'hbbd9accb),
	.w7(32'h3b92e56b),
	.w8(32'hba7f50ef),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31150e),
	.w1(32'h3a5c3208),
	.w2(32'hbb9e3e04),
	.w3(32'h3aadb884),
	.w4(32'hb961b3e8),
	.w5(32'hb9d51e47),
	.w6(32'hba89f49a),
	.w7(32'hbafe082a),
	.w8(32'hbb3a2e48),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98d0a5),
	.w1(32'hbb28e7e3),
	.w2(32'h3b7edb58),
	.w3(32'hba20cc9f),
	.w4(32'h3b751f65),
	.w5(32'h3b18acd5),
	.w6(32'h3b4a7343),
	.w7(32'h3b817701),
	.w8(32'hb9456a5c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad1f7c),
	.w1(32'h3b1a5007),
	.w2(32'h3ba9e3c4),
	.w3(32'h3c167632),
	.w4(32'h3b7611b6),
	.w5(32'hba3e8e1c),
	.w6(32'h39c2a84d),
	.w7(32'h3ace97bd),
	.w8(32'hbbb14042),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e745d),
	.w1(32'hbb242951),
	.w2(32'hb9ca3c99),
	.w3(32'h3b7b79f9),
	.w4(32'h3b29db5e),
	.w5(32'h3b0c866b),
	.w6(32'hba2ee8f6),
	.w7(32'h3916b97f),
	.w8(32'h3b2c3e79),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4066c1),
	.w1(32'h3c2daf97),
	.w2(32'h3b0ebcf0),
	.w3(32'h3bc05294),
	.w4(32'h3a133376),
	.w5(32'h3afbcec7),
	.w6(32'hbb07a093),
	.w7(32'hbacfb444),
	.w8(32'h3a517fa9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ed502),
	.w1(32'h3a43cd96),
	.w2(32'hbb4cce92),
	.w3(32'h3a7cf1c4),
	.w4(32'hbb342f53),
	.w5(32'h3b8ea8a6),
	.w6(32'h3957795c),
	.w7(32'hbb9eb313),
	.w8(32'h3bc57ead),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34b744),
	.w1(32'hb9bbc877),
	.w2(32'h3baf2449),
	.w3(32'hb94aaaa3),
	.w4(32'h3b66873f),
	.w5(32'h3b3fc661),
	.w6(32'hbac88cbb),
	.w7(32'h3bbda9bb),
	.w8(32'h3a2cf6d9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27b74e),
	.w1(32'h3bd5d0d6),
	.w2(32'h39ff4d7e),
	.w3(32'h3c0e0c70),
	.w4(32'h39ca6f6a),
	.w5(32'h3b93a618),
	.w6(32'h3c5bc3ee),
	.w7(32'hb9d4c3f2),
	.w8(32'h3b505dc8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ae068),
	.w1(32'hbb7bbea9),
	.w2(32'h3b372507),
	.w3(32'hbb11ef50),
	.w4(32'h3b3b3e43),
	.w5(32'hbb44337e),
	.w6(32'hbc1fa33f),
	.w7(32'h39432933),
	.w8(32'h39b2d435),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0997e),
	.w1(32'hbbc26845),
	.w2(32'hbbbcd9f4),
	.w3(32'hbc185c19),
	.w4(32'hbb94f7dd),
	.w5(32'hba2f03f2),
	.w6(32'hbbf70c80),
	.w7(32'hbbc1a8c7),
	.w8(32'h3b2a2e6c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c6646),
	.w1(32'hbb405bfe),
	.w2(32'h3b48987a),
	.w3(32'hb8d69bea),
	.w4(32'h3b65a3c9),
	.w5(32'hbad68df9),
	.w6(32'hbadb9c8b),
	.w7(32'h3a11a325),
	.w8(32'hba5150e0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a1408),
	.w1(32'hbab873dc),
	.w2(32'hb701c060),
	.w3(32'h3ab63645),
	.w4(32'h3a0ed384),
	.w5(32'hbbf0e3bf),
	.w6(32'hbb155a46),
	.w7(32'hbb2a77a5),
	.w8(32'h3abf816f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b711957),
	.w1(32'hbb277ffb),
	.w2(32'h3b810dc8),
	.w3(32'hbb04f291),
	.w4(32'h3b7004cf),
	.w5(32'h3b1b42e6),
	.w6(32'hbbeba579),
	.w7(32'h3bcac5c6),
	.w8(32'h3b1ec4e2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2d0fd),
	.w1(32'hbaec3434),
	.w2(32'hbb7ec4e5),
	.w3(32'h3aa75ced),
	.w4(32'h3a1b9cf2),
	.w5(32'h3a809bac),
	.w6(32'h3a603ff6),
	.w7(32'hbae6ee18),
	.w8(32'h3ba0a537),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83c646),
	.w1(32'hbb5d95fa),
	.w2(32'hbb1663ac),
	.w3(32'hbb537e94),
	.w4(32'h38d750b5),
	.w5(32'h3bb33517),
	.w6(32'h3b64b3a1),
	.w7(32'h3ae42a93),
	.w8(32'h3beb970f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc71f0),
	.w1(32'h3a98ac47),
	.w2(32'h3b5d9ad8),
	.w3(32'h3ae53796),
	.w4(32'h398d46fb),
	.w5(32'h3a341b68),
	.w6(32'h3a391a76),
	.w7(32'h3b8255c8),
	.w8(32'h3aaed6f1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb099863),
	.w1(32'hbb006676),
	.w2(32'h3b4d7d62),
	.w3(32'hbb41ad87),
	.w4(32'h389c5181),
	.w5(32'h3b322067),
	.w6(32'h3a47a406),
	.w7(32'h3be72091),
	.w8(32'h3b68e567),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b986275),
	.w1(32'hbb5142d0),
	.w2(32'h3aeb864d),
	.w3(32'hba55744c),
	.w4(32'h3b89edaa),
	.w5(32'h3c109501),
	.w6(32'hbbc168dc),
	.w7(32'hb82ac797),
	.w8(32'hba9b0522),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cd5e05),
	.w1(32'hbc69e684),
	.w2(32'h3be02c89),
	.w3(32'hba8516d9),
	.w4(32'h3c592f2a),
	.w5(32'hbb2c96fc),
	.w6(32'hbca061b1),
	.w7(32'h3b871d1e),
	.w8(32'hba85aed5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b718160),
	.w1(32'hbb9c1847),
	.w2(32'hbb7b4da9),
	.w3(32'h3c06acb1),
	.w4(32'h398d78ef),
	.w5(32'hb94f4774),
	.w6(32'hbb3b3121),
	.w7(32'hbb4627bd),
	.w8(32'hb9caf9ce),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c56fe),
	.w1(32'h3b0efb9c),
	.w2(32'h3a8ced9c),
	.w3(32'h3a7d764e),
	.w4(32'hbaadb09e),
	.w5(32'hba180bcd),
	.w6(32'h3c06a625),
	.w7(32'hbb6c8b02),
	.w8(32'hba90c157),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac438e2),
	.w1(32'hbba75de5),
	.w2(32'hb9510956),
	.w3(32'hbaf2b27c),
	.w4(32'hbb26f4d9),
	.w5(32'h3b043297),
	.w6(32'h38c62ba0),
	.w7(32'h3b86eabf),
	.w8(32'h399d159c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5099d8),
	.w1(32'hbbcedded),
	.w2(32'hba52d338),
	.w3(32'hbb5c9050),
	.w4(32'h3a12e9c3),
	.w5(32'h3b481bd9),
	.w6(32'hbb67999b),
	.w7(32'h3ac64f5d),
	.w8(32'h39a0cfe7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad959f),
	.w1(32'hbbabe681),
	.w2(32'hbb5277f0),
	.w3(32'hbb111df9),
	.w4(32'h3a324602),
	.w5(32'h3b78027b),
	.w6(32'h39dd3618),
	.w7(32'hbb184c4e),
	.w8(32'h3b80c227),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb674cb),
	.w1(32'hbbbe5857),
	.w2(32'h392aab31),
	.w3(32'h3b4d052e),
	.w4(32'hb9c6a537),
	.w5(32'hbaac2746),
	.w6(32'hbb612da3),
	.w7(32'h3a8d11d9),
	.w8(32'h3adc0eb9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83aec5),
	.w1(32'h3be5133e),
	.w2(32'hba8fbfff),
	.w3(32'hbb856122),
	.w4(32'h3b990bd8),
	.w5(32'hbaf95b1b),
	.w6(32'hbb8aefe3),
	.w7(32'h3be8f1a1),
	.w8(32'h3b0a5b60),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea04bb),
	.w1(32'h3c99fc91),
	.w2(32'h3b776e97),
	.w3(32'h3c653ae2),
	.w4(32'h3c0aa466),
	.w5(32'h3b6b829f),
	.w6(32'h3c6a0b53),
	.w7(32'h3b9b629c),
	.w8(32'h3ba0fa07),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd57255),
	.w1(32'h3b3d9145),
	.w2(32'hbb62b09e),
	.w3(32'hbb2ba4fa),
	.w4(32'hb75d2ac6),
	.w5(32'hbbccf36b),
	.w6(32'h3b6d8d24),
	.w7(32'hbacd42fa),
	.w8(32'hbba90555),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf447ee),
	.w1(32'hba12c561),
	.w2(32'h380baf4d),
	.w3(32'hb9f84c3c),
	.w4(32'hbbcf70d1),
	.w5(32'h3a45fc2b),
	.w6(32'h3b84de2c),
	.w7(32'hbb85835d),
	.w8(32'h3baf1ee3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02529a),
	.w1(32'hbabf5728),
	.w2(32'h3a7940bb),
	.w3(32'hbaddc02a),
	.w4(32'h3b30ed5d),
	.w5(32'hbc1d55dd),
	.w6(32'hbb904089),
	.w7(32'hb97b84f5),
	.w8(32'hbbfca4a9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edbc29),
	.w1(32'h3c0e1e9f),
	.w2(32'hbc2de099),
	.w3(32'h3bcb0037),
	.w4(32'hba13c534),
	.w5(32'hbbebb8d3),
	.w6(32'h3cb6bd0f),
	.w7(32'hbc45c02e),
	.w8(32'h3b6c8966),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c69c0),
	.w1(32'hbc5b8a20),
	.w2(32'hbbd83598),
	.w3(32'hbbb8f3c6),
	.w4(32'h3b77cab7),
	.w5(32'hbb2c1e45),
	.w6(32'h3c504d91),
	.w7(32'h3b215273),
	.w8(32'hbbe1867a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4b7a6),
	.w1(32'hbc089d00),
	.w2(32'h3a3a9cef),
	.w3(32'h3b5add46),
	.w4(32'hbc0bd13c),
	.w5(32'hbb8f369e),
	.w6(32'h3be3f3d9),
	.w7(32'h3b7a2d24),
	.w8(32'h3ac6fd86),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae83623),
	.w1(32'h3b9545f2),
	.w2(32'h3b067355),
	.w3(32'hbb32c9eb),
	.w4(32'h3ae2e818),
	.w5(32'hb95f998a),
	.w6(32'hbb8685fd),
	.w7(32'h3c0c9e3a),
	.w8(32'hba0e4881),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd411b3),
	.w1(32'h3b542f55),
	.w2(32'h3a7d53af),
	.w3(32'h3b0d4c15),
	.w4(32'hbb0b0175),
	.w5(32'h3bd9d26a),
	.w6(32'h3c3a3317),
	.w7(32'h390a3f76),
	.w8(32'h3c2228a1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb353bac),
	.w1(32'h3b034cc7),
	.w2(32'h3c078958),
	.w3(32'h3b8a5002),
	.w4(32'h3b8ecb42),
	.w5(32'h3a28958b),
	.w6(32'hbc074568),
	.w7(32'h3a965714),
	.w8(32'hbac0f5d2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba27a7),
	.w1(32'hbbc877e1),
	.w2(32'hb98bb56e),
	.w3(32'hbb4bd48a),
	.w4(32'h3b31fd34),
	.w5(32'h3b4b2385),
	.w6(32'hbbabdab8),
	.w7(32'hbaea9e65),
	.w8(32'h3bafc23c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1998d4),
	.w1(32'h3b91132c),
	.w2(32'h3b4957a9),
	.w3(32'h3ae0ba34),
	.w4(32'h3bbbed9e),
	.w5(32'hbb54ea81),
	.w6(32'h3ba5119d),
	.w7(32'h3bb66d56),
	.w8(32'h3a58ea80),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917421c),
	.w1(32'h3c137fd6),
	.w2(32'hbaaae100),
	.w3(32'h3a88c18c),
	.w4(32'hb9c6cc77),
	.w5(32'h3b54dce5),
	.w6(32'h3ba44311),
	.w7(32'h3b766561),
	.w8(32'hbac21a98),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc23109),
	.w1(32'h3aa06317),
	.w2(32'h3b812369),
	.w3(32'h3c412f98),
	.w4(32'h3bb8dcb5),
	.w5(32'h39270a58),
	.w6(32'h3b994510),
	.w7(32'h3b851eab),
	.w8(32'hbb177ab2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d3b42),
	.w1(32'hbb17cb17),
	.w2(32'h3ab82a8e),
	.w3(32'h3b2e5613),
	.w4(32'hbb08f321),
	.w5(32'h3b48168c),
	.w6(32'h3bfb5a3c),
	.w7(32'h3b32364c),
	.w8(32'h3a882636),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f4f4b),
	.w1(32'hbaa67c32),
	.w2(32'hb995e19f),
	.w3(32'hbb4bf16e),
	.w4(32'h3b3baf38),
	.w5(32'h3bfddfaa),
	.w6(32'hbb89edaf),
	.w7(32'hbaf08a72),
	.w8(32'h3c3624d7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37b180),
	.w1(32'h3c3ce30f),
	.w2(32'h3c35526e),
	.w3(32'h3c76a99c),
	.w4(32'h3c2477fe),
	.w5(32'h39f96f39),
	.w6(32'h3c7cd7d7),
	.w7(32'h3c013363),
	.w8(32'h3a30f2e5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23584a),
	.w1(32'h3a8bc765),
	.w2(32'h38b59dc7),
	.w3(32'hbae88833),
	.w4(32'h3aff7878),
	.w5(32'h3b20b100),
	.w6(32'hbaa07aab),
	.w7(32'h3abafbfe),
	.w8(32'hba333f5d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5327fc),
	.w1(32'h3be9677d),
	.w2(32'hbb765e6a),
	.w3(32'h3b931994),
	.w4(32'h3b6da907),
	.w5(32'hbb954472),
	.w6(32'hbbd77a08),
	.w7(32'hba76bb9f),
	.w8(32'hba934bcd),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395572fb),
	.w1(32'h38c7245e),
	.w2(32'hb9a686ee),
	.w3(32'hbba09fb2),
	.w4(32'h3b7bf134),
	.w5(32'h3b9258cf),
	.w6(32'hbb16d660),
	.w7(32'h3b5ea34c),
	.w8(32'h3b0f13d6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8714f3),
	.w1(32'hbbae6f5f),
	.w2(32'h3a236e57),
	.w3(32'h3b85555c),
	.w4(32'hb99af33f),
	.w5(32'h3b0be139),
	.w6(32'hbb215801),
	.w7(32'hb823bc3f),
	.w8(32'h3b803629),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9f625),
	.w1(32'h3bc336a2),
	.w2(32'h39a37d08),
	.w3(32'h3b83df33),
	.w4(32'h3ad51c6e),
	.w5(32'hbacde25b),
	.w6(32'hb9d10f48),
	.w7(32'hbb4c0441),
	.w8(32'hbb786139),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e4d5d),
	.w1(32'h3c89cb53),
	.w2(32'hbc6d6c3d),
	.w3(32'hbb3ebf1f),
	.w4(32'hbc8a53b4),
	.w5(32'hbbb426c3),
	.w6(32'h3c953eec),
	.w7(32'hbc2dbcc1),
	.w8(32'h3c47c5b1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f1c9d),
	.w1(32'hba3bf398),
	.w2(32'hbbc41f0f),
	.w3(32'hbbd30d67),
	.w4(32'hbbb23cf1),
	.w5(32'hbb5536de),
	.w6(32'hbb66e667),
	.w7(32'hba2151b7),
	.w8(32'hb98d0226),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b917014),
	.w1(32'h3c09c914),
	.w2(32'hbaa5a513),
	.w3(32'hbadc2c79),
	.w4(32'hbb6a33f3),
	.w5(32'hbb45f51d),
	.w6(32'h3b836a88),
	.w7(32'hbb927b1d),
	.w8(32'h3b409d99),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02fec9),
	.w1(32'hbadaec98),
	.w2(32'hbb98b396),
	.w3(32'hbc101c7d),
	.w4(32'hbac3333d),
	.w5(32'h3b0f1cc3),
	.w6(32'hbb8bf29d),
	.w7(32'hbb80eff8),
	.w8(32'h3b17cea4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee4070),
	.w1(32'hbaf99bdc),
	.w2(32'h3a4f9b2e),
	.w3(32'hb94f2041),
	.w4(32'h3aea9a91),
	.w5(32'hbbc43ecb),
	.w6(32'hbb014e79),
	.w7(32'h398a5529),
	.w8(32'hbb9b8aaa),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaef89),
	.w1(32'h39c30082),
	.w2(32'hbb9f23e9),
	.w3(32'h3a139ce4),
	.w4(32'h3a14901e),
	.w5(32'hb9c4cd88),
	.w6(32'h3c0e3b17),
	.w7(32'hbbebe87a),
	.w8(32'h3af83bcc),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f1f81),
	.w1(32'h3b49f175),
	.w2(32'h3a9a96c8),
	.w3(32'hbbdd4940),
	.w4(32'h3b2d414f),
	.w5(32'h3ac1c295),
	.w6(32'hbbe4c265),
	.w7(32'hb98387e9),
	.w8(32'h3bc0c997),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac266b1),
	.w1(32'hbb36325d),
	.w2(32'h3c1fba48),
	.w3(32'h39e8632e),
	.w4(32'h3b9b864c),
	.w5(32'h3b9b7f6b),
	.w6(32'h3a031a1d),
	.w7(32'h3c19d881),
	.w8(32'h3c031c5e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c518636),
	.w1(32'h3962e8a9),
	.w2(32'h3b3cf87d),
	.w3(32'h3c2067e8),
	.w4(32'hbb089542),
	.w5(32'h3b01cc1c),
	.w6(32'hbba16f36),
	.w7(32'hbbe2dbdc),
	.w8(32'hb97d5952),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf92a79),
	.w1(32'hba2df75d),
	.w2(32'hbba7df6a),
	.w3(32'hbb290e92),
	.w4(32'hbb8e1ac6),
	.w5(32'hbbc66caf),
	.w6(32'hbb8a2ad7),
	.w7(32'hbb738ec8),
	.w8(32'hba320753),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2a30b),
	.w1(32'h3a5976ff),
	.w2(32'hbb05691f),
	.w3(32'hbbef75b4),
	.w4(32'h3926101e),
	.w5(32'h3c004f01),
	.w6(32'h3b36e378),
	.w7(32'hbb11163e),
	.w8(32'h39c04c56),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c116da0),
	.w1(32'hba13cc4b),
	.w2(32'h3be869e6),
	.w3(32'h3c822de5),
	.w4(32'hbb4aab78),
	.w5(32'h3b56ffb9),
	.w6(32'h3baf5d45),
	.w7(32'hba9fc7a8),
	.w8(32'hbb52e85c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedeed0),
	.w1(32'h3b757973),
	.w2(32'h3bb0650c),
	.w3(32'h3c071a0a),
	.w4(32'h3b643a18),
	.w5(32'h3c248eae),
	.w6(32'h3baeca80),
	.w7(32'hbb8ca03e),
	.w8(32'h3b81d4fc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c9896),
	.w1(32'h3b20ca6f),
	.w2(32'hbb1f0281),
	.w3(32'h3a9ee988),
	.w4(32'hb90200d2),
	.w5(32'h3b01819a),
	.w6(32'h3b22fdc0),
	.w7(32'h39b388b6),
	.w8(32'hbae65b22),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38887986),
	.w1(32'hbb46902b),
	.w2(32'h38dd21e2),
	.w3(32'h3b93d831),
	.w4(32'hbaed8d54),
	.w5(32'h3b0aab20),
	.w6(32'hbab0f3f7),
	.w7(32'hbb02afcd),
	.w8(32'hbc4a7f4a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02c964),
	.w1(32'h3c5866c9),
	.w2(32'h3b5bbbd5),
	.w3(32'h3bd7aa89),
	.w4(32'h3b3dc285),
	.w5(32'h3a642c56),
	.w6(32'hbc3b4476),
	.w7(32'hbc7ea4a1),
	.w8(32'hbadb9f73),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4beb59),
	.w1(32'hb99a4bec),
	.w2(32'h3ab13917),
	.w3(32'hbaf33b3d),
	.w4(32'hb92270fc),
	.w5(32'h3bb6e953),
	.w6(32'h3b8db5be),
	.w7(32'h3abb17e4),
	.w8(32'hbb89df2e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb94e70),
	.w1(32'hb982a089),
	.w2(32'hbba51d11),
	.w3(32'hba93e6fe),
	.w4(32'hbb3d32d8),
	.w5(32'h3b693d18),
	.w6(32'h3b2ce051),
	.w7(32'h3a4c0f2c),
	.w8(32'h3bcb47cc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24f219),
	.w1(32'hbb5501d9),
	.w2(32'hbacaf0b5),
	.w3(32'hba1a6c22),
	.w4(32'h3aa55601),
	.w5(32'h3b87d539),
	.w6(32'h3b57c3ac),
	.w7(32'h3a74cfca),
	.w8(32'hba7ad3b4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f73328),
	.w1(32'hbb238b64),
	.w2(32'hbbc39ba4),
	.w3(32'h3be86076),
	.w4(32'hb9e9ac03),
	.w5(32'hbb2b221c),
	.w6(32'hbb341c7b),
	.w7(32'hbbc1fe84),
	.w8(32'h3c07f008),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be75781),
	.w1(32'h3b8624be),
	.w2(32'h3b4a3a96),
	.w3(32'h3b8f1fc9),
	.w4(32'h3b1381b6),
	.w5(32'hbb4c93a5),
	.w6(32'h3c10eb72),
	.w7(32'hb9e24cdf),
	.w8(32'h3b424d25),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9884cb),
	.w1(32'hbb897beb),
	.w2(32'hba1f206d),
	.w3(32'hbb3d9865),
	.w4(32'h3a87fef5),
	.w5(32'h3b0efc3a),
	.w6(32'h3c2b91c3),
	.w7(32'hba0ae296),
	.w8(32'h3ab64592),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b131376),
	.w1(32'hbaf35a91),
	.w2(32'hbb1df233),
	.w3(32'h3b98568f),
	.w4(32'h3a4ac559),
	.w5(32'h3b458949),
	.w6(32'h3af2129e),
	.w7(32'hbb28a17b),
	.w8(32'hb9c86017),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb209b1),
	.w1(32'h3c017681),
	.w2(32'h3ab26f84),
	.w3(32'hba12c9c4),
	.w4(32'h3aba7b22),
	.w5(32'h3b92854d),
	.w6(32'h3a3af022),
	.w7(32'hba76e579),
	.w8(32'hbb33ce18),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7539e),
	.w1(32'h3b7c90b0),
	.w2(32'h3b4e4bb6),
	.w3(32'h3b827371),
	.w4(32'h3b2b5eb6),
	.w5(32'hbb0e09ef),
	.w6(32'h3b93ac03),
	.w7(32'h3b2a4731),
	.w8(32'h3b4a7f8d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb1e85),
	.w1(32'hbb912252),
	.w2(32'hbb492a1f),
	.w3(32'h3b6e1afc),
	.w4(32'h3b4474a8),
	.w5(32'hbabb9ba2),
	.w6(32'hbb9e7ecc),
	.w7(32'hbba443b1),
	.w8(32'hbac329fa),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25305d),
	.w1(32'hbb92d01e),
	.w2(32'hbac0fcdf),
	.w3(32'hbb7c203e),
	.w4(32'hba43d39b),
	.w5(32'h3b8b2dec),
	.w6(32'h3b76c4ba),
	.w7(32'h3a903c19),
	.w8(32'h3ae355a8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0373a8),
	.w1(32'hb9369d76),
	.w2(32'h3bb2de0e),
	.w3(32'h3b46cb35),
	.w4(32'h3b245fd1),
	.w5(32'h3af9f100),
	.w6(32'hbc230f55),
	.w7(32'hbb24d2b1),
	.w8(32'hbc0d85f5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ae2ac),
	.w1(32'hbb6d0e1d),
	.w2(32'hbbf92f34),
	.w3(32'h3b422edb),
	.w4(32'h3aae84ec),
	.w5(32'h3ad036a7),
	.w6(32'hbba2f950),
	.w7(32'hbb1383c3),
	.w8(32'hbae90708),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c4def),
	.w1(32'hbafc8dc9),
	.w2(32'hbb4ee5b5),
	.w3(32'h3b02909a),
	.w4(32'hbaecf005),
	.w5(32'hba7d6bf8),
	.w6(32'hbbb90f98),
	.w7(32'hbb406b8a),
	.w8(32'hbbab289d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab8a6e),
	.w1(32'hbbbb2cfa),
	.w2(32'hbc09e279),
	.w3(32'h3b2646cd),
	.w4(32'hbbecffce),
	.w5(32'hbb67d433),
	.w6(32'hbc3483ed),
	.w7(32'hbbe6b1be),
	.w8(32'hbac1e676),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5f387),
	.w1(32'h3b1d6bc5),
	.w2(32'hba93aeae),
	.w3(32'hbb46dd5e),
	.w4(32'hbbaddc66),
	.w5(32'h3b104b65),
	.w6(32'hbabb020f),
	.w7(32'hbb9f8e27),
	.w8(32'hbabfc8ce),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c0b50),
	.w1(32'hbad06cbf),
	.w2(32'hbc0e7e7f),
	.w3(32'hbbdf6e12),
	.w4(32'h3a98ef66),
	.w5(32'hbc779da7),
	.w6(32'hbaae0bbb),
	.w7(32'hbbcad88a),
	.w8(32'hbc3a3e9d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0b29b),
	.w1(32'hba898c00),
	.w2(32'h3bf63938),
	.w3(32'hbc52655b),
	.w4(32'hbc5321ef),
	.w5(32'h3985b176),
	.w6(32'h3cf4fea6),
	.w7(32'h3c39015e),
	.w8(32'h3be86f3a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c7ac6),
	.w1(32'h3bace97f),
	.w2(32'hbbac75f4),
	.w3(32'hbac7b8ba),
	.w4(32'h3bb8a394),
	.w5(32'hbc7a6c52),
	.w6(32'h3b32f2d9),
	.w7(32'h3b186d7c),
	.w8(32'h3a4f069c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aa36b),
	.w1(32'hba60f4eb),
	.w2(32'h3b261310),
	.w3(32'hbc930e38),
	.w4(32'hbc40d8bf),
	.w5(32'h3997f1f2),
	.w6(32'h3d12fae5),
	.w7(32'h3c4c4b5a),
	.w8(32'hbb9a1720),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d8f59),
	.w1(32'hb9d973f6),
	.w2(32'hb90e0fa6),
	.w3(32'hba6c1f8f),
	.w4(32'hba53fab7),
	.w5(32'hba2407e7),
	.w6(32'h39bc8f17),
	.w7(32'hbaef2331),
	.w8(32'h3b2ef146),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6e84e),
	.w1(32'hbb9f0579),
	.w2(32'hbbbca4d4),
	.w3(32'hbb145855),
	.w4(32'hbbb61269),
	.w5(32'hbae0f955),
	.w6(32'h3c4fe5e7),
	.w7(32'h3b4ce931),
	.w8(32'h39cf0612),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb178d70),
	.w1(32'hbb01bc12),
	.w2(32'hbb013363),
	.w3(32'hbb0610e4),
	.w4(32'hb98a4976),
	.w5(32'h3bbf78ad),
	.w6(32'hbb777041),
	.w7(32'hbb46fa84),
	.w8(32'h3ad091ea),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be393d5),
	.w1(32'h3bae3b5a),
	.w2(32'h3b2fb3a6),
	.w3(32'h3ac1cf79),
	.w4(32'hbb09d888),
	.w5(32'h3b32c996),
	.w6(32'h3be2c275),
	.w7(32'h3b0cc4bd),
	.w8(32'hbb3affcc),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9f0b3),
	.w1(32'hbba0e75d),
	.w2(32'hbb7415ee),
	.w3(32'hba80ae23),
	.w4(32'h3af41eb4),
	.w5(32'h3b6665d6),
	.w6(32'h3b6168e7),
	.w7(32'hbb5ec4e6),
	.w8(32'hba3b3a16),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93d333),
	.w1(32'h3b043ccf),
	.w2(32'hbb0d1641),
	.w3(32'h398f5fa1),
	.w4(32'hba3f8aef),
	.w5(32'hbb3591a4),
	.w6(32'h3b3e43f4),
	.w7(32'h3ba194c7),
	.w8(32'h393f0e9c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba380dfd),
	.w1(32'h39e3c6a2),
	.w2(32'h3b851441),
	.w3(32'h3b49002a),
	.w4(32'h3b72c4ff),
	.w5(32'hbb2f4ed8),
	.w6(32'hb9b5bdb4),
	.w7(32'h3b84c3fa),
	.w8(32'hbc296b90),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc522b),
	.w1(32'h3a9a4983),
	.w2(32'h3b8cd9f4),
	.w3(32'h3ac2f893),
	.w4(32'hbb011adb),
	.w5(32'hbba00c9d),
	.w6(32'h3a3ea98a),
	.w7(32'hbaac9529),
	.w8(32'h3a308400),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d4f07),
	.w1(32'h3ae9a76f),
	.w2(32'h3be00a19),
	.w3(32'hbbb27eb0),
	.w4(32'hbadff4e0),
	.w5(32'h3b6835e4),
	.w6(32'h3c2f5e9d),
	.w7(32'h3b718cd0),
	.w8(32'h3925965d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f1581),
	.w1(32'h38d8d340),
	.w2(32'h3a95c4d7),
	.w3(32'hbab77c0f),
	.w4(32'hbb3d5b05),
	.w5(32'h3b1d4dbe),
	.w6(32'h39d84610),
	.w7(32'h3ba55611),
	.w8(32'hbbaaa394),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cba7e),
	.w1(32'hbc1ffe3e),
	.w2(32'h3a0c8a70),
	.w3(32'h3be4ed84),
	.w4(32'h3b12ff38),
	.w5(32'h3b52ae31),
	.w6(32'hbb8efc70),
	.w7(32'hbc01c19a),
	.w8(32'h3b17525b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4f48e),
	.w1(32'h3b740a0f),
	.w2(32'h3bfbfd0b),
	.w3(32'h3acda235),
	.w4(32'h3b690f66),
	.w5(32'hbab25787),
	.w6(32'hb8ba2e59),
	.w7(32'h3b1645af),
	.w8(32'h3b6b5c92),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30418b),
	.w1(32'h3b58cab5),
	.w2(32'h3baa1ee3),
	.w3(32'hbaf6f586),
	.w4(32'hbac5fbc2),
	.w5(32'hbb190490),
	.w6(32'h3c1f6ce3),
	.w7(32'h3bdb979b),
	.w8(32'hbabe49cb),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34e272),
	.w1(32'h3aaff5d8),
	.w2(32'h3b8b8acb),
	.w3(32'hbbc204d3),
	.w4(32'hbb7bcd1e),
	.w5(32'h394647bc),
	.w6(32'h3be92a07),
	.w7(32'h3be45510),
	.w8(32'h399219a0),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf985d),
	.w1(32'h3c0f7267),
	.w2(32'hbb7d2597),
	.w3(32'h3bf34808),
	.w4(32'h3b800e18),
	.w5(32'hbafba6db),
	.w6(32'h3b405ea3),
	.w7(32'h3c036e90),
	.w8(32'h3a50d9f5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f861c),
	.w1(32'h3b598e43),
	.w2(32'hbb3fc48a),
	.w3(32'hbbcc2b05),
	.w4(32'hba2894db),
	.w5(32'h3b567cc4),
	.w6(32'h3bcb7256),
	.w7(32'h3b325f6c),
	.w8(32'hbb5b9e6e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f9f94),
	.w1(32'hb91c7ffb),
	.w2(32'h39c5b792),
	.w3(32'h3abf8427),
	.w4(32'hba81c3d4),
	.w5(32'hbb8a855b),
	.w6(32'hba518424),
	.w7(32'hbb83c145),
	.w8(32'h3b58e684),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1503bc),
	.w1(32'hba676f64),
	.w2(32'h3ad2545e),
	.w3(32'hbba13a28),
	.w4(32'hba524c1f),
	.w5(32'h39e237b3),
	.w6(32'h3b9cfcc9),
	.w7(32'hbad2174e),
	.w8(32'hbb5d058d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b5d88),
	.w1(32'hbbc0da33),
	.w2(32'hbbde25fa),
	.w3(32'h3a9bb883),
	.w4(32'hbbbf4012),
	.w5(32'h3af1bbec),
	.w6(32'h39f69a3c),
	.w7(32'hbb0b57c9),
	.w8(32'hb9936183),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba298fea),
	.w1(32'h3ac71b2c),
	.w2(32'h3a762ad5),
	.w3(32'hbaede5bb),
	.w4(32'h3ba9e806),
	.w5(32'hb973c5fe),
	.w6(32'h3b09e1f2),
	.w7(32'hbb70070f),
	.w8(32'hbb83b32f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a3e2b),
	.w1(32'hb98221c1),
	.w2(32'hba434baf),
	.w3(32'hb92ce65f),
	.w4(32'hba366ef2),
	.w5(32'h3a4b9f26),
	.w6(32'hb8ca01ca),
	.w7(32'hb90a0564),
	.w8(32'hbbc52738),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb830daf),
	.w1(32'hba91638a),
	.w2(32'hba901988),
	.w3(32'h3bb94ee9),
	.w4(32'h3b16cb02),
	.w5(32'h3b089cd9),
	.w6(32'hbb809ca3),
	.w7(32'hbc0c94a1),
	.w8(32'h3a4168e0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba728c9d),
	.w1(32'hba75861f),
	.w2(32'h3b00cf86),
	.w3(32'h3b193df4),
	.w4(32'h3b1bda7e),
	.w5(32'h3b22a303),
	.w6(32'hbb0181b6),
	.w7(32'h37b4a263),
	.w8(32'h3b372a99),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a4397),
	.w1(32'hbc27d7b8),
	.w2(32'hbbff5728),
	.w3(32'hbb4c05ce),
	.w4(32'hbbf17311),
	.w5(32'h3baaf534),
	.w6(32'hbaa945d1),
	.w7(32'hba8e087a),
	.w8(32'h3a0f8c8b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393030b1),
	.w1(32'h3ae1ec12),
	.w2(32'h3ba2acce),
	.w3(32'h3b9f52e9),
	.w4(32'h3bc1c738),
	.w5(32'h3c0e5531),
	.w6(32'hbb1c2712),
	.w7(32'hbb2f7513),
	.w8(32'h3a9324db),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86d466),
	.w1(32'h3b92e731),
	.w2(32'h3b192dd4),
	.w3(32'hba5739e5),
	.w4(32'h3b0d94d7),
	.w5(32'h3a7c39d8),
	.w6(32'hbb15c7e8),
	.w7(32'h3b276ffa),
	.w8(32'hbc0d2a45),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8aa5e),
	.w1(32'hbb412e35),
	.w2(32'hbb983848),
	.w3(32'hbba888f1),
	.w4(32'hbc0901da),
	.w5(32'h3965a487),
	.w6(32'hbbcabac1),
	.w7(32'h3b82608b),
	.w8(32'hbb7a1308),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b595729),
	.w1(32'hbbc8ba1a),
	.w2(32'hbb8bdf1d),
	.w3(32'h3b3bd4a6),
	.w4(32'hbba4b437),
	.w5(32'h3ad00afd),
	.w6(32'h3c2ca06e),
	.w7(32'hbb23d676),
	.w8(32'h3b465fe4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b37094),
	.w1(32'hbb003d6d),
	.w2(32'h3b342337),
	.w3(32'h3c12190c),
	.w4(32'h3bb1abcf),
	.w5(32'h3b8c7607),
	.w6(32'hbc0ddb34),
	.w7(32'hbb5a79e3),
	.w8(32'hbaf2eddb),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9554ee),
	.w1(32'hbb083d07),
	.w2(32'h3966db8f),
	.w3(32'h3b837834),
	.w4(32'hbb0ea3ed),
	.w5(32'hb967d662),
	.w6(32'hbc1525d5),
	.w7(32'hbbc1e0e2),
	.w8(32'h3ba3c4ee),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06cdab),
	.w1(32'h3b1d3f20),
	.w2(32'hba303ad7),
	.w3(32'h3b8e4527),
	.w4(32'h3ad01487),
	.w5(32'h3b581dd1),
	.w6(32'h3c1a2455),
	.w7(32'h3b85b73f),
	.w8(32'hbb6a42fa),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee6ed1),
	.w1(32'hbaf19cbf),
	.w2(32'h3a6defc4),
	.w3(32'h3b994b73),
	.w4(32'hbb567ef6),
	.w5(32'h3abadb6a),
	.w6(32'hbafb8190),
	.w7(32'hbb0a36b2),
	.w8(32'hbb41438a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcccbbc),
	.w1(32'hbb886f20),
	.w2(32'hbc11c352),
	.w3(32'hbbf70595),
	.w4(32'hbb5aad41),
	.w5(32'hbb219305),
	.w6(32'hbc2547df),
	.w7(32'hbbb00719),
	.w8(32'h3ad42a74),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56533e),
	.w1(32'hbb53de76),
	.w2(32'hbb7d71cc),
	.w3(32'h3b94e398),
	.w4(32'h3b35c628),
	.w5(32'hbc1de26a),
	.w6(32'hbb3ee79b),
	.w7(32'hbbd04d68),
	.w8(32'h3b3cafbc),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9caa46),
	.w1(32'h3ad4bc07),
	.w2(32'h3a247355),
	.w3(32'hb917b922),
	.w4(32'hbc01b639),
	.w5(32'h39fa4d08),
	.w6(32'h3b134ec1),
	.w7(32'hbadb061d),
	.w8(32'h3ba13da8),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a893a3b),
	.w1(32'hbaac97bc),
	.w2(32'h3b8f4291),
	.w3(32'h3c43b1a5),
	.w4(32'h3ba6e7cc),
	.w5(32'h3b5519c0),
	.w6(32'hbbfc1c21),
	.w7(32'hbbb801bf),
	.w8(32'hbb9e774a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ac719),
	.w1(32'hbb01a02a),
	.w2(32'h39fa8390),
	.w3(32'hbb5f5ba9),
	.w4(32'h3b3a0ca9),
	.w5(32'hbad1607c),
	.w6(32'h3b19abbb),
	.w7(32'h3ac069c9),
	.w8(32'hbac5ff48),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f74cf),
	.w1(32'h3aa33dff),
	.w2(32'hba788704),
	.w3(32'h3ba6be2f),
	.w4(32'h3b155c44),
	.w5(32'hbbc40873),
	.w6(32'h3b040772),
	.w7(32'hba88fa75),
	.w8(32'hbbacc3bc),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afee126),
	.w1(32'h3be33e29),
	.w2(32'hba646842),
	.w3(32'hbaf7ebd3),
	.w4(32'hbb261f8f),
	.w5(32'hbb135681),
	.w6(32'hba806f9a),
	.w7(32'h3b0937ab),
	.w8(32'hbc198697),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9b257),
	.w1(32'h3b30e3b3),
	.w2(32'hba7f8285),
	.w3(32'h3bcc3dd7),
	.w4(32'h3b2a4708),
	.w5(32'hba34d1f5),
	.w6(32'hbc0d9750),
	.w7(32'hbbd739bb),
	.w8(32'h3baf1eb0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb1847),
	.w1(32'h3afef729),
	.w2(32'h3bdb5f39),
	.w3(32'hba7bbcc5),
	.w4(32'hbacdb8c8),
	.w5(32'hbbc7d8c0),
	.w6(32'hbb619b42),
	.w7(32'hb949362d),
	.w8(32'h3b221dc7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ec0e9),
	.w1(32'h3b5dd9a3),
	.w2(32'hb9a0357c),
	.w3(32'hbc1fa38a),
	.w4(32'hbad13649),
	.w5(32'h3c81a75c),
	.w6(32'h3ca4e6f1),
	.w7(32'h3c33368a),
	.w8(32'h3a978733),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82c3bf),
	.w1(32'h3ad1b6db),
	.w2(32'h3b5d9533),
	.w3(32'h3c1af9bf),
	.w4(32'h3bb71596),
	.w5(32'hbb17b52d),
	.w6(32'hbbaa40c2),
	.w7(32'h3a39e808),
	.w8(32'hbb86986a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b1e4e),
	.w1(32'h3bf0e939),
	.w2(32'hbb197703),
	.w3(32'h3b44421d),
	.w4(32'h3b01cf65),
	.w5(32'h3babf380),
	.w6(32'h3a9313be),
	.w7(32'hbb91371b),
	.w8(32'h3b5820d0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7ad0b),
	.w1(32'hbb234a72),
	.w2(32'h39b63dbf),
	.w3(32'h3b5c18c5),
	.w4(32'hba84906d),
	.w5(32'hbbbc2375),
	.w6(32'hbbe3bb57),
	.w7(32'hbac8e867),
	.w8(32'h3ab67723),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10d5a8),
	.w1(32'h3ba5bd90),
	.w2(32'h3b57e17f),
	.w3(32'h3b31de5f),
	.w4(32'hbafe1d60),
	.w5(32'hbae50cb4),
	.w6(32'h3b2a3d7f),
	.w7(32'h3b983a6b),
	.w8(32'hbb83443b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b39202),
	.w1(32'h37e8ae57),
	.w2(32'hbb9136af),
	.w3(32'hbb7603af),
	.w4(32'hbb898757),
	.w5(32'hb9b8492d),
	.w6(32'h3afc1de2),
	.w7(32'hbb469d71),
	.w8(32'hbb39c6a0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b727885),
	.w1(32'hba9025da),
	.w2(32'hbb0ecb56),
	.w3(32'h3c2735af),
	.w4(32'hbac5c19a),
	.w5(32'hbae830dc),
	.w6(32'hbbc97f2f),
	.w7(32'hbb9867de),
	.w8(32'h3b97eebe),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51ddc5),
	.w1(32'hbb80eccc),
	.w2(32'hbb448ba5),
	.w3(32'hbac4bb52),
	.w4(32'hbb27b185),
	.w5(32'hbb17552a),
	.w6(32'h3c8bd56c),
	.w7(32'h3b88f971),
	.w8(32'hbb9e9735),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c197a),
	.w1(32'hbb4ca695),
	.w2(32'hbbc5e35b),
	.w3(32'h3b9423d1),
	.w4(32'hbb7ff285),
	.w5(32'h3b86a37d),
	.w6(32'hbb3c5f22),
	.w7(32'hbbe2ad20),
	.w8(32'h3b650f41),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4094e),
	.w1(32'h3c1d474e),
	.w2(32'h3c3f9f5e),
	.w3(32'h39cd3525),
	.w4(32'h3bc31e5a),
	.w5(32'hbb0ddad4),
	.w6(32'h3a722d9d),
	.w7(32'h3b7de733),
	.w8(32'h3b0395da),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ed420),
	.w1(32'hbb2c3265),
	.w2(32'hbb62e15b),
	.w3(32'hbbadfdf2),
	.w4(32'hbb100030),
	.w5(32'h3bd43616),
	.w6(32'h3c3cbb46),
	.w7(32'h3bf1fd43),
	.w8(32'h3a16b73d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989e15c),
	.w1(32'h3bb6445a),
	.w2(32'h3be155ac),
	.w3(32'h3baa35f2),
	.w4(32'h3b76772f),
	.w5(32'h3b4a16da),
	.w6(32'hbbd80d27),
	.w7(32'hbb1c3182),
	.w8(32'h3b226bfd),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96df8f8),
	.w1(32'hbbd14e09),
	.w2(32'hb881694e),
	.w3(32'h3afd29c7),
	.w4(32'h39a7cb92),
	.w5(32'hbae90901),
	.w6(32'hbac12495),
	.w7(32'hba4e4bcc),
	.w8(32'hbb6098af),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fd278),
	.w1(32'hbad0af39),
	.w2(32'hbb3144dd),
	.w3(32'h39921b1e),
	.w4(32'hba15d1dd),
	.w5(32'hbbb51727),
	.w6(32'hbb7c01d0),
	.w7(32'hbb06078c),
	.w8(32'hbb07b8e8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbaab78),
	.w1(32'h3bcbc124),
	.w2(32'h39db22d8),
	.w3(32'hbb1daeac),
	.w4(32'hb9dc8b5f),
	.w5(32'h3b1c0047),
	.w6(32'h3b91bd1e),
	.w7(32'h3b967e75),
	.w8(32'hbb037981),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d28de),
	.w1(32'h3b681ebd),
	.w2(32'hbc11cb9c),
	.w3(32'h3a88d92e),
	.w4(32'hbbcb9338),
	.w5(32'h3b025349),
	.w6(32'hbc0100c4),
	.w7(32'h3a675e67),
	.w8(32'h3b61c764),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18cd3b),
	.w1(32'hbb117d2a),
	.w2(32'hba6b53b8),
	.w3(32'h3b4d1abb),
	.w4(32'h39a5b979),
	.w5(32'hbac9726d),
	.w6(32'h3bb2154a),
	.w7(32'h3acefb92),
	.w8(32'h3a611d1b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae18d39),
	.w1(32'hbb010dfb),
	.w2(32'h39b2615e),
	.w3(32'h3aded40c),
	.w4(32'hbb9dd8d9),
	.w5(32'hbb4e8655),
	.w6(32'h3bb68031),
	.w7(32'h3ac5a857),
	.w8(32'h3b020e92),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2f49b),
	.w1(32'h3b74a83d),
	.w2(32'h3ba2ff74),
	.w3(32'h3b05431f),
	.w4(32'h39c7dd8d),
	.w5(32'h38c0fa41),
	.w6(32'h3a88b78c),
	.w7(32'hbb3c3962),
	.w8(32'hbb8313fa),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc109d95),
	.w1(32'hb8040a1b),
	.w2(32'hbb679871),
	.w3(32'hbb114b04),
	.w4(32'hbbb1eaf6),
	.w5(32'h3be9d100),
	.w6(32'hbb7c0927),
	.w7(32'h3ab18ef8),
	.w8(32'h39954633),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b124bc9),
	.w1(32'h3b891558),
	.w2(32'h3bf6651f),
	.w3(32'h3bd92245),
	.w4(32'h3b43f508),
	.w5(32'hbbcf2bef),
	.w6(32'hbc39829f),
	.w7(32'h37f90479),
	.w8(32'hbc21f796),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a25c7),
	.w1(32'h3c979140),
	.w2(32'h3c640281),
	.w3(32'h3c605743),
	.w4(32'h3c29ad9b),
	.w5(32'h3acc0ef5),
	.w6(32'h3c7e5c83),
	.w7(32'h3bae1db8),
	.w8(32'h3b2837a2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82447a),
	.w1(32'h3978576d),
	.w2(32'h3b7c608f),
	.w3(32'hb99c0c5f),
	.w4(32'hbb180f60),
	.w5(32'hba996a18),
	.w6(32'h3c449658),
	.w7(32'h3aeb0ad2),
	.w8(32'h3b8d3cfe),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00db22),
	.w1(32'hbb846dc4),
	.w2(32'hbb476e0a),
	.w3(32'h3bf56ede),
	.w4(32'h3af01e03),
	.w5(32'hbbd4c00f),
	.w6(32'h3bd3fb3d),
	.w7(32'hba9b49e4),
	.w8(32'hbbc4a008),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f08e4),
	.w1(32'hbbdeaa70),
	.w2(32'hbb9403d6),
	.w3(32'hbbcac659),
	.w4(32'hbbc3c224),
	.w5(32'h39b8a193),
	.w6(32'hbae458d4),
	.w7(32'hbbbbe62c),
	.w8(32'hbac7780f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab88a5f),
	.w1(32'h39ce7d3c),
	.w2(32'h39d6799c),
	.w3(32'h3b62e45a),
	.w4(32'h3a1de8e2),
	.w5(32'hba92426f),
	.w6(32'hbb80181f),
	.w7(32'hbaa80e7c),
	.w8(32'h3b3cb347),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3929a9f0),
	.w1(32'hbb7133a2),
	.w2(32'hbbc44a1f),
	.w3(32'hbac85f7c),
	.w4(32'hbad5f33c),
	.w5(32'hbb4d6af0),
	.w6(32'hbb68e815),
	.w7(32'hbb7e302b),
	.w8(32'hbba58de9),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab61d60),
	.w1(32'h3b004d63),
	.w2(32'h39bfcf4f),
	.w3(32'hbbaf867c),
	.w4(32'hbbdd0283),
	.w5(32'hbbd5914c),
	.w6(32'h3be29a7f),
	.w7(32'h3b0c49be),
	.w8(32'hbbdeb07a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4fcef),
	.w1(32'hbb850367),
	.w2(32'hba8560e1),
	.w3(32'hbbfe41f2),
	.w4(32'h3b121462),
	.w5(32'hbbe1b25e),
	.w6(32'h3c4527b0),
	.w7(32'h39a5176b),
	.w8(32'h3bc3f45f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf487f),
	.w1(32'h3b9f16b6),
	.w2(32'h3b559eb4),
	.w3(32'h3a8cfb15),
	.w4(32'h3a725516),
	.w5(32'hbae54604),
	.w6(32'h3bd252aa),
	.w7(32'hba01de1e),
	.w8(32'h3a52b568),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36bb30),
	.w1(32'hbb6e1f60),
	.w2(32'hbb118d58),
	.w3(32'hbae2891b),
	.w4(32'hbb56864f),
	.w5(32'h3b8f7d68),
	.w6(32'hbbc4ec31),
	.w7(32'hbba44b4e),
	.w8(32'h3b11a6a3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93c6d1),
	.w1(32'h3b9b3e01),
	.w2(32'h3b6d3602),
	.w3(32'hb9c7424b),
	.w4(32'h3b835123),
	.w5(32'h3c061a68),
	.w6(32'h3b898b40),
	.w7(32'h3ae4deab),
	.w8(32'h3b002224),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ed2be),
	.w1(32'h3b764a36),
	.w2(32'h3bb85f80),
	.w3(32'h3c3dc02a),
	.w4(32'h3c13e393),
	.w5(32'h3c472b64),
	.w6(32'hbb90b8a8),
	.w7(32'hbacdadcd),
	.w8(32'h38ce52c1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc156216),
	.w1(32'hbc0b7fd7),
	.w2(32'h3bd47ed2),
	.w3(32'h3bd4f0a2),
	.w4(32'hbb93f00b),
	.w5(32'h3b2fd763),
	.w6(32'hbc46062c),
	.w7(32'h3aded81a),
	.w8(32'hbc51c4aa),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea4ce8),
	.w1(32'h3cd11382),
	.w2(32'h3c3bc07b),
	.w3(32'h3cb920e9),
	.w4(32'h3b2b9ebc),
	.w5(32'hba94c5bb),
	.w6(32'hbcb1e45f),
	.w7(32'hbbc1cc64),
	.w8(32'hbb136aac),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf4643),
	.w1(32'hbb22260c),
	.w2(32'hbba8bfab),
	.w3(32'hbc05769c),
	.w4(32'hba1aee9f),
	.w5(32'hbbcb1f03),
	.w6(32'h3a800a35),
	.w7(32'hbb6f5770),
	.w8(32'hbb2197d9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ffea41),
	.w1(32'h3b5a6c40),
	.w2(32'h3a0e4304),
	.w3(32'hbc1cb278),
	.w4(32'hbb88f209),
	.w5(32'hbb55001a),
	.w6(32'h3c34327f),
	.w7(32'hb9b9019a),
	.w8(32'h3a65321d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34943),
	.w1(32'h3b28ef20),
	.w2(32'h3a94bb1f),
	.w3(32'hbc3c9bd4),
	.w4(32'hbc1d51c3),
	.w5(32'h3b259c1a),
	.w6(32'h3bd59706),
	.w7(32'h3b98789a),
	.w8(32'hbbe91219),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a645f),
	.w1(32'h3b80165b),
	.w2(32'h3adc1c9d),
	.w3(32'hbb23bcc8),
	.w4(32'hba31eab1),
	.w5(32'hbb029031),
	.w6(32'hbb1b2a3b),
	.w7(32'hbb077d6b),
	.w8(32'hbb9a6ddf),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb800eac),
	.w1(32'hbabc33ae),
	.w2(32'hbb4050a4),
	.w3(32'h3ace0a09),
	.w4(32'h3ab708ce),
	.w5(32'h3ad15a65),
	.w6(32'hbb685a54),
	.w7(32'hbb27113b),
	.w8(32'hba349b9e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7a893),
	.w1(32'h3a39253d),
	.w2(32'h3b21290b),
	.w3(32'h3be3cd2c),
	.w4(32'h3b883870),
	.w5(32'h3b3b6f5b),
	.w6(32'h3c24f01f),
	.w7(32'h3a8cc141),
	.w8(32'hba0d81c4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d09cd),
	.w1(32'h3b749627),
	.w2(32'h3b9c6bb5),
	.w3(32'h3aa77bcd),
	.w4(32'h3be95276),
	.w5(32'h3be682a6),
	.w6(32'h3c897e4c),
	.w7(32'h3a8e6c36),
	.w8(32'h3bea59e1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c206e2a),
	.w1(32'h3a2c8667),
	.w2(32'h3c08549f),
	.w3(32'h3a0a798c),
	.w4(32'h3a27e9e5),
	.w5(32'h3aa3bb50),
	.w6(32'hbb92cf7e),
	.w7(32'hbb438f3a),
	.w8(32'hbb031013),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83ec78),
	.w1(32'h398077b7),
	.w2(32'hba9d0050),
	.w3(32'hbb47b005),
	.w4(32'hbaba18a3),
	.w5(32'h38940f02),
	.w6(32'h3b9c4c38),
	.w7(32'h3a4ed5e7),
	.w8(32'hb9e71fed),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4d0f3),
	.w1(32'hb9997537),
	.w2(32'hbb6f688f),
	.w3(32'hbbd52506),
	.w4(32'hbb7ab380),
	.w5(32'h3a8b3bde),
	.w6(32'hba8822c1),
	.w7(32'hb987343b),
	.w8(32'h3c009797),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0abe74),
	.w1(32'h3b302ca5),
	.w2(32'h3b470656),
	.w3(32'hbbf4d320),
	.w4(32'h38b55f4d),
	.w5(32'h3adfe936),
	.w6(32'h3c190469),
	.w7(32'h3c472127),
	.w8(32'h395bdfbe),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d853d),
	.w1(32'h3b697499),
	.w2(32'h3a1c5961),
	.w3(32'hbaa52f3d),
	.w4(32'hb95c1c60),
	.w5(32'hbc298a8b),
	.w6(32'hbad58396),
	.w7(32'hba8ff7e5),
	.w8(32'h3c00c56d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf63b3c),
	.w1(32'hbaee3e04),
	.w2(32'h3b1dd459),
	.w3(32'hbc22bb46),
	.w4(32'hbc3797f6),
	.w5(32'h3c4f3797),
	.w6(32'h3cc7b6ea),
	.w7(32'h3c51c538),
	.w8(32'h3aadd72f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae22263),
	.w1(32'h3b7f1621),
	.w2(32'hbba405b0),
	.w3(32'h3bde2acc),
	.w4(32'hba990cec),
	.w5(32'h3b2de289),
	.w6(32'hbadac6a7),
	.w7(32'h3b0fbc06),
	.w8(32'hbbf80a83),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73bbf7),
	.w1(32'hbb9add6d),
	.w2(32'hbb85b4a8),
	.w3(32'h3a7170f3),
	.w4(32'h391d4f54),
	.w5(32'hbad8dd4f),
	.w6(32'h37356ea5),
	.w7(32'hbb984241),
	.w8(32'hbb2aef9d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cb42f),
	.w1(32'h3a977774),
	.w2(32'h3b2e2934),
	.w3(32'hbb5f537b),
	.w4(32'hba0d19fc),
	.w5(32'h3af87519),
	.w6(32'hbaa0e92c),
	.w7(32'hbb633593),
	.w8(32'h3bdba7c9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1807a7),
	.w1(32'hbad4b692),
	.w2(32'h3a80e0e6),
	.w3(32'hbc179c1a),
	.w4(32'h3b926301),
	.w5(32'h3c5bfe45),
	.w6(32'hbbf02716),
	.w7(32'hba192b18),
	.w8(32'h3b2a0230),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c043e51),
	.w1(32'hbb0c068c),
	.w2(32'h3b31fa39),
	.w3(32'h3a6b2089),
	.w4(32'h3b86e981),
	.w5(32'h3ba987b2),
	.w6(32'h3b699d1c),
	.w7(32'h372950d8),
	.w8(32'h3bc86841),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d1c56),
	.w1(32'hbb96c5d9),
	.w2(32'hbbbf7921),
	.w3(32'h39a84a3c),
	.w4(32'hbba145de),
	.w5(32'hbbbd95e6),
	.w6(32'hbc52eaa1),
	.w7(32'hbb761375),
	.w8(32'hbbdc511e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9863ce),
	.w1(32'hb98f7a14),
	.w2(32'hbaa12622),
	.w3(32'h3bafaefe),
	.w4(32'h39e35573),
	.w5(32'h3a59549f),
	.w6(32'hbb69f143),
	.w7(32'hbb8ddf98),
	.w8(32'h3ad39ebc),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b881058),
	.w1(32'h3a7809f5),
	.w2(32'hbb43b61f),
	.w3(32'h3be5eab6),
	.w4(32'hbbbb1fdb),
	.w5(32'h3b0837b8),
	.w6(32'h3b7468d2),
	.w7(32'hba8b9a26),
	.w8(32'h3c19d2ee),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09b6a9),
	.w1(32'hba8ea3bd),
	.w2(32'h3b99a0a5),
	.w3(32'h3be491eb),
	.w4(32'h3a9d8bec),
	.w5(32'hbc1b2352),
	.w6(32'hbbf59de3),
	.w7(32'hbb58c073),
	.w8(32'hbafdfa0d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aceb960),
	.w1(32'h3c0c7d7c),
	.w2(32'h3c16dfaa),
	.w3(32'hbad42c9d),
	.w4(32'hbb1e618c),
	.w5(32'hbb4b82bb),
	.w6(32'h3a9bc344),
	.w7(32'h3beca4db),
	.w8(32'h397269b0),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1074ff),
	.w1(32'hba41fe1d),
	.w2(32'hbba5c38c),
	.w3(32'hba6db56c),
	.w4(32'hb92d364a),
	.w5(32'h3a6a08e6),
	.w6(32'h3c2d9c14),
	.w7(32'h3bd51716),
	.w8(32'h3ba767b5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fc401),
	.w1(32'hbbdce335),
	.w2(32'hba8f73bf),
	.w3(32'h3b91aa88),
	.w4(32'h3c0650b1),
	.w5(32'hb9ef4f96),
	.w6(32'hbc218557),
	.w7(32'hbc03efe9),
	.w8(32'hb97ab2bc),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaccb6),
	.w1(32'hbac3ca3f),
	.w2(32'hba9037c6),
	.w3(32'hbb4aae52),
	.w4(32'hbadc0405),
	.w5(32'hbb14843c),
	.w6(32'hbb312ed7),
	.w7(32'hbaa0cfd2),
	.w8(32'hb9cc2b88),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b030d),
	.w1(32'h3b6e146b),
	.w2(32'h390025f3),
	.w3(32'h3b00b54f),
	.w4(32'hb95fecea),
	.w5(32'h399ba7aa),
	.w6(32'h3b9b3d11),
	.w7(32'hb9d6e876),
	.w8(32'hba6a9bc4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95149f),
	.w1(32'h3a556ea7),
	.w2(32'h3b325f83),
	.w3(32'h39f5b30e),
	.w4(32'h399ef342),
	.w5(32'hba895ad4),
	.w6(32'hbac088c4),
	.w7(32'hba9a1085),
	.w8(32'h3b3e88bb),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c37f3),
	.w1(32'h3b7142e7),
	.w2(32'h3b871880),
	.w3(32'hbb096d12),
	.w4(32'hba750a51),
	.w5(32'hb9bc75d9),
	.w6(32'h3b2f5bd9),
	.w7(32'h3b4bf784),
	.w8(32'hb9b428cc),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9da195),
	.w1(32'h3a5ed4de),
	.w2(32'hbb17ecd0),
	.w3(32'hbb423af2),
	.w4(32'h3a5dcdd2),
	.w5(32'h3a1d138a),
	.w6(32'h3920f2dd),
	.w7(32'h39714b67),
	.w8(32'h3b1668e1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ddd7e),
	.w1(32'h3b1f5f31),
	.w2(32'hb80e142e),
	.w3(32'h3ac3c947),
	.w4(32'hba9382f5),
	.w5(32'hba9b1fe1),
	.w6(32'h3a44d6cc),
	.w7(32'h3b00e37b),
	.w8(32'hbb133817),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b46f44),
	.w1(32'hba95d043),
	.w2(32'h3981925b),
	.w3(32'hbaaf2f5e),
	.w4(32'h390ea1f6),
	.w5(32'h38f9ab7c),
	.w6(32'hba54d1a4),
	.w7(32'hba55f94b),
	.w8(32'h3a33aee2),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f52775),
	.w1(32'h3ade0b72),
	.w2(32'h3a195d58),
	.w3(32'h393660ee),
	.w4(32'h3a692edd),
	.w5(32'hbab55844),
	.w6(32'h3a097ab7),
	.w7(32'h3a75ebb4),
	.w8(32'hba867d68),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084385),
	.w1(32'hbb0d15e3),
	.w2(32'hbaa6eac0),
	.w3(32'hbb07df9e),
	.w4(32'hbb15bba6),
	.w5(32'hba621e95),
	.w6(32'hb9a7d7a4),
	.w7(32'hba9bab20),
	.w8(32'hbabe8443),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdd770),
	.w1(32'hba199206),
	.w2(32'hbae05bb1),
	.w3(32'h38891b9b),
	.w4(32'hba1869db),
	.w5(32'h396bc250),
	.w6(32'h3a6e1767),
	.w7(32'hba64cc62),
	.w8(32'h3a079e59),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b4bda),
	.w1(32'h39271972),
	.w2(32'h3927478e),
	.w3(32'hba18b521),
	.w4(32'hba1af253),
	.w5(32'hbad4b114),
	.w6(32'hba37c82c),
	.w7(32'h39182de9),
	.w8(32'hba904878),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b934c),
	.w1(32'hba9d1fee),
	.w2(32'hbabbb344),
	.w3(32'hbac32098),
	.w4(32'hba33dc90),
	.w5(32'hba5797de),
	.w6(32'hba874572),
	.w7(32'hba987372),
	.w8(32'hb7ff13e0),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ad44d),
	.w1(32'h3a0886c8),
	.w2(32'h39202ff6),
	.w3(32'h3a9a358e),
	.w4(32'h39a83852),
	.w5(32'hba9b2335),
	.w6(32'h3b1bfa11),
	.w7(32'h39d9aaa3),
	.w8(32'hb9328ed9),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69a276),
	.w1(32'h3ab2dc52),
	.w2(32'h3acdea1a),
	.w3(32'h3b949bcf),
	.w4(32'h3a2d0b56),
	.w5(32'h3b0ae312),
	.w6(32'h3b4de661),
	.w7(32'hb88c0d2e),
	.w8(32'h3a3cda15),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75e3fe),
	.w1(32'h3a87a894),
	.w2(32'h3a0352cb),
	.w3(32'h3b1b8f75),
	.w4(32'h3a853607),
	.w5(32'h3a31d456),
	.w6(32'hbaa50309),
	.w7(32'hbaeee0cf),
	.w8(32'h39b4ce7d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb35153),
	.w1(32'h3b6b7a7e),
	.w2(32'h3b48bbb6),
	.w3(32'h3b725654),
	.w4(32'h3ad14bd1),
	.w5(32'h3ab5d25c),
	.w6(32'h3ae3319c),
	.w7(32'h38b098dc),
	.w8(32'hba149d44),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cee7f),
	.w1(32'h3aee024d),
	.w2(32'h3ae8c426),
	.w3(32'h3a5b0963),
	.w4(32'h3a54ba84),
	.w5(32'hba7d72c4),
	.w6(32'h3ab84e6d),
	.w7(32'h3abb20a1),
	.w8(32'h3a49a888),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06293c),
	.w1(32'h3acb317c),
	.w2(32'h3aae389a),
	.w3(32'hb7948cee),
	.w4(32'h3a4505a1),
	.w5(32'h3a3fcd2c),
	.w6(32'h3ae0679a),
	.w7(32'h3acdd980),
	.w8(32'h3a0ff66f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b1a88),
	.w1(32'h3a398be0),
	.w2(32'h39f15024),
	.w3(32'h39ad95c5),
	.w4(32'h3a1c7426),
	.w5(32'hba87b8a9),
	.w6(32'h39c4428e),
	.w7(32'h39b4db7a),
	.w8(32'hba427727),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab69b1a),
	.w1(32'hb8092dc3),
	.w2(32'hb98a0c11),
	.w3(32'hba17f289),
	.w4(32'hbb028d54),
	.w5(32'hbae6e961),
	.w6(32'h3a7ca0a9),
	.w7(32'h3a82563d),
	.w8(32'hbb01abad),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb654d),
	.w1(32'hbad037dc),
	.w2(32'hbacc9bed),
	.w3(32'h3a691944),
	.w4(32'hba60eda4),
	.w5(32'hbabcab66),
	.w6(32'hba85c4ac),
	.w7(32'hbab7d675),
	.w8(32'hba179ce3),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba103baf),
	.w1(32'hbae7823b),
	.w2(32'hbad6e044),
	.w3(32'hbb3858f2),
	.w4(32'hbad10370),
	.w5(32'h3a975788),
	.w6(32'hbb98b40f),
	.w7(32'hbaf3f092),
	.w8(32'h3a292f8a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9347bde),
	.w1(32'h3b3117ef),
	.w2(32'h3aa5dc9c),
	.w3(32'hb9415639),
	.w4(32'h3aa3587b),
	.w5(32'hbab06a2a),
	.w6(32'hb9521afe),
	.w7(32'h3a272c14),
	.w8(32'h39d3fb91),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa40610),
	.w1(32'hb9237f35),
	.w2(32'h395c8138),
	.w3(32'hb9faeeb2),
	.w4(32'hba8fdb7f),
	.w5(32'h3a96c023),
	.w6(32'hb9ba9ecb),
	.w7(32'hb989c746),
	.w8(32'h3b23e23e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb841aa4d),
	.w1(32'hb83daabf),
	.w2(32'h3a3f2b55),
	.w3(32'h39e0c1bc),
	.w4(32'h3a69de57),
	.w5(32'hba2801a5),
	.w6(32'h3adafef7),
	.w7(32'h3a7583f3),
	.w8(32'hbaee4878),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba875d98),
	.w1(32'hba070d8d),
	.w2(32'hbaa30a46),
	.w3(32'hba8c625a),
	.w4(32'h3924f013),
	.w5(32'h3b2cef9e),
	.w6(32'hbb01d79a),
	.w7(32'hba7275a9),
	.w8(32'h3b586411),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4222f9),
	.w1(32'h3b00dbae),
	.w2(32'h3a34b730),
	.w3(32'h3a115cf7),
	.w4(32'h3ab0d326),
	.w5(32'hba4977c5),
	.w6(32'h3a809a99),
	.w7(32'hb868e278),
	.w8(32'h3ad93d2a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf71f52),
	.w1(32'h3b6d2717),
	.w2(32'h3b1e88ee),
	.w3(32'h3ba44f2f),
	.w4(32'hb98e8f8f),
	.w5(32'h39f65272),
	.w6(32'h3bd43859),
	.w7(32'h3b087b04),
	.w8(32'hba48fc9c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade7c62),
	.w1(32'hb8cfabf5),
	.w2(32'hba3737e3),
	.w3(32'h3a755d02),
	.w4(32'hba063e5a),
	.w5(32'hb8cfedfe),
	.w6(32'h3b0718e7),
	.w7(32'hb8b6589f),
	.w8(32'h378f0d28),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27c140),
	.w1(32'h3b186d29),
	.w2(32'h37ecb8a6),
	.w3(32'hb99825ec),
	.w4(32'hba97ff87),
	.w5(32'hb9bc3169),
	.w6(32'hbb349f61),
	.w7(32'hba613e48),
	.w8(32'h38b12e6d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule