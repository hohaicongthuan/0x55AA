module layer_10_featuremap_397(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93c797),
	.w1(32'hbbd54028),
	.w2(32'hbba40122),
	.w3(32'h3a194314),
	.w4(32'hbbe7d09c),
	.w5(32'hbbce6a76),
	.w6(32'hbbeddb56),
	.w7(32'h3bc36d74),
	.w8(32'hbbd7ea2f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e2150),
	.w1(32'hb92fd78e),
	.w2(32'h3c225cac),
	.w3(32'hbb2608fe),
	.w4(32'h3b9a303e),
	.w5(32'h3c5a52d7),
	.w6(32'h3a894e05),
	.w7(32'h3b8c4cf5),
	.w8(32'h3c36fcb8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b94ef),
	.w1(32'hbb197dc4),
	.w2(32'hbc11d19a),
	.w3(32'hbbfd1ec8),
	.w4(32'hbc161263),
	.w5(32'hbaa3cd8d),
	.w6(32'h3c201faa),
	.w7(32'hbb0ca74f),
	.w8(32'hbc063739),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9971cb),
	.w1(32'hbc016b44),
	.w2(32'hbc259219),
	.w3(32'h3862150a),
	.w4(32'hbbbdfe8e),
	.w5(32'hba055e30),
	.w6(32'h3a493caa),
	.w7(32'hbc4e0c33),
	.w8(32'hbcaef7ee),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddf854),
	.w1(32'h3be42828),
	.w2(32'h3b9158ba),
	.w3(32'hbc2bf5d0),
	.w4(32'hbb232cf1),
	.w5(32'hbbaf1ccb),
	.w6(32'hbc91954a),
	.w7(32'hb9050265),
	.w8(32'hbbed16be),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae51ee3),
	.w1(32'h3a94f7ef),
	.w2(32'hbad4b907),
	.w3(32'hbba2d35e),
	.w4(32'h3bae3c40),
	.w5(32'h3b9b05aa),
	.w6(32'hbb07bde5),
	.w7(32'h3b136a98),
	.w8(32'hbb3908f9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af52a32),
	.w1(32'h3cb51b08),
	.w2(32'h3bd29262),
	.w3(32'h3a36f3b1),
	.w4(32'h3cc66655),
	.w5(32'h3c62cb19),
	.w6(32'h3bddf0db),
	.w7(32'h3c6204b7),
	.w8(32'h3bdaf84c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd1ff7),
	.w1(32'hbabe1549),
	.w2(32'hbc475b2b),
	.w3(32'h3c4b2e1b),
	.w4(32'h3c14e9eb),
	.w5(32'hbb522241),
	.w6(32'h3c938cdd),
	.w7(32'h3badc8ab),
	.w8(32'h3a3347e8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b707024),
	.w1(32'h3982dbc2),
	.w2(32'h3ad445ba),
	.w3(32'h3aa31d53),
	.w4(32'hbbe03fc8),
	.w5(32'hbbf7eef0),
	.w6(32'h3b0c6c31),
	.w7(32'hbc15d9c1),
	.w8(32'hbbc7cbc9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb6040),
	.w1(32'hbb85348e),
	.w2(32'hbb83ece7),
	.w3(32'hbc652bc2),
	.w4(32'hbb97670f),
	.w5(32'hbb90c20f),
	.w6(32'hbc575937),
	.w7(32'hbbb44686),
	.w8(32'hbc5e16d6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac5b93),
	.w1(32'hbc02c708),
	.w2(32'hbbcf645f),
	.w3(32'h39e8371a),
	.w4(32'hbb9bd207),
	.w5(32'hba2ca458),
	.w6(32'h3b8d69b1),
	.w7(32'hbb4d772b),
	.w8(32'hbb7560ff),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef3bdb),
	.w1(32'hbb186c8c),
	.w2(32'hbc31ca2b),
	.w3(32'h3b766482),
	.w4(32'h3b071251),
	.w5(32'hbb1fb350),
	.w6(32'hba89fa64),
	.w7(32'h3b4052fa),
	.w8(32'h3c0394c2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5e93d),
	.w1(32'h3c45c3ca),
	.w2(32'h3c8097ba),
	.w3(32'h3b613f03),
	.w4(32'h3acc530c),
	.w5(32'hbc1a0195),
	.w6(32'h3bc8d2a8),
	.w7(32'hbb958dc5),
	.w8(32'h3c779634),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969ffb9),
	.w1(32'h3b1e1ee8),
	.w2(32'h3b8a269f),
	.w3(32'h389eaf22),
	.w4(32'hbbb1c999),
	.w5(32'hbb00b093),
	.w6(32'h3c9d0ef2),
	.w7(32'hbb5c5e87),
	.w8(32'hb9cb06e3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79c7b5),
	.w1(32'hbc050bac),
	.w2(32'hbbf1f5dc),
	.w3(32'hbad1ad4f),
	.w4(32'hbbebcd43),
	.w5(32'hba8519a1),
	.w6(32'hbb6a4ce7),
	.w7(32'hbc101e8c),
	.w8(32'hbc68756d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0615e1),
	.w1(32'hb994f7f6),
	.w2(32'hbb66556d),
	.w3(32'h3985f37f),
	.w4(32'hbb2b3a6e),
	.w5(32'hbc09df53),
	.w6(32'h38b42e99),
	.w7(32'hbc4f45f1),
	.w8(32'hbc3a4afa),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb694ed0),
	.w1(32'h3bcff7b8),
	.w2(32'h3be24002),
	.w3(32'h3b873a8b),
	.w4(32'h3aeb96c0),
	.w5(32'h3b597c58),
	.w6(32'h3b11e9ba),
	.w7(32'hba8d0f24),
	.w8(32'h3aeaf10e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf18463),
	.w1(32'hbbe87892),
	.w2(32'hbc529bdc),
	.w3(32'hbb2aeeb6),
	.w4(32'hbbfdd54a),
	.w5(32'hbc56079f),
	.w6(32'hba94fbf4),
	.w7(32'hbb293c92),
	.w8(32'hbc15347a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0fa0a),
	.w1(32'hbbd5b42a),
	.w2(32'hbc56e318),
	.w3(32'hbb2ab8cc),
	.w4(32'hbb6712d0),
	.w5(32'hbc0728d1),
	.w6(32'hba734089),
	.w7(32'hbc0f99de),
	.w8(32'hbbf3a93c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4d106),
	.w1(32'hbb1d2bbf),
	.w2(32'h3b0695bc),
	.w3(32'hbb4d1dd0),
	.w4(32'h3ac3c0e8),
	.w5(32'h3b9d49c4),
	.w6(32'hbb99168d),
	.w7(32'hba9a4243),
	.w8(32'hbc4afaae),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba18339),
	.w1(32'hbbcbea4f),
	.w2(32'hbbb6a18e),
	.w3(32'h3b832c50),
	.w4(32'hbb599cd0),
	.w5(32'hbbca0967),
	.w6(32'h39a90c9b),
	.w7(32'hbbc65374),
	.w8(32'hbb75f181),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb1521),
	.w1(32'hbb5cce7f),
	.w2(32'hb9ae758e),
	.w3(32'hba323f63),
	.w4(32'h3ba4a513),
	.w5(32'hbc22aa16),
	.w6(32'hbaf60faa),
	.w7(32'h3b65abb8),
	.w8(32'hbc09fc6b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ef297),
	.w1(32'hbb839c38),
	.w2(32'hbc19b46f),
	.w3(32'h3b97743c),
	.w4(32'h3aa9bf8b),
	.w5(32'h3b50472b),
	.w6(32'hbb52e6a7),
	.w7(32'h39f8287b),
	.w8(32'hbc1a88f1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25ed5a),
	.w1(32'h3b197d8e),
	.w2(32'hbbb6b8fd),
	.w3(32'hbc2c0bc0),
	.w4(32'h39cd9c89),
	.w5(32'hbb54ab28),
	.w6(32'hbb4e9d61),
	.w7(32'hbbb456bf),
	.w8(32'hbc009749),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94ea34),
	.w1(32'hbb8f4156),
	.w2(32'h3bae877e),
	.w3(32'h38eab279),
	.w4(32'h3ab69bbc),
	.w5(32'hbb9eebcc),
	.w6(32'hbc2037cd),
	.w7(32'hbb7636bd),
	.w8(32'hb8dbc83a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02333c),
	.w1(32'h3bf79257),
	.w2(32'hbad46282),
	.w3(32'hbb9431aa),
	.w4(32'h3bb124de),
	.w5(32'hb938c4c5),
	.w6(32'hbc194a68),
	.w7(32'h3a1e60e6),
	.w8(32'hbb62e590),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf54fa5),
	.w1(32'hbb847856),
	.w2(32'h3bb0d9ef),
	.w3(32'hbabe4082),
	.w4(32'h3bbd1130),
	.w5(32'h3c9abea5),
	.w6(32'hbb0cddee),
	.w7(32'h3b1d8e2c),
	.w8(32'hb98de9c1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb94d6),
	.w1(32'hbacf1207),
	.w2(32'hba9f816f),
	.w3(32'h3bb2ff93),
	.w4(32'hbaaefd24),
	.w5(32'h3bfed1cd),
	.w6(32'hbc200cc4),
	.w7(32'h397fb4e8),
	.w8(32'h3b99fdeb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c059362),
	.w1(32'h3bd9b0c9),
	.w2(32'h3b9d3f13),
	.w3(32'h3c558425),
	.w4(32'h3b23b796),
	.w5(32'h3acd2358),
	.w6(32'h3c2f2f07),
	.w7(32'h3b8783c8),
	.w8(32'hba85d2ec),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb525c92),
	.w1(32'hbb22d69e),
	.w2(32'hbb00eec5),
	.w3(32'hbc214118),
	.w4(32'h3a56db9b),
	.w5(32'h3a0baffc),
	.w6(32'hbb4baf43),
	.w7(32'h3b56952b),
	.w8(32'h3bba2023),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadeab7),
	.w1(32'h3b3e1f72),
	.w2(32'h3a74a6c9),
	.w3(32'h3b13ef0d),
	.w4(32'h3b8e9b06),
	.w5(32'h3c08e3b0),
	.w6(32'h3c0f304b),
	.w7(32'hbad809ba),
	.w8(32'hbba6d950),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac09619),
	.w1(32'h3c1d00aa),
	.w2(32'h3bde03ab),
	.w3(32'h3ae3d7fd),
	.w4(32'hb9616150),
	.w5(32'h3a0a331b),
	.w6(32'hbb96bd45),
	.w7(32'hbb070bd8),
	.w8(32'hbb52cccc),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2e9dd),
	.w1(32'h3b4f0fb1),
	.w2(32'h3b6249eb),
	.w3(32'h3be8e81a),
	.w4(32'h3b49e81b),
	.w5(32'hbc2207f5),
	.w6(32'h399bdda7),
	.w7(32'h3c9c478c),
	.w8(32'h3cf8dbad),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e686f3),
	.w1(32'h3c75f508),
	.w2(32'h3b93c527),
	.w3(32'h3b8bf759),
	.w4(32'h3c850edb),
	.w5(32'h3cd22f79),
	.w6(32'h3c591866),
	.w7(32'h3c5b9f79),
	.w8(32'h3c39d6d3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e4a7b),
	.w1(32'hbb73e13d),
	.w2(32'hbc0c8356),
	.w3(32'h3c7d4712),
	.w4(32'h3bcec038),
	.w5(32'h3c260e77),
	.w6(32'h3b84df35),
	.w7(32'h39a2ee3e),
	.w8(32'h3a5034c9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e5ad1),
	.w1(32'h3b13decf),
	.w2(32'h398b3526),
	.w3(32'h3ba8f365),
	.w4(32'h3a4797df),
	.w5(32'hbaa57a32),
	.w6(32'h3ba39ec2),
	.w7(32'h3bd78699),
	.w8(32'h3b2311cf),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb440e7e),
	.w1(32'hbc18c4de),
	.w2(32'hbc4fe9f1),
	.w3(32'h3b4f686c),
	.w4(32'hbaef4baf),
	.w5(32'h3cb90ac6),
	.w6(32'hba3910fe),
	.w7(32'h3b690c7e),
	.w8(32'h3ae53210),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0589e),
	.w1(32'h3c481ec2),
	.w2(32'h3cb65c4b),
	.w3(32'hbb801adb),
	.w4(32'h3c5c2430),
	.w5(32'h3c8ac2fa),
	.w6(32'hbb595567),
	.w7(32'hbb0a8de4),
	.w8(32'h3bd1164d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2ed63),
	.w1(32'h3b92aebb),
	.w2(32'h3c8bc238),
	.w3(32'h3b9d714d),
	.w4(32'h3c22dd4d),
	.w5(32'h3bbf2690),
	.w6(32'h3c866832),
	.w7(32'h3bcec46d),
	.w8(32'h3c2528cf),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c349df5),
	.w1(32'h3be24a40),
	.w2(32'h3c561b26),
	.w3(32'h3b8fdfe2),
	.w4(32'h3b84a116),
	.w5(32'hbb3d174f),
	.w6(32'h3bfe8f0d),
	.w7(32'hbc28a484),
	.w8(32'hbc161fac),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45cb94),
	.w1(32'h3b978636),
	.w2(32'h3c25077d),
	.w3(32'hbb7f8e0c),
	.w4(32'hba6785ea),
	.w5(32'hbba4d51b),
	.w6(32'hbbac7fe8),
	.w7(32'hbc0ad6e0),
	.w8(32'h3bbad779),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3a629),
	.w1(32'hb90f18ef),
	.w2(32'h3bf9fdf9),
	.w3(32'hba215120),
	.w4(32'hbb0f4957),
	.w5(32'h3aa28e5c),
	.w6(32'h3b6b71b9),
	.w7(32'hbae2dfe5),
	.w8(32'hbc0c000b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34ad94),
	.w1(32'h3c064057),
	.w2(32'h3c0c5cc8),
	.w3(32'hbb869e57),
	.w4(32'hb9caefdb),
	.w5(32'h3b0da4a3),
	.w6(32'hbba081dc),
	.w7(32'hbb4dedc1),
	.w8(32'h3c7d1b97),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0669f7),
	.w1(32'hbc41b431),
	.w2(32'hbc872c77),
	.w3(32'hbbde4cef),
	.w4(32'hbc01ad46),
	.w5(32'hbb639c65),
	.w6(32'h3bb6da9b),
	.w7(32'h3b2ca172),
	.w8(32'hbc6be2c6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb090869),
	.w1(32'hbbca8482),
	.w2(32'hbb16d119),
	.w3(32'hbc1b666b),
	.w4(32'hbbc014af),
	.w5(32'h3aa786d1),
	.w6(32'hbc4efd04),
	.w7(32'hbb326bb5),
	.w8(32'h3c0f2164),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39918dcd),
	.w1(32'h3bbb7459),
	.w2(32'h38923d93),
	.w3(32'h3b2d7030),
	.w4(32'hbbe275b7),
	.w5(32'hba8c69a9),
	.w6(32'hba2a827b),
	.w7(32'hbba1406e),
	.w8(32'h3ba9f04b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9694c),
	.w1(32'h3b83d262),
	.w2(32'h3b943116),
	.w3(32'hbb3b8189),
	.w4(32'hbc0906f6),
	.w5(32'hbcfb03a7),
	.w6(32'hbb9b4b35),
	.w7(32'h3baf7f9b),
	.w8(32'h3c809ce6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37f2f4),
	.w1(32'hbb75c826),
	.w2(32'hbc8d9e79),
	.w3(32'h39dbabcd),
	.w4(32'h3b3654ab),
	.w5(32'hbc88dc6d),
	.w6(32'h3c0384f5),
	.w7(32'hbbbc4ca3),
	.w8(32'hbc80ba4f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51c4f4),
	.w1(32'h3b1cd2d7),
	.w2(32'h3b3bb842),
	.w3(32'hbbc8db14),
	.w4(32'h3ace98d6),
	.w5(32'hbb1df4a1),
	.w6(32'hbc1c0928),
	.w7(32'h3b985f30),
	.w8(32'h3bfc1b2c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07f78),
	.w1(32'h3870a291),
	.w2(32'hbb16a2f4),
	.w3(32'h3b853080),
	.w4(32'h3c0b081b),
	.w5(32'hbaaf4282),
	.w6(32'h3c09469c),
	.w7(32'h3c693994),
	.w8(32'h3bbddfb2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2bf36),
	.w1(32'h3a7eacf5),
	.w2(32'h3b05bb2c),
	.w3(32'h3c861619),
	.w4(32'hba293fd7),
	.w5(32'hbbdca68f),
	.w6(32'h3c590998),
	.w7(32'hbbc2c760),
	.w8(32'hbbdd42e1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdabab),
	.w1(32'h3b48498b),
	.w2(32'hbb81af83),
	.w3(32'hbb8a0277),
	.w4(32'hbae2a545),
	.w5(32'hbb309923),
	.w6(32'h3a9b68c2),
	.w7(32'h3aa0fb63),
	.w8(32'hbbb36a1e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0949b7),
	.w1(32'h3c3e9873),
	.w2(32'hbb9c39cc),
	.w3(32'hbbda3dd6),
	.w4(32'h3c210f1b),
	.w5(32'h3b535c6e),
	.w6(32'hbc0614f2),
	.w7(32'h3b0142e0),
	.w8(32'hba80dbad),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c221d55),
	.w1(32'hbb368a17),
	.w2(32'hbbd84241),
	.w3(32'h3b6167df),
	.w4(32'h3b8ce66d),
	.w5(32'h3aa982bd),
	.w6(32'h3c126e2a),
	.w7(32'hbbb5e11b),
	.w8(32'hbbb59f1e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfe0eb),
	.w1(32'h3bc0a850),
	.w2(32'h3bf608d0),
	.w3(32'hbae02266),
	.w4(32'hbb28a026),
	.w5(32'hbb85f73a),
	.w6(32'hbb340ece),
	.w7(32'hbc81bae6),
	.w8(32'hbc3c7601),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadc5af),
	.w1(32'h3b88dc48),
	.w2(32'h3b03ef68),
	.w3(32'h3ba1bd96),
	.w4(32'h3bddc163),
	.w5(32'h3c2cdea4),
	.w6(32'h3bcd7eaf),
	.w7(32'hba16d183),
	.w8(32'h3c38f30f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8a4b6),
	.w1(32'h3a69f50b),
	.w2(32'h3b477e19),
	.w3(32'h3bf40da5),
	.w4(32'h3b3d1b28),
	.w5(32'h3bba4554),
	.w6(32'h3c578b4d),
	.w7(32'h3ac4a336),
	.w8(32'h393a60ff),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8309a3),
	.w1(32'h3b3085cc),
	.w2(32'hbb18f0cd),
	.w3(32'h3b37df10),
	.w4(32'hbaec2efb),
	.w5(32'h3be1aeab),
	.w6(32'h3b2abb93),
	.w7(32'h3b1e0f85),
	.w8(32'h3c485f77),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb109650),
	.w1(32'h3ac8d4d4),
	.w2(32'h3bf3c642),
	.w3(32'hbc0f9b25),
	.w4(32'hbb6c631f),
	.w5(32'h3c8b2212),
	.w6(32'hbb85150e),
	.w7(32'hba4433ef),
	.w8(32'h3c1a461e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59cc3f),
	.w1(32'hbb4f0ba0),
	.w2(32'hbbd070f6),
	.w3(32'hbb9a18aa),
	.w4(32'hba14d338),
	.w5(32'hbc722d5f),
	.w6(32'h3c3c0026),
	.w7(32'hbc7b2771),
	.w8(32'hbc1be319),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5f35f),
	.w1(32'hbaa83d4c),
	.w2(32'hbbc6d4fb),
	.w3(32'hbbb44ae7),
	.w4(32'h3950d6a3),
	.w5(32'hbb54ef7e),
	.w6(32'hbb9c3e09),
	.w7(32'hbb653164),
	.w8(32'hbb554f9a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab44ea),
	.w1(32'hbaaaa633),
	.w2(32'h3b7380f1),
	.w3(32'h3aae0962),
	.w4(32'hbb34f3ce),
	.w5(32'h3bc8abc3),
	.w6(32'hbb4b17c8),
	.w7(32'hba5a907c),
	.w8(32'h3ba5a8ca),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c5f1f),
	.w1(32'hbc04e86e),
	.w2(32'hbc499347),
	.w3(32'h3b14120a),
	.w4(32'hb88511ff),
	.w5(32'hbc34cf48),
	.w6(32'h3ba5aac2),
	.w7(32'hbbd9fa0f),
	.w8(32'hbbd3724e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c1f59),
	.w1(32'h3a1d1afb),
	.w2(32'h3a732253),
	.w3(32'hbb38346c),
	.w4(32'hbbaed6aa),
	.w5(32'hbbd98d5a),
	.w6(32'h3ad32ea5),
	.w7(32'hbad4fcf3),
	.w8(32'h3adf1e35),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba70751),
	.w1(32'hbbaf2b94),
	.w2(32'h396ed1d6),
	.w3(32'hba116abb),
	.w4(32'h3b75f1bd),
	.w5(32'h3a8b8f8a),
	.w6(32'h3bc96f95),
	.w7(32'hba9cd908),
	.w8(32'hbba232ca),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf7f1b),
	.w1(32'h3b03569a),
	.w2(32'h3b63f851),
	.w3(32'h3b96785c),
	.w4(32'h3c425ce6),
	.w5(32'h3c1e588a),
	.w6(32'h3b55cbed),
	.w7(32'h3c601e26),
	.w8(32'h3c380272),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c638750),
	.w1(32'hbc69889b),
	.w2(32'hbcae6e58),
	.w3(32'h3c8ab73c),
	.w4(32'hbb7a5824),
	.w5(32'hbc8f0d73),
	.w6(32'h3b7303ca),
	.w7(32'hbb9da759),
	.w8(32'hba70a441),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd6ffa),
	.w1(32'h3c17ffb7),
	.w2(32'hbc3231bd),
	.w3(32'hbc189472),
	.w4(32'h3b490730),
	.w5(32'hbaee08fa),
	.w6(32'h3c05cb97),
	.w7(32'hbad14af5),
	.w8(32'h3c10b13e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4ae80),
	.w1(32'hbbf42942),
	.w2(32'hbc4130aa),
	.w3(32'h3c449db4),
	.w4(32'h3a4dd33e),
	.w5(32'hbc5dda52),
	.w6(32'h3c27c0e1),
	.w7(32'hbb0dac12),
	.w8(32'hbc85e59c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2acd51),
	.w1(32'h3ae20da8),
	.w2(32'h3bea5f12),
	.w3(32'hbc10b679),
	.w4(32'hbb529ec6),
	.w5(32'h3b0eb601),
	.w6(32'hbc4c4ac4),
	.w7(32'hbb758a6f),
	.w8(32'h3961a1fe),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb9cd2),
	.w1(32'hba952c1e),
	.w2(32'hba9e5ab4),
	.w3(32'h3b7b1b31),
	.w4(32'hbb0516a0),
	.w5(32'h3ab848af),
	.w6(32'h3b4bea35),
	.w7(32'hb72e27ff),
	.w8(32'hb8cd854b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacddb9c),
	.w1(32'hbaa419c1),
	.w2(32'h391e5af8),
	.w3(32'hba971754),
	.w4(32'h3ae94944),
	.w5(32'h3aab1cbd),
	.w6(32'hbaa50789),
	.w7(32'h3aa33105),
	.w8(32'h3a5988ba),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf7b1e),
	.w1(32'h3b389ec4),
	.w2(32'h3a88f844),
	.w3(32'hbb24cbba),
	.w4(32'h3a82be8d),
	.w5(32'h3ac32109),
	.w6(32'h3aeec2dc),
	.w7(32'hba22e0e9),
	.w8(32'h3a98c494),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a976d94),
	.w1(32'h3972f9e6),
	.w2(32'hbaf4cef4),
	.w3(32'h3aa5cf03),
	.w4(32'hba50809f),
	.w5(32'hbafe4109),
	.w6(32'h3b0fe9a1),
	.w7(32'hbb0df13b),
	.w8(32'hbb216154),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395e5977),
	.w1(32'hbaa0c0ef),
	.w2(32'hbb16c10f),
	.w3(32'hb825d02b),
	.w4(32'hbb1cf688),
	.w5(32'hbb075d07),
	.w6(32'h39cce47b),
	.w7(32'hbb33b578),
	.w8(32'h38564ffe),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8866b78),
	.w1(32'h38936304),
	.w2(32'hbb49dff4),
	.w3(32'hba9ffbdc),
	.w4(32'h3a606fcc),
	.w5(32'h39ecabe7),
	.w6(32'h39e27161),
	.w7(32'hba405386),
	.w8(32'hba50f1d2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7d84b),
	.w1(32'h3b2738f4),
	.w2(32'hbabd3a52),
	.w3(32'h3b5c82e0),
	.w4(32'h3b33e111),
	.w5(32'hbabacd07),
	.w6(32'h3b9442f5),
	.w7(32'h399827b5),
	.w8(32'hbb37930a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb029fb4),
	.w1(32'h3af0be5d),
	.w2(32'h38c8104a),
	.w3(32'hba5bc5a3),
	.w4(32'h37e7f9e1),
	.w5(32'hbb399a8d),
	.w6(32'hba0aaa22),
	.w7(32'h39443fe9),
	.w8(32'h38fe272d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf595e4),
	.w1(32'h3a07eeec),
	.w2(32'hbb3fd3e9),
	.w3(32'hbabbadfc),
	.w4(32'h3b146e41),
	.w5(32'hbad8ab09),
	.w6(32'h39632f88),
	.w7(32'h3b023b9c),
	.w8(32'hba5545f0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50a3c7),
	.w1(32'hbaaf1245),
	.w2(32'hbb949f3e),
	.w3(32'h3ae25fcd),
	.w4(32'h3aeab987),
	.w5(32'hbaec9ce8),
	.w6(32'h3b514236),
	.w7(32'h3a13d19a),
	.w8(32'hbb26d282),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53c620),
	.w1(32'h3b8fd956),
	.w2(32'h3b969022),
	.w3(32'hbafcac8a),
	.w4(32'h3ba7996c),
	.w5(32'h3a791cf3),
	.w6(32'hba956639),
	.w7(32'h3b9d8130),
	.w8(32'h3b71b96f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c112937),
	.w1(32'hba464c5d),
	.w2(32'hbb20f04f),
	.w3(32'h3c0230f7),
	.w4(32'hb822bae9),
	.w5(32'hbab09dd0),
	.w6(32'h3bdb30b4),
	.w7(32'hba43296b),
	.w8(32'hbb1dbd7d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94af68),
	.w1(32'h3921c488),
	.w2(32'hba9305f2),
	.w3(32'h3a27b71e),
	.w4(32'h3aa3bf60),
	.w5(32'hba85f5fa),
	.w6(32'h38fafe43),
	.w7(32'h3a2075eb),
	.w8(32'hbad63b40),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9294a66),
	.w1(32'h3b1b8300),
	.w2(32'h3b0bdc0c),
	.w3(32'hb90c5b3a),
	.w4(32'h3a5099b1),
	.w5(32'h3b945c39),
	.w6(32'h3a08c902),
	.w7(32'h3adb803f),
	.w8(32'h3b921526),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f8b63),
	.w1(32'hbb032fbf),
	.w2(32'hbb18ddf4),
	.w3(32'h3baaf982),
	.w4(32'hbb1d27e4),
	.w5(32'h392b3f3b),
	.w6(32'h3a480cb5),
	.w7(32'hbaf0c711),
	.w8(32'hbae7fcbd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4e256),
	.w1(32'hbb6e8fd0),
	.w2(32'hb9015855),
	.w3(32'hbb00d5a9),
	.w4(32'hb9d2acb8),
	.w5(32'h3ba1e1fe),
	.w6(32'hba873643),
	.w7(32'hba93df41),
	.w8(32'hbb2bf476),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80fe8f),
	.w1(32'h3a53aa86),
	.w2(32'hba7d412c),
	.w3(32'hbbaa94bc),
	.w4(32'hba254a2e),
	.w5(32'hba938023),
	.w6(32'hbb91c575),
	.w7(32'h39d09a3a),
	.w8(32'h38018a66),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb169f0c),
	.w1(32'h3a3f7f8a),
	.w2(32'hba84b5da),
	.w3(32'hbac39354),
	.w4(32'hba800100),
	.w5(32'hba50c90d),
	.w6(32'hbaa08456),
	.w7(32'hba8ad7be),
	.w8(32'hb899c544),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf65ed6),
	.w1(32'h3ad7b14c),
	.w2(32'hba538870),
	.w3(32'hbb143304),
	.w4(32'hba87d673),
	.w5(32'h3b082822),
	.w6(32'hba117239),
	.w7(32'h3b641732),
	.w8(32'h3b375a30),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babcb64),
	.w1(32'h3b186cf8),
	.w2(32'hbb269d8b),
	.w3(32'h3bea9b75),
	.w4(32'h3b22ad70),
	.w5(32'hbb15cd43),
	.w6(32'h3b99688a),
	.w7(32'hbb3cbc27),
	.w8(32'hbb811cd9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7db660),
	.w1(32'hb9ecaeb6),
	.w2(32'h3a89e393),
	.w3(32'hba8577fe),
	.w4(32'hb9f985cd),
	.w5(32'h3b88ed82),
	.w6(32'hbae40ec7),
	.w7(32'hbb2a7de0),
	.w8(32'hba5ad60e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84cef1),
	.w1(32'hba892ac8),
	.w2(32'hbc57d28d),
	.w3(32'h3beb55e6),
	.w4(32'h3b79086e),
	.w5(32'hbbaeedc8),
	.w6(32'h3bab0a54),
	.w7(32'h3a8b0afc),
	.w8(32'hbc096b8e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc83f4),
	.w1(32'hb9030a66),
	.w2(32'h3aae1f3d),
	.w3(32'hba19fe69),
	.w4(32'hbaae2e32),
	.w5(32'h3a4e3c0b),
	.w6(32'hbb5a7184),
	.w7(32'hba78b14c),
	.w8(32'h3aca6506),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f5d1b),
	.w1(32'hbb4ae9c7),
	.w2(32'hbbb91825),
	.w3(32'h3b01bde8),
	.w4(32'h3a235fa2),
	.w5(32'hbba7151f),
	.w6(32'h3b25c2f4),
	.w7(32'hbabb1a4e),
	.w8(32'hbbcc507f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37c698),
	.w1(32'hba4ad36a),
	.w2(32'hbb696365),
	.w3(32'h3b99a269),
	.w4(32'h3b889e4b),
	.w5(32'h3a16e56d),
	.w6(32'h3b17730d),
	.w7(32'h3b78a352),
	.w8(32'hb98642d7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c29f3),
	.w1(32'hbaa1fb9b),
	.w2(32'h3aaae6e6),
	.w3(32'hb941fdf3),
	.w4(32'hbb49ca4a),
	.w5(32'h3aa59bba),
	.w6(32'hbb5b896c),
	.w7(32'hbb8893fe),
	.w8(32'hbb2f2545),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fe18f),
	.w1(32'hb8f11a42),
	.w2(32'hbb101a36),
	.w3(32'hbb090594),
	.w4(32'hbab9a2c3),
	.w5(32'h3b580a79),
	.w6(32'h3b0064a1),
	.w7(32'h39998b7b),
	.w8(32'hb9a5692e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab10cc9),
	.w1(32'h3a71be0f),
	.w2(32'hbad58c12),
	.w3(32'h3a7e502b),
	.w4(32'h3b52ea32),
	.w5(32'hba5b8423),
	.w6(32'h3b2d59ff),
	.w7(32'h3987b1b5),
	.w8(32'hbb903e34),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ab7ef),
	.w1(32'h39bd9ea5),
	.w2(32'hbab33e61),
	.w3(32'h3b6ad296),
	.w4(32'h3bb89794),
	.w5(32'h3ac3cf82),
	.w6(32'hba64c292),
	.w7(32'hbb091ce2),
	.w8(32'hbbe3bda4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c6e6f),
	.w1(32'h3c082335),
	.w2(32'h3ab36a52),
	.w3(32'hba5dc497),
	.w4(32'h3ad74e1e),
	.w5(32'hbb4f53e1),
	.w6(32'h3b5e76fd),
	.w7(32'h3c22f2a7),
	.w8(32'h3bc5b952),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ca6d5),
	.w1(32'h3b114a48),
	.w2(32'h3ab52cab),
	.w3(32'hbc02fbba),
	.w4(32'h3b60d1ba),
	.w5(32'h3bf958f2),
	.w6(32'hbc2fdec5),
	.w7(32'h3a6587d4),
	.w8(32'h3b9d1dc4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04e5f5),
	.w1(32'h3aee151c),
	.w2(32'h3b2259f8),
	.w3(32'hbaeefcc5),
	.w4(32'hb920e909),
	.w5(32'h39d71830),
	.w6(32'hbb49d007),
	.w7(32'h3a7c6571),
	.w8(32'hbaca2bfc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a95b0f),
	.w1(32'hba67b024),
	.w2(32'hbbe903a7),
	.w3(32'hbaaf3839),
	.w4(32'h3b8f1586),
	.w5(32'h3a9f8d52),
	.w6(32'hba3eb4fb),
	.w7(32'h3aac5e47),
	.w8(32'hbb97cce1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926e6ea),
	.w1(32'h3b103bd5),
	.w2(32'hb80fbbc4),
	.w3(32'hbb451e09),
	.w4(32'hba01c446),
	.w5(32'h3a97d6ae),
	.w6(32'h3a9b5382),
	.w7(32'h3b1013de),
	.w8(32'h3acb469a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec477d),
	.w1(32'hba7af27c),
	.w2(32'hbbc4c0eb),
	.w3(32'hbb8d4f4d),
	.w4(32'h382dcee5),
	.w5(32'hbb0b33d1),
	.w6(32'hba8dc194),
	.w7(32'h3bb15cb2),
	.w8(32'h3b105d52),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e5527),
	.w1(32'hba90dec7),
	.w2(32'hbb4f4a23),
	.w3(32'hb96acbe9),
	.w4(32'hb95987cc),
	.w5(32'hba931e12),
	.w6(32'hbb240e0a),
	.w7(32'h3ac7179e),
	.w8(32'hb9cdf46c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31af4d),
	.w1(32'h3b35073a),
	.w2(32'h3a0be3b8),
	.w3(32'h3aaabcaf),
	.w4(32'h3b55301b),
	.w5(32'hb95915b5),
	.w6(32'h3b25a06c),
	.w7(32'h3b1b87e8),
	.w8(32'hb9119d45),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aea51a),
	.w1(32'hba9e7a49),
	.w2(32'hbb393e6e),
	.w3(32'h393855cc),
	.w4(32'hba2ed697),
	.w5(32'hbb42c397),
	.w6(32'hba4dd0c6),
	.w7(32'hba8179aa),
	.w8(32'hbb983fd7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67c78b),
	.w1(32'hb78d50c5),
	.w2(32'hbb666178),
	.w3(32'h3ba190e4),
	.w4(32'hba1e10ed),
	.w5(32'hbb80e642),
	.w6(32'h3b1c70eb),
	.w7(32'hbb8a4cc3),
	.w8(32'hbbb49939),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9279c6),
	.w1(32'h3b24852e),
	.w2(32'h3b52c9d2),
	.w3(32'hba1a5979),
	.w4(32'h3b4d9edb),
	.w5(32'h3ae8986a),
	.w6(32'h3a8b0a42),
	.w7(32'h3b05af98),
	.w8(32'h382def34),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc617c),
	.w1(32'hbbaac7dd),
	.w2(32'hb9ed498b),
	.w3(32'hbb771b6c),
	.w4(32'hba51e2c8),
	.w5(32'hb974909b),
	.w6(32'hbac713e0),
	.w7(32'hbb71621f),
	.w8(32'hbb2de073),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4744df),
	.w1(32'h39294fca),
	.w2(32'h3ae220c0),
	.w3(32'hbb899139),
	.w4(32'h39573b54),
	.w5(32'h3b150bb5),
	.w6(32'hba4d3abc),
	.w7(32'h3a603939),
	.w8(32'h391c32ae),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add52e6),
	.w1(32'h3ba387eb),
	.w2(32'h3b2391be),
	.w3(32'hbb8dad48),
	.w4(32'h3a7e7cd6),
	.w5(32'h3ac01930),
	.w6(32'hba0b0fef),
	.w7(32'h3bae19bd),
	.w8(32'h3ae5b6e6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafae113),
	.w1(32'hbb8ebcd6),
	.w2(32'hbbfaeb32),
	.w3(32'hbb28cd7b),
	.w4(32'hbafd7419),
	.w5(32'hbb7e78f6),
	.w6(32'hbae72467),
	.w7(32'hbaf0300a),
	.w8(32'hbb654841),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f0fdf),
	.w1(32'h3ab8c9ba),
	.w2(32'h3ab07ba7),
	.w3(32'hbaa8e166),
	.w4(32'h3a7d8419),
	.w5(32'h3a8c7078),
	.w6(32'hbb322224),
	.w7(32'h3ad14360),
	.w8(32'hb871980e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5339a7),
	.w1(32'hb97ffd86),
	.w2(32'hbaa92640),
	.w3(32'h3a623770),
	.w4(32'hb9f86eb8),
	.w5(32'hba9e9d3d),
	.w6(32'h3acae1f0),
	.w7(32'hba19e073),
	.w8(32'hbab7fba3),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3755e),
	.w1(32'hbb0d2ab3),
	.w2(32'hba30f2f9),
	.w3(32'hb92aa66d),
	.w4(32'hba471ff1),
	.w5(32'h3a87d580),
	.w6(32'h391a0f08),
	.w7(32'hba7382e6),
	.w8(32'hba5bd008),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab771e1),
	.w1(32'h396b0921),
	.w2(32'hba908553),
	.w3(32'h3b1f8cb8),
	.w4(32'h38ba1990),
	.w5(32'hbb143814),
	.w6(32'h3a7c4b36),
	.w7(32'hbac87449),
	.w8(32'hbb185ce7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7105ce),
	.w1(32'h3abb9b7b),
	.w2(32'hb8a25132),
	.w3(32'h39802c6c),
	.w4(32'hb855829c),
	.w5(32'h3abc5917),
	.w6(32'hb94469bb),
	.w7(32'hb9c5d09b),
	.w8(32'h3b06e718),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5166c8),
	.w1(32'hba8a17bd),
	.w2(32'h3a060ad9),
	.w3(32'hbadac504),
	.w4(32'hba098fba),
	.w5(32'h3b09fa0e),
	.w6(32'h3a63ffd2),
	.w7(32'h3996173f),
	.w8(32'h384b283b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f3f74),
	.w1(32'h3b17a07f),
	.w2(32'h3872d8a6),
	.w3(32'hba8e3851),
	.w4(32'h3aa5aece),
	.w5(32'h3a836607),
	.w6(32'hbab2651d),
	.w7(32'h3b1bb63f),
	.w8(32'h3a8a0562),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b915c39),
	.w1(32'hb9df00c6),
	.w2(32'hbb91a7ab),
	.w3(32'h3ba02a0b),
	.w4(32'hba3d89a6),
	.w5(32'hba467a06),
	.w6(32'h3ae0bc4d),
	.w7(32'hbba1c888),
	.w8(32'hbb4a1b8c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d5afb),
	.w1(32'hba13a091),
	.w2(32'h3aedc7ee),
	.w3(32'h35fca818),
	.w4(32'hbb3cd797),
	.w5(32'h3b0665a0),
	.w6(32'hbb195e69),
	.w7(32'hbac88d1d),
	.w8(32'h3a67761b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab72d56),
	.w1(32'hba3981c5),
	.w2(32'h3a73e365),
	.w3(32'hbacd9644),
	.w4(32'h39df750e),
	.w5(32'h3b076c19),
	.w6(32'hb8a819ca),
	.w7(32'h3739e026),
	.w8(32'h3a4256fe),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14fb1d),
	.w1(32'hbb32469b),
	.w2(32'hbb268e0a),
	.w3(32'h388922e8),
	.w4(32'hbb2cd097),
	.w5(32'hbb290a14),
	.w6(32'hba4bc8dc),
	.w7(32'hbb39c577),
	.w8(32'hbafa3730),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba919e33),
	.w1(32'h39a2e3aa),
	.w2(32'hba8fd252),
	.w3(32'hbb4ff466),
	.w4(32'hb8a77d0a),
	.w5(32'h39a69186),
	.w6(32'hbb047997),
	.w7(32'hba99fa92),
	.w8(32'hbb132018),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa88fa3),
	.w1(32'h3995a2c9),
	.w2(32'h3a904589),
	.w3(32'hbb33547f),
	.w4(32'hb9e543bf),
	.w5(32'h3b5d029d),
	.w6(32'hbaac0814),
	.w7(32'h39bb6829),
	.w8(32'hb987f1d5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8284b),
	.w1(32'hba451096),
	.w2(32'hbb74cef0),
	.w3(32'hbb858e33),
	.w4(32'hbba84fee),
	.w5(32'hbba18f8a),
	.w6(32'h3b37158a),
	.w7(32'hbab1f674),
	.w8(32'hbb68bd6f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba754af1),
	.w1(32'hbaa5f7a5),
	.w2(32'hbbd61bb7),
	.w3(32'hb9c2989b),
	.w4(32'h3976c016),
	.w5(32'hbb9556f9),
	.w6(32'hb973cce2),
	.w7(32'hbb6502d0),
	.w8(32'hbb8e2171),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9821f95),
	.w1(32'hba499522),
	.w2(32'hba8d1bbc),
	.w3(32'h3a3dca73),
	.w4(32'h39a0d83f),
	.w5(32'h3a28a5a3),
	.w6(32'h3a87e435),
	.w7(32'hba6af8af),
	.w8(32'hbb138312),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafef7da),
	.w1(32'hba0f04fe),
	.w2(32'hbb210afa),
	.w3(32'hbb48c47a),
	.w4(32'hbaa526d2),
	.w5(32'hbb6afaa9),
	.w6(32'hbac39c73),
	.w7(32'h39224b9b),
	.w8(32'hbac52bac),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71bd34),
	.w1(32'h3aa7b661),
	.w2(32'hbab5aa0d),
	.w3(32'hbb029024),
	.w4(32'hb940038f),
	.w5(32'hb83fd244),
	.w6(32'hbb3f8fb0),
	.w7(32'hbab49806),
	.w8(32'hbb419a2b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9daf148),
	.w1(32'hba4ec7c1),
	.w2(32'hbac78d71),
	.w3(32'hba6846b4),
	.w4(32'h3ab192e4),
	.w5(32'hbadc4b6a),
	.w6(32'h3abeb101),
	.w7(32'hba08e6a2),
	.w8(32'hbb10cf76),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca62d1),
	.w1(32'hba00da7d),
	.w2(32'hba209a9f),
	.w3(32'h3a9e5519),
	.w4(32'h3a667054),
	.w5(32'h3ab83277),
	.w6(32'h3b36783f),
	.w7(32'h3a8715cd),
	.w8(32'hbad58a9c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ac236),
	.w1(32'h3970558b),
	.w2(32'hbbde6fd3),
	.w3(32'h3a972002),
	.w4(32'h3b0e2bdc),
	.w5(32'hbb30698d),
	.w6(32'hba79b0ee),
	.w7(32'hbb7af15b),
	.w8(32'hbbb060ff),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5084bd),
	.w1(32'h3b654c9a),
	.w2(32'h3b96701a),
	.w3(32'hbb478a61),
	.w4(32'h3adec4af),
	.w5(32'h3b0e0686),
	.w6(32'hbac8dc17),
	.w7(32'h3b10d886),
	.w8(32'h3b151bee),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46e524),
	.w1(32'hba66aacc),
	.w2(32'hbb833966),
	.w3(32'h3ba63c71),
	.w4(32'h3ac9cb8b),
	.w5(32'hbaa7eda1),
	.w6(32'h3ac46077),
	.w7(32'h3aa926af),
	.w8(32'hbb4bcf6d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74eef1),
	.w1(32'h3a6f763a),
	.w2(32'hbbde1769),
	.w3(32'h3acd3fe3),
	.w4(32'h3ae02687),
	.w5(32'hbb28766c),
	.w6(32'h3b2ac6fc),
	.w7(32'hba626f73),
	.w8(32'hbbaf8053),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56d4a6),
	.w1(32'h3a9ffa2a),
	.w2(32'hba25f399),
	.w3(32'hbb134d5e),
	.w4(32'h3a871e1c),
	.w5(32'hb935a048),
	.w6(32'hba754236),
	.w7(32'h3a8f0f9f),
	.w8(32'hba906b93),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ba842),
	.w1(32'hbaa5bbbc),
	.w2(32'hbb4a85fe),
	.w3(32'hba42d0c7),
	.w4(32'h3ac3418c),
	.w5(32'hb9f7ee33),
	.w6(32'h39c15c87),
	.w7(32'h3b1ee4f4),
	.w8(32'h38bb9c64),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0871c2),
	.w1(32'hba6945e8),
	.w2(32'hbb20b102),
	.w3(32'h3b08dfca),
	.w4(32'hbb317476),
	.w5(32'hbae2ec08),
	.w6(32'h3ac4fc48),
	.w7(32'hba874aca),
	.w8(32'hbb1b4cc1),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0f6f1),
	.w1(32'hbb32cc68),
	.w2(32'h3a8f5a74),
	.w3(32'hbb0c35c1),
	.w4(32'hbb8f95a5),
	.w5(32'hbaa68b53),
	.w6(32'hbb663c6e),
	.w7(32'hbbb17a39),
	.w8(32'hbb43905c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36fe61),
	.w1(32'h388c36f0),
	.w2(32'hba9abd79),
	.w3(32'hb9b2a51e),
	.w4(32'hbb08f693),
	.w5(32'hba3e180d),
	.w6(32'hb8489a50),
	.w7(32'hbadfb23a),
	.w8(32'hbb108929),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9773093),
	.w1(32'hbb34ef19),
	.w2(32'hba72b4fe),
	.w3(32'hbb364439),
	.w4(32'hbb182c4b),
	.w5(32'hbacc95e5),
	.w6(32'hbad6c6c2),
	.w7(32'hba9c4c2b),
	.w8(32'hbaaf27a0),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e38a51),
	.w1(32'h3979a1e0),
	.w2(32'h3a2ef302),
	.w3(32'hb95759a1),
	.w4(32'h3b094f9f),
	.w5(32'h3afa8a08),
	.w6(32'h361c076d),
	.w7(32'h3b336dc8),
	.w8(32'h3b62e430),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a457f2f),
	.w1(32'h3ab83d52),
	.w2(32'h39bf75c9),
	.w3(32'h3a645ce3),
	.w4(32'h3b2eaf8e),
	.w5(32'h3aa451ec),
	.w6(32'h3afbf3d9),
	.w7(32'h3ae2a672),
	.w8(32'h387c223a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5d8d1),
	.w1(32'h3acc56cf),
	.w2(32'h3a377609),
	.w3(32'hb8130969),
	.w4(32'hba84e6f5),
	.w5(32'h3b20a88d),
	.w6(32'hbb088214),
	.w7(32'hbae9a475),
	.w8(32'h3805b201),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3eac9a),
	.w1(32'h3a9044c7),
	.w2(32'h39e78694),
	.w3(32'h3a310f5b),
	.w4(32'hba0af2c2),
	.w5(32'hb9a9acbe),
	.w6(32'hb94dfb62),
	.w7(32'hb921e3e6),
	.w8(32'hbad2d32c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb714c),
	.w1(32'hb9d269d6),
	.w2(32'h3a6c07c2),
	.w3(32'hba659836),
	.w4(32'h39331de8),
	.w5(32'h3a8334de),
	.w6(32'hb9356a07),
	.w7(32'h397d7d0f),
	.w8(32'h388529e7),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34e30c),
	.w1(32'hbb09d9be),
	.w2(32'hbaf61bd3),
	.w3(32'h3723fc87),
	.w4(32'hbadcd51c),
	.w5(32'hba8af36c),
	.w6(32'hbaf132f2),
	.w7(32'hbb897d6b),
	.w8(32'hbb4387b3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b788ad0),
	.w1(32'h3a837818),
	.w2(32'h3aa62a27),
	.w3(32'h3b1d9844),
	.w4(32'hba1530ea),
	.w5(32'hb9b91048),
	.w6(32'h3ac04514),
	.w7(32'hb84e5701),
	.w8(32'hba262961),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c11fd),
	.w1(32'hbb7ff0bd),
	.w2(32'hbc1c83f5),
	.w3(32'h3b04e6f1),
	.w4(32'hba9e76ef),
	.w5(32'hbc08b3d8),
	.w6(32'h3b176571),
	.w7(32'hbba069a7),
	.w8(32'hbc295dcc),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59b17c),
	.w1(32'hbb9df4ce),
	.w2(32'h3b391fb5),
	.w3(32'hbaa74974),
	.w4(32'hbbaaab28),
	.w5(32'hb98eebec),
	.w6(32'hbb616ce8),
	.w7(32'hbbf5b9ef),
	.w8(32'hbc072f5d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2ba58),
	.w1(32'h3bc5d713),
	.w2(32'h3b89ec70),
	.w3(32'h3b85915d),
	.w4(32'h3b804878),
	.w5(32'h3a9de5d9),
	.w6(32'h3b824c07),
	.w7(32'h3a94efb4),
	.w8(32'hbac837d9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5b8e7),
	.w1(32'hb9afbd1e),
	.w2(32'h3a672edc),
	.w3(32'h3bea5ed2),
	.w4(32'h3abebf5c),
	.w5(32'h3b8f6138),
	.w6(32'h3bc43eb1),
	.w7(32'h3b520246),
	.w8(32'h3b8c75fa),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb889319),
	.w1(32'hba92a492),
	.w2(32'hbb40dc40),
	.w3(32'hbc0acf09),
	.w4(32'hbb8f6086),
	.w5(32'hbb59a2ea),
	.w6(32'hbbb90000),
	.w7(32'hbbaf1507),
	.w8(32'hbb510105),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81569b),
	.w1(32'hbabeb015),
	.w2(32'h3b439df7),
	.w3(32'hba828b12),
	.w4(32'h3b0e6f1f),
	.w5(32'h3bbba60e),
	.w6(32'hbb1951e6),
	.w7(32'h39fdea26),
	.w8(32'h3aae2b45),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cbd68),
	.w1(32'h3b3c27a2),
	.w2(32'h3bb23b8c),
	.w3(32'hb970f73b),
	.w4(32'h3b4f4507),
	.w5(32'h3b65af5d),
	.w6(32'h3a8294df),
	.w7(32'h3b1bc840),
	.w8(32'h3b5edaac),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b357676),
	.w1(32'h389c362c),
	.w2(32'h383b6a09),
	.w3(32'h3b3a068c),
	.w4(32'h3ace05bb),
	.w5(32'h39a8bd4f),
	.w6(32'h3aa8d8e9),
	.w7(32'h3a599f08),
	.w8(32'h3a831bff),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac99bdc),
	.w1(32'hba26e9aa),
	.w2(32'hbab99038),
	.w3(32'h3abe7a90),
	.w4(32'hb9ea0acb),
	.w5(32'hba4fa570),
	.w6(32'h3b2c30a6),
	.w7(32'hb9f753c6),
	.w8(32'hbac96ae2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86944e),
	.w1(32'hbb0c390d),
	.w2(32'hbb36a681),
	.w3(32'hb936ebc7),
	.w4(32'hb9d18384),
	.w5(32'hbafe532e),
	.w6(32'h398bda75),
	.w7(32'hba827e47),
	.w8(32'hb97e2af8),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8ad3e),
	.w1(32'h3a1760fc),
	.w2(32'hba72e4be),
	.w3(32'hbb2ea502),
	.w4(32'hbaa1d927),
	.w5(32'h387cec42),
	.w6(32'hba810a84),
	.w7(32'hba9d84a5),
	.w8(32'h3822090b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02217e),
	.w1(32'h3b13f52d),
	.w2(32'h3ad74391),
	.w3(32'hbb5fff6e),
	.w4(32'hba3f4ed0),
	.w5(32'hbb18e292),
	.w6(32'hba90d5ab),
	.w7(32'h39a460fc),
	.w8(32'hba548969),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad44b84),
	.w1(32'h3ad3568d),
	.w2(32'h39bd2958),
	.w3(32'h39fd6ac8),
	.w4(32'h3b346ea7),
	.w5(32'h3acf0b03),
	.w6(32'h3ab91aae),
	.w7(32'h3b16cce6),
	.w8(32'h3b130197),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08b295),
	.w1(32'h3b7b0e11),
	.w2(32'h3ad0b3ef),
	.w3(32'h3bb5da26),
	.w4(32'h3a5b74a1),
	.w5(32'h3b1a7bc1),
	.w6(32'h3bdc992a),
	.w7(32'hbad74e66),
	.w8(32'hbb174eaa),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4874a3),
	.w1(32'h3b53aacf),
	.w2(32'h39efbf67),
	.w3(32'h39c8a323),
	.w4(32'h3b0062cc),
	.w5(32'h3a97f394),
	.w6(32'h39948f7c),
	.w7(32'h3addaa0f),
	.w8(32'h3af4c082),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55f170),
	.w1(32'h3a212b50),
	.w2(32'h3aa19703),
	.w3(32'h3a985175),
	.w4(32'h3ad9380a),
	.w5(32'h3ae55f5e),
	.w6(32'h3a984a98),
	.w7(32'h3a64f0ee),
	.w8(32'hba508a95),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade6326),
	.w1(32'h3b2fe079),
	.w2(32'hba8e92fe),
	.w3(32'hbb2fa2d4),
	.w4(32'h3934ff35),
	.w5(32'h3a05f712),
	.w6(32'hba805802),
	.w7(32'h3b52a29a),
	.w8(32'h3afe14fc),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b452c9e),
	.w1(32'hba7d64ba),
	.w2(32'hbb18f9e4),
	.w3(32'hba13bcd8),
	.w4(32'hbb5a2d94),
	.w5(32'hba602d59),
	.w6(32'hbab6c7dc),
	.w7(32'hbae3c495),
	.w8(32'hbb3ff954),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d4fa2),
	.w1(32'h3a0ae6a3),
	.w2(32'hb88609b6),
	.w3(32'h3a9d9699),
	.w4(32'h3ab1f50d),
	.w5(32'h3b24a9a7),
	.w6(32'h39c99bd2),
	.w7(32'h3aedf01b),
	.w8(32'h3a1b6664),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9724a),
	.w1(32'h3a671c12),
	.w2(32'hba6e7aac),
	.w3(32'hbaaeb976),
	.w4(32'h39d58ceb),
	.w5(32'hba51d206),
	.w6(32'hba9b4ff2),
	.w7(32'h3a86a09e),
	.w8(32'hbb826591),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c2472),
	.w1(32'h3b00f8d6),
	.w2(32'h39276198),
	.w3(32'hbaf0ab37),
	.w4(32'h3b038d70),
	.w5(32'hbb1a629d),
	.w6(32'hbb17a677),
	.w7(32'h39b0fdd1),
	.w8(32'hbb2762ef),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc47755),
	.w1(32'hbb84edc1),
	.w2(32'hbbe0f729),
	.w3(32'hbaaca247),
	.w4(32'hbbc41ee8),
	.w5(32'hbb5c8ff6),
	.w6(32'hbb5273e8),
	.w7(32'hbbe3912e),
	.w8(32'hbbb206f2),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba472e9a),
	.w1(32'hbb8c3b62),
	.w2(32'hbba73ea1),
	.w3(32'hba08ea93),
	.w4(32'hb9f32b2f),
	.w5(32'hbb0532e3),
	.w6(32'hba4689f8),
	.w7(32'hbac99f41),
	.w8(32'hbb3bc4cd),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20c8f6),
	.w1(32'hbb5a409c),
	.w2(32'hbbbae741),
	.w3(32'hbb4634f3),
	.w4(32'h38ca8d2b),
	.w5(32'hbb398424),
	.w6(32'hbaaff9d4),
	.w7(32'hbac7a663),
	.w8(32'hbbce7a3d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939f653),
	.w1(32'h39459374),
	.w2(32'h3a5b4a94),
	.w3(32'hbabeb9d6),
	.w4(32'h3acb979a),
	.w5(32'h3b8ff4f4),
	.w6(32'hb6f2fd68),
	.w7(32'h3b071ff4),
	.w8(32'h3b68be0e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafd87e),
	.w1(32'hbb689324),
	.w2(32'hba95edd5),
	.w3(32'hba2464c7),
	.w4(32'hbb1d9a8c),
	.w5(32'hbb285ebe),
	.w6(32'hba0cb323),
	.w7(32'h398f9132),
	.w8(32'hba107851),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29b951),
	.w1(32'h3a4b3c14),
	.w2(32'h3aca4b16),
	.w3(32'hba983813),
	.w4(32'h3b35c451),
	.w5(32'h3a959da7),
	.w6(32'hba65acb6),
	.w7(32'h3b8c4f01),
	.w8(32'h3b3e352f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd3bfe),
	.w1(32'h3a16929f),
	.w2(32'h39a8b4dc),
	.w3(32'h3ae860e6),
	.w4(32'h3aa90d19),
	.w5(32'h3a79cebe),
	.w6(32'h39d13d72),
	.w7(32'h3af93b3a),
	.w8(32'hb9e56b5a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a71d4),
	.w1(32'hbaa6c5be),
	.w2(32'h39f55332),
	.w3(32'hb9a92eba),
	.w4(32'hb9e6dbd1),
	.w5(32'h3acf8e26),
	.w6(32'h3a4d2632),
	.w7(32'h392a1805),
	.w8(32'h3a8e236d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cfb31),
	.w1(32'hba786204),
	.w2(32'hbb0fa7b5),
	.w3(32'hb9ee7c55),
	.w4(32'h3b079730),
	.w5(32'hba8ff74b),
	.w6(32'hb825a96b),
	.w7(32'h3ac94928),
	.w8(32'h3a89268e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b175e2b),
	.w1(32'h3ad35269),
	.w2(32'h3a3102ed),
	.w3(32'h3b4a6c29),
	.w4(32'h3a9e15bd),
	.w5(32'h38e07f3e),
	.w6(32'h3b2bfddb),
	.w7(32'h3b46989a),
	.w8(32'h3b144572),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ad1d2),
	.w1(32'h3b73d197),
	.w2(32'hba594572),
	.w3(32'h3a828a81),
	.w4(32'h3b0c9473),
	.w5(32'h39a74e8c),
	.w6(32'h3af554dd),
	.w7(32'h3aff048e),
	.w8(32'hba6db801),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb685560d),
	.w1(32'h3a6dd898),
	.w2(32'hb7e39fb7),
	.w3(32'hbacad051),
	.w4(32'hb91076ec),
	.w5(32'hb9e8d9e0),
	.w6(32'hb9eb33b4),
	.w7(32'hba8026cb),
	.w8(32'hbaf3cb00),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e934d),
	.w1(32'hbaca528c),
	.w2(32'hbbb729d9),
	.w3(32'hbb49c0f7),
	.w4(32'h3b4915c6),
	.w5(32'hbb45f7ab),
	.w6(32'hbb601243),
	.w7(32'h3b097e9d),
	.w8(32'hbbc943d1),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a34de5),
	.w1(32'h3b54921d),
	.w2(32'hbae4654b),
	.w3(32'hbb1232f2),
	.w4(32'h3acba959),
	.w5(32'hb9ff76b9),
	.w6(32'hbb49276a),
	.w7(32'h3ad24a67),
	.w8(32'h39fe3bec),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7dd26),
	.w1(32'hba30eca4),
	.w2(32'hbb65a824),
	.w3(32'h3a64a42b),
	.w4(32'hba790a46),
	.w5(32'hbb7df70a),
	.w6(32'hba09927f),
	.w7(32'hba960768),
	.w8(32'hbb673fcd),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b6ccdc),
	.w1(32'hba0a34f7),
	.w2(32'hbbd5ed68),
	.w3(32'h3aa3d683),
	.w4(32'hb9f1b88a),
	.w5(32'hbbb4d1d8),
	.w6(32'h3a934347),
	.w7(32'hb9c3fc14),
	.w8(32'hbc091e5e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba4ca9),
	.w1(32'hbba63577),
	.w2(32'hbbd35149),
	.w3(32'h3b3d989b),
	.w4(32'hba29b310),
	.w5(32'hbb214d63),
	.w6(32'h3a3285a9),
	.w7(32'hbaf45fb3),
	.w8(32'hbbf91410),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dad6e),
	.w1(32'hbac40216),
	.w2(32'hbb7f8762),
	.w3(32'hba2ea102),
	.w4(32'hb9d39b3f),
	.w5(32'hba501e95),
	.w6(32'h3a1f1bc0),
	.w7(32'hbae0f5cb),
	.w8(32'hbb7ad6f8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8256e),
	.w1(32'h3a2474b9),
	.w2(32'hbb2c479d),
	.w3(32'hbb056c21),
	.w4(32'hba381e2b),
	.w5(32'hbb06e279),
	.w6(32'hbb0b3a0b),
	.w7(32'hb9f3965f),
	.w8(32'hbb8db191),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c776e),
	.w1(32'h3a9f44fc),
	.w2(32'hb8bd94c0),
	.w3(32'hbacf27b0),
	.w4(32'h3ae757fe),
	.w5(32'h389476ef),
	.w6(32'hba912896),
	.w7(32'h3aab0d54),
	.w8(32'h3947dc71),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a012e4e),
	.w1(32'h3b82cf77),
	.w2(32'h3aff0a14),
	.w3(32'h3a518c35),
	.w4(32'h3b53e9f0),
	.w5(32'hba072d1f),
	.w6(32'h3aad1cd1),
	.w7(32'h3b35a511),
	.w8(32'h3ad8cc46),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcc3fb),
	.w1(32'h3b036e4d),
	.w2(32'hb9a6b8af),
	.w3(32'h3b1bb363),
	.w4(32'h3afcadd5),
	.w5(32'h3af217e3),
	.w6(32'h3b784f3f),
	.w7(32'h3a961452),
	.w8(32'hb9b3300d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07f278),
	.w1(32'hba860fb0),
	.w2(32'hba32c31d),
	.w3(32'h3b534acf),
	.w4(32'hb82636c8),
	.w5(32'hb978b9d4),
	.w6(32'h3b2562be),
	.w7(32'h3a95f714),
	.w8(32'hba47df0b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88ed3f),
	.w1(32'hba3e51e3),
	.w2(32'h3a8fb458),
	.w3(32'hbb611df5),
	.w4(32'hba7cd98d),
	.w5(32'h3a983a35),
	.w6(32'hbb412f45),
	.w7(32'h39e943af),
	.w8(32'hba80ab5e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb861b52),
	.w1(32'h3af5dfb8),
	.w2(32'h3a0619fd),
	.w3(32'hbbc515b2),
	.w4(32'h3acefb9d),
	.w5(32'h3ac137c0),
	.w6(32'hbb9a5d95),
	.w7(32'h3b07ed6f),
	.w8(32'hba73a6fa),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f7eb4),
	.w1(32'hbb020434),
	.w2(32'hbb95f8af),
	.w3(32'hb893e0a4),
	.w4(32'hbaf2a29f),
	.w5(32'hbc20e7b2),
	.w6(32'hba5d53ab),
	.w7(32'h3abe7492),
	.w8(32'hbbe1d76c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09994e),
	.w1(32'hbb1197f0),
	.w2(32'hbbc30b64),
	.w3(32'hbadcc79e),
	.w4(32'hbb2a5486),
	.w5(32'h3a891e91),
	.w6(32'hbb78bde4),
	.w7(32'hbb94f1f4),
	.w8(32'hbb5aa879),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90c429),
	.w1(32'hbb11ae77),
	.w2(32'h3be1a6c4),
	.w3(32'hbb0dff20),
	.w4(32'hbab1237c),
	.w5(32'h3c80fc19),
	.w6(32'hbad92c0f),
	.w7(32'hbb7b154d),
	.w8(32'hbc468a6c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6f6ed),
	.w1(32'hbc23c919),
	.w2(32'hbb1e8069),
	.w3(32'hba962c19),
	.w4(32'hbbc9fd48),
	.w5(32'h3b815c51),
	.w6(32'h3bba5a3f),
	.w7(32'hbc0f37cc),
	.w8(32'hbbc195e4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c25cf),
	.w1(32'hbba914b9),
	.w2(32'hba306d50),
	.w3(32'hbb3963db),
	.w4(32'h3b5f37c2),
	.w5(32'h3ba734ea),
	.w6(32'hbbc0d44b),
	.w7(32'h3ac1022a),
	.w8(32'hbaa6fcb5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375b4e8a),
	.w1(32'hbb467383),
	.w2(32'hbc059354),
	.w3(32'h398350f7),
	.w4(32'h3b9010e2),
	.w5(32'hbca02cfd),
	.w6(32'hba008ae5),
	.w7(32'hbb447c0c),
	.w8(32'hbc3401ce),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc356a56),
	.w1(32'hbb7733e7),
	.w2(32'h3ae5c8eb),
	.w3(32'hbc21799a),
	.w4(32'hbb007b44),
	.w5(32'hbb983007),
	.w6(32'hbc0fea6e),
	.w7(32'hbb24051b),
	.w8(32'hbb6f7de0),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b796c6c),
	.w1(32'h3abe38b7),
	.w2(32'h3bca2f83),
	.w3(32'hba9f1ce3),
	.w4(32'h3915268a),
	.w5(32'h3c139171),
	.w6(32'h3ad3ca8f),
	.w7(32'hbbc9ff81),
	.w8(32'h3a8b7950),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ca185),
	.w1(32'hbbb0a7c1),
	.w2(32'hbb181617),
	.w3(32'h3baf589d),
	.w4(32'hbaf4c817),
	.w5(32'h3bb5dd0e),
	.w6(32'h3b20dba2),
	.w7(32'hbb7bd280),
	.w8(32'hbb50082b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53b86f),
	.w1(32'hbb650523),
	.w2(32'h3aa05a82),
	.w3(32'hbc0652d0),
	.w4(32'hbb81d390),
	.w5(32'hbb85f9a9),
	.w6(32'hbc1eb5f1),
	.w7(32'hbb2efb56),
	.w8(32'h39eca619),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a37b6),
	.w1(32'hbb3146de),
	.w2(32'hbb1499ed),
	.w3(32'hbc507544),
	.w4(32'hbb199fe5),
	.w5(32'hbb2cba94),
	.w6(32'hb9ee7ae4),
	.w7(32'h3b6c4eae),
	.w8(32'h3b4231ae),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a9304),
	.w1(32'hbc3f15c6),
	.w2(32'hbbb44bcd),
	.w3(32'h39e1d983),
	.w4(32'hbc0e1408),
	.w5(32'hbc1a4125),
	.w6(32'hbc74e4d0),
	.w7(32'hbc4cf49a),
	.w8(32'hbc6f209e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba19b4d),
	.w1(32'hbb314ff1),
	.w2(32'hbb1a000d),
	.w3(32'hbc1cef9d),
	.w4(32'hb9f83c85),
	.w5(32'hba927948),
	.w6(32'hbb18fc1c),
	.w7(32'hba215cae),
	.w8(32'hbabb611e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396ce002),
	.w1(32'hbad40a98),
	.w2(32'h3b840845),
	.w3(32'h3a8f40b3),
	.w4(32'hbb7c49f0),
	.w5(32'h3ae4e855),
	.w6(32'h39c8ea43),
	.w7(32'hbb88db9a),
	.w8(32'hbbaa1a45),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85b26d),
	.w1(32'h3a10dd59),
	.w2(32'hbc15afcc),
	.w3(32'hb908dc20),
	.w4(32'h3b1f80a5),
	.w5(32'h3b2a50b2),
	.w6(32'hbad101f2),
	.w7(32'hb9651924),
	.w8(32'h3bc4eb07),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5e135),
	.w1(32'hbbb5733c),
	.w2(32'hbbd045d5),
	.w3(32'h3bd6903f),
	.w4(32'hbb23ee12),
	.w5(32'hba9c53ff),
	.w6(32'h3bbc3df4),
	.w7(32'hbb3f7761),
	.w8(32'hbba84d2e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ed5f3),
	.w1(32'h3bc69110),
	.w2(32'h3bd14771),
	.w3(32'hbb8da16d),
	.w4(32'h3c196e1c),
	.w5(32'h3c177e94),
	.w6(32'hbbe25485),
	.w7(32'h3ac7c732),
	.w8(32'hbb6e5f90),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ff4b4),
	.w1(32'hbc140513),
	.w2(32'hbc32bc30),
	.w3(32'hb92d998b),
	.w4(32'hba917187),
	.w5(32'h3bd3f54f),
	.w6(32'h3c27baf3),
	.w7(32'hbc46e008),
	.w8(32'hbb5e7202),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc951b3),
	.w1(32'h39aa07e4),
	.w2(32'hb9bb5bb2),
	.w3(32'hbbd1bfdd),
	.w4(32'hba5d3cd8),
	.w5(32'h3ba453cc),
	.w6(32'hba59955d),
	.w7(32'hbbf86a2a),
	.w8(32'hbc76f1b6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f107d),
	.w1(32'h3a0ee8d7),
	.w2(32'h3b0202b5),
	.w3(32'hbb57d1b2),
	.w4(32'hba4adb0a),
	.w5(32'h3b469c3e),
	.w6(32'h3b7a7303),
	.w7(32'hbc1394d5),
	.w8(32'hb9cc77a5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae4dca),
	.w1(32'h3b8fabd0),
	.w2(32'hbbefa194),
	.w3(32'h3a9acce4),
	.w4(32'hbad76c97),
	.w5(32'hbba096b6),
	.w6(32'h3b53be11),
	.w7(32'h3a91b666),
	.w8(32'h389a1488),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0e317),
	.w1(32'hbc0bdf3a),
	.w2(32'hbbe177e1),
	.w3(32'hba7abfa9),
	.w4(32'h3b9fdec8),
	.w5(32'hba3c5359),
	.w6(32'hbb47bfc3),
	.w7(32'hbac4f252),
	.w8(32'hbbeb1939),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c459d),
	.w1(32'h3c85f6c8),
	.w2(32'h3aab7be4),
	.w3(32'hba562155),
	.w4(32'h3c0f9449),
	.w5(32'hbb301dc9),
	.w6(32'hbb97273c),
	.w7(32'h3bcd44a8),
	.w8(32'hba170b89),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9b2b8),
	.w1(32'hbae3b31d),
	.w2(32'hbbe8a5eb),
	.w3(32'h3a670ee9),
	.w4(32'hbb70c92f),
	.w5(32'h3ab7a26b),
	.w6(32'h3af0ab0d),
	.w7(32'hba70fc4d),
	.w8(32'hbc6b3cbc),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0add46),
	.w1(32'hbb1ee3b7),
	.w2(32'hbbaece92),
	.w3(32'hbc5b4554),
	.w4(32'h3b865f5b),
	.w5(32'h3c29d343),
	.w6(32'hbb87e77a),
	.w7(32'hbbbb81f4),
	.w8(32'hbbdc3555),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39387f43),
	.w1(32'h3ad9ca56),
	.w2(32'h3b14d44b),
	.w3(32'hb9af3d21),
	.w4(32'hbaedc684),
	.w5(32'h3c070bca),
	.w6(32'h3b175afd),
	.w7(32'hbb19240f),
	.w8(32'h3b6b2187),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2d2e7),
	.w1(32'hbbcaac02),
	.w2(32'hbaae9080),
	.w3(32'hbaf0361f),
	.w4(32'hbb87d1ba),
	.w5(32'h3c5d9942),
	.w6(32'hbbd45763),
	.w7(32'hbb821b4c),
	.w8(32'h3a43b6db),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33e289),
	.w1(32'hbb6eca34),
	.w2(32'hbb064f53),
	.w3(32'hbb74ab65),
	.w4(32'h3b089613),
	.w5(32'h3bb3c29e),
	.w6(32'hbb242c64),
	.w7(32'hbbce769f),
	.w8(32'hbbc66667),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bd55b),
	.w1(32'h3c16e0af),
	.w2(32'h3b62db3f),
	.w3(32'hbbc12668),
	.w4(32'h3c222471),
	.w5(32'hbb65233b),
	.w6(32'h3a5cf677),
	.w7(32'h3c3763a8),
	.w8(32'h3aa3d8b1),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d861b),
	.w1(32'hbb3a6229),
	.w2(32'hbb4a9d13),
	.w3(32'h3ad75c68),
	.w4(32'hbb971d01),
	.w5(32'hbbce3e72),
	.w6(32'hbb694323),
	.w7(32'hba86e085),
	.w8(32'h3b9ec6c3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb550c95),
	.w1(32'h39ec329a),
	.w2(32'h3b6767bc),
	.w3(32'h3b5f85f4),
	.w4(32'hbb01457c),
	.w5(32'hbb2d3ef4),
	.w6(32'hbc081a98),
	.w7(32'h3bfc370a),
	.w8(32'hb92488ec),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba081f90),
	.w1(32'hbbb96ad2),
	.w2(32'hbbae689b),
	.w3(32'hbb4d4706),
	.w4(32'h3aef03ce),
	.w5(32'hb92230be),
	.w6(32'hbbbb8a97),
	.w7(32'hbb928cdf),
	.w8(32'h3b00b9e8),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb207525),
	.w1(32'hbc0dc241),
	.w2(32'hbbcd8fd9),
	.w3(32'hbb0bb9e9),
	.w4(32'hbbb8d8a6),
	.w5(32'h3b879348),
	.w6(32'h3aa0a5c2),
	.w7(32'hbaf0e56f),
	.w8(32'hbbc40f55),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97910f),
	.w1(32'h3b75a7af),
	.w2(32'h3b622859),
	.w3(32'hbb445b95),
	.w4(32'h3bb360f2),
	.w5(32'h3b7d48e5),
	.w6(32'h3909e218),
	.w7(32'hbb135637),
	.w8(32'hbc6ad0a2),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f723d),
	.w1(32'hbb5556d4),
	.w2(32'hbaa676b0),
	.w3(32'hba4055e0),
	.w4(32'hbb2f3ff5),
	.w5(32'h3bef7e9f),
	.w6(32'hbb5a2a17),
	.w7(32'hbc32c696),
	.w8(32'hbbf0c948),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb7f4d),
	.w1(32'h3ac5456a),
	.w2(32'hbb9075e7),
	.w3(32'hbac8b670),
	.w4(32'hbb05b786),
	.w5(32'hb9d0a03b),
	.w6(32'hbb0744cc),
	.w7(32'hba2cfa56),
	.w8(32'h3b62b55f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb905c99),
	.w1(32'h3aae7853),
	.w2(32'hb97e548a),
	.w3(32'h3af63e8d),
	.w4(32'h3b5b3daa),
	.w5(32'h398027f3),
	.w6(32'h3ba04b54),
	.w7(32'h383393cf),
	.w8(32'hbaa416e7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb113c8f),
	.w1(32'hba57fb94),
	.w2(32'h3bd477b8),
	.w3(32'hbb09ed13),
	.w4(32'h3af9288c),
	.w5(32'h3c29626b),
	.w6(32'hbac33c9b),
	.w7(32'hbb8e8a18),
	.w8(32'h3a78e649),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b6cd9),
	.w1(32'hbb3f9f26),
	.w2(32'h3b4cede9),
	.w3(32'h3af015c8),
	.w4(32'hba047dd1),
	.w5(32'h3c148149),
	.w6(32'h3b08476a),
	.w7(32'h3bc9056b),
	.w8(32'h3bcecfc9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb87e7d),
	.w1(32'hb9c0ec73),
	.w2(32'hbb9b100c),
	.w3(32'h3b88b9d9),
	.w4(32'h3a02574e),
	.w5(32'h3ab9875a),
	.w6(32'hbbc5f74f),
	.w7(32'h3c252f01),
	.w8(32'h3bab4d5d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d2e9d),
	.w1(32'hbb52aac2),
	.w2(32'hbb9fdac3),
	.w3(32'h3c1e91b2),
	.w4(32'hbacc58e3),
	.w5(32'h3c195603),
	.w6(32'h3b536351),
	.w7(32'h3b3551c1),
	.w8(32'hbb38b122),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6ae73),
	.w1(32'h3c05b7b5),
	.w2(32'h3c457b87),
	.w3(32'hbb52fcd7),
	.w4(32'h3b4b6352),
	.w5(32'h38a052f1),
	.w6(32'hb91e2d4b),
	.w7(32'hbb2d4687),
	.w8(32'hb8ac60b0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbc2f0),
	.w1(32'hbbd86017),
	.w2(32'hbc1055b4),
	.w3(32'hbb848b38),
	.w4(32'h3b480a7b),
	.w5(32'hbb4c4e13),
	.w6(32'h3ba63e1e),
	.w7(32'hbb292631),
	.w8(32'hbc0af5fb),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc013137),
	.w1(32'hbbaf1d34),
	.w2(32'hbb5ab6ac),
	.w3(32'hbbe296f4),
	.w4(32'hbbabdbfe),
	.w5(32'hbb82a5dc),
	.w6(32'hbb08d230),
	.w7(32'h3b3f31e2),
	.w8(32'hbb1777f5),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01ca35),
	.w1(32'hba8ca4e7),
	.w2(32'hbc50f280),
	.w3(32'h3b70a990),
	.w4(32'hbaac0c30),
	.w5(32'hbc2863e3),
	.w6(32'hbbcbe930),
	.w7(32'h39bb4fcf),
	.w8(32'hbc509f2e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084cef),
	.w1(32'h3b33b339),
	.w2(32'h3ac41ffe),
	.w3(32'hbbfa7002),
	.w4(32'hb9dc7480),
	.w5(32'h3b7fca74),
	.w6(32'h3b2fce9a),
	.w7(32'h3aa0e52b),
	.w8(32'hbb21b8fc),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1512b0),
	.w1(32'hbab09fea),
	.w2(32'hbba941f3),
	.w3(32'hbbb95bfd),
	.w4(32'h39773c3f),
	.w5(32'hbb331582),
	.w6(32'hbb5db444),
	.w7(32'hb9282784),
	.w8(32'hbbd1e455),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84c60e),
	.w1(32'h3b890fb5),
	.w2(32'h3bf2c86b),
	.w3(32'hbac8016b),
	.w4(32'h3c0e3462),
	.w5(32'h3b65ad15),
	.w6(32'hbbc3e604),
	.w7(32'h3bb03d29),
	.w8(32'h3a096ee5),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9606bc6),
	.w1(32'hbc31e52e),
	.w2(32'hbada7dec),
	.w3(32'hb90504fc),
	.w4(32'h3986dc2b),
	.w5(32'h3bdf8864),
	.w6(32'h3a843994),
	.w7(32'hbb9a9a8f),
	.w8(32'hbc1f7541),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55e87b),
	.w1(32'hbba94c3b),
	.w2(32'hbc425f51),
	.w3(32'h3a42e284),
	.w4(32'hbb2ff0fd),
	.w5(32'hbb332775),
	.w6(32'hbc314fcd),
	.w7(32'hbb42bca2),
	.w8(32'hbb931e33),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe16163),
	.w1(32'hbb7fab8b),
	.w2(32'hba8ccd3c),
	.w3(32'hbabb2e83),
	.w4(32'hbb1b5ff4),
	.w5(32'hbbc4e678),
	.w6(32'hb772542d),
	.w7(32'hb99f4a7c),
	.w8(32'hbbce5bb7),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a21757),
	.w1(32'hbafab46a),
	.w2(32'h3a4cb246),
	.w3(32'h3b0380f5),
	.w4(32'hba8eab6f),
	.w5(32'h3baa0218),
	.w6(32'hba9ddfbc),
	.w7(32'hb9b06a86),
	.w8(32'hbb4176f5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06e6ae),
	.w1(32'h3be87466),
	.w2(32'h3ba7ee22),
	.w3(32'h3b215636),
	.w4(32'hba87db8b),
	.w5(32'hba9a2b9b),
	.w6(32'h3bb057b5),
	.w7(32'h3bba38f3),
	.w8(32'hbad382e8),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca4893),
	.w1(32'hbb91822b),
	.w2(32'hbb2fb5bd),
	.w3(32'h395cfecf),
	.w4(32'hba7367da),
	.w5(32'h3bb16ab7),
	.w6(32'hbb37035c),
	.w7(32'hbbcb60fe),
	.w8(32'hbbb9f891),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ecf99),
	.w1(32'h3a467e73),
	.w2(32'h3b9a3d51),
	.w3(32'h3abb558f),
	.w4(32'hb9de4ead),
	.w5(32'hbb1431df),
	.w6(32'hb9994301),
	.w7(32'hbb051f4f),
	.w8(32'hbbbe1cfc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe662f4),
	.w1(32'hbb83f4f6),
	.w2(32'hba6229ff),
	.w3(32'hbcab6c8d),
	.w4(32'hbb86a3d7),
	.w5(32'h3bf7a649),
	.w6(32'hbb863ae4),
	.w7(32'hbbb3ba44),
	.w8(32'hbc2c80b5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28281a),
	.w1(32'hbc1c9295),
	.w2(32'hbbfd8eeb),
	.w3(32'h3b54f012),
	.w4(32'h3afcf03d),
	.w5(32'h3c1d8b62),
	.w6(32'h3b4875a4),
	.w7(32'hbb94f79c),
	.w8(32'hbbf9b21a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22127a),
	.w1(32'hbaea1778),
	.w2(32'h3bbb2518),
	.w3(32'hbbb60710),
	.w4(32'h3baed5c1),
	.w5(32'h3c21e10d),
	.w6(32'h3b11cef9),
	.w7(32'hbbbec753),
	.w8(32'hbbde6935),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf3f96),
	.w1(32'h3c07dee7),
	.w2(32'hbbe86606),
	.w3(32'hbc00bb76),
	.w4(32'hbbc84d0d),
	.w5(32'hbc507317),
	.w6(32'hbc592d7d),
	.w7(32'h3962a345),
	.w8(32'h3c41c977),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule