module layer_10_featuremap_102(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d09c660),
	.w1(32'h3b0a6adc),
	.w2(32'hbc8ac260),
	.w3(32'h3c81b578),
	.w4(32'h389180da),
	.w5(32'hbbb95e72),
	.w6(32'hbaf240e7),
	.w7(32'hbbb8efa8),
	.w8(32'hba0ac348),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b983a5a),
	.w1(32'h3b995e19),
	.w2(32'h3b9a9e55),
	.w3(32'h3959435a),
	.w4(32'hbb9cf6b6),
	.w5(32'h3b0c6b48),
	.w6(32'hbae5ab3c),
	.w7(32'hbb71d9c5),
	.w8(32'hb8c24b2d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7f104),
	.w1(32'h3b6f1c6a),
	.w2(32'h38f348df),
	.w3(32'h3ac22dbf),
	.w4(32'hbbc103e6),
	.w5(32'hbbe816fb),
	.w6(32'hba9d281e),
	.w7(32'hbba76a0b),
	.w8(32'hbba76ba0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc7652),
	.w1(32'h3bdd076b),
	.w2(32'h3c1c3047),
	.w3(32'hbb8d6e16),
	.w4(32'hbbe876c8),
	.w5(32'hbb89459a),
	.w6(32'hbb107ee8),
	.w7(32'h3b12ab33),
	.w8(32'h3be33317),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d2f8f),
	.w1(32'hbc0cd1de),
	.w2(32'h3c467387),
	.w3(32'h3b602752),
	.w4(32'hbaa86984),
	.w5(32'h3ad27ebb),
	.w6(32'hbb2d1042),
	.w7(32'hb9b0bf75),
	.w8(32'hbc15102b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20911e),
	.w1(32'hbcd2af13),
	.w2(32'hba6ba63a),
	.w3(32'hbc0aebb4),
	.w4(32'hbc6a47cc),
	.w5(32'hbb0c97fa),
	.w6(32'hbcb61463),
	.w7(32'hbb031e45),
	.w8(32'h3c25c457),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d11f4f0),
	.w1(32'h3bd3f9ef),
	.w2(32'h3c2b4a3a),
	.w3(32'h3c777cb3),
	.w4(32'hbabc2a9f),
	.w5(32'h3bcf70ac),
	.w6(32'hbad676c3),
	.w7(32'hbb12c801),
	.w8(32'hba6e3fb1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4bda5),
	.w1(32'hbcf0a4f9),
	.w2(32'h3b1e588b),
	.w3(32'h3b0bd61e),
	.w4(32'hbc5442f1),
	.w5(32'h3b65e302),
	.w6(32'hbcf98e96),
	.w7(32'h38a430be),
	.w8(32'h3c8cce35),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d15feb9),
	.w1(32'hbc8c0d8e),
	.w2(32'h3b821989),
	.w3(32'h3c89d9b0),
	.w4(32'hbbe782b4),
	.w5(32'h3ab8e1e6),
	.w6(32'hbbfe3744),
	.w7(32'h3b250942),
	.w8(32'h3b2ac27d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c441f07),
	.w1(32'h3ced55bf),
	.w2(32'hb92e0610),
	.w3(32'h3b34cf3b),
	.w4(32'h3aa17486),
	.w5(32'hbbeb8cd0),
	.w6(32'h3c3116ac),
	.w7(32'hbc6fbb19),
	.w8(32'hbc90a57d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd23ccd5),
	.w1(32'hbc143105),
	.w2(32'h3b8f3176),
	.w3(32'hbc94971a),
	.w4(32'hbbe5cf11),
	.w5(32'hbaa1c22e),
	.w6(32'hbb656538),
	.w7(32'h3b6b78cc),
	.w8(32'h3c1ec9a1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ced5630),
	.w1(32'hbc182234),
	.w2(32'hbbb15130),
	.w3(32'h3c01bb16),
	.w4(32'hba174d19),
	.w5(32'h3becd7c6),
	.w6(32'hbc2482e2),
	.w7(32'hbb26d6c0),
	.w8(32'h3c24d4e3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c436a29),
	.w1(32'hbca37945),
	.w2(32'hb9da1195),
	.w3(32'h3c00eacb),
	.w4(32'hbc4c2a6e),
	.w5(32'hb924aca0),
	.w6(32'hbc9fc2c1),
	.w7(32'hbba6dcea),
	.w8(32'h3bc8d019),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ab9c3),
	.w1(32'hbd154955),
	.w2(32'hbb6783f8),
	.w3(32'h3c086061),
	.w4(32'hbbdd54d9),
	.w5(32'h3bd00b94),
	.w6(32'hbcb092ad),
	.w7(32'h3be04f41),
	.w8(32'h3cc5444e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4f6650),
	.w1(32'hba0a6877),
	.w2(32'hbaccbb7f),
	.w3(32'h3cc3659f),
	.w4(32'hbb5be25f),
	.w5(32'h3ba7a838),
	.w6(32'hbb05e84c),
	.w7(32'hbb5c6679),
	.w8(32'h3a2c3bb7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9557005),
	.w1(32'hbc6e2785),
	.w2(32'h3c021617),
	.w3(32'hba3c5ed7),
	.w4(32'hbbd0f935),
	.w5(32'h3b646eed),
	.w6(32'hbc1704ac),
	.w7(32'h3bb6ef6c),
	.w8(32'h3b74861a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4aa398),
	.w1(32'hbb82abeb),
	.w2(32'hba3e61dd),
	.w3(32'h3afabe04),
	.w4(32'hba84b235),
	.w5(32'hbb19744c),
	.w6(32'hbbe71df0),
	.w7(32'hb9190c60),
	.w8(32'hbaa4623b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eeb0b2),
	.w1(32'h3c8fd5b2),
	.w2(32'h3b692a19),
	.w3(32'hbb0f14e2),
	.w4(32'hb8568975),
	.w5(32'hbb26d677),
	.w6(32'h3af4dd15),
	.w7(32'hbc3b0896),
	.w8(32'hbc73097e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdab9f0),
	.w1(32'hbb3cfd57),
	.w2(32'hbac0e44f),
	.w3(32'hbc36e036),
	.w4(32'hbc005629),
	.w5(32'hbb1cca45),
	.w6(32'hbc2dc670),
	.w7(32'hbbd96113),
	.w8(32'hbab4862e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb802a9b),
	.w1(32'hbc8882aa),
	.w2(32'h3a3f1620),
	.w3(32'h3a50fc0c),
	.w4(32'hbc203675),
	.w5(32'hba8af6a7),
	.w6(32'hbc30447e),
	.w7(32'hbb0857ea),
	.w8(32'hbb051f74),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c010ac4),
	.w1(32'hbce97be3),
	.w2(32'hbb61151c),
	.w3(32'h39de174d),
	.w4(32'hbc5c22f1),
	.w5(32'hb8c3661b),
	.w6(32'hbc8a6afa),
	.w7(32'h3b8a5338),
	.w8(32'h3bf983ad),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8be72),
	.w1(32'hbbb81e75),
	.w2(32'hbb3abb08),
	.w3(32'h3bba3a09),
	.w4(32'hbc38a70f),
	.w5(32'hbbe4cb0b),
	.w6(32'h3b972dfd),
	.w7(32'h3aaac355),
	.w8(32'h3b9d3634),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf22e16),
	.w1(32'hbb137f4f),
	.w2(32'h3c1cd67d),
	.w3(32'h3c07ab7c),
	.w4(32'hbb9cea6a),
	.w5(32'h3c1085c7),
	.w6(32'hbb0d63bb),
	.w7(32'h3b67b5b6),
	.w8(32'hbab84a33),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75e831),
	.w1(32'hbce3bc9f),
	.w2(32'h3bbb4909),
	.w3(32'h3b61b2fa),
	.w4(32'hbc2fa0c9),
	.w5(32'h3bd1069d),
	.w6(32'hbcaa3eb6),
	.w7(32'h3b9f01ed),
	.w8(32'h3c90877e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d142d84),
	.w1(32'h3b99c4df),
	.w2(32'h3ad99ea1),
	.w3(32'h3c8160ca),
	.w4(32'hbb19ef6d),
	.w5(32'h3a293612),
	.w6(32'h3b30510e),
	.w7(32'h390d9579),
	.w8(32'hbb2e7d36),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47dc3c),
	.w1(32'hbb333a74),
	.w2(32'h3bcd689d),
	.w3(32'hb9f87788),
	.w4(32'hbb84bdc5),
	.w5(32'hbb802081),
	.w6(32'hbbfba18a),
	.w7(32'hbb5f6244),
	.w8(32'h3b36271a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56cdbf),
	.w1(32'hbcb9d194),
	.w2(32'hbb9765ad),
	.w3(32'h3ba71a43),
	.w4(32'hbc5575e0),
	.w5(32'hbb3bca8d),
	.w6(32'hbc898326),
	.w7(32'hbb8232ee),
	.w8(32'h3adbd8ab),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a3d00),
	.w1(32'h3c0686b5),
	.w2(32'h3b8f972e),
	.w3(32'h3bdac941),
	.w4(32'hbaaf3956),
	.w5(32'hbaf8f5e7),
	.w6(32'h3c15ee60),
	.w7(32'h3baef69c),
	.w8(32'h397f0ce6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99048cd),
	.w1(32'hbaefe1bc),
	.w2(32'hbc24355f),
	.w3(32'hbb3048d4),
	.w4(32'h3b216746),
	.w5(32'hbc170d87),
	.w6(32'hbb39fcc0),
	.w7(32'hbc20aa8c),
	.w8(32'hbbcdfd2e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1088ee),
	.w1(32'hba4baa0f),
	.w2(32'hbb63813b),
	.w3(32'h3b04ae68),
	.w4(32'h3aa2e7ba),
	.w5(32'hbacf67b0),
	.w6(32'h3be22788),
	.w7(32'h3a802180),
	.w8(32'h3ab25ef6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d8d72),
	.w1(32'hbcaa2f9c),
	.w2(32'hbb82c7cd),
	.w3(32'hbb7d292c),
	.w4(32'hbc3c75e8),
	.w5(32'hbb0b533e),
	.w6(32'hbc785f84),
	.w7(32'hba936063),
	.w8(32'h3ba09965),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64b2e7),
	.w1(32'hbcbacc7e),
	.w2(32'hbb620783),
	.w3(32'h3b653aad),
	.w4(32'hbc448362),
	.w5(32'hba45a95c),
	.w6(32'hbc976e9e),
	.w7(32'hbb051c70),
	.w8(32'h3be9e5b0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c955179),
	.w1(32'hbb8afb1b),
	.w2(32'hbbbf9169),
	.w3(32'h3bd57dcd),
	.w4(32'h3a6b47d3),
	.w5(32'hbabbcd0e),
	.w6(32'hbaeabad6),
	.w7(32'hbb82b87e),
	.w8(32'h3be43ee9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91e9cc),
	.w1(32'hbc4863b8),
	.w2(32'hbb21784a),
	.w3(32'h3c020fc6),
	.w4(32'hbbd9077f),
	.w5(32'hba4e6287),
	.w6(32'hbc23fa04),
	.w7(32'hbc1a6b30),
	.w8(32'hbaa6ede3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91bcfb),
	.w1(32'h3c79b677),
	.w2(32'hbbf88290),
	.w3(32'h3c3465b4),
	.w4(32'h3ac05312),
	.w5(32'hbc12b45f),
	.w6(32'h3be13543),
	.w7(32'hbc542859),
	.w8(32'hbcb866e9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0a502f),
	.w1(32'hbc870e9c),
	.w2(32'h3ad8cecb),
	.w3(32'hbca980aa),
	.w4(32'hbc2cf61b),
	.w5(32'hba267601),
	.w6(32'hbc93d516),
	.w7(32'hbb0940e0),
	.w8(32'h3bd9fb91),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54d0e8),
	.w1(32'h3b84e843),
	.w2(32'h3bc14ebd),
	.w3(32'hbc0f31eb),
	.w4(32'hbc2e8add),
	.w5(32'h3acee6c7),
	.w6(32'hba9a10eb),
	.w7(32'hbc405265),
	.w8(32'hbb721947),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d746d),
	.w1(32'h3b46327a),
	.w2(32'h3b473df4),
	.w3(32'h37be0f33),
	.w4(32'hbbdf7d81),
	.w5(32'hbadd17c6),
	.w6(32'h3a855fbf),
	.w7(32'hbb93fc5f),
	.w8(32'hbba23672),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ef6da),
	.w1(32'hbcc4d755),
	.w2(32'h3bbd30d9),
	.w3(32'hba04af0b),
	.w4(32'hbc41d303),
	.w5(32'h3b878d64),
	.w6(32'hbc28efc3),
	.w7(32'h3c08db82),
	.w8(32'h3c6b80b8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d06e00d),
	.w1(32'hbb12475f),
	.w2(32'h3b2713e0),
	.w3(32'h3c6453c4),
	.w4(32'hbc14355d),
	.w5(32'hb9893b2a),
	.w6(32'hbbb8d536),
	.w7(32'hbb57a8d9),
	.w8(32'hba617d88),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c2b15),
	.w1(32'h3b60fd62),
	.w2(32'hbafcd908),
	.w3(32'h3ac917e7),
	.w4(32'h3a888728),
	.w5(32'hbb12e105),
	.w6(32'h3a0a589a),
	.w7(32'h3a0f9856),
	.w8(32'h3af9b39c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add176f),
	.w1(32'hbbb94e4a),
	.w2(32'h3a6cf3c0),
	.w3(32'h3a8eff85),
	.w4(32'hbc22b40d),
	.w5(32'hbb55fb5f),
	.w6(32'hbbfbc4c3),
	.w7(32'hbb1660cd),
	.w8(32'hbb6ebd00),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52d6da),
	.w1(32'hbcb07565),
	.w2(32'h39a248a2),
	.w3(32'hbac69ad2),
	.w4(32'hbc4b05cf),
	.w5(32'h3b00b679),
	.w6(32'hbc7cfb76),
	.w7(32'h3b04fe6f),
	.w8(32'h3c2ca4c2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf82bf),
	.w1(32'h3d5b9b37),
	.w2(32'h3b9aa2c5),
	.w3(32'h3c52cd3b),
	.w4(32'h3c587f05),
	.w5(32'hbbc53083),
	.w6(32'h3cbee2cd),
	.w7(32'hbc7eb8b2),
	.w8(32'hbc9917b6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2d18bb),
	.w1(32'h3c8bf9e0),
	.w2(32'h3c00e824),
	.w3(32'hbc86d56c),
	.w4(32'h3bbae439),
	.w5(32'h3b283b90),
	.w6(32'h3c6d84ea),
	.w7(32'h3ab2d5ae),
	.w8(32'h3c159e0a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafce5de),
	.w1(32'h3c6555f8),
	.w2(32'h3bf0c4eb),
	.w3(32'h3b999c98),
	.w4(32'h39df8f45),
	.w5(32'hbb0781a1),
	.w6(32'h3bc623bd),
	.w7(32'hbaac317e),
	.w8(32'hbb2ea57f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb0d02),
	.w1(32'hba9e8a5e),
	.w2(32'h3b39ffdb),
	.w3(32'hbb065737),
	.w4(32'hbbfba063),
	.w5(32'h3b65f1e1),
	.w6(32'h39684806),
	.w7(32'h39dab37c),
	.w8(32'hbb001297),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1fef5),
	.w1(32'h3907108c),
	.w2(32'hbb4e63b0),
	.w3(32'h3a2c6daf),
	.w4(32'h3ac56367),
	.w5(32'h38f85a23),
	.w6(32'hbc3556b4),
	.w7(32'hbc302496),
	.w8(32'hbb024dce),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc3acf),
	.w1(32'hbc8dac48),
	.w2(32'h3781b9b7),
	.w3(32'hbaed45aa),
	.w4(32'hbc1897fc),
	.w5(32'h3a715d86),
	.w6(32'hbc7453f2),
	.w7(32'hb8f11d77),
	.w8(32'h3c080372),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96e192),
	.w1(32'hbcd4039b),
	.w2(32'h3b3b303b),
	.w3(32'h3c44456c),
	.w4(32'hbc1cc0c1),
	.w5(32'h3b833d2d),
	.w6(32'hbc8bbe06),
	.w7(32'h3b905a46),
	.w8(32'h3c69a51e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d06eb36),
	.w1(32'h3c9c95ff),
	.w2(32'h3bf337a9),
	.w3(32'h3c85c79c),
	.w4(32'h3c0ef88c),
	.w5(32'h3b890158),
	.w6(32'h3c326f91),
	.w7(32'hba55ed49),
	.w8(32'hbbcb5306),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc301242),
	.w1(32'h3bb2211a),
	.w2(32'hbc3777d3),
	.w3(32'hbb827875),
	.w4(32'h3bbdf1c7),
	.w5(32'hbc1d9f32),
	.w6(32'h3b6239f8),
	.w7(32'hbb9b58b8),
	.w8(32'hbc02cd96),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6bc78),
	.w1(32'hbc723c58),
	.w2(32'h3c113555),
	.w3(32'hba9481bb),
	.w4(32'hbc376db7),
	.w5(32'h3c0b48ce),
	.w6(32'hbc6a6e90),
	.w7(32'h3c0b21a2),
	.w8(32'h3c262b03),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d06e0dd),
	.w1(32'h3b8568f6),
	.w2(32'h3b103db2),
	.w3(32'h3c834d36),
	.w4(32'h3bf24dc3),
	.w5(32'hb9c3ed05),
	.w6(32'hbb6349e2),
	.w7(32'hbb11c930),
	.w8(32'h3ab250e1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2b966),
	.w1(32'h3bb0fe6b),
	.w2(32'hb9d044fd),
	.w3(32'hba5a4008),
	.w4(32'h3a9fcf86),
	.w5(32'hbb7aec31),
	.w6(32'hba84a8f3),
	.w7(32'hbb7bb67c),
	.w8(32'hbbd5c8b6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc245518),
	.w1(32'h39d12a3f),
	.w2(32'hbb14eaa7),
	.w3(32'hbb978a6f),
	.w4(32'hb82c90e4),
	.w5(32'hbb17a7c1),
	.w6(32'h38d3f546),
	.w7(32'h3abf2190),
	.w8(32'hbafbec73),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02d71c),
	.w1(32'hba3df32c),
	.w2(32'hbb10248c),
	.w3(32'hbaca3ff3),
	.w4(32'h3ad0f319),
	.w5(32'h3b09ba39),
	.w6(32'hba92f7af),
	.w7(32'h3a0ff0d3),
	.w8(32'h3bf3b62b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0e8d5),
	.w1(32'hbc07437c),
	.w2(32'hbcd76b08),
	.w3(32'h3c029f6d),
	.w4(32'hbb13fc58),
	.w5(32'hbc6d67dd),
	.w6(32'hbc11643b),
	.w7(32'hbc583a52),
	.w8(32'hba897ae7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba959927),
	.w1(32'h3bb732c8),
	.w2(32'h385c4a5a),
	.w3(32'hbb7d0d00),
	.w4(32'hbc212715),
	.w5(32'hbbc5cf43),
	.w6(32'hbb0de79b),
	.w7(32'hbbf7cf77),
	.w8(32'hbb0710c5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc214154),
	.w1(32'hbcd3cce4),
	.w2(32'h3b9bd285),
	.w3(32'hbb329ccb),
	.w4(32'hbc41c25a),
	.w5(32'h3b662d0b),
	.w6(32'hbc97c09b),
	.w7(32'h3b92b700),
	.w8(32'h3c5e2e32),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0fc9de),
	.w1(32'hbc2e3ec6),
	.w2(32'hbb47f620),
	.w3(32'h3c81d60c),
	.w4(32'hbc956d86),
	.w5(32'hbbebe572),
	.w6(32'hbc8b37d0),
	.w7(32'hbc4972bd),
	.w8(32'hbbe4ccce),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fc41a),
	.w1(32'hbcb987d5),
	.w2(32'hba10fc45),
	.w3(32'hba7e8b9a),
	.w4(32'hbc289b46),
	.w5(32'hba8f9381),
	.w6(32'hbc21d6b9),
	.w7(32'h3b9f82eb),
	.w8(32'h3bc9fd85),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4c8bb),
	.w1(32'hbc57d374),
	.w2(32'hbc2d08b9),
	.w3(32'h3c1ae93f),
	.w4(32'hbb3be529),
	.w5(32'hbc526ca9),
	.w6(32'h3b42a109),
	.w7(32'hbc54c8d1),
	.w8(32'hbba24abb),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1965e8),
	.w1(32'h3d0ac047),
	.w2(32'hb8302e6c),
	.w3(32'hba4b62f2),
	.w4(32'h3bc48a74),
	.w5(32'hbbde8dd3),
	.w6(32'h3c7c3b65),
	.w7(32'hbc555e73),
	.w8(32'hbc691b8c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01d36d),
	.w1(32'hbb9b476e),
	.w2(32'hbb0b10ab),
	.w3(32'hbc4fac08),
	.w4(32'hbc1459a6),
	.w5(32'hbbda7d34),
	.w6(32'hbbb04b52),
	.w7(32'hbbafbeb5),
	.w8(32'hbaf64727),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffd727),
	.w1(32'hbc012ed8),
	.w2(32'hbc553d43),
	.w3(32'h3a2164ae),
	.w4(32'hbbe288c0),
	.w5(32'hbc8570d5),
	.w6(32'hbc0d2b63),
	.w7(32'hbc14b8c6),
	.w8(32'h3a847274),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fda2e),
	.w1(32'hbb21e37b),
	.w2(32'hbc009f5e),
	.w3(32'hba8d0191),
	.w4(32'hbb89ca9a),
	.w5(32'hbc033a17),
	.w6(32'h3b043599),
	.w7(32'h3c24bf2d),
	.w8(32'h3bbbcf67),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb5ffb),
	.w1(32'hba93c3ca),
	.w2(32'h3b035e2e),
	.w3(32'hbc420359),
	.w4(32'hbb0f3f2b),
	.w5(32'h3aca0f3a),
	.w6(32'hbc0dc255),
	.w7(32'hba40b039),
	.w8(32'h3b3c458b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66b341),
	.w1(32'hbc826618),
	.w2(32'h3bf46bff),
	.w3(32'h3bc1bcda),
	.w4(32'hbbb42436),
	.w5(32'h3bf23d6c),
	.w6(32'hbc2f54b4),
	.w7(32'h3be672f4),
	.w8(32'h3bc9f15c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd212d1),
	.w1(32'h3cb88fad),
	.w2(32'hba63116f),
	.w3(32'h3bde061f),
	.w4(32'h3c87e4be),
	.w5(32'hbb54de53),
	.w6(32'h3c87f9c7),
	.w7(32'hbba95f38),
	.w8(32'hbc25cf5a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc887c9f),
	.w1(32'h3c212c95),
	.w2(32'hbb127590),
	.w3(32'hbc0dcd47),
	.w4(32'hbaa7f537),
	.w5(32'hbbc965d6),
	.w6(32'h3b3c50c3),
	.w7(32'hbc050ee8),
	.w8(32'hbc390bff),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb35ac1),
	.w1(32'hbce09d6f),
	.w2(32'hb8842ae0),
	.w3(32'hbc2eefb9),
	.w4(32'hbc4e4f37),
	.w5(32'h38c9a778),
	.w6(32'hbc9393e2),
	.w7(32'hb8fc0b57),
	.w8(32'h3c14622e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd59eb5),
	.w1(32'hbcb5e9d9),
	.w2(32'h3ba4dae2),
	.w3(32'h3c2d9482),
	.w4(32'hbc269e16),
	.w5(32'h3b58cdb9),
	.w6(32'hbc7f222f),
	.w7(32'h3ba2a64b),
	.w8(32'h3c486316),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d00a10e),
	.w1(32'hbcb6465e),
	.w2(32'hb97f23a6),
	.w3(32'h3c5cbd74),
	.w4(32'hbc28e573),
	.w5(32'h3b34516d),
	.w6(32'hbcb822f9),
	.w7(32'hba1beca0),
	.w8(32'h3c2ab37c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbefe66),
	.w1(32'h3b35422d),
	.w2(32'h398ac980),
	.w3(32'h3bbda0d2),
	.w4(32'hbc0126bf),
	.w5(32'hbb471fe2),
	.w6(32'hbb72db4c),
	.w7(32'hbb9f2434),
	.w8(32'hba83074a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba02b95),
	.w1(32'hbad28007),
	.w2(32'h3b99cab1),
	.w3(32'h3b16129c),
	.w4(32'hbb814979),
	.w5(32'hbb8fb623),
	.w6(32'hbc04ee69),
	.w7(32'h3b064312),
	.w8(32'h3b54898b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12b3f5),
	.w1(32'hbce9ca8b),
	.w2(32'h3aed8030),
	.w3(32'h3b70fed7),
	.w4(32'hbc13cfb3),
	.w5(32'h3ac5aba9),
	.w6(32'hbcbfbec8),
	.w7(32'h3947e251),
	.w8(32'h3c9dd497),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d279762),
	.w1(32'hbc7b9b46),
	.w2(32'hbc5c1de7),
	.w3(32'h3c9684f9),
	.w4(32'hbcbc201e),
	.w5(32'hbc946087),
	.w6(32'hbc7b41a4),
	.w7(32'hbc881f68),
	.w8(32'hbc14a1b4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84de38),
	.w1(32'h3ab634fb),
	.w2(32'h3b8c52c4),
	.w3(32'hbbe0cdaa),
	.w4(32'h3a9e829f),
	.w5(32'h3b65f2a0),
	.w6(32'hbbe402c0),
	.w7(32'h3a660892),
	.w8(32'h3b495565),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3b397),
	.w1(32'hbd038042),
	.w2(32'hbbe26827),
	.w3(32'h3c1509b0),
	.w4(32'hbc7c1b84),
	.w5(32'hbb704cc1),
	.w6(32'hbc90db1c),
	.w7(32'h3b1e7d18),
	.w8(32'h3b884755),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64f0a5),
	.w1(32'hbaa90af4),
	.w2(32'hbadd22b1),
	.w3(32'h3a995cfd),
	.w4(32'hbb313e0b),
	.w5(32'hb683a50c),
	.w6(32'hbaca8795),
	.w7(32'h3b26ee87),
	.w8(32'h3b67e7a0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f2abf),
	.w1(32'hbb990fb8),
	.w2(32'h3b99529d),
	.w3(32'h3b8eb2f2),
	.w4(32'hbc37dd02),
	.w5(32'h3b3866fe),
	.w6(32'hbc1b6bcd),
	.w7(32'hbb8e13be),
	.w8(32'hbb125bae),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3a251),
	.w1(32'h3abc7623),
	.w2(32'hba09fe01),
	.w3(32'hb99fe41e),
	.w4(32'hbb0d4dd8),
	.w5(32'hbb37a21d),
	.w6(32'hbb245000),
	.w7(32'hbb0b6f85),
	.w8(32'hbba83a0b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9f54b),
	.w1(32'hbbb7b387),
	.w2(32'hbaac2d0b),
	.w3(32'hbb39c9e2),
	.w4(32'hbc52bb3d),
	.w5(32'hbba185bf),
	.w6(32'hbc16012a),
	.w7(32'hbba76028),
	.w8(32'hba391e1e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0127a9),
	.w1(32'hbb919eb9),
	.w2(32'h3b1caae0),
	.w3(32'hbb96648c),
	.w4(32'hb95db279),
	.w5(32'h3ba60054),
	.w6(32'hbbaa717b),
	.w7(32'h3b8d0d61),
	.w8(32'h3bad60e5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b279b91),
	.w1(32'hbb84580d),
	.w2(32'hbb187be8),
	.w3(32'h3b870f45),
	.w4(32'hbbe1014f),
	.w5(32'hbb0d77b2),
	.w6(32'hbb901344),
	.w7(32'hbad3c79f),
	.w8(32'h3a5d413c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74e94f),
	.w1(32'h3a9a9dff),
	.w2(32'hbbb65040),
	.w3(32'hbada864c),
	.w4(32'h38554781),
	.w5(32'hb98dc42f),
	.w6(32'h3a87b6c5),
	.w7(32'hbab98a96),
	.w8(32'h3c1456c1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4133fa),
	.w1(32'hbc97fe06),
	.w2(32'hbb46ddaa),
	.w3(32'h3b90ecb0),
	.w4(32'hbc190026),
	.w5(32'hba5c8162),
	.w6(32'hbc51c4b0),
	.w7(32'h3a8f6a12),
	.w8(32'h3b944915),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c521c),
	.w1(32'h3b9cc0f9),
	.w2(32'h3aabe3f5),
	.w3(32'h3a794e08),
	.w4(32'hba81f8c9),
	.w5(32'h3a9a6380),
	.w6(32'hbb27ffa4),
	.w7(32'hbb340813),
	.w8(32'hba907802),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45b0f4),
	.w1(32'hbce7b28c),
	.w2(32'hbb8e473d),
	.w3(32'h3a9ad02f),
	.w4(32'hbc5bf2b7),
	.w5(32'hb5c74516),
	.w6(32'hbcb96985),
	.w7(32'h3a797e51),
	.w8(32'h3bfdde9c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9cc747),
	.w1(32'hbc919c2d),
	.w2(32'h39ee42b5),
	.w3(32'h3bb96f06),
	.w4(32'hbc2542ca),
	.w5(32'h3a81c6b4),
	.w6(32'hbc5226bb),
	.w7(32'h3af4a4fe),
	.w8(32'h3c049fe2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb45dfe),
	.w1(32'h3c380851),
	.w2(32'h3b56c7dd),
	.w3(32'h3c042e5b),
	.w4(32'h3ab234a5),
	.w5(32'h3a82ee3e),
	.w6(32'h3bc290ac),
	.w7(32'hbb8e470f),
	.w8(32'hbbce4304),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca7f12),
	.w1(32'h3b5805d4),
	.w2(32'hbb3c6cea),
	.w3(32'hbc1202d7),
	.w4(32'hbb1b1031),
	.w5(32'hbb90c2b4),
	.w6(32'h390b8903),
	.w7(32'hbb962d34),
	.w8(32'hbc0eb4b6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc734c29),
	.w1(32'h3ab7e1eb),
	.w2(32'h3b9b7c67),
	.w3(32'hbc18ac9d),
	.w4(32'h3a1ef8b5),
	.w5(32'h3baac68b),
	.w6(32'hbb70206c),
	.w7(32'h3be7a195),
	.w8(32'h3bc0f93d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a762428),
	.w1(32'hbaa645e7),
	.w2(32'h39fde4a0),
	.w3(32'h3b6c7612),
	.w4(32'hbbea4c1c),
	.w5(32'hbb8c8c87),
	.w6(32'h3af8bef4),
	.w7(32'h3a3d9159),
	.w8(32'hbab9cf0c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4c7cd),
	.w1(32'hbbb1acca),
	.w2(32'h3bbc6cd6),
	.w3(32'hbb961bd1),
	.w4(32'hbbcd9ec5),
	.w5(32'h3a3d535b),
	.w6(32'hbb42fab9),
	.w7(32'h3be9e04c),
	.w8(32'h3b9b1647),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be56e25),
	.w1(32'hbbd9be8a),
	.w2(32'hbbc4e125),
	.w3(32'h3be92d5e),
	.w4(32'hbb8339f2),
	.w5(32'hbb8483a7),
	.w6(32'hbbb6a16b),
	.w7(32'hbba5e459),
	.w8(32'hbb8488f4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8d96d),
	.w1(32'h391d57d3),
	.w2(32'hbc308f64),
	.w3(32'h3a5ffc74),
	.w4(32'hba80fda2),
	.w5(32'hbc3baeda),
	.w6(32'hbb52ef5e),
	.w7(32'hbc389f82),
	.w8(32'hbbf23534),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd63781),
	.w1(32'hbc3d273f),
	.w2(32'hb910f980),
	.w3(32'hba572380),
	.w4(32'hbcb4bed2),
	.w5(32'hbbc49019),
	.w6(32'hbc3930c6),
	.w7(32'hbb8c700e),
	.w8(32'hbac9ffcd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f6676),
	.w1(32'h3b9fa99b),
	.w2(32'h3bfaef8b),
	.w3(32'hbc19f954),
	.w4(32'hbb9ab12d),
	.w5(32'h3bf2b1a4),
	.w6(32'hbbcd6ff3),
	.w7(32'hbbdcdb79),
	.w8(32'hbbf72bd0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5ec54),
	.w1(32'h3af24fa3),
	.w2(32'hbc396555),
	.w3(32'hbb02a0ed),
	.w4(32'h3b4a2a36),
	.w5(32'hbc49eaad),
	.w6(32'h3c0337f2),
	.w7(32'hbc1845db),
	.w8(32'hbb6c96b6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8081ae),
	.w1(32'hbc00f4c4),
	.w2(32'h3cef2e4c),
	.w3(32'h3a099ae7),
	.w4(32'hbb886106),
	.w5(32'hbc2396d3),
	.w6(32'hbbce43ab),
	.w7(32'h3b44df9c),
	.w8(32'hbc39fffc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc10e3b),
	.w1(32'hbd3ed923),
	.w2(32'h39105335),
	.w3(32'hbc8ca4eb),
	.w4(32'hbc5d0305),
	.w5(32'h3ac1d8a9),
	.w6(32'hbcdac04c),
	.w7(32'h3b93a543),
	.w8(32'h3ce8c287),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d81ffc0),
	.w1(32'hbcdc69a7),
	.w2(32'hbb7a1b0d),
	.w3(32'h3ceca3fa),
	.w4(32'hbc422175),
	.w5(32'hbac77124),
	.w6(32'hbc8e691a),
	.w7(32'h371391db),
	.w8(32'h3c000a00),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd9159f),
	.w1(32'hbcc0a8b1),
	.w2(32'hbadfc69c),
	.w3(32'h3b6192e2),
	.w4(32'hbc1f944b),
	.w5(32'h38d68ef2),
	.w6(32'hbca103ee),
	.w7(32'hbb8c3f26),
	.w8(32'h3c6268f8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d07d350),
	.w1(32'hbc7943c5),
	.w2(32'hbb4c2b88),
	.w3(32'h3c8198da),
	.w4(32'hbbd8ace9),
	.w5(32'hb92bd390),
	.w6(32'hbc3a3bfb),
	.w7(32'h3948f3b4),
	.w8(32'h3b76d079),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c483dab),
	.w1(32'hbb4f66ae),
	.w2(32'h39f34743),
	.w3(32'h3b719ada),
	.w4(32'hbc2b5960),
	.w5(32'hbbfd3747),
	.w6(32'hbb555b84),
	.w7(32'hba9dd6e4),
	.w8(32'hba97401a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc180335),
	.w1(32'hbca8762a),
	.w2(32'h3b424123),
	.w3(32'hbc10934c),
	.w4(32'hbc2cbd72),
	.w5(32'h3b5b1eef),
	.w6(32'hbc8a279a),
	.w7(32'h3b91a705),
	.w8(32'h3c07e2d8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd1752a),
	.w1(32'hbcbac8e6),
	.w2(32'h3ac2e08f),
	.w3(32'h3c31a945),
	.w4(32'hbbda40eb),
	.w5(32'h3a729acf),
	.w6(32'hbc8c10f9),
	.w7(32'h3adadc80),
	.w8(32'h3c702241),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0a08ef),
	.w1(32'h3bd81ed1),
	.w2(32'h3c21a3b7),
	.w3(32'h3c74fadb),
	.w4(32'hbb08a14e),
	.w5(32'h3bc347c2),
	.w6(32'h3b57c07d),
	.w7(32'hb9eec37f),
	.w8(32'h3b958205),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d19ee),
	.w1(32'hbc6398b0),
	.w2(32'h3c0b6361),
	.w3(32'h3beb299e),
	.w4(32'hbbc8421e),
	.w5(32'h3bcb3ea6),
	.w6(32'hbc292aeb),
	.w7(32'h3c1e7ad8),
	.w8(32'h3c23ddf6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce8079b),
	.w1(32'hbbb5fc70),
	.w2(32'h3b928d68),
	.w3(32'h3c40429c),
	.w4(32'hbb3ef537),
	.w5(32'hbad36740),
	.w6(32'h3c087fb4),
	.w7(32'h3b4160b1),
	.w8(32'h3aef0ab3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08ff33),
	.w1(32'hbc6dbec2),
	.w2(32'h3b9b4451),
	.w3(32'h3ad2ae67),
	.w4(32'hbbfdb094),
	.w5(32'h3b8d1381),
	.w6(32'hbc88b29e),
	.w7(32'hb9dda7dd),
	.w8(32'h3bc831dc),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf30ce),
	.w1(32'h3c1384d4),
	.w2(32'h3b06a437),
	.w3(32'h3be066a9),
	.w4(32'h39fc568c),
	.w5(32'h3aabf6cc),
	.w6(32'h3b1d0971),
	.w7(32'hbb66f0af),
	.w8(32'hbba594ac),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffb198),
	.w1(32'hbcad96c0),
	.w2(32'hbaa52911),
	.w3(32'hba94721f),
	.w4(32'hbc1dea34),
	.w5(32'h3b000e5f),
	.w6(32'hbc57fbd5),
	.w7(32'h3b5860d6),
	.w8(32'h3c10b57a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc41bcc),
	.w1(32'hbd0672a7),
	.w2(32'hba96e5f4),
	.w3(32'h3c3a91a5),
	.w4(32'hbc30a2f8),
	.w5(32'hbad83558),
	.w6(32'hbca7e6cf),
	.w7(32'h3b38f7cc),
	.w8(32'h3c9ff925),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d410444),
	.w1(32'hbcd0a61f),
	.w2(32'h39d21389),
	.w3(32'h3caff87e),
	.w4(32'hbc2a331f),
	.w5(32'h3a183f5f),
	.w6(32'hbc83b9d4),
	.w7(32'h3b41d100),
	.w8(32'h3c5c1ad8),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf9e01a),
	.w1(32'hbccdaba6),
	.w2(32'h3a9b6e9e),
	.w3(32'h3c74b084),
	.w4(32'hbc26a540),
	.w5(32'h39a3d83d),
	.w6(32'hbc85744d),
	.w7(32'h3b04ae75),
	.w8(32'h3c5e097f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d07c0da),
	.w1(32'hbbc44584),
	.w2(32'hbb41e9a0),
	.w3(32'h3c6fd0fe),
	.w4(32'hbc439fbd),
	.w5(32'hbc3927dc),
	.w6(32'hbbd95521),
	.w7(32'hbb456e53),
	.w8(32'hb98523c2),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b600880),
	.w1(32'h3b155cda),
	.w2(32'hbb8b3d80),
	.w3(32'h3bdc31a5),
	.w4(32'hbbb994db),
	.w5(32'hbbb494bc),
	.w6(32'hbbb8a0af),
	.w7(32'hbbe2a440),
	.w8(32'h3aa6d4be),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03586d),
	.w1(32'hbcb5a71a),
	.w2(32'hba96d75c),
	.w3(32'h3be08efa),
	.w4(32'hbc4b0cda),
	.w5(32'h3a5d06d5),
	.w6(32'hbc9f9d89),
	.w7(32'hbbac6392),
	.w8(32'h3c07653f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc7c014),
	.w1(32'hbc8b5a56),
	.w2(32'h3c06a586),
	.w3(32'h3c4866c6),
	.w4(32'hbc2b678b),
	.w5(32'h3bb1b2b1),
	.w6(32'hbc606b0b),
	.w7(32'h3a34f2ba),
	.w8(32'h3b8e01c3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8574f2),
	.w1(32'hbcf32a03),
	.w2(32'h3b0223ad),
	.w3(32'h3c05dbfb),
	.w4(32'hbc644a7b),
	.w5(32'h3b452ab1),
	.w6(32'hbc9f96fd),
	.w7(32'h3b85f4ca),
	.w8(32'h3c772b44),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d13c0ff),
	.w1(32'h3bccc34f),
	.w2(32'h3c04e0db),
	.w3(32'h3c8af80e),
	.w4(32'hbb4cd1ff),
	.w5(32'hbc285a13),
	.w6(32'hbb87dae2),
	.w7(32'h3b6072aa),
	.w8(32'hbb30cfac),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd73af),
	.w1(32'hbc561732),
	.w2(32'h3c01f7a1),
	.w3(32'hbb0aaed7),
	.w4(32'hbc1d619d),
	.w5(32'h3b652dfd),
	.w6(32'hbc44e30f),
	.w7(32'h3be85079),
	.w8(32'h3c1bcec6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce30059),
	.w1(32'hbccfe05a),
	.w2(32'hba0f6c5c),
	.w3(32'h3c582799),
	.w4(32'hbc677aa6),
	.w5(32'hbaac3f56),
	.w6(32'hbca6073c),
	.w7(32'hbb03bf91),
	.w8(32'h3bbd9a6f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab240b),
	.w1(32'hb91cbaab),
	.w2(32'hb80b82b0),
	.w3(32'h3b67900b),
	.w4(32'hba02623a),
	.w5(32'hb9b8f9a0),
	.w6(32'hb9946a00),
	.w7(32'hb9d30c7a),
	.w8(32'hb94a4fd9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b438ebc),
	.w1(32'h3b42dcae),
	.w2(32'h3b88884d),
	.w3(32'hbb5ae798),
	.w4(32'hbabd69c9),
	.w5(32'h3b52a19c),
	.w6(32'hbbcaa6c3),
	.w7(32'hbba2ce04),
	.w8(32'hba6c09aa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b046c58),
	.w1(32'h3b067001),
	.w2(32'h3b211a4c),
	.w3(32'h39ef6b5c),
	.w4(32'h3add3be3),
	.w5(32'h3b2a96f0),
	.w6(32'hbb096408),
	.w7(32'h3a7b56b2),
	.w8(32'h3b1327cf),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9235dd2),
	.w1(32'hb982f23f),
	.w2(32'h39ae4237),
	.w3(32'h39416993),
	.w4(32'h38e30a2d),
	.w5(32'h39998662),
	.w6(32'hb6f91764),
	.w7(32'h398dec4f),
	.w8(32'h39b3e4e1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e58a6e),
	.w1(32'hb9710da2),
	.w2(32'h39ed47d6),
	.w3(32'hb959dceb),
	.w4(32'hb9c86101),
	.w5(32'h393d3cda),
	.w6(32'hb9f3ebf3),
	.w7(32'hba7fa1c4),
	.w8(32'h380c27eb),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7861a02),
	.w1(32'hb9890872),
	.w2(32'hb99ec389),
	.w3(32'h394e5dcd),
	.w4(32'hb9b9fcb5),
	.w5(32'hb9a2e18e),
	.w6(32'h3a3bcfb9),
	.w7(32'h392a2228),
	.w8(32'h3946aa05),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918e10b),
	.w1(32'h3988ff34),
	.w2(32'h3a21ac82),
	.w3(32'h399d8dc7),
	.w4(32'h39665589),
	.w5(32'h39e25665),
	.w6(32'hb80f98d1),
	.w7(32'hb74e6d48),
	.w8(32'h396d0842),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e749e),
	.w1(32'hb9e926da),
	.w2(32'h389700d8),
	.w3(32'h390e38e4),
	.w4(32'hba890895),
	.w5(32'hba89b5ff),
	.w6(32'h3b0b2af0),
	.w7(32'h3a5e24f4),
	.w8(32'h398746a8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2eddff),
	.w1(32'h3a238238),
	.w2(32'h3b0f1f95),
	.w3(32'h39830a6f),
	.w4(32'h3af2061c),
	.w5(32'h3b33b667),
	.w6(32'hbb381fd4),
	.w7(32'h3a38f68d),
	.w8(32'h3aec7ff5),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90cc32b),
	.w1(32'hb9380592),
	.w2(32'hb921228c),
	.w3(32'hb93a668b),
	.w4(32'hb9d66160),
	.w5(32'h3a0876c6),
	.w6(32'h3a942f92),
	.w7(32'h3a540dde),
	.w8(32'h3a5f46bf),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82ead0),
	.w1(32'hb90284e0),
	.w2(32'h3ab163f1),
	.w3(32'hba8c41d6),
	.w4(32'hba0fd654),
	.w5(32'h3a39e4bd),
	.w6(32'hb9a5e1f5),
	.w7(32'hba1212b7),
	.w8(32'h3a4823ea),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a445ac7),
	.w1(32'h3a868ac3),
	.w2(32'h3ae61aa7),
	.w3(32'h3a3ccf84),
	.w4(32'h39fc6a41),
	.w5(32'h3abe860e),
	.w6(32'hbacb1ebb),
	.w7(32'hbaa2c1be),
	.w8(32'h3a54b68e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946ee45),
	.w1(32'h391fe0d0),
	.w2(32'h38b91a9a),
	.w3(32'hbb18913a),
	.w4(32'hbaf397f9),
	.w5(32'hb99931a8),
	.w6(32'hbb05f172),
	.w7(32'hbb0809fb),
	.w8(32'hba171f75),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e47fe),
	.w1(32'h39a29ebd),
	.w2(32'h3af77ad2),
	.w3(32'h3a13df68),
	.w4(32'h3a532ef8),
	.w5(32'h3b21569a),
	.w6(32'hb955363f),
	.w7(32'h3ac863f0),
	.w8(32'h3b5beb05),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b0c21),
	.w1(32'h394388e3),
	.w2(32'h39cc904e),
	.w3(32'h383f28ae),
	.w4(32'h388219ab),
	.w5(32'h39cd0ed2),
	.w6(32'hb86faccf),
	.w7(32'hb79c22e1),
	.w8(32'h39ae889e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6e29d),
	.w1(32'hba14c287),
	.w2(32'h39cbbccc),
	.w3(32'h3adcb276),
	.w4(32'h39d23bd5),
	.w5(32'h3b1fedf8),
	.w6(32'h3bb033eb),
	.w7(32'h3b753458),
	.w8(32'h3b9e5c1f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d76190),
	.w1(32'h3ab4a88c),
	.w2(32'h3aafafce),
	.w3(32'h395a0d1a),
	.w4(32'h3a6e716e),
	.w5(32'h3ad34579),
	.w6(32'hb8cd9223),
	.w7(32'h3a6f5897),
	.w8(32'h3aa44d4f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90417f0),
	.w1(32'h38079fe0),
	.w2(32'h38a9e469),
	.w3(32'hb7e42968),
	.w4(32'h38ee94b6),
	.w5(32'h38ee1102),
	.w6(32'hb9161175),
	.w7(32'hb779c45b),
	.w8(32'hb66b9376),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80773e5),
	.w1(32'hb83fc670),
	.w2(32'h37b3ab8e),
	.w3(32'hb89b0dd0),
	.w4(32'hb8ee5da2),
	.w5(32'hb8dc156e),
	.w6(32'h386291b5),
	.w7(32'hb884700e),
	.w8(32'hb7ba2a7c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e93455),
	.w1(32'hb989415e),
	.w2(32'hba2dc86a),
	.w3(32'hb9b20db4),
	.w4(32'hb8a2a5ae),
	.w5(32'h393a755e),
	.w6(32'hb9a948a6),
	.w7(32'h3a5049ae),
	.w8(32'hb9329779),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49f5cc),
	.w1(32'h3a103473),
	.w2(32'hb953bacf),
	.w3(32'hba2b7e77),
	.w4(32'hb909f7b2),
	.w5(32'h3a69e40e),
	.w6(32'h3ac690c8),
	.w7(32'h3abab35b),
	.w8(32'h3ac7603f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f9bd1),
	.w1(32'h3a8c3067),
	.w2(32'h39fa572a),
	.w3(32'h3a709fd1),
	.w4(32'h3a62d4e9),
	.w5(32'h3a315968),
	.w6(32'hbab6a24e),
	.w7(32'hb9fa8d21),
	.w8(32'hb9c3ca76),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb767116b),
	.w1(32'h35e6380e),
	.w2(32'h3752ff63),
	.w3(32'h37531540),
	.w4(32'h371c3d57),
	.w5(32'hb6ea6b44),
	.w6(32'h38345118),
	.w7(32'h37b74e3f),
	.w8(32'hb62b4a79),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3bd4b),
	.w1(32'h3ad3f166),
	.w2(32'h3b3d536a),
	.w3(32'h3ae1f152),
	.w4(32'h3b1022f9),
	.w5(32'h3b375c39),
	.w6(32'hb9f9555d),
	.w7(32'h3b12e4c3),
	.w8(32'h3b3fa062),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391caa42),
	.w1(32'h3a4af458),
	.w2(32'h3ad5fb65),
	.w3(32'hb9c157ac),
	.w4(32'h39b041c6),
	.w5(32'h3ab600ea),
	.w6(32'hb8ffc31c),
	.w7(32'h39107a60),
	.w8(32'h3a8b2229),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77d514),
	.w1(32'hbac03fe6),
	.w2(32'h3ab01a59),
	.w3(32'h3a2963d0),
	.w4(32'hb960d9ad),
	.w5(32'h3a9e8221),
	.w6(32'hbab93cd0),
	.w7(32'hba202971),
	.w8(32'h3957d463),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6cc81),
	.w1(32'hba0ef879),
	.w2(32'h3b7cfb0f),
	.w3(32'h3bb56ddb),
	.w4(32'hbac8688a),
	.w5(32'h3ab4d732),
	.w6(32'h3bc2e8c9),
	.w7(32'h3b27b769),
	.w8(32'h3a22b627),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a396b8a),
	.w1(32'h3a292faa),
	.w2(32'hb962e273),
	.w3(32'h3a341ef9),
	.w4(32'h3a1e8850),
	.w5(32'h399bc9ed),
	.w6(32'h3a975ddb),
	.w7(32'h3a872e60),
	.w8(32'h3a39c3f8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e8f5a),
	.w1(32'hb966db51),
	.w2(32'hb8b1b915),
	.w3(32'hb9c1afc3),
	.w4(32'hb98b6d18),
	.w5(32'hb9295a35),
	.w6(32'hb9687bff),
	.w7(32'hb90ed330),
	.w8(32'h3890345f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df4803),
	.w1(32'h39abe637),
	.w2(32'h3a487d51),
	.w3(32'h39e6359c),
	.w4(32'hb7a643e6),
	.w5(32'h3995631e),
	.w6(32'h3a8d228b),
	.w7(32'h395532ee),
	.w8(32'h39e39ede),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb85d0),
	.w1(32'h3a835e57),
	.w2(32'h3962322a),
	.w3(32'h3ad4fbb4),
	.w4(32'h3a916a35),
	.w5(32'h3a263897),
	.w6(32'h3b5933b4),
	.w7(32'h3b245410),
	.w8(32'h3ae5f244),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac6ac6),
	.w1(32'hba917432),
	.w2(32'hba631eae),
	.w3(32'hba756a96),
	.w4(32'hba9a17d7),
	.w5(32'hba59e66d),
	.w6(32'h39d16712),
	.w7(32'hb770b169),
	.w8(32'hb92abd44),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89acf5f),
	.w1(32'hb8573ad1),
	.w2(32'h39a990d7),
	.w3(32'h3912bfc3),
	.w4(32'h39a62657),
	.w5(32'h39b9e5ae),
	.w6(32'hb9d9fb29),
	.w7(32'hb73783df),
	.w8(32'h395e7c35),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915e503),
	.w1(32'hb932f4ac),
	.w2(32'hb9a9e4be),
	.w3(32'hb868327a),
	.w4(32'hb8cee21a),
	.w5(32'hb97f97b7),
	.w6(32'h38bbe123),
	.w7(32'hb70b50ac),
	.w8(32'hb9580e2f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfc05c),
	.w1(32'h3adbe615),
	.w2(32'h3b277120),
	.w3(32'h3811224e),
	.w4(32'h3a2bd65d),
	.w5(32'h3b0d7ede),
	.w6(32'hbaf4c0a4),
	.w7(32'hba33b23e),
	.w8(32'h3aade61b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39764818),
	.w1(32'h3a0f2b66),
	.w2(32'h390eda35),
	.w3(32'h37f87256),
	.w4(32'hb9a9ba25),
	.w5(32'hb86c4d9c),
	.w6(32'hb92ef591),
	.w7(32'h39ab95a3),
	.w8(32'h37f53aaa),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69184f),
	.w1(32'h391b2264),
	.w2(32'h3a570745),
	.w3(32'h3aa26d50),
	.w4(32'h394098ea),
	.w5(32'hb959751f),
	.w6(32'h3ad7ce62),
	.w7(32'hba9dceee),
	.w8(32'hba81b881),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eab8c7),
	.w1(32'hb9147916),
	.w2(32'hb9894324),
	.w3(32'hb77fbaff),
	.w4(32'hb8b4d31a),
	.w5(32'hb94dba91),
	.w6(32'h38cbff6d),
	.w7(32'hb8323ef1),
	.w8(32'hb8bff36c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e15427),
	.w1(32'h39499007),
	.w2(32'hb8eb7464),
	.w3(32'hbaf4a328),
	.w4(32'h3920af82),
	.w5(32'h3a08399e),
	.w6(32'hbb58831a),
	.w7(32'hbb0373d3),
	.w8(32'hb8b34d67),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c257c0),
	.w1(32'h39002d6e),
	.w2(32'h38eb7c8b),
	.w3(32'h38ef1ad8),
	.w4(32'h38e3b1f7),
	.w5(32'h3884090b),
	.w6(32'h3822d459),
	.w7(32'h383c43d3),
	.w8(32'h38918bd8),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a8bb8),
	.w1(32'h38829a1d),
	.w2(32'hb8f4f06e),
	.w3(32'h39229447),
	.w4(32'h38af61f9),
	.w5(32'hb8f5f6ad),
	.w6(32'h39b1f119),
	.w7(32'h398b9bb8),
	.w8(32'h389f6e7d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39487e22),
	.w1(32'h3a1cbc4f),
	.w2(32'h3a91017b),
	.w3(32'hb97c9db0),
	.w4(32'h388e5b1c),
	.w5(32'h3a703581),
	.w6(32'h3aaf0341),
	.w7(32'h3ab62b04),
	.w8(32'h3aa92a3d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b835f10),
	.w1(32'h3aead375),
	.w2(32'h3b8a0f74),
	.w3(32'hba36bb8e),
	.w4(32'h3b098225),
	.w5(32'h3b9d0394),
	.w6(32'hbb67c3b3),
	.w7(32'hbb0899c0),
	.w8(32'h3b2b5e3a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a8e42),
	.w1(32'hba1fd673),
	.w2(32'hba159edf),
	.w3(32'hba1e196a),
	.w4(32'hba3128d0),
	.w5(32'hba2f422b),
	.w6(32'hba0f1c6e),
	.w7(32'hba311933),
	.w8(32'hb9f80a6e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a9a38),
	.w1(32'hb91a18bf),
	.w2(32'h3940d57b),
	.w3(32'hb9de005d),
	.w4(32'hba5a8d20),
	.w5(32'h3a22d2b0),
	.w6(32'h3a059442),
	.w7(32'hb8daec36),
	.w8(32'h3a89dd4d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fe978),
	.w1(32'hba1a8cbf),
	.w2(32'hb8814821),
	.w3(32'h3a0512a2),
	.w4(32'hba4e2456),
	.w5(32'h39a2167f),
	.w6(32'h3b04cec8),
	.w7(32'h3b10232f),
	.w8(32'h3a809c00),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4350b),
	.w1(32'h3b2452ef),
	.w2(32'h3b27b800),
	.w3(32'h3a55ad58),
	.w4(32'h3b613e35),
	.w5(32'h3b254300),
	.w6(32'h3b2f9484),
	.w7(32'h3b57e556),
	.w8(32'hbaddaed9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33baad),
	.w1(32'h399cb15e),
	.w2(32'h3a91fee0),
	.w3(32'h3a62cef9),
	.w4(32'h3a44d1eb),
	.w5(32'h3a84c793),
	.w6(32'h38d92ffd),
	.w7(32'h3aca687e),
	.w8(32'h3aa59553),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9e455),
	.w1(32'h3ae45d41),
	.w2(32'h3b344f52),
	.w3(32'h3a58f920),
	.w4(32'h3aad3e7d),
	.w5(32'h3b1edeed),
	.w6(32'hbb061863),
	.w7(32'hba31a114),
	.w8(32'h3add5781),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385a3422),
	.w1(32'h373452a2),
	.w2(32'h3982e35b),
	.w3(32'hb8f50e34),
	.w4(32'hb8ea5b24),
	.w5(32'h386d8ff8),
	.w6(32'h3886be72),
	.w7(32'h38ead81b),
	.w8(32'h39403df7),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38122b2f),
	.w1(32'h39c93fa0),
	.w2(32'h39c9ae86),
	.w3(32'h3a94b277),
	.w4(32'h3a4ed2f0),
	.w5(32'h396d5ca5),
	.w6(32'h3b0497fc),
	.w7(32'h3b4f4d8b),
	.w8(32'h3ae02828),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bd630b),
	.w1(32'hb7844e76),
	.w2(32'hb8219ad4),
	.w3(32'hb78b6943),
	.w4(32'hb716b9f1),
	.w5(32'hb7f38e71),
	.w6(32'hb7aaee9c),
	.w7(32'hb747f99e),
	.w8(32'hb8386685),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992d23d),
	.w1(32'h39277453),
	.w2(32'h383ce9cf),
	.w3(32'h395590f5),
	.w4(32'hb595d120),
	.w5(32'hb8c000b1),
	.w6(32'h391894a1),
	.w7(32'hb79d0784),
	.w8(32'h38aec7e3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a92939),
	.w1(32'hb99453d2),
	.w2(32'hb9c83e54),
	.w3(32'hb90e4ef2),
	.w4(32'hb9afb546),
	.w5(32'hb95f7dd2),
	.w6(32'h396eabc4),
	.w7(32'hb7ba795f),
	.w8(32'hb912b0a9),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb004b9b),
	.w1(32'hb9acd832),
	.w2(32'h3a9aac0a),
	.w3(32'h38bb2172),
	.w4(32'h39813d0c),
	.w5(32'h3936452d),
	.w6(32'h39991c4c),
	.w7(32'h3b0454a4),
	.w8(32'h39ed80c4),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a58154),
	.w1(32'hb795f863),
	.w2(32'hb7c28093),
	.w3(32'hb6a0c27c),
	.w4(32'hb79bd434),
	.w5(32'hb7c7c11d),
	.w6(32'h3630197a),
	.w7(32'hb7500896),
	.w8(32'hb7ed664a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3854cadc),
	.w1(32'h38c68c1d),
	.w2(32'h38e64ed6),
	.w3(32'h383357ca),
	.w4(32'h389cc61c),
	.w5(32'h38e0639e),
	.w6(32'h388cbe0b),
	.w7(32'h38576942),
	.w8(32'h38edf098),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad84b2),
	.w1(32'hb92d81df),
	.w2(32'hb9de6579),
	.w3(32'h392be04d),
	.w4(32'hb9f63e21),
	.w5(32'hba81214b),
	.w6(32'hba089f23),
	.w7(32'hb9d55b71),
	.w8(32'hbaa37377),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3941e2ed),
	.w1(32'hbaeb534f),
	.w2(32'hba758799),
	.w3(32'h39d405cd),
	.w4(32'hb92f9d2f),
	.w5(32'hba94ee5b),
	.w6(32'h3b24e1b7),
	.w7(32'h3a8f6859),
	.w8(32'hbb0e5936),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c92748),
	.w1(32'hbb148815),
	.w2(32'hba7aff83),
	.w3(32'hbb055929),
	.w4(32'hbb0585ca),
	.w5(32'h3a76a855),
	.w6(32'hbb46e504),
	.w7(32'hbb6a14a8),
	.w8(32'h3a5c511a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943736b),
	.w1(32'hb9917c6d),
	.w2(32'hb88833ba),
	.w3(32'hb919d7b7),
	.w4(32'hb91d469b),
	.w5(32'hb8b9378e),
	.w6(32'hb8f85de7),
	.w7(32'hb8f73c63),
	.w8(32'hb8193870),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aceb933),
	.w1(32'h3b8ca282),
	.w2(32'h3b8ec30b),
	.w3(32'h3a4f735c),
	.w4(32'h3b76f0cb),
	.w5(32'h3bafaf25),
	.w6(32'hbb774ab5),
	.w7(32'h3a74b1bf),
	.w8(32'h3b55f799),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0bce4),
	.w1(32'hba431d42),
	.w2(32'h3b50db44),
	.w3(32'h3ad00fb2),
	.w4(32'hbb3fa6c2),
	.w5(32'h39c4b192),
	.w6(32'h3bfdb8b3),
	.w7(32'h3bd63b06),
	.w8(32'h3b5b0224),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9a5ae),
	.w1(32'hba5d62c8),
	.w2(32'h36f0c4b4),
	.w3(32'hb918ab85),
	.w4(32'hb99b6e4d),
	.w5(32'hb9a2eed1),
	.w6(32'hbaa2c70a),
	.w7(32'hba061a2c),
	.w8(32'h3a919105),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cb6c36),
	.w1(32'hb6ca0135),
	.w2(32'hb8274a50),
	.w3(32'hb7be2de0),
	.w4(32'hb6893a6c),
	.w5(32'hb878d896),
	.w6(32'hb6d25da0),
	.w7(32'hb7843de7),
	.w8(32'hb7aed1ec),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3861d0b7),
	.w1(32'h38e590b7),
	.w2(32'h390951bc),
	.w3(32'h3892e5a8),
	.w4(32'h38c10fcc),
	.w5(32'h391f0532),
	.w6(32'h3879caa2),
	.w7(32'h38ff0f43),
	.w8(32'h3943daa4),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c46809),
	.w1(32'hb723a08d),
	.w2(32'hb7a3a589),
	.w3(32'h35765a01),
	.w4(32'hb633cc64),
	.w5(32'hb780ceca),
	.w6(32'hb7067baa),
	.w7(32'hb7620526),
	.w8(32'hb7c1b2e4),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6fd22),
	.w1(32'h3a3d7964),
	.w2(32'h3aa092d2),
	.w3(32'h39cf2428),
	.w4(32'h3a37db45),
	.w5(32'h3b15e96a),
	.w6(32'hbad34915),
	.w7(32'hbaa3d1a8),
	.w8(32'h3ac16126),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaaa914),
	.w1(32'h3a9597f4),
	.w2(32'h3a7b0fdd),
	.w3(32'h39b21639),
	.w4(32'h3a18cb04),
	.w5(32'h39e52d04),
	.w6(32'hb9a23427),
	.w7(32'hba03571f),
	.w8(32'h398ee908),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a8488),
	.w1(32'hb9cb40ea),
	.w2(32'hbab1386d),
	.w3(32'hb92cfb71),
	.w4(32'hbae7227d),
	.w5(32'hba8c5ab8),
	.w6(32'h3a8aa462),
	.w7(32'h38dd427d),
	.w8(32'hb9193fa7),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bda80f),
	.w1(32'h3a2243db),
	.w2(32'h39cd9374),
	.w3(32'h38af756c),
	.w4(32'h38ffa53f),
	.w5(32'hb814d14b),
	.w6(32'hb848cf2f),
	.w7(32'hb99648dd),
	.w8(32'hb99b6927),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c1f1d),
	.w1(32'h3a6c98c7),
	.w2(32'h3af1a064),
	.w3(32'hb9ab09c1),
	.w4(32'h3a38dc05),
	.w5(32'h3b0eabc5),
	.w6(32'hbb159fe4),
	.w7(32'hba837f7d),
	.w8(32'h3a1d0a21),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e23a6),
	.w1(32'hb9836f80),
	.w2(32'hba990093),
	.w3(32'h39e1c6e3),
	.w4(32'hba0d78f6),
	.w5(32'hba642e8f),
	.w6(32'h391135f7),
	.w7(32'hb98fe744),
	.w8(32'hba90b77b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d0fa33),
	.w1(32'hb7b8469a),
	.w2(32'hb8271754),
	.w3(32'hb725e9d9),
	.w4(32'hb7959126),
	.w5(32'hb81e8a02),
	.w6(32'hb79ef6b1),
	.w7(32'hb7d98eba),
	.w8(32'hb84d8449),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2b461),
	.w1(32'h3a058092),
	.w2(32'h3aa6a360),
	.w3(32'hba154294),
	.w4(32'h3a437dd5),
	.w5(32'h3b260f19),
	.w6(32'hb90615fb),
	.w7(32'h382cf5ab),
	.w8(32'h3a8522a5),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb849a5e9),
	.w1(32'hb7e7e41e),
	.w2(32'hb87e3a42),
	.w3(32'hb7bee6e0),
	.w4(32'h36e939c2),
	.w5(32'hb8334629),
	.w6(32'hb7adaa92),
	.w7(32'hb7555bb0),
	.w8(32'hb88f06ef),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73291e),
	.w1(32'h3a9b8356),
	.w2(32'h3a8ff8a4),
	.w3(32'h3971d4ff),
	.w4(32'h3a2b39f6),
	.w5(32'h3a79b7ed),
	.w6(32'hba07560d),
	.w7(32'hb8e69e01),
	.w8(32'h392ea788),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c1473),
	.w1(32'h3a306be4),
	.w2(32'h3a8afa94),
	.w3(32'h3a66a5bf),
	.w4(32'hba2542ef),
	.w5(32'hb8dcfffd),
	.w6(32'h3aeec15c),
	.w7(32'h3a34b1b5),
	.w8(32'h3a20d011),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b0577),
	.w1(32'h37fc4c04),
	.w2(32'h3a781970),
	.w3(32'h3960490a),
	.w4(32'hb9457506),
	.w5(32'h3a3f49b8),
	.w6(32'h3a8f31f2),
	.w7(32'h39bf8db8),
	.w8(32'h3a49e37f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9065ad6),
	.w1(32'hb965d14d),
	.w2(32'hb9980e60),
	.w3(32'hb9451230),
	.w4(32'hb95d8c5d),
	.w5(32'hb9b87428),
	.w6(32'hb84b730e),
	.w7(32'hb77b32bf),
	.w8(32'hb8fac2de),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43ba48),
	.w1(32'hba17d32f),
	.w2(32'h39822689),
	.w3(32'h3993f87b),
	.w4(32'hbac2d107),
	.w5(32'hbaa2be99),
	.w6(32'h3b17cc48),
	.w7(32'h39cd5cec),
	.w8(32'hb96f8557),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e60823),
	.w1(32'h3a1f3999),
	.w2(32'h3af0dbb8),
	.w3(32'h37b0ac4a),
	.w4(32'h3a4f7001),
	.w5(32'h3afcb95e),
	.w6(32'hb9a76963),
	.w7(32'h399e9406),
	.w8(32'h3b16088f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a011e47),
	.w1(32'h3a9362c3),
	.w2(32'h3aa73d6c),
	.w3(32'hb9063d40),
	.w4(32'h3a4a0d53),
	.w5(32'h3ab655ac),
	.w6(32'hbad64c6e),
	.w7(32'hb6cca898),
	.w8(32'h3a005c73),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8673ddd),
	.w1(32'hb7be2600),
	.w2(32'h36c85f3c),
	.w3(32'hb7e6377e),
	.w4(32'hb68ae4b4),
	.w5(32'h366db7ec),
	.w6(32'h3675d78c),
	.w7(32'h37a37754),
	.w8(32'h3808258c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc7787),
	.w1(32'hb86950b7),
	.w2(32'h374c00dd),
	.w3(32'hb16d114c),
	.w4(32'hb8ac38d0),
	.w5(32'hb811fd90),
	.w6(32'h378f399e),
	.w7(32'h38d47c23),
	.w8(32'h38a0d150),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb30aa),
	.w1(32'h3a16a1d8),
	.w2(32'h3aec1f33),
	.w3(32'hbb2ad1b9),
	.w4(32'hbaceb835),
	.w5(32'h3931b063),
	.w6(32'hbb71e7a7),
	.w7(32'hbb603e25),
	.w8(32'hba37837f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d5a35),
	.w1(32'h3b0e9c84),
	.w2(32'h3b8788ee),
	.w3(32'h391a6739),
	.w4(32'h3af2bdfa),
	.w5(32'h3b7870cd),
	.w6(32'hba630aaf),
	.w7(32'h393a88f8),
	.w8(32'h3b0c3319),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0aff91),
	.w1(32'h393779fc),
	.w2(32'h3a26bbc1),
	.w3(32'h39f7fd8a),
	.w4(32'hba831464),
	.w5(32'hb865d804),
	.w6(32'h39c87eba),
	.w7(32'hba03a451),
	.w8(32'hb9a77d4e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb087398),
	.w1(32'hbb11e2ef),
	.w2(32'hba3c3536),
	.w3(32'h3aa53e49),
	.w4(32'hbb0ce6c6),
	.w5(32'hb94df271),
	.w6(32'h3b23d7b2),
	.w7(32'h3bbcc683),
	.w8(32'h3b72cab6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0aba10),
	.w1(32'h39a4527f),
	.w2(32'h39d28fd5),
	.w3(32'hb9c2ab8f),
	.w4(32'h3a1aaeba),
	.w5(32'h398b48d0),
	.w6(32'hba0c1cde),
	.w7(32'h397adddd),
	.w8(32'h3813f07f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9231ac0),
	.w1(32'h3a016db5),
	.w2(32'h3a64ee78),
	.w3(32'hb96df12b),
	.w4(32'h39a25bb3),
	.w5(32'h3a85da6b),
	.w6(32'hb9e329a6),
	.w7(32'h38cb9272),
	.w8(32'h3a4c771a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad59c0),
	.w1(32'h3b28c521),
	.w2(32'h3b21b8fa),
	.w3(32'hb8ba5cb3),
	.w4(32'h385aaf09),
	.w5(32'h3be3076e),
	.w6(32'hbb8caa2d),
	.w7(32'hbbcfc0b6),
	.w8(32'h3b16f869),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b219a80),
	.w1(32'h3b1cf246),
	.w2(32'h3b022121),
	.w3(32'h3a1e478a),
	.w4(32'h3ae25df7),
	.w5(32'h3b2d883e),
	.w6(32'hbb65d655),
	.w7(32'hbaba377f),
	.w8(32'hb88d0477),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17e556),
	.w1(32'hbab8f299),
	.w2(32'h39dc17da),
	.w3(32'hba8de864),
	.w4(32'hba1afe9a),
	.w5(32'h3aa276d9),
	.w6(32'hbb774a25),
	.w7(32'hbb622fc2),
	.w8(32'hba8f3e90),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38af278c),
	.w1(32'hb9fcab03),
	.w2(32'hb9a526b7),
	.w3(32'h3a1c36ce),
	.w4(32'hb99f6b7a),
	.w5(32'h390434ef),
	.w6(32'h3abaff12),
	.w7(32'h39c90626),
	.w8(32'hb929a922),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c1bc3),
	.w1(32'h39776d36),
	.w2(32'h3a0193c4),
	.w3(32'h3a58ab01),
	.w4(32'hba81c8f6),
	.w5(32'hba00d79e),
	.w6(32'h3b5fbbbb),
	.w7(32'h3ae3e608),
	.w8(32'h3a4ad708),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e52ae1),
	.w1(32'hb793b98d),
	.w2(32'hb80133ac),
	.w3(32'hb7aa097b),
	.w4(32'hb772868f),
	.w5(32'hb7e0e124),
	.w6(32'hb757369d),
	.w7(32'hb78101d2),
	.w8(32'hb8006020),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a66905),
	.w1(32'hb68730c9),
	.w2(32'hb77c2e9a),
	.w3(32'hb75fa41b),
	.w4(32'hb6bae4f5),
	.w5(32'hb79d1671),
	.w6(32'hb766e831),
	.w7(32'hb765b3bf),
	.w8(32'hb7c1aa6e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ea23d),
	.w1(32'h3995cfd9),
	.w2(32'hba026631),
	.w3(32'hb6e7ac28),
	.w4(32'h39b7444b),
	.w5(32'hb99e4d24),
	.w6(32'hbabe75c5),
	.w7(32'hba381738),
	.w8(32'hb990dd34),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79821bd),
	.w1(32'hb58a2129),
	.w2(32'hb7f8c6dd),
	.w3(32'hb7b5cf89),
	.w4(32'h36afb397),
	.w5(32'hb7f559bb),
	.w6(32'hb7ae3a8a),
	.w7(32'hb7d6661f),
	.w8(32'hb7c2b6b0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69f470),
	.w1(32'h39d7b1db),
	.w2(32'hba48af26),
	.w3(32'h3a71a9ec),
	.w4(32'h39e0e69e),
	.w5(32'h39f53bf7),
	.w6(32'hba8224a9),
	.w7(32'h3903e64a),
	.w8(32'h3a484143),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0992af),
	.w1(32'h3a96349d),
	.w2(32'h3b503db9),
	.w3(32'hbafe051b),
	.w4(32'hba5ee572),
	.w5(32'h3b495ae7),
	.w6(32'hbad4206c),
	.w7(32'hbaaded75),
	.w8(32'h3ae4bb6a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0df483),
	.w1(32'h3a08a01b),
	.w2(32'h3a931dba),
	.w3(32'h39294a0f),
	.w4(32'h39e20ebd),
	.w5(32'h3a7bca4a),
	.w6(32'hb91b644f),
	.w7(32'h38c684cd),
	.w8(32'h3a007350),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74f681c),
	.w1(32'hb74a1dc2),
	.w2(32'hb7f08602),
	.w3(32'h37320fc9),
	.w4(32'hb7b06b06),
	.w5(32'hb80d11d1),
	.w6(32'h371a4dc2),
	.w7(32'hb75acbcc),
	.w8(32'hb7cce761),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b100517),
	.w1(32'hba9ba28b),
	.w2(32'h3b0c85cf),
	.w3(32'hba405702),
	.w4(32'h3a90efb5),
	.w5(32'h3b3eac58),
	.w6(32'hbbedd5f7),
	.w7(32'hbbc72a81),
	.w8(32'hbacab10a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55caca),
	.w1(32'h3a05d370),
	.w2(32'h3aa8a2e9),
	.w3(32'hb96f1d1c),
	.w4(32'h39692e0d),
	.w5(32'h3a97f4a0),
	.w6(32'hbb061045),
	.w7(32'hba9bac45),
	.w8(32'h3986ee7e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39382b38),
	.w1(32'h37d84e39),
	.w2(32'hb8bc8314),
	.w3(32'h3887f8eb),
	.w4(32'h3803111f),
	.w5(32'hb849cb17),
	.w6(32'hb7282206),
	.w7(32'h372f521c),
	.w8(32'hb7f1fa0e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34df8d),
	.w1(32'h39b59aa0),
	.w2(32'h3a8b407a),
	.w3(32'hb9660eb0),
	.w4(32'h3a0eef52),
	.w5(32'h3a92297c),
	.w6(32'hbb190453),
	.w7(32'hbad65a72),
	.w8(32'h375e14d6),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb878aefc),
	.w1(32'h387651da),
	.w2(32'h38fa641b),
	.w3(32'hb881ca8a),
	.w4(32'h383d0882),
	.w5(32'h392e0aca),
	.w6(32'h37bf4352),
	.w7(32'h38d9dfa5),
	.w8(32'h39438c41),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3803f91f),
	.w1(32'hb61c6515),
	.w2(32'h39db9507),
	.w3(32'hb94c35da),
	.w4(32'hb98a33ff),
	.w5(32'h38e8203f),
	.w6(32'hb935ee3b),
	.w7(32'hb91bac69),
	.w8(32'h385bbba6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378ea0d3),
	.w1(32'h3761680b),
	.w2(32'hb8320f21),
	.w3(32'h37a9f484),
	.w4(32'h3782fddc),
	.w5(32'hb822202c),
	.w6(32'h37b50f13),
	.w7(32'h370b0d4b),
	.w8(32'hb8188b2b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bfb690),
	.w1(32'hb75eb96a),
	.w2(32'hb7fa4c38),
	.w3(32'hb738b958),
	.w4(32'hb74ebd13),
	.w5(32'hb81b65ec),
	.w6(32'hb7a562a7),
	.w7(32'hb6f07d4e),
	.w8(32'hb7098382),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77c720),
	.w1(32'hba188d12),
	.w2(32'hb9fb0901),
	.w3(32'h3a69b77b),
	.w4(32'hb9a3e7c1),
	.w5(32'hb9b9dd86),
	.w6(32'h3b003db8),
	.w7(32'h39a38cba),
	.w8(32'hb8e1c8f8),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fba68),
	.w1(32'h39d37377),
	.w2(32'h3b480af0),
	.w3(32'h3ab939a2),
	.w4(32'h3ab96583),
	.w5(32'h3b0a55ce),
	.w6(32'h3b3b5b02),
	.w7(32'h3b915182),
	.w8(32'h3b4b4d1e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34b1db),
	.w1(32'h3aff1eaa),
	.w2(32'h3b0e0c60),
	.w3(32'h3abec814),
	.w4(32'h3ac1db8a),
	.w5(32'h3af912d8),
	.w6(32'hbaa8ba78),
	.w7(32'hb9d0e89d),
	.w8(32'h3a9bb6b3),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e69b1),
	.w1(32'h3a9ed912),
	.w2(32'h3ae698cd),
	.w3(32'h39e22cd0),
	.w4(32'h3ab44f16),
	.w5(32'h3af77d5a),
	.w6(32'h39443c74),
	.w7(32'h3b0d24a3),
	.w8(32'h3ae95779),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3742c55c),
	.w1(32'hb9230805),
	.w2(32'hb9ac170a),
	.w3(32'hb6b51d48),
	.w4(32'hb98ced39),
	.w5(32'hb9c3328c),
	.w6(32'h383bc5d1),
	.w7(32'hb95c2843),
	.w8(32'hb96f886d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904531a),
	.w1(32'hb7b4ec9c),
	.w2(32'h39460e81),
	.w3(32'hb96a44af),
	.w4(32'hb7f0b1f8),
	.w5(32'h39c629ee),
	.w6(32'hb9bf9366),
	.w7(32'h38b271fe),
	.w8(32'h39b89e2c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67dd280),
	.w1(32'hb728d890),
	.w2(32'hb769eed1),
	.w3(32'hb6b5a917),
	.w4(32'hb73d3f8c),
	.w5(32'hb7bb7e61),
	.w6(32'hb6e1f88d),
	.w7(32'hb7103dd6),
	.w8(32'hb76b603a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cabea8),
	.w1(32'hb79b2be0),
	.w2(32'h3684ed34),
	.w3(32'hb841f09a),
	.w4(32'hb817a899),
	.w5(32'hb7eb8fb6),
	.w6(32'hb8106df7),
	.w7(32'hb8189ab7),
	.w8(32'hb72d63cd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e2b02),
	.w1(32'h3a209106),
	.w2(32'h397ff35b),
	.w3(32'h3a8b254f),
	.w4(32'h3a2819d4),
	.w5(32'hb7516acc),
	.w6(32'hba03fa54),
	.w7(32'h3a2e6334),
	.w8(32'hb9f5876b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ad83fa),
	.w1(32'h38f9c2e2),
	.w2(32'h38f02ce4),
	.w3(32'h390ada6b),
	.w4(32'h39003f5d),
	.w5(32'h3907a1c1),
	.w6(32'h3910acb0),
	.w7(32'h390f5975),
	.w8(32'h39192475),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d73d96),
	.w1(32'hb98dfa7f),
	.w2(32'hb9f14562),
	.w3(32'hb9925354),
	.w4(32'hb96ac94c),
	.w5(32'hba1f058a),
	.w6(32'hb84fe80e),
	.w7(32'hb8dfcc96),
	.w8(32'hb9ae9695),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ca973),
	.w1(32'hb91d38c5),
	.w2(32'hb9d01850),
	.w3(32'hb99e6e8a),
	.w4(32'h399c8275),
	.w5(32'hb781f04b),
	.w6(32'hb9923500),
	.w7(32'h3a008a8a),
	.w8(32'hb9095286),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4ffccfc),
	.w1(32'hb6321132),
	.w2(32'hb7756831),
	.w3(32'hb7b23c93),
	.w4(32'h35c7d95a),
	.w5(32'hb7329377),
	.w6(32'hb7376bff),
	.w7(32'hb68a76f1),
	.w8(32'hb6d470b9),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3772a458),
	.w1(32'h398760cb),
	.w2(32'h3982d217),
	.w3(32'h384f12fc),
	.w4(32'h39c4d0b4),
	.w5(32'h39cd7e2f),
	.w6(32'hba4b5d61),
	.w7(32'hb9632f92),
	.w8(32'hb90c2046),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3898325c),
	.w1(32'h388b7c0a),
	.w2(32'h39160233),
	.w3(32'h3824af93),
	.w4(32'h38e44e46),
	.w5(32'h38cfbdcd),
	.w6(32'h38a451cb),
	.w7(32'h3914700a),
	.w8(32'h395e5e96),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d93d8),
	.w1(32'h3a101279),
	.w2(32'h3b2e194a),
	.w3(32'h3ab267c2),
	.w4(32'h3ad3e8ec),
	.w5(32'hba0ff0c4),
	.w6(32'h3b208a98),
	.w7(32'h3ba1e4cd),
	.w8(32'h3a3ed17d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab3474),
	.w1(32'hb8afe4e4),
	.w2(32'hb9660986),
	.w3(32'hb8b1d48f),
	.w4(32'hb88df854),
	.w5(32'hb90dce1b),
	.w6(32'h33345e08),
	.w7(32'hb706a87c),
	.w8(32'hb821a9ce),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f63cd),
	.w1(32'hb92ab822),
	.w2(32'hbaa8fc5b),
	.w3(32'h3988a80a),
	.w4(32'hb9d263a7),
	.w5(32'hbb21505d),
	.w6(32'hba927532),
	.w7(32'hbb2fcd71),
	.w8(32'hbb351585),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule