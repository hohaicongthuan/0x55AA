module layer_8_featuremap_61(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69bb05),
	.w1(32'h39e03ebf),
	.w2(32'h397294ab),
	.w3(32'hbc348d01),
	.w4(32'hbb971d8c),
	.w5(32'hba7d8426),
	.w6(32'hbb1e4851),
	.w7(32'h3a32c174),
	.w8(32'h3b8ebda2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2ffe3),
	.w1(32'h3b5e99ab),
	.w2(32'hba96bde0),
	.w3(32'h3ba849fd),
	.w4(32'h3b007eb7),
	.w5(32'hb891fd2b),
	.w6(32'h3b0b2e3a),
	.w7(32'h3a147a80),
	.w8(32'h3b341095),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b042bc8),
	.w1(32'h39e7c6cd),
	.w2(32'hbaa8d275),
	.w3(32'h3ad4852d),
	.w4(32'h39ffe41d),
	.w5(32'hba137407),
	.w6(32'h3acb9001),
	.w7(32'h3a02a6b8),
	.w8(32'hbb6fa58d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fc2d9),
	.w1(32'h3bb04783),
	.w2(32'h3b47fcc1),
	.w3(32'h3c105c68),
	.w4(32'h3bc29c41),
	.w5(32'h3b938f09),
	.w6(32'h3beab30e),
	.w7(32'h3c5c304a),
	.w8(32'h3bcbb395),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd73de5),
	.w1(32'h3b070399),
	.w2(32'hbbbd488c),
	.w3(32'h3b48191f),
	.w4(32'h3a0d262a),
	.w5(32'hbb6782d5),
	.w6(32'h3b9939e3),
	.w7(32'hbb12a2be),
	.w8(32'h3cf41d9a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7ea051),
	.w1(32'h3acaec9d),
	.w2(32'hbd4fd12b),
	.w3(32'h3d1fda09),
	.w4(32'hbae606f4),
	.w5(32'hbd0b384b),
	.w6(32'hbb81f2da),
	.w7(32'hbd17a862),
	.w8(32'hbc136c71),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2d846),
	.w1(32'h3985c91e),
	.w2(32'hbb833677),
	.w3(32'hba627920),
	.w4(32'hba6a94af),
	.w5(32'hba755eae),
	.w6(32'h3ab34a00),
	.w7(32'hb9ee84a7),
	.w8(32'hb9087397),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b126678),
	.w1(32'h3bbbb290),
	.w2(32'h3b392e9e),
	.w3(32'hbafa2ef5),
	.w4(32'h3bb1a5eb),
	.w5(32'h3c0238fc),
	.w6(32'h3b81b8d4),
	.w7(32'h3aa22736),
	.w8(32'h3b0025a2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba326880),
	.w1(32'hba2cb492),
	.w2(32'hbb844d0a),
	.w3(32'hbb6e8121),
	.w4(32'hbb4edea5),
	.w5(32'hbb2b3c68),
	.w6(32'hb8661410),
	.w7(32'hba8e874d),
	.w8(32'hbc6e9cf7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98a7ed),
	.w1(32'hbb8e8fee),
	.w2(32'h3ce0949f),
	.w3(32'hbb15ca05),
	.w4(32'hbb825311),
	.w5(32'hbc12fcb9),
	.w6(32'hbbe226de),
	.w7(32'h3c89caf4),
	.w8(32'h3b120e26),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3eccb7),
	.w1(32'hbb82bb87),
	.w2(32'hbb9d52a7),
	.w3(32'hbc69e792),
	.w4(32'hbba04932),
	.w5(32'hb821a70e),
	.w6(32'h3a519c2a),
	.w7(32'h39fd01dc),
	.w8(32'h3ba4613d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6156a9),
	.w1(32'h391be9f5),
	.w2(32'h3a1aa07c),
	.w3(32'hbba9aefc),
	.w4(32'hbbb4a349),
	.w5(32'h3af34ecc),
	.w6(32'hbb4848db),
	.w7(32'hba2880b3),
	.w8(32'hbb4ffbcd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b023bf7),
	.w1(32'h3a0238ab),
	.w2(32'hbad4ff9e),
	.w3(32'hba09bd04),
	.w4(32'hba09bd03),
	.w5(32'h39b44e32),
	.w6(32'h3b7c34e2),
	.w7(32'h3b008b69),
	.w8(32'h3d1e11d2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7e8c49),
	.w1(32'h38c22e41),
	.w2(32'hbd5d2a43),
	.w3(32'h3d1dd4b9),
	.w4(32'hbb061b1c),
	.w5(32'hbd060535),
	.w6(32'hbc0da1ce),
	.w7(32'hbd24d2e5),
	.w8(32'h3c89a063),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d02efda),
	.w1(32'h3abe40e2),
	.w2(32'hbd07e24b),
	.w3(32'h3ca2b82e),
	.w4(32'h3b26e46f),
	.w5(32'hbc9b53bb),
	.w6(32'hbb31f533),
	.w7(32'hbcbac111),
	.w8(32'h3b2f01c0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80fe5a),
	.w1(32'hba599002),
	.w2(32'hb97bcd22),
	.w3(32'h3abb8f06),
	.w4(32'hba855823),
	.w5(32'h3a813929),
	.w6(32'hba2e37e9),
	.w7(32'hb8bebb4d),
	.w8(32'hbb3d8fa0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc389cd9),
	.w1(32'h399c231f),
	.w2(32'h3cc4cc28),
	.w3(32'h3bf7e3cc),
	.w4(32'hb980bf39),
	.w5(32'hbbcfd10e),
	.w6(32'hbb92fd2b),
	.w7(32'h3b277457),
	.w8(32'h3a91f718),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4d956),
	.w1(32'h3bcb2968),
	.w2(32'h3c1719cb),
	.w3(32'hbbfcc09a),
	.w4(32'hbac57f06),
	.w5(32'h3b69589d),
	.w6(32'h3b4bacde),
	.w7(32'h3b810c73),
	.w8(32'hbbe56b78),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfac8d4),
	.w1(32'h3a2bb647),
	.w2(32'h3bb4666f),
	.w3(32'hbcc87281),
	.w4(32'h3b9ae51d),
	.w5(32'h3cbde8a1),
	.w6(32'hbbbd5e1a),
	.w7(32'hbacb8538),
	.w8(32'h3c44a53e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fbc93d),
	.w1(32'h3c22a3bc),
	.w2(32'h3c86cc5a),
	.w3(32'hbc7141fa),
	.w4(32'hbc3fc775),
	.w5(32'hbc003777),
	.w6(32'h3ad0e202),
	.w7(32'hbb8d51a6),
	.w8(32'hbc45b3fb),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8aa1ac),
	.w1(32'h3b9d4af8),
	.w2(32'h3c8c92b4),
	.w3(32'hbc974bc4),
	.w4(32'hbb861935),
	.w5(32'h3b1b1245),
	.w6(32'h3aaef922),
	.w7(32'h3c07d5b9),
	.w8(32'hbac7bc5e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a9631),
	.w1(32'h3bbf4bd6),
	.w2(32'hbb12a033),
	.w3(32'h3c15b71d),
	.w4(32'h3be3d373),
	.w5(32'h3adfbb53),
	.w6(32'h3c0bc875),
	.w7(32'h3a3f8bfc),
	.w8(32'hbc978ce0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8357c8),
	.w1(32'hbb8f7677),
	.w2(32'h3d631ac7),
	.w3(32'hbd7277ba),
	.w4(32'hbc6351e8),
	.w5(32'h3d06b28c),
	.w6(32'hbcdb6cbd),
	.w7(32'h3cc8cdb8),
	.w8(32'hbba35910),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab92a5e),
	.w1(32'h3ba13580),
	.w2(32'hbabdacae),
	.w3(32'hbbc32fc9),
	.w4(32'hbb4fa9ad),
	.w5(32'hbb1950d8),
	.w6(32'hbae99268),
	.w7(32'h3aef5bd6),
	.w8(32'hbbacbd1f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c179a),
	.w1(32'h3ae72b4a),
	.w2(32'h3cdb16c3),
	.w3(32'hbc2834f8),
	.w4(32'hbb6a656d),
	.w5(32'h3c6311ed),
	.w6(32'h3aba64ca),
	.w7(32'h3c288d22),
	.w8(32'hbc9bae5e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0845b4),
	.w1(32'h3b138767),
	.w2(32'h3d49a9c0),
	.w3(32'hbcc9472a),
	.w4(32'hbb5fe2c9),
	.w5(32'h3cf8b531),
	.w6(32'hbc2c53bb),
	.w7(32'h3cc49a8c),
	.w8(32'hbc8d5875),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc927c7),
	.w1(32'h3a55bc9f),
	.w2(32'h3d1ab006),
	.w3(32'hbc772c0f),
	.w4(32'hbb95d015),
	.w5(32'h3caf2de1),
	.w6(32'hbb5cd226),
	.w7(32'h3ca22730),
	.w8(32'hbc8a821f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf25fc3),
	.w1(32'h3d50d1ef),
	.w2(32'h3daee55e),
	.w3(32'hbd142894),
	.w4(32'h3d02b49c),
	.w5(32'h3d8fb858),
	.w6(32'hbc71bf1c),
	.w7(32'h3cbbc783),
	.w8(32'h3c983f35),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6dba63),
	.w1(32'hbb2a21be),
	.w2(32'h3c32fd1e),
	.w3(32'hbc723994),
	.w4(32'hbc273495),
	.w5(32'h3b83e564),
	.w6(32'hbc44d4c1),
	.w7(32'hbb295130),
	.w8(32'h3b982785),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a3cd1),
	.w1(32'hb909c3ef),
	.w2(32'hbb86dcd1),
	.w3(32'h3b450202),
	.w4(32'h3ab27338),
	.w5(32'hba3afc9e),
	.w6(32'h3ace127f),
	.w7(32'hb95d5ace),
	.w8(32'h3c2a2c35),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36d60e),
	.w1(32'h399b3e3a),
	.w2(32'h3c084b6c),
	.w3(32'hbcc8da6e),
	.w4(32'h3b8c6ce4),
	.w5(32'h3caf40c2),
	.w6(32'h3ba089b0),
	.w7(32'hbbc2eaa0),
	.w8(32'hbcb48f46),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd13e3bf),
	.w1(32'h3bb28210),
	.w2(32'h3d181c27),
	.w3(32'hbc9c2669),
	.w4(32'h3be6a1ee),
	.w5(32'h3cd9992b),
	.w6(32'h3bca2121),
	.w7(32'h3cbaa560),
	.w8(32'hbb32cc69),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba6d10),
	.w1(32'h3b0803c2),
	.w2(32'hbc4ca779),
	.w3(32'hbbbbc441),
	.w4(32'hbbf230f6),
	.w5(32'hbb401dfe),
	.w6(32'hbac13728),
	.w7(32'h3ab8c58c),
	.w8(32'h3b96f9e9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bf35f),
	.w1(32'h3c491478),
	.w2(32'h3c80a197),
	.w3(32'hbb06a730),
	.w4(32'hba6c10f3),
	.w5(32'hbb182671),
	.w6(32'h3b529a82),
	.w7(32'h3a0a9646),
	.w8(32'h3d047159),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d72442b),
	.w1(32'hb8954c20),
	.w2(32'hbd4a59b3),
	.w3(32'h3d162730),
	.w4(32'hbbb8d530),
	.w5(32'hbd10f0bb),
	.w6(32'hbbbc42bb),
	.w7(32'hbd158f76),
	.w8(32'hbbe5e2cf),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ed6b1),
	.w1(32'h3bbcd717),
	.w2(32'h3bf4665f),
	.w3(32'hbb7bdc6f),
	.w4(32'h3b98f14a),
	.w5(32'h3c444a40),
	.w6(32'hba470ad4),
	.w7(32'h3b2b8cdc),
	.w8(32'hbc6f07f0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd1e453),
	.w1(32'h3b7f14ec),
	.w2(32'h3cc36031),
	.w3(32'hbc9630ba),
	.w4(32'hbb11ddc3),
	.w5(32'h3bcf6af7),
	.w6(32'h3b17b7d7),
	.w7(32'h3c53d19e),
	.w8(32'h3b45d2a6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93713e),
	.w1(32'h3a87dfbc),
	.w2(32'hbb53dda4),
	.w3(32'h3b79cfba),
	.w4(32'h3b4015f7),
	.w5(32'hb9fa41ae),
	.w6(32'h3b2c1c9b),
	.w7(32'h3af93404),
	.w8(32'h3cd3838f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5c8f6f),
	.w1(32'h3b8351d8),
	.w2(32'hbd7710d7),
	.w3(32'h3cfe9585),
	.w4(32'h3bbbae82),
	.w5(32'hbd0b5427),
	.w6(32'hbba18465),
	.w7(32'hbd29baa9),
	.w8(32'hbc8ea7b3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb837f9),
	.w1(32'h3b85d1bf),
	.w2(32'h3cbae140),
	.w3(32'hbc7c309a),
	.w4(32'h3a073ebc),
	.w5(32'h3c53cb54),
	.w6(32'hba515a5c),
	.w7(32'h3c5a33ff),
	.w8(32'hbc0c2bad),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc913a66),
	.w1(32'h3ad6e128),
	.w2(32'h3ce2a20d),
	.w3(32'hbc93cab3),
	.w4(32'hbbb18426),
	.w5(32'h3c41c878),
	.w6(32'h3a30eb9a),
	.w7(32'h3c9b10d6),
	.w8(32'h3b57bd03),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8035b3),
	.w1(32'hba6e7e2b),
	.w2(32'h3b62540b),
	.w3(32'h38e5744b),
	.w4(32'hb92cfd7a),
	.w5(32'h3bec3fee),
	.w6(32'hb9c0724a),
	.w7(32'hbc10bb52),
	.w8(32'hbc8d7456),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd205d3),
	.w1(32'hbaea6e58),
	.w2(32'h3bda53e8),
	.w3(32'h3c5079fd),
	.w4(32'h3b92e765),
	.w5(32'hbc2cf194),
	.w6(32'hbcac77eb),
	.w7(32'h3c002111),
	.w8(32'h3a8017c9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f85a2),
	.w1(32'hbbc649c9),
	.w2(32'h3b35da26),
	.w3(32'hbc4ab31e),
	.w4(32'hbc1014c2),
	.w5(32'hb907b182),
	.w6(32'h3a5b3f05),
	.w7(32'hbb328f71),
	.w8(32'hbaabf9e0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b2066),
	.w1(32'hbbeab5e8),
	.w2(32'h3990729d),
	.w3(32'hbc7a9893),
	.w4(32'hbb184eb2),
	.w5(32'h3c0f56fd),
	.w6(32'hbbb745dd),
	.w7(32'hbc28e939),
	.w8(32'h3b17fe11),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9e540),
	.w1(32'h3833d339),
	.w2(32'h3b6cfaf2),
	.w3(32'h3c3401cd),
	.w4(32'h3bf2bcea),
	.w5(32'h3c89259f),
	.w6(32'hbb21fd20),
	.w7(32'hbc3fa0a2),
	.w8(32'h362c4e70),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd875c8),
	.w1(32'hbc28d696),
	.w2(32'hbade7094),
	.w3(32'h3c211dc8),
	.w4(32'hbce5c113),
	.w5(32'h3b8f62ad),
	.w6(32'hbc4eb885),
	.w7(32'hbc3f1f52),
	.w8(32'hbbbe2575),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca506b9),
	.w1(32'hbc802d44),
	.w2(32'hbc23bf76),
	.w3(32'hbb3fbf78),
	.w4(32'hbc48859b),
	.w5(32'hbb9225c6),
	.w6(32'hbc45e963),
	.w7(32'hbc43b366),
	.w8(32'h3b96ca9f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cda9c73),
	.w1(32'h3ae4d79b),
	.w2(32'hbc571cbb),
	.w3(32'h3ccfa0ff),
	.w4(32'h3cb35622),
	.w5(32'h3bf29c23),
	.w6(32'hbca640c7),
	.w7(32'hbc5cb588),
	.w8(32'h3a4a9f55),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d02c9),
	.w1(32'hbc2a0286),
	.w2(32'h3b182bc3),
	.w3(32'hbc00f996),
	.w4(32'hbc0db681),
	.w5(32'h3be1a1e1),
	.w6(32'h39ceb0b6),
	.w7(32'hbc34830c),
	.w8(32'h3b7f1037),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08c324),
	.w1(32'h3bccc9f3),
	.w2(32'h3b801d88),
	.w3(32'h3c002522),
	.w4(32'h3bc87cc2),
	.w5(32'hbb09cf09),
	.w6(32'h3c4ced9b),
	.w7(32'h3c201fa7),
	.w8(32'h3a856f34),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0be11),
	.w1(32'h3b358a07),
	.w2(32'h3c1b621a),
	.w3(32'hbcc71c16),
	.w4(32'h3bc9557f),
	.w5(32'h3c868b21),
	.w6(32'h3b14573f),
	.w7(32'hbb4abe29),
	.w8(32'h3be282a8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a4038),
	.w1(32'h3c09b518),
	.w2(32'hbc5445d7),
	.w3(32'hbd0e51a7),
	.w4(32'h3c513411),
	.w5(32'h3b3c8e5d),
	.w6(32'hbd1eb6e6),
	.w7(32'hbc0cfd8e),
	.w8(32'h3bcfa552),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca24aae),
	.w1(32'h3c167301),
	.w2(32'hbb197469),
	.w3(32'h3c42bf56),
	.w4(32'h3c858e31),
	.w5(32'h3b84c9b3),
	.w6(32'hbbff34ba),
	.w7(32'hbc9f8944),
	.w8(32'hbc9c707a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bbe58),
	.w1(32'hbb005777),
	.w2(32'h3ba53386),
	.w3(32'h3d0b243d),
	.w4(32'hbc9c4d33),
	.w5(32'hbc2bd959),
	.w6(32'hbb4afe2a),
	.w7(32'h3ca486b6),
	.w8(32'h3c528708),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2462d6),
	.w1(32'hbbe33d7b),
	.w2(32'h3cc23aef),
	.w3(32'hbc3dfc3f),
	.w4(32'hbab8d6fc),
	.w5(32'h3ca30af0),
	.w6(32'hbc033fd9),
	.w7(32'h3bdc2a6f),
	.w8(32'h3c8ad146),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92e327),
	.w1(32'hbc0aebed),
	.w2(32'h3bca891c),
	.w3(32'hbc139919),
	.w4(32'hba65d303),
	.w5(32'hbbb8f779),
	.w6(32'h3bbc7fb4),
	.w7(32'h3b8851ba),
	.w8(32'hbb90b7ae),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dad42),
	.w1(32'hbb8dacc8),
	.w2(32'hbc3984cc),
	.w3(32'h39e82e04),
	.w4(32'hbb0bd285),
	.w5(32'h3a6247ba),
	.w6(32'hbc27d860),
	.w7(32'h3b1e99d4),
	.w8(32'h3c3c40da),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc697311),
	.w1(32'hbbff971f),
	.w2(32'h3c621799),
	.w3(32'hbc7e1969),
	.w4(32'hbbed8b73),
	.w5(32'h3c2a9612),
	.w6(32'h3bd688dd),
	.w7(32'h3ca6666c),
	.w8(32'h3b348d2b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0c900),
	.w1(32'hbbbb6662),
	.w2(32'hbc32a45a),
	.w3(32'h3c0c1599),
	.w4(32'hba9b9721),
	.w5(32'hbb9a6370),
	.w6(32'hbc62176a),
	.w7(32'hbc5da274),
	.w8(32'h3b3ef994),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5b114),
	.w1(32'h3bc27fa3),
	.w2(32'h3c8efe2b),
	.w3(32'h3cd2ad87),
	.w4(32'h3b7a0c08),
	.w5(32'h3b7a5842),
	.w6(32'hbc8f2cb1),
	.w7(32'hbc25265b),
	.w8(32'h3b16799b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9f246),
	.w1(32'hbc00a14a),
	.w2(32'hbba45937),
	.w3(32'h3c3b88b7),
	.w4(32'h3bfddd36),
	.w5(32'hba8e3b42),
	.w6(32'h3c0460d8),
	.w7(32'hba1791df),
	.w8(32'h3bbf6469),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1fd44),
	.w1(32'h3bbf1762),
	.w2(32'h3ccf8641),
	.w3(32'hbc864037),
	.w4(32'hbb4daf72),
	.w5(32'h3c8a4bae),
	.w6(32'h3b3a9532),
	.w7(32'h3c0982cb),
	.w8(32'h3b963390),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99799b),
	.w1(32'hb98c4155),
	.w2(32'hbc4fc20d),
	.w3(32'h3b5dd56b),
	.w4(32'hbabc6b40),
	.w5(32'h3bfb22dc),
	.w6(32'hbcd87dc1),
	.w7(32'hbb6a51a2),
	.w8(32'h3bb91d76),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a4484),
	.w1(32'hbbafa729),
	.w2(32'h3a18b99e),
	.w3(32'h3a4f9d04),
	.w4(32'hbbb67ced),
	.w5(32'h3abe418a),
	.w6(32'hbb7931e9),
	.w7(32'hbb86f7f4),
	.w8(32'h3a75da4c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941b67),
	.w1(32'h3ac1f1d2),
	.w2(32'h3b81b03d),
	.w3(32'hbb3b48e3),
	.w4(32'h38aac517),
	.w5(32'h3b055d73),
	.w6(32'h3b204d34),
	.w7(32'hbafc152c),
	.w8(32'h3b09538b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95a8ed),
	.w1(32'hba3cd6e2),
	.w2(32'h3b2fa1bd),
	.w3(32'h38f88d2d),
	.w4(32'h3b0f6299),
	.w5(32'h3b25e8dd),
	.w6(32'h3b94393e),
	.w7(32'h3a69f954),
	.w8(32'hbbf1e898),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca7b3b6),
	.w1(32'hbc27129a),
	.w2(32'h3a91e31e),
	.w3(32'h3c0a5e81),
	.w4(32'h3ba524e8),
	.w5(32'h3c52d16a),
	.w6(32'hbc20b0e0),
	.w7(32'hbc5c7bab),
	.w8(32'hbb04114b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95c25b),
	.w1(32'hbb8f6a57),
	.w2(32'hbac6bbca),
	.w3(32'hbb196e56),
	.w4(32'hbaad8be3),
	.w5(32'h3b1e01e9),
	.w6(32'hbb096d53),
	.w7(32'hbc0449b9),
	.w8(32'h3c448d0a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd70b09f),
	.w1(32'hbc86f910),
	.w2(32'h3cfe7e1c),
	.w3(32'hbd5b5196),
	.w4(32'hbd12ad41),
	.w5(32'h3b82cc09),
	.w6(32'h3d29db4e),
	.w7(32'h3d59c77e),
	.w8(32'hbbd6d4a7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95afdc),
	.w1(32'hbb79402c),
	.w2(32'hbb097164),
	.w3(32'hbb2ffd96),
	.w4(32'hbb0bd37c),
	.w5(32'h3ab28c24),
	.w6(32'hbb9edac3),
	.w7(32'hbc20e225),
	.w8(32'hbb05577d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6db7b7),
	.w1(32'hbafa923a),
	.w2(32'hbadd417a),
	.w3(32'hbb4fe768),
	.w4(32'hbb0cee58),
	.w5(32'h3a364445),
	.w6(32'hbb10f2f1),
	.w7(32'hbbdca408),
	.w8(32'h3b8e88ef),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb932960),
	.w1(32'hbb39b0c8),
	.w2(32'hbb91ac15),
	.w3(32'hbb2f52db),
	.w4(32'hb9f6150b),
	.w5(32'h3a5a3a1c),
	.w6(32'hbb8f0fb4),
	.w7(32'hbc5a6561),
	.w8(32'hbc07f5be),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce44a3a),
	.w1(32'hb98537d7),
	.w2(32'hbd12cfd5),
	.w3(32'hbd0cdcff),
	.w4(32'hbd171e61),
	.w5(32'h3a9395a8),
	.w6(32'hbd1b5c07),
	.w7(32'hbcf0a963),
	.w8(32'h3af4f5eb),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa54f8a),
	.w1(32'hbb904ba1),
	.w2(32'hbc16ed0e),
	.w3(32'h3bcba716),
	.w4(32'h3b08c1d4),
	.w5(32'h3acc2741),
	.w6(32'hbbf93b2e),
	.w7(32'hbc494617),
	.w8(32'hb9411864),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9043d5),
	.w1(32'hbb6c2d71),
	.w2(32'h3989cd53),
	.w3(32'hbbe2446c),
	.w4(32'hbba4586b),
	.w5(32'hb939840b),
	.w6(32'hbb312b73),
	.w7(32'hbbfcbbda),
	.w8(32'hbad6d047),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab2018),
	.w1(32'hbb8ca34a),
	.w2(32'hbb87329b),
	.w3(32'h3b0b03d0),
	.w4(32'h3af5cf71),
	.w5(32'h3a1744ad),
	.w6(32'hbb96d316),
	.w7(32'hbc1f8847),
	.w8(32'h3c743c6f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd60fb0a),
	.w1(32'hbc073808),
	.w2(32'h3d49b349),
	.w3(32'hbd522ab8),
	.w4(32'hbd12751f),
	.w5(32'h3c32750b),
	.w6(32'h3d404c03),
	.w7(32'h3d8388e6),
	.w8(32'h3b8981a8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec24b2),
	.w1(32'h3b735f29),
	.w2(32'h3d2b444d),
	.w3(32'hbd114c9a),
	.w4(32'hbcb3d0ab),
	.w5(32'h3c95122a),
	.w6(32'h3cc11f36),
	.w7(32'h3d022c04),
	.w8(32'h3c6d658a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97d0ff),
	.w1(32'hbbf3767d),
	.w2(32'hbb81de19),
	.w3(32'h3a037a3b),
	.w4(32'hbbdc9175),
	.w5(32'hbb3c6c8a),
	.w6(32'hbb64ecb3),
	.w7(32'hbb02d39c),
	.w8(32'h3bfd835c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f6a26),
	.w1(32'hbb177eba),
	.w2(32'hbd09d217),
	.w3(32'hbc5ef294),
	.w4(32'hbc804230),
	.w5(32'hbcbd19d2),
	.w6(32'hbb62b01a),
	.w7(32'hbb610819),
	.w8(32'h3b897735),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b368076),
	.w1(32'hba8011ec),
	.w2(32'hbaef1736),
	.w3(32'hb9e86402),
	.w4(32'h3b2a7419),
	.w5(32'hbb7c82de),
	.w6(32'hbaaea099),
	.w7(32'hbb73fa0d),
	.w8(32'h3b379455),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf2b49),
	.w1(32'hbb966117),
	.w2(32'hbbdb05e4),
	.w3(32'hbb07a344),
	.w4(32'h3af1385c),
	.w5(32'hb9da44c9),
	.w6(32'hbc19d2e2),
	.w7(32'hbc93b7c1),
	.w8(32'h3bf3b4fd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66a728),
	.w1(32'h3afe7c19),
	.w2(32'hbcddc6c8),
	.w3(32'h3d033626),
	.w4(32'h3d4b8228),
	.w5(32'hbb425da8),
	.w6(32'h3d18414d),
	.w7(32'hbc0dd15a),
	.w8(32'h3c06524b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beaf0cf),
	.w1(32'h3bddd8cf),
	.w2(32'hbbb25829),
	.w3(32'h3b2b758a),
	.w4(32'h3c8c31f7),
	.w5(32'h3b7c1536),
	.w6(32'hbc76a899),
	.w7(32'hbca8ef84),
	.w8(32'hbb9fa6d4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90fc57),
	.w1(32'hbac9ce0e),
	.w2(32'h39e987b4),
	.w3(32'hbc759475),
	.w4(32'hbb7bff0c),
	.w5(32'h3b899d5f),
	.w6(32'hbb936306),
	.w7(32'hbbac9593),
	.w8(32'h3c02ace0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d7fcf),
	.w1(32'hb9992c08),
	.w2(32'hbc9f05ae),
	.w3(32'h3d052a75),
	.w4(32'h3ce3c79a),
	.w5(32'h3c0c70b0),
	.w6(32'hbcefd97d),
	.w7(32'hbc9db00d),
	.w8(32'h3b9f94d3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96d8b7),
	.w1(32'hbb1a539a),
	.w2(32'hbba31e9b),
	.w3(32'h3b925a10),
	.w4(32'hbbb40d05),
	.w5(32'hbbb29727),
	.w6(32'hb999f4db),
	.w7(32'hbc39402d),
	.w8(32'hbbbca4ca),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c143869),
	.w1(32'h3abd3932),
	.w2(32'hbcbc35b4),
	.w3(32'h3c64598e),
	.w4(32'h3cb13a24),
	.w5(32'hbb89d246),
	.w6(32'hbc12b1cd),
	.w7(32'hbc8cca59),
	.w8(32'h3b202189),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d06be35),
	.w1(32'h39b2ff67),
	.w2(32'hbc959fd5),
	.w3(32'h3cfc4445),
	.w4(32'h3cda56c8),
	.w5(32'h3c115af9),
	.w6(32'hbce0146b),
	.w7(32'hbc91f148),
	.w8(32'h3b3baf25),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d02fd40),
	.w1(32'h3b631c60),
	.w2(32'hbc5a9a3d),
	.w3(32'h3cc3c27f),
	.w4(32'h3ca740ae),
	.w5(32'h3bba1765),
	.w6(32'hbcc6d6cb),
	.w7(32'hbc54ba91),
	.w8(32'hbb9113d4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c502331),
	.w1(32'h3acab7f8),
	.w2(32'hbc78918b),
	.w3(32'h3bc6604f),
	.w4(32'h3c35f8b0),
	.w5(32'hbb2ccfa6),
	.w6(32'hbc53d3a4),
	.w7(32'hbcd31ed0),
	.w8(32'hbbfa74ed),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbefd7c),
	.w1(32'hbcaba691),
	.w2(32'hbcfedddf),
	.w3(32'hbcabca78),
	.w4(32'hbd106ee9),
	.w5(32'hbcaaf60e),
	.w6(32'hbd1f9f1e),
	.w7(32'hbd0a27c0),
	.w8(32'h3a418f41),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941c61),
	.w1(32'h3b1b428e),
	.w2(32'h3bba2a40),
	.w3(32'hbbb7310b),
	.w4(32'hbaabe40a),
	.w5(32'h3b226985),
	.w6(32'h3b358033),
	.w7(32'h3aa4d3f4),
	.w8(32'hbc157def),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb869505),
	.w1(32'hbb1a2f6d),
	.w2(32'hbbbe5127),
	.w3(32'h3d2f7c1c),
	.w4(32'h3ca681ad),
	.w5(32'hbcca0fb9),
	.w6(32'hba5714fb),
	.w7(32'h3bc9a655),
	.w8(32'hba4f3c18),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf490a6),
	.w1(32'h3b0cccb1),
	.w2(32'hbc98a50e),
	.w3(32'h3c87de2d),
	.w4(32'h3cd455f4),
	.w5(32'h3a49f832),
	.w6(32'hbcf027cf),
	.w7(32'hbd241452),
	.w8(32'hbbeabb1a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd2c3c),
	.w1(32'hbc55c5a7),
	.w2(32'h3c1e54b0),
	.w3(32'hbabe27eb),
	.w4(32'h3ad8ed0c),
	.w5(32'hbb8decba),
	.w6(32'h3aeb798a),
	.w7(32'h3bd75e0a),
	.w8(32'hbace0729),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8757b0),
	.w1(32'h3c12a162),
	.w2(32'hbc2cdf27),
	.w3(32'h3c7eb2ca),
	.w4(32'h3aad281b),
	.w5(32'hbb752667),
	.w6(32'h3bd543e5),
	.w7(32'h3c2cc783),
	.w8(32'h3c552037),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1fd2a2),
	.w1(32'hbbdb2fdc),
	.w2(32'h3d2b8409),
	.w3(32'hbd20de9d),
	.w4(32'hbd0763ef),
	.w5(32'h3c17d572),
	.w6(32'h3d2dc076),
	.w7(32'h3d5c8f6a),
	.w8(32'h3b863b29),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b3763),
	.w1(32'hbb5a1816),
	.w2(32'h3a879e44),
	.w3(32'h3af8d63d),
	.w4(32'hbb0797ec),
	.w5(32'h3a2f5b9a),
	.w6(32'hba811cb8),
	.w7(32'hbc120761),
	.w8(32'h3a750c1d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c6ea5),
	.w1(32'hbc363705),
	.w2(32'hbcaeda47),
	.w3(32'h3ca962fe),
	.w4(32'h3b8fa84c),
	.w5(32'hbbaf2340),
	.w6(32'hbca94b56),
	.w7(32'hbca3de8d),
	.w8(32'h3b70298e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b9efb),
	.w1(32'h3b2df4a6),
	.w2(32'h3bb3e4f7),
	.w3(32'hba463659),
	.w4(32'h3a423e95),
	.w5(32'h3b246099),
	.w6(32'h3bae509e),
	.w7(32'h3a600b99),
	.w8(32'h3ba9c162),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd56ed0b),
	.w1(32'hbc3bfbbf),
	.w2(32'h3d2de539),
	.w3(32'hbd68358d),
	.w4(32'hbd582db5),
	.w5(32'h39fd855c),
	.w6(32'h3d4ce173),
	.w7(32'h3d3fcfc7),
	.w8(32'hbbbdb9f7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a1f67),
	.w1(32'h3af9bd32),
	.w2(32'hbc97d720),
	.w3(32'h3c1b7a85),
	.w4(32'h3c3b4902),
	.w5(32'hbc3c53e9),
	.w6(32'hbc6d0347),
	.w7(32'hbcd719f9),
	.w8(32'h3af2dafb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87942a),
	.w1(32'h3886224f),
	.w2(32'hbc108bf1),
	.w3(32'h3c73ffa4),
	.w4(32'h3c212d86),
	.w5(32'h3a956c94),
	.w6(32'hbc2a81dd),
	.w7(32'hbc0c80f3),
	.w8(32'hb7b6b52c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe60c83),
	.w1(32'hb96f368a),
	.w2(32'h3aa59086),
	.w3(32'hbbd36c23),
	.w4(32'h3ac09aa6),
	.w5(32'h3b88b96f),
	.w6(32'hba6f8f10),
	.w7(32'h3a6ecf70),
	.w8(32'hbaa76a91),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8733d8),
	.w1(32'h3aaa8611),
	.w2(32'h3a3e587f),
	.w3(32'h3a857523),
	.w4(32'h3aba7d0c),
	.w5(32'h3a7cedbb),
	.w6(32'h3a8ee406),
	.w7(32'h3a7ac8cf),
	.w8(32'h39eeb6f0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b0deb),
	.w1(32'hb85aa142),
	.w2(32'hb9ee2dc9),
	.w3(32'h3b033f77),
	.w4(32'hba5f05fa),
	.w5(32'hbaff769f),
	.w6(32'h3b230d54),
	.w7(32'h3a7a725d),
	.w8(32'h394b994d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabe1ed),
	.w1(32'hb9c94ace),
	.w2(32'hba19af2b),
	.w3(32'h3a819d34),
	.w4(32'hba039e61),
	.w5(32'hba55848f),
	.w6(32'h3a0166dd),
	.w7(32'h399614cd),
	.w8(32'h3a3c8310),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b092907),
	.w1(32'h3b0d5aab),
	.w2(32'hb9d2d1ba),
	.w3(32'h3a04f47b),
	.w4(32'h3b1c3abd),
	.w5(32'h3a0788a0),
	.w6(32'hba8b62be),
	.w7(32'h3a789f29),
	.w8(32'h3a4fa972),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27784f),
	.w1(32'h3b3363bc),
	.w2(32'h3b92d940),
	.w3(32'h3a8ed5a1),
	.w4(32'hb946131a),
	.w5(32'hba2b5f45),
	.w6(32'h3b044351),
	.w7(32'h3ab09321),
	.w8(32'h3ae9fbf0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3570bd),
	.w1(32'h3b1c1264),
	.w2(32'h3b2727c4),
	.w3(32'h3b6bcf83),
	.w4(32'h3afa78fd),
	.w5(32'h3b247605),
	.w6(32'h3b75cc8a),
	.w7(32'h39abf570),
	.w8(32'h3b2fc232),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a6178),
	.w1(32'hb83ccab2),
	.w2(32'hbb10eb57),
	.w3(32'h3b32221e),
	.w4(32'hbac822dd),
	.w5(32'hbb249f44),
	.w6(32'h3b08c91d),
	.w7(32'hba281cb9),
	.w8(32'hb92e0364),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38110aa2),
	.w1(32'hb900b46c),
	.w2(32'hb9a5c6b3),
	.w3(32'h392c5538),
	.w4(32'h39020fe8),
	.w5(32'hb9981ac8),
	.w6(32'hb91e0411),
	.w7(32'hb989b9cc),
	.w8(32'hb9d9e53a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf470a5),
	.w1(32'hba67f64d),
	.w2(32'h3ac2c3c0),
	.w3(32'hbaf56dd1),
	.w4(32'h3884425a),
	.w5(32'h3af67786),
	.w6(32'hba9bd6a6),
	.w7(32'hba11029e),
	.w8(32'h3b2b00ee),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98baffe),
	.w1(32'hb96933f9),
	.w2(32'hba2f081d),
	.w3(32'hb9ef1277),
	.w4(32'hb92393e5),
	.w5(32'hba0c549d),
	.w6(32'hb738082b),
	.w7(32'hb891c3e2),
	.w8(32'hb9bc8830),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9dbde6),
	.w1(32'hb6be1040),
	.w2(32'hb9709904),
	.w3(32'hba1dc51b),
	.w4(32'hbadd5efa),
	.w5(32'hbaa8843b),
	.w6(32'h3a4a8a47),
	.w7(32'h39035ecd),
	.w8(32'h3a8f3659),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb999899),
	.w1(32'hbb1d7eb1),
	.w2(32'h3b1767f3),
	.w3(32'hbb960b65),
	.w4(32'hbacc7421),
	.w5(32'h3b7dd5de),
	.w6(32'hbb1e179b),
	.w7(32'hb9a2eb9c),
	.w8(32'hb9b54c30),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7146e3b),
	.w1(32'hb804c4d7),
	.w2(32'hb87f1959),
	.w3(32'hb7482870),
	.w4(32'hb7c893c2),
	.w5(32'hb839aa57),
	.w6(32'hb7c0a636),
	.w7(32'hb7ad0377),
	.w8(32'hb8214de3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c6fce),
	.w1(32'h39ab1634),
	.w2(32'h3a7ecb63),
	.w3(32'hba6c96a0),
	.w4(32'hba41c802),
	.w5(32'h39fb424d),
	.w6(32'hb982b425),
	.w7(32'h3a0428e8),
	.w8(32'h3a54f547),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96c870),
	.w1(32'h3b39170d),
	.w2(32'h3b2681f8),
	.w3(32'hbbbe2bbe),
	.w4(32'hbc000ded),
	.w5(32'hbbd18ed4),
	.w6(32'h39d06d77),
	.w7(32'h3b7bb82b),
	.w8(32'h3bc20156),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5eb8b),
	.w1(32'h3b157a6c),
	.w2(32'h3b0a7487),
	.w3(32'h3a6bb3fa),
	.w4(32'h3b6724ff),
	.w5(32'h3b14ee3f),
	.w6(32'hba2201a4),
	.w7(32'h39cf7b07),
	.w8(32'hba607639),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aed2c0),
	.w1(32'h381983b6),
	.w2(32'h37079d4b),
	.w3(32'h39b76733),
	.w4(32'hb878a6da),
	.w5(32'hb9312aad),
	.w6(32'h396af790),
	.w7(32'hb7caca81),
	.w8(32'hb91e19c5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dc794c),
	.w1(32'hb9d15356),
	.w2(32'hb9f1ead9),
	.w3(32'hb914a7d3),
	.w4(32'hba3a5261),
	.w5(32'hba435b7b),
	.w6(32'h38b00b53),
	.w7(32'hb99452f7),
	.w8(32'hb8df8259),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aceca6),
	.w1(32'h38facb2b),
	.w2(32'h381c60f2),
	.w3(32'hb8bc55af),
	.w4(32'h39f81ed3),
	.w5(32'h38c48376),
	.w6(32'hb903b02d),
	.w7(32'h3961156c),
	.w8(32'hb755e0bf),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b363777),
	.w1(32'hbaaa61a9),
	.w2(32'hb9bf4d14),
	.w3(32'h3ad63827),
	.w4(32'hb9bae9ab),
	.w5(32'hba8465b1),
	.w6(32'h3a93f02a),
	.w7(32'hbb14ac3c),
	.w8(32'h3adcb8a2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af65744),
	.w1(32'h3b362235),
	.w2(32'h3bd18bae),
	.w3(32'h3a19ef48),
	.w4(32'hb99a7dde),
	.w5(32'h3b3875f5),
	.w6(32'h3adf18e9),
	.w7(32'h3b1c86c9),
	.w8(32'h3b1b097a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c5ede),
	.w1(32'hbb4e5c19),
	.w2(32'h3b706644),
	.w3(32'hbb7eb10f),
	.w4(32'hbad1c06a),
	.w5(32'h3b8a80c1),
	.w6(32'h3891beaa),
	.w7(32'h39cd9141),
	.w8(32'h3bad559e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule