module layer_10_featuremap_211(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb591476a),
	.w1(32'h36a895bb),
	.w2(32'h3683fc6f),
	.w3(32'hb6943e7b),
	.w4(32'h36dd223b),
	.w5(32'hb5840a05),
	.w6(32'h36b4c660),
	.w7(32'hb5be9887),
	.w8(32'h371c40e6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7860757),
	.w1(32'hb97e8bc7),
	.w2(32'hb9e7450f),
	.w3(32'h38807c11),
	.w4(32'hb9176b00),
	.w5(32'h397e31fc),
	.w6(32'h3a13d5ab),
	.w7(32'h39be9e23),
	.w8(32'h3a1dc753),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d0bf83),
	.w1(32'h36a2538e),
	.w2(32'h37061a61),
	.w3(32'h3625fbcc),
	.w4(32'h36395f20),
	.w5(32'h36a17fbd),
	.w6(32'hb61e18d2),
	.w7(32'hb68c99f7),
	.w8(32'hb5cf0cfb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913e016),
	.w1(32'h3810a489),
	.w2(32'h393cbe78),
	.w3(32'h39575fdd),
	.w4(32'h390c6ae0),
	.w5(32'h39115f53),
	.w6(32'h3911f0c6),
	.w7(32'h38f80f95),
	.w8(32'hb7d3380b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a89173),
	.w1(32'hb6f76fe2),
	.w2(32'h3746c792),
	.w3(32'hb68efabf),
	.w4(32'hb7a6e4c4),
	.w5(32'h33703c70),
	.w6(32'h35e5e4ad),
	.w7(32'hb74e1644),
	.w8(32'h3587728a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61ef2a8),
	.w1(32'hb608029b),
	.w2(32'h369d882c),
	.w3(32'h36e4ead5),
	.w4(32'h358fd7c6),
	.w5(32'h360736ad),
	.w6(32'h37730e41),
	.w7(32'h369465a3),
	.w8(32'h36a7dae8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf3d70),
	.w1(32'hb9b85b25),
	.w2(32'hba12734c),
	.w3(32'hb9fd854f),
	.w4(32'hba2d9bed),
	.w5(32'hba69801b),
	.w6(32'hba5cba29),
	.w7(32'hba50dec2),
	.w8(32'hba3f3d3c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d707d),
	.w1(32'hb8a9c870),
	.w2(32'h39a042b0),
	.w3(32'hb6e0f798),
	.w4(32'h3a194359),
	.w5(32'hb924c5d9),
	.w6(32'h3a9a31c5),
	.w7(32'hb88910a6),
	.w8(32'h3a133e19),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb98ff),
	.w1(32'hba82cdd7),
	.w2(32'hba8cdd5a),
	.w3(32'hb9d0d679),
	.w4(32'hba0fc7e4),
	.w5(32'hba8fb223),
	.w6(32'hb92da674),
	.w7(32'hba21f6eb),
	.w8(32'hbaa25902),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba697e74),
	.w1(32'hb98cde75),
	.w2(32'hb9676f21),
	.w3(32'h3a79d746),
	.w4(32'h3a8511a3),
	.w5(32'hbaba37b7),
	.w6(32'h3a8c0942),
	.w7(32'h3a40226c),
	.w8(32'hbac82eb6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e2d97),
	.w1(32'hb9ac3476),
	.w2(32'hb9d76c2d),
	.w3(32'h383abb35),
	.w4(32'hb9b929b7),
	.w5(32'hba1866ca),
	.w6(32'hb940e081),
	.w7(32'hba139469),
	.w8(32'hba21af4e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ffa314),
	.w1(32'hba770b08),
	.w2(32'hbaa99b6a),
	.w3(32'hba0c2f68),
	.w4(32'hba1ebb50),
	.w5(32'hbac7edc1),
	.w6(32'hba8d7a9c),
	.w7(32'hb90c090f),
	.w8(32'hb9f7edba),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91da0c7),
	.w1(32'hb9845c0f),
	.w2(32'hb924f579),
	.w3(32'h3a7092fe),
	.w4(32'h3a1ba250),
	.w5(32'hba65e2ae),
	.w6(32'h3a48c71c),
	.w7(32'h39c49595),
	.w8(32'hba9adcc0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ea2be),
	.w1(32'h35c0680e),
	.w2(32'hb94d99b4),
	.w3(32'h398b363a),
	.w4(32'h3a07d17e),
	.w5(32'h38cef6bb),
	.w6(32'h394dc703),
	.w7(32'h39ea5d77),
	.w8(32'h38f55493),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba946286),
	.w1(32'hba064016),
	.w2(32'hba1e1071),
	.w3(32'h38eb1523),
	.w4(32'hb89395d7),
	.w5(32'hb9a9f11b),
	.w6(32'hba20214d),
	.w7(32'hb9919bd4),
	.w8(32'hba19178d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e826a),
	.w1(32'h39e371ff),
	.w2(32'h3a9907a8),
	.w3(32'h3a0c71ce),
	.w4(32'h3a2c04a3),
	.w5(32'h3a1eef73),
	.w6(32'h39b11dce),
	.w7(32'h3a4c1eec),
	.w8(32'h390d238f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb777b287),
	.w1(32'hb8e5ce6f),
	.w2(32'hb8bb04f3),
	.w3(32'hb8a0f797),
	.w4(32'hb967c048),
	.w5(32'hb86b69e8),
	.w6(32'hb8e2c5ab),
	.w7(32'hb97f2d9a),
	.w8(32'hb877f0c3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad159c8),
	.w1(32'hba7e2195),
	.w2(32'hb93b1c65),
	.w3(32'hb949442b),
	.w4(32'hb7cd710c),
	.w5(32'hba43d404),
	.w6(32'hba0e72ad),
	.w7(32'hb9b69823),
	.w8(32'hb9da8354),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f7ec9e),
	.w1(32'h38cd06db),
	.w2(32'hb9c86695),
	.w3(32'h3a86e79d),
	.w4(32'h3927387a),
	.w5(32'hba7e4a6d),
	.w6(32'h3a0b86ac),
	.w7(32'hb9b9c9ac),
	.w8(32'hba92b53d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h359dd6b1),
	.w1(32'h36904446),
	.w2(32'h36105427),
	.w3(32'h371f0741),
	.w4(32'hb7fdce70),
	.w5(32'h34231095),
	.w6(32'hb7168697),
	.w7(32'hb7b53072),
	.w8(32'h3763e9ea),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5628f78),
	.w1(32'h36bbbe59),
	.w2(32'h3819be1e),
	.w3(32'h37e163fc),
	.w4(32'h37c3a9ad),
	.w5(32'h383b69a1),
	.w6(32'h37a46ac9),
	.w7(32'h37994091),
	.w8(32'h384d8d54),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947cb66),
	.w1(32'h39d40960),
	.w2(32'h39964983),
	.w3(32'hb71915d9),
	.w4(32'h39afb5e9),
	.w5(32'h39d7a0ad),
	.w6(32'h37ef08a6),
	.w7(32'h39aba471),
	.w8(32'h3a08692d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7f477),
	.w1(32'hbad3e55b),
	.w2(32'hbad74397),
	.w3(32'hba0d45ea),
	.w4(32'hb940d588),
	.w5(32'hbad5a539),
	.w6(32'hba25ce46),
	.w7(32'h3a9d69d5),
	.w8(32'hbb014003),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8caf1),
	.w1(32'h398762ae),
	.w2(32'hb9d3d795),
	.w3(32'h3a2fb961),
	.w4(32'h3a89d7ce),
	.w5(32'hba44c1e3),
	.w6(32'h3a55cd19),
	.w7(32'h3a57305f),
	.w8(32'hb9f28dfa),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaceb0cc),
	.w1(32'hba4c0a2d),
	.w2(32'hbab8159b),
	.w3(32'hba213405),
	.w4(32'hb94a5308),
	.w5(32'hba1d99a4),
	.w6(32'h397e2410),
	.w7(32'h3a2880cd),
	.w8(32'h3954d39f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d45580),
	.w1(32'h39ffd373),
	.w2(32'h3a27210e),
	.w3(32'h398eecb7),
	.w4(32'h3a0cfa21),
	.w5(32'h391b1ae8),
	.w6(32'hb97d2bb5),
	.w7(32'h393fb35e),
	.w8(32'hb8d77d14),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c36e6e),
	.w1(32'hb7ec197c),
	.w2(32'hb7f7469b),
	.w3(32'hb5dfba41),
	.w4(32'hb855a6df),
	.w5(32'hb7922a9d),
	.w6(32'h37d7f355),
	.w7(32'hb81d6b71),
	.w8(32'h37691efc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef8e5a),
	.w1(32'h39bc6195),
	.w2(32'hb9198757),
	.w3(32'hb92893ab),
	.w4(32'hb90049d7),
	.w5(32'hb9f8aee6),
	.w6(32'hb8c55e3f),
	.w7(32'hb9af388f),
	.w8(32'hb97286ac),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885ff18),
	.w1(32'h39850e35),
	.w2(32'h39926980),
	.w3(32'hb855a258),
	.w4(32'h392106ab),
	.w5(32'h39da637c),
	.w6(32'hb65bfc69),
	.w7(32'h398120be),
	.w8(32'h3a43eb94),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec9583),
	.w1(32'h3a907da2),
	.w2(32'h3a4dc75d),
	.w3(32'h3aad83aa),
	.w4(32'h3b06bc48),
	.w5(32'h397484d5),
	.w6(32'h3aa76a7c),
	.w7(32'h3abde1c9),
	.w8(32'hb9b81d2a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37567dc9),
	.w1(32'h36112594),
	.w2(32'h3715299d),
	.w3(32'h36fbb01c),
	.w4(32'hb45e81d6),
	.w5(32'h36ea6e09),
	.w6(32'h36977d64),
	.w7(32'hb6955a0c),
	.w8(32'h3669b2c5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85febcd),
	.w1(32'hb8530cf0),
	.w2(32'hb5e03ecc),
	.w3(32'hb8525936),
	.w4(32'hb8128392),
	.w5(32'h37fbda68),
	.w6(32'hb7fcbea5),
	.w7(32'hb7cef22b),
	.w8(32'h381bcb1c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d85c37),
	.w1(32'hb98eafb0),
	.w2(32'hb98d425d),
	.w3(32'h39418e75),
	.w4(32'h3965d3ce),
	.w5(32'hb9eda94c),
	.w6(32'h39292379),
	.w7(32'h3997dedf),
	.w8(32'hb9465920),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0f81e),
	.w1(32'hb9a5eb1a),
	.w2(32'hb9d8e24f),
	.w3(32'hb73a3568),
	.w4(32'hb88486c7),
	.w5(32'hb934790a),
	.w6(32'h398dac02),
	.w7(32'h39061829),
	.w8(32'hb8223a13),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ca72ec),
	.w1(32'hb8ee831c),
	.w2(32'hb8733aff),
	.w3(32'hb8319f23),
	.w4(32'hb8641104),
	.w5(32'hb923a72d),
	.w6(32'hb91bb222),
	.w7(32'hb8daec2d),
	.w8(32'h37a0f193),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04fb2b),
	.w1(32'hba361485),
	.w2(32'hb9a790b7),
	.w3(32'hb98c1870),
	.w4(32'hba15332a),
	.w5(32'hb99e47bf),
	.w6(32'hb9bb2372),
	.w7(32'hb99b7f0f),
	.w8(32'hb859fac4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05ebcd),
	.w1(32'hbb03fa8e),
	.w2(32'hb98fa1dc),
	.w3(32'hbaac5334),
	.w4(32'hb9eb45f1),
	.w5(32'h39f50942),
	.w6(32'hbac4ffe9),
	.w7(32'h3a068be7),
	.w8(32'h396e30f5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb380906),
	.w1(32'hb9fee87a),
	.w2(32'hbacd518f),
	.w3(32'hbb123c68),
	.w4(32'h397b349e),
	.w5(32'h392f7719),
	.w6(32'hbac2a66b),
	.w7(32'h39c2479b),
	.w8(32'h3a850ae0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2c8bc),
	.w1(32'hba8abd59),
	.w2(32'hbb12a57c),
	.w3(32'hbaeb4996),
	.w4(32'hb90119b3),
	.w5(32'hb8d4f765),
	.w6(32'h38d1e2e1),
	.w7(32'h3acc3bf3),
	.w8(32'h3adf9aa6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b255a3),
	.w1(32'hb8c354c0),
	.w2(32'hb97af2ac),
	.w3(32'h37a7312e),
	.w4(32'hb7c6156a),
	.w5(32'hb9077d9f),
	.w6(32'h395b8ec9),
	.w7(32'h38e7bf89),
	.w8(32'h35a176af),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381fb918),
	.w1(32'h37423c67),
	.w2(32'h375a36d3),
	.w3(32'h37e39cb2),
	.w4(32'hb7b744a2),
	.w5(32'hb7f00821),
	.w6(32'hb60bb2ac),
	.w7(32'hb82b7716),
	.w8(32'hb7ea0554),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cac8ea),
	.w1(32'h37e5d631),
	.w2(32'h37d59cb7),
	.w3(32'h38a60af9),
	.w4(32'h371b9df6),
	.w5(32'h3851af97),
	.w6(32'h38ed513d),
	.w7(32'hb78d744a),
	.w8(32'hb77372b9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb934057c),
	.w1(32'hb8a5e5bc),
	.w2(32'hb8ac4231),
	.w3(32'hb8612e66),
	.w4(32'h3990f33b),
	.w5(32'h39dadc34),
	.w6(32'h38e95127),
	.w7(32'h3a242d83),
	.w8(32'h3a575dbe),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7def1),
	.w1(32'h3a5394d3),
	.w2(32'h3973f2a0),
	.w3(32'h3aa51f82),
	.w4(32'h3ab0b5f8),
	.w5(32'hba987c5c),
	.w6(32'h3ab0167e),
	.w7(32'h3a288966),
	.w8(32'hba8610bf),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1aa477),
	.w1(32'h39397510),
	.w2(32'hb9d18111),
	.w3(32'h3a1b65de),
	.w4(32'h3a92139e),
	.w5(32'hb9e6da8e),
	.w6(32'h3a5cfd82),
	.w7(32'h3a3dfdad),
	.w8(32'hba1d10cc),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90eb9e0),
	.w1(32'h3a0cedd2),
	.w2(32'h3785df46),
	.w3(32'h3a735099),
	.w4(32'h3ad539cd),
	.w5(32'hb9e115bd),
	.w6(32'h3a9b514c),
	.w7(32'h3a8548a3),
	.w8(32'hba24582e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26e325),
	.w1(32'h386354aa),
	.w2(32'hba5fb45c),
	.w3(32'hb77bbec9),
	.w4(32'h3a2f130a),
	.w5(32'hb900a534),
	.w6(32'h3a0ce44a),
	.w7(32'h3aa0c440),
	.w8(32'h39b5c692),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a0246),
	.w1(32'h39d1d6a3),
	.w2(32'h3a8543b3),
	.w3(32'h3ab87c65),
	.w4(32'h3a99df28),
	.w5(32'hb9b9e871),
	.w6(32'h3a17123c),
	.w7(32'hb8b4e222),
	.w8(32'hb9d9436a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a3a3ee),
	.w1(32'h36a7fe82),
	.w2(32'hb7e82d2b),
	.w3(32'hb829a13a),
	.w4(32'h382853b3),
	.w5(32'hb7e37f16),
	.w6(32'h371dd9cd),
	.w7(32'hb6aa60bf),
	.w8(32'hb839fc7c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8be7ecc),
	.w1(32'hb84c8b83),
	.w2(32'hb907da6b),
	.w3(32'h3a188245),
	.w4(32'h390d73fa),
	.w5(32'hb98d5dcc),
	.w6(32'h39d69726),
	.w7(32'hb91d7a21),
	.w8(32'hba0d6704),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce0a0f),
	.w1(32'hb8cb14b1),
	.w2(32'hb7d0c572),
	.w3(32'h38b63584),
	.w4(32'hb8e6a088),
	.w5(32'hb8737923),
	.w6(32'h38ba883d),
	.w7(32'hb7564920),
	.w8(32'hb8036c0b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39374f18),
	.w1(32'h3a0dd87b),
	.w2(32'h3a028a9c),
	.w3(32'h3a9612d3),
	.w4(32'h3a7b432e),
	.w5(32'h3a1c4f5c),
	.w6(32'h3a1051d1),
	.w7(32'h3a4a7eff),
	.w8(32'h38c314a2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9097492),
	.w1(32'hb931995d),
	.w2(32'hb9b04654),
	.w3(32'hb6f556ae),
	.w4(32'h3805fd4b),
	.w5(32'hb93890a7),
	.w6(32'h39818732),
	.w7(32'h393eb8a4),
	.w8(32'h3844958f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f038a),
	.w1(32'hbb0fe7d4),
	.w2(32'hbacbc8ad),
	.w3(32'h3a4115b0),
	.w4(32'hb9ff13c3),
	.w5(32'hbb233c88),
	.w6(32'h3adbffee),
	.w7(32'hb92464e9),
	.w8(32'hbac164cc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cff439),
	.w1(32'hb9de92de),
	.w2(32'hba0fa1a0),
	.w3(32'hb9aec20e),
	.w4(32'hb98aea23),
	.w5(32'hb9ca387d),
	.w6(32'h37a63310),
	.w7(32'hb8e82633),
	.w8(32'h3912ffa3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c9bb0),
	.w1(32'h3951cdc1),
	.w2(32'h394b43b1),
	.w3(32'h392a51e3),
	.w4(32'h39489225),
	.w5(32'h388db576),
	.w6(32'h389d2406),
	.w7(32'h38a99285),
	.w8(32'h36b60989),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3701d62b),
	.w1(32'h36cd4284),
	.w2(32'h370a5bc0),
	.w3(32'hb633f5cd),
	.w4(32'h369ae423),
	.w5(32'h370b13ff),
	.w6(32'h36100793),
	.w7(32'hb609c16a),
	.w8(32'hb5adff29),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ac4f99),
	.w1(32'hb87cc1ba),
	.w2(32'hb85ca877),
	.w3(32'hb87bc130),
	.w4(32'hb767e908),
	.w5(32'hb866b9f3),
	.w6(32'hb874c891),
	.w7(32'hb75b2991),
	.w8(32'hb887bf91),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88511c9),
	.w1(32'h394d20c7),
	.w2(32'h38d8fb78),
	.w3(32'hb8bf0448),
	.w4(32'h395e806f),
	.w5(32'h3900a67c),
	.w6(32'hb818934d),
	.w7(32'h39411e6e),
	.w8(32'h392f6e77),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81367da),
	.w1(32'h37e60603),
	.w2(32'hb87541c6),
	.w3(32'h3772ced9),
	.w4(32'h371d8a02),
	.w5(32'hb9817165),
	.w6(32'h37c1635f),
	.w7(32'hb8cb8e6a),
	.w8(32'hb8f05b65),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a88bdc),
	.w1(32'hb838c6b9),
	.w2(32'hb81664b0),
	.w3(32'h39860a3d),
	.w4(32'hb954312c),
	.w5(32'hb9b2a411),
	.w6(32'h39bf8bd3),
	.w7(32'hb8cee5cb),
	.w8(32'hb9808a01),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba437855),
	.w1(32'h3814220e),
	.w2(32'h3a629bc2),
	.w3(32'hb9c60f16),
	.w4(32'h39008dc1),
	.w5(32'h3a1b3c82),
	.w6(32'hb9a404e6),
	.w7(32'h3a03ac25),
	.w8(32'h3a18f18e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b14083),
	.w1(32'h359b86a9),
	.w2(32'h366c2ea2),
	.w3(32'h378832bb),
	.w4(32'hb6ac5d7c),
	.w5(32'hb68459cf),
	.w6(32'h370f059d),
	.w7(32'hb7358b6b),
	.w8(32'hb6342f0b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3776b588),
	.w1(32'hb30bbcd6),
	.w2(32'hb6a49f66),
	.w3(32'h379bf623),
	.w4(32'hb6b57c6c),
	.w5(32'hb73284b7),
	.w6(32'h366d3c47),
	.w7(32'hb72e7a72),
	.w8(32'hb7584a0a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7282159),
	.w1(32'hb7ef5e21),
	.w2(32'hb7471e25),
	.w3(32'h37935486),
	.w4(32'hb739d89d),
	.w5(32'h36b87cd5),
	.w6(32'hb63a0728),
	.w7(32'hb7a43fb3),
	.w8(32'hb769dbfe),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370fac32),
	.w1(32'hb78960d6),
	.w2(32'h362b1342),
	.w3(32'hb64d3761),
	.w4(32'hb7cbcf01),
	.w5(32'h3731e356),
	.w6(32'h368920eb),
	.w7(32'hb734a96a),
	.w8(32'h3730fff7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabadec),
	.w1(32'hb9f61528),
	.w2(32'h3a46ea25),
	.w3(32'hba77a1b4),
	.w4(32'hba31825f),
	.w5(32'hb98562af),
	.w6(32'hba7cff3f),
	.w7(32'hb9bbc0ed),
	.w8(32'h38e22b32),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab958fb),
	.w1(32'hba8c35da),
	.w2(32'hbaf40663),
	.w3(32'hba27f978),
	.w4(32'h37a43c69),
	.w5(32'hba82bbcb),
	.w6(32'h39bebcd9),
	.w7(32'h3a3b5298),
	.w8(32'h3a0b3049),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15b86e),
	.w1(32'hbac47ea0),
	.w2(32'hbab30ee7),
	.w3(32'hbaced210),
	.w4(32'hba87ea74),
	.w5(32'hb9f85651),
	.w6(32'hb9cd391f),
	.w7(32'h39a44f0f),
	.w8(32'h3a6fce53),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb537b5b),
	.w1(32'hbb3938c5),
	.w2(32'hbb81392c),
	.w3(32'hba1ed1d6),
	.w4(32'hba800e7d),
	.w5(32'hbaf888df),
	.w6(32'h3a1ae031),
	.w7(32'h3a0e3463),
	.w8(32'hba722f77),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c7be51),
	.w1(32'h376c27c6),
	.w2(32'h3801496b),
	.w3(32'h37b31ef0),
	.w4(32'h341ad82f),
	.w5(32'h379bebef),
	.w6(32'h358a0870),
	.w7(32'hb779d20d),
	.w8(32'h351eea91),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383a2930),
	.w1(32'h37ce95e3),
	.w2(32'h384df77f),
	.w3(32'h37ad502d),
	.w4(32'hb494eb85),
	.w5(32'h3808cefb),
	.w6(32'h3694e064),
	.w7(32'hb7b68b91),
	.w8(32'h371738b2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3882348f),
	.w1(32'h387fc809),
	.w2(32'h389504e3),
	.w3(32'h3866861b),
	.w4(32'h3788f3f2),
	.w5(32'h378b8376),
	.w6(32'h37be1c1f),
	.w7(32'hb81fc459),
	.w8(32'hb803f4a7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d352c),
	.w1(32'hba42f4ab),
	.w2(32'hba5af020),
	.w3(32'hb935d15f),
	.w4(32'hb9c0b69d),
	.w5(32'hba59641e),
	.w6(32'h38956ad8),
	.w7(32'hb98f48ce),
	.w8(32'hba2056ae),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386a7633),
	.w1(32'h37de45a4),
	.w2(32'h341badfe),
	.w3(32'h38509e4b),
	.w4(32'h37c55ec5),
	.w5(32'h37be73d9),
	.w6(32'h38683899),
	.w7(32'h36164582),
	.w8(32'hb748ffcf),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2c5df),
	.w1(32'hba2bc686),
	.w2(32'hb9cece2d),
	.w3(32'hb8b76477),
	.w4(32'hb9c298fa),
	.w5(32'hba1b1f75),
	.w6(32'hb98ce110),
	.w7(32'hb9e5824f),
	.w8(32'hba0be4ef),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3634a6),
	.w1(32'hb9dc46bb),
	.w2(32'hba46a0e6),
	.w3(32'hb99a65e5),
	.w4(32'hbab5ce59),
	.w5(32'hbabc5c3b),
	.w6(32'hb9edb23e),
	.w7(32'hba7541a2),
	.w8(32'hb9bcc475),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1197b8),
	.w1(32'h3a5456f3),
	.w2(32'h3a664de3),
	.w3(32'h3a6b476c),
	.w4(32'h3aa1331b),
	.w5(32'h39c2fade),
	.w6(32'h3a1412f5),
	.w7(32'h3a361a0a),
	.w8(32'h386fe162),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb8d4d),
	.w1(32'hbabd5557),
	.w2(32'hbad11df5),
	.w3(32'hb9a72a4a),
	.w4(32'hba498946),
	.w5(32'hbaad7922),
	.w6(32'h39432fbd),
	.w7(32'hb8c4ca8d),
	.w8(32'hba8004e3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e4ad1),
	.w1(32'hba0baf0a),
	.w2(32'hb83eac5e),
	.w3(32'h384885ac),
	.w4(32'hb91fae7e),
	.w5(32'hb9a1f085),
	.w6(32'hb9bd57a1),
	.w7(32'hb9834855),
	.w8(32'hb990e07a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901face),
	.w1(32'h39fbb52d),
	.w2(32'h395075c7),
	.w3(32'h3a1e225d),
	.w4(32'h3a4e22a8),
	.w5(32'h38c2bc96),
	.w6(32'h39db4ae4),
	.w7(32'h39e7913c),
	.w8(32'hb8e614cf),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88aeaab),
	.w1(32'hb8cfafdf),
	.w2(32'h397adcd4),
	.w3(32'hb8742079),
	.w4(32'h39564839),
	.w5(32'hb990d32d),
	.w6(32'hb9d53bf9),
	.w7(32'hb96a664b),
	.w8(32'hb9c94ffa),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6eb9055),
	.w1(32'hb6b6a258),
	.w2(32'h36c61597),
	.w3(32'hb70fa8ab),
	.w4(32'hb6ad3128),
	.w5(32'h36cd5b86),
	.w6(32'hb6e0c37a),
	.w7(32'hb64d96fb),
	.w8(32'h36e00c8e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7757379),
	.w1(32'hb7330f1b),
	.w2(32'h363ba9e7),
	.w3(32'h3680e785),
	.w4(32'h36d4446b),
	.w5(32'h376e2de5),
	.w6(32'h370c705d),
	.w7(32'h3787ba82),
	.w8(32'h37c92647),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370bc5a4),
	.w1(32'h35ee1e94),
	.w2(32'h371d7c13),
	.w3(32'h36b54bf3),
	.w4(32'hb6e9156f),
	.w5(32'h36692b75),
	.w6(32'hb60cf551),
	.w7(32'hb6a68e7f),
	.w8(32'hb64d39dc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7341d76),
	.w1(32'hb845b97b),
	.w2(32'hb8e2380d),
	.w3(32'hb7a1bda4),
	.w4(32'hb62cd273),
	.w5(32'hb878260d),
	.w6(32'h368475f5),
	.w7(32'h385af1d2),
	.w8(32'hb798d9d0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdadcd),
	.w1(32'hba78718c),
	.w2(32'hba24ef33),
	.w3(32'hba3a37a7),
	.w4(32'hb98faaed),
	.w5(32'hb83f172b),
	.w6(32'h39cbaa0f),
	.w7(32'h37b2189d),
	.w8(32'hb89ab180),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382f036a),
	.w1(32'h394c75c9),
	.w2(32'h3894a242),
	.w3(32'hb8e195af),
	.w4(32'h39191a90),
	.w5(32'h392711b6),
	.w6(32'hb91ac081),
	.w7(32'h398b551e),
	.w8(32'h39cb1371),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2b7f0),
	.w1(32'hba6c5176),
	.w2(32'hb9c810f6),
	.w3(32'h39088bdf),
	.w4(32'hb89e01c7),
	.w5(32'hba58b24e),
	.w6(32'h3aa6f697),
	.w7(32'h398837b7),
	.w8(32'hba5af6c8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5d2ee),
	.w1(32'hb9bb1553),
	.w2(32'h38c66f6b),
	.w3(32'hb97ac804),
	.w4(32'h38cce8f3),
	.w5(32'h3680424c),
	.w6(32'hb9dfd36a),
	.w7(32'hb71df624),
	.w8(32'h39f16caf),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a9258),
	.w1(32'h38eef3e6),
	.w2(32'hba2ba94f),
	.w3(32'hba836c77),
	.w4(32'h38ccc486),
	.w5(32'hb8f97f77),
	.w6(32'hb8e80cf1),
	.w7(32'h3a22006a),
	.w8(32'h3a020eb4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c8a65),
	.w1(32'hbb45c91e),
	.w2(32'hba81262f),
	.w3(32'hb9e0d319),
	.w4(32'hb8f8237e),
	.w5(32'hba2016e5),
	.w6(32'hba0b1f02),
	.w7(32'h39ee208c),
	.w8(32'hba465e2d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf26dc3),
	.w1(32'hba92cfb6),
	.w2(32'hbacc4a60),
	.w3(32'hbaa99760),
	.w4(32'hb9d6ac24),
	.w5(32'hba2ec091),
	.w6(32'hba4c8e15),
	.w7(32'hb888bacc),
	.w8(32'hb8241d61),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97eb0b),
	.w1(32'hbb958968),
	.w2(32'hbb98b1ce),
	.w3(32'hba38773e),
	.w4(32'hbb14ec42),
	.w5(32'hbb9b1b45),
	.w6(32'h3b0e705c),
	.w7(32'h389b8fdd),
	.w8(32'hbb2ad9d1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c92bd),
	.w1(32'hb909269a),
	.w2(32'h384e08d7),
	.w3(32'h37f9e2a4),
	.w4(32'h3a0dd028),
	.w5(32'hb89fec70),
	.w6(32'h399e98ff),
	.w7(32'h39436cd3),
	.w8(32'hb9a7b455),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba867155),
	.w1(32'hba264408),
	.w2(32'hba86bb3c),
	.w3(32'hb9a22d4e),
	.w4(32'hb925bb1b),
	.w5(32'hba1219b2),
	.w6(32'h399a172a),
	.w7(32'h397b7d58),
	.w8(32'hb8bd6e5d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb725c1a3),
	.w1(32'hb8b5efbd),
	.w2(32'hb7cd118a),
	.w3(32'hb7aa0e9e),
	.w4(32'hb90dcc4c),
	.w5(32'hb9052669),
	.w6(32'hb9206475),
	.w7(32'hb9720625),
	.w8(32'hb8daa4e6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb600d),
	.w1(32'hb922442f),
	.w2(32'hba366c98),
	.w3(32'h3a2983f8),
	.w4(32'h3a8911fa),
	.w5(32'hba969289),
	.w6(32'h3a10f219),
	.w7(32'h3a645d7d),
	.w8(32'hba59b9ef),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb207e98),
	.w1(32'hbb0ecf79),
	.w2(32'hbad725f8),
	.w3(32'hbae0292d),
	.w4(32'hbadec7b0),
	.w5(32'hbad543e9),
	.w6(32'hba10fe61),
	.w7(32'hba570f8b),
	.w8(32'hba53ea91),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1a59d),
	.w1(32'hba909cfe),
	.w2(32'hb948784d),
	.w3(32'hb9a6bfcc),
	.w4(32'hba420101),
	.w5(32'h39774a9f),
	.w6(32'hba9b5fc5),
	.w7(32'h39018b42),
	.w8(32'h3a1beba0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbece3fa),
	.w1(32'hbbc0ca96),
	.w2(32'hbb965b72),
	.w3(32'hbb897089),
	.w4(32'hbae10928),
	.w5(32'hbaa002c0),
	.w6(32'h3a4428a7),
	.w7(32'h3a8112e1),
	.w8(32'hb8dd3dbe),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5042bc),
	.w1(32'h3a975b61),
	.w2(32'h3a81547a),
	.w3(32'h3abcd975),
	.w4(32'h3b0318ff),
	.w5(32'hba275934),
	.w6(32'h3a70d02b),
	.w7(32'h3a128d04),
	.w8(32'hbaa0e45a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32dbbe),
	.w1(32'hbb369be1),
	.w2(32'hbb16fe6d),
	.w3(32'hbaed7fb1),
	.w4(32'hbae79bd8),
	.w5(32'hbb07d3f9),
	.w6(32'hbac3fcf3),
	.w7(32'hba78c30a),
	.w8(32'hbb1f3bdb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd5431),
	.w1(32'hb92a01b9),
	.w2(32'hb771b0d5),
	.w3(32'hb8a74bb9),
	.w4(32'hb80ab84d),
	.w5(32'h3842dc3d),
	.w6(32'h38b57b05),
	.w7(32'h38dc9a19),
	.w8(32'h388afdaf),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a31e4),
	.w1(32'hbb66121d),
	.w2(32'hbb31045c),
	.w3(32'hbabd6666),
	.w4(32'hbb3d5036),
	.w5(32'hbaa3ac5d),
	.w6(32'hb8ab16d6),
	.w7(32'hbab0d17b),
	.w8(32'hbac16953),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f21544),
	.w1(32'hba3acad4),
	.w2(32'hb99e2244),
	.w3(32'hb9f4a328),
	.w4(32'hb900bf99),
	.w5(32'h39a87b5a),
	.w6(32'hba0cb76d),
	.w7(32'hb98751d9),
	.w8(32'h3a270e05),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fc7c40),
	.w1(32'h37cf273b),
	.w2(32'h351c1866),
	.w3(32'h379ee7fa),
	.w4(32'h382737ce),
	.w5(32'h3796dd4c),
	.w6(32'h38ddec1e),
	.w7(32'h38e7432c),
	.w8(32'h38af004d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981ea33),
	.w1(32'hb8970167),
	.w2(32'h39592cbe),
	.w3(32'hb8b7a087),
	.w4(32'hb7e91060),
	.w5(32'h39a8adbc),
	.w6(32'hb9050214),
	.w7(32'h39698275),
	.w8(32'h39be443a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bbcb3),
	.w1(32'h3aae4bac),
	.w2(32'h3a8b43e4),
	.w3(32'h3ac2e275),
	.w4(32'h3af5210a),
	.w5(32'h398fd5c6),
	.w6(32'h3a43a28f),
	.w7(32'h3a35e0d5),
	.w8(32'hba082051),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395aa29c),
	.w1(32'h3a4b28f2),
	.w2(32'h394a40c7),
	.w3(32'h3a5dbcc2),
	.w4(32'h3aa396f2),
	.w5(32'hb91df90c),
	.w6(32'h39b94c3e),
	.w7(32'h3a7b0e3c),
	.w8(32'hb982a97e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3079a),
	.w1(32'hba9a3831),
	.w2(32'hbab8ae5a),
	.w3(32'hba44b223),
	.w4(32'h375b7802),
	.w5(32'hba0182d0),
	.w6(32'h381f82b7),
	.w7(32'h3a34ab95),
	.w8(32'h39504424),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6b6ed),
	.w1(32'hbadadefd),
	.w2(32'hbb00f81d),
	.w3(32'hb99d37c0),
	.w4(32'hba31d295),
	.w5(32'hbabff21d),
	.w6(32'h3a03b77f),
	.w7(32'hb958a418),
	.w8(32'hba98822a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f338f2),
	.w1(32'hb99d8d7e),
	.w2(32'hb9488022),
	.w3(32'h39b0be26),
	.w4(32'h388b0b79),
	.w5(32'h3a089897),
	.w6(32'h3984264b),
	.w7(32'h3a316952),
	.w8(32'h3abf4f3c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3726601c),
	.w1(32'h3a8db15c),
	.w2(32'h3addf502),
	.w3(32'h39ea38a4),
	.w4(32'h3a537f35),
	.w5(32'h3a0414e0),
	.w6(32'h3a9aa2d8),
	.w7(32'h3a2b744f),
	.w8(32'h3a09d2ed),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6cf2b),
	.w1(32'h38a76dc6),
	.w2(32'h3935c852),
	.w3(32'h39bce071),
	.w4(32'h3a0f9a16),
	.w5(32'hba0d1c66),
	.w6(32'h3a1bab54),
	.w7(32'h3a033a7e),
	.w8(32'hb9dc4627),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80ed631),
	.w1(32'hb80d193b),
	.w2(32'hb72d039b),
	.w3(32'hb8384917),
	.w4(32'hb805dce3),
	.w5(32'hb6c51e8c),
	.w6(32'hb7ec1ed2),
	.w7(32'hb7f888a0),
	.w8(32'hb7511636),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89ba6a1),
	.w1(32'h37af3996),
	.w2(32'h3915cb02),
	.w3(32'h3850ab2b),
	.w4(32'h378a49dd),
	.w5(32'h39177947),
	.w6(32'h388b76c2),
	.w7(32'h38504aca),
	.w8(32'h38dcb771),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h351383fb),
	.w1(32'h36a85f4b),
	.w2(32'h37160558),
	.w3(32'h36fa26df),
	.w4(32'h36fe72b7),
	.w5(32'h371bd596),
	.w6(32'hb6a2267a),
	.w7(32'hb6b2e5f3),
	.w8(32'h34ad4a5d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9927353),
	.w1(32'hb9c14254),
	.w2(32'hb9aa93ae),
	.w3(32'hb90d338e),
	.w4(32'hb94ac908),
	.w5(32'hb934260f),
	.w6(32'h379f63eb),
	.w7(32'hb92d3eeb),
	.w8(32'hb9355748),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ad555),
	.w1(32'h3946951b),
	.w2(32'h38ab87cf),
	.w3(32'h3a0fcf31),
	.w4(32'h3a75fddc),
	.w5(32'h382f624f),
	.w6(32'h3a305c85),
	.w7(32'h3a0fb74f),
	.w8(32'hb8ef5fab),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84f852),
	.w1(32'hba9b022e),
	.w2(32'hba6674f2),
	.w3(32'hb967c762),
	.w4(32'hba1bf027),
	.w5(32'hba466268),
	.w6(32'h398594d3),
	.w7(32'hb9dd3ab4),
	.w8(32'hba72cf4f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c91a15),
	.w1(32'hb9e7f868),
	.w2(32'hb90cd6a4),
	.w3(32'hb9784d75),
	.w4(32'hb87e7912),
	.w5(32'hb9f13630),
	.w6(32'hb9b1ec14),
	.w7(32'hb939ad34),
	.w8(32'hb9e29c45),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6cb202),
	.w1(32'hb9a5bf2a),
	.w2(32'hb961f9a5),
	.w3(32'hb9ca9c7d),
	.w4(32'h390df9d9),
	.w5(32'h3a220a30),
	.w6(32'h37f65633),
	.w7(32'h3a2c41e2),
	.w8(32'h3a6f40a8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3786b164),
	.w1(32'h37032710),
	.w2(32'h37aee02b),
	.w3(32'h3760b9ad),
	.w4(32'h3678357b),
	.w5(32'h37af1946),
	.w6(32'h370e6bd4),
	.w7(32'hb6f7e59f),
	.w8(32'h37274f3c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bb21c6),
	.w1(32'h390dab04),
	.w2(32'h38bdb8d8),
	.w3(32'hb81125a0),
	.w4(32'h38b6f645),
	.w5(32'h39438057),
	.w6(32'h38140701),
	.w7(32'h395a473f),
	.w8(32'h3978e896),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36827ad9),
	.w1(32'hb6c854e3),
	.w2(32'h37621e99),
	.w3(32'hb4873a27),
	.w4(32'hb66cccf7),
	.w5(32'h37989ed4),
	.w6(32'h36b907a9),
	.w7(32'hb616b637),
	.w8(32'h379e534e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f12fa),
	.w1(32'h3a59c5ba),
	.w2(32'h3a151ce0),
	.w3(32'hb9856cef),
	.w4(32'hbac126bf),
	.w5(32'hb899cf6e),
	.w6(32'hba901bd4),
	.w7(32'h3a96cb60),
	.w8(32'hb70ad8e0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab32ade),
	.w1(32'h398829dc),
	.w2(32'h3a8f3dae),
	.w3(32'h3a3f5cdf),
	.w4(32'hb924ac51),
	.w5(32'hb9cfcc9d),
	.w6(32'hbaa60328),
	.w7(32'hba1e7905),
	.w8(32'hb8ffeb87),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4721c6),
	.w1(32'h3a8310c7),
	.w2(32'hbb9a2f5b),
	.w3(32'h3af9fa74),
	.w4(32'h3af9b4d4),
	.w5(32'hbb81f588),
	.w6(32'hbaff1385),
	.w7(32'hbafcb4bc),
	.w8(32'hbab28bb0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8c01e),
	.w1(32'hb9e04d63),
	.w2(32'hb815733b),
	.w3(32'h3a10afbb),
	.w4(32'hb9747ce0),
	.w5(32'hba4ad0f1),
	.w6(32'h38554527),
	.w7(32'hba0cc3c0),
	.w8(32'hb9e0a668),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa8699),
	.w1(32'hb9935390),
	.w2(32'h3b45b79e),
	.w3(32'hbaa6f243),
	.w4(32'h38b46ecb),
	.w5(32'h3a3429fe),
	.w6(32'hba28de68),
	.w7(32'hb9b9a4f5),
	.w8(32'h370b7208),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb359acf),
	.w1(32'h3b848516),
	.w2(32'h39b4913c),
	.w3(32'h39a565b2),
	.w4(32'h3b6ea932),
	.w5(32'h3b7d738d),
	.w6(32'h3a320809),
	.w7(32'hbaa17a15),
	.w8(32'hbb422ec1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d479e),
	.w1(32'hbaff831d),
	.w2(32'hbaec1a45),
	.w3(32'h3a080f54),
	.w4(32'hb9b78c28),
	.w5(32'hbb640265),
	.w6(32'hba19069b),
	.w7(32'h38ae0e1a),
	.w8(32'hb8dd9c83),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39199132),
	.w1(32'hba40f4f2),
	.w2(32'h399b764b),
	.w3(32'hb9bc418a),
	.w4(32'hbb27ccf0),
	.w5(32'hbab8f6ed),
	.w6(32'h3a237f66),
	.w7(32'h3aa64154),
	.w8(32'hb7d9c812),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385bd425),
	.w1(32'hb9ccc74e),
	.w2(32'h3a4f1094),
	.w3(32'h3a4389d8),
	.w4(32'hba7bfe6f),
	.w5(32'hbac51d42),
	.w6(32'h3a4e8ceb),
	.w7(32'h39f0b67e),
	.w8(32'hba0019ad),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24b27d),
	.w1(32'hba01b171),
	.w2(32'hba0bb824),
	.w3(32'hbae8f63c),
	.w4(32'h38b3c7d6),
	.w5(32'h3803c83b),
	.w6(32'hbac8ac46),
	.w7(32'hba67a614),
	.w8(32'hba93f118),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba113219),
	.w1(32'hb979e73f),
	.w2(32'h3ab314ab),
	.w3(32'h3a1535c5),
	.w4(32'hb9c2e647),
	.w5(32'h393a7b05),
	.w6(32'h3a75ba1a),
	.w7(32'h3ae375aa),
	.w8(32'h3a0b8755),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbe125),
	.w1(32'hba9d8713),
	.w2(32'hbaffaf8c),
	.w3(32'hba1de7bd),
	.w4(32'hbb1f71e3),
	.w5(32'hbb69b339),
	.w6(32'h3a10e813),
	.w7(32'h39ce3d7e),
	.w8(32'hbab9f5e8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31bf8d),
	.w1(32'hbaac529f),
	.w2(32'hb9f7197d),
	.w3(32'hbb01a7de),
	.w4(32'hbb6471b6),
	.w5(32'hbb0e2d51),
	.w6(32'h3bade944),
	.w7(32'h3b5c0491),
	.w8(32'h3b3a0814),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a0929),
	.w1(32'hbaa58152),
	.w2(32'h3aa80a52),
	.w3(32'hbb3a8fa3),
	.w4(32'h3985b612),
	.w5(32'h3a677570),
	.w6(32'hbaf1cf59),
	.w7(32'hbacab408),
	.w8(32'hbafc782c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39725851),
	.w1(32'h39a521fa),
	.w2(32'h3a6a8b25),
	.w3(32'h3ac3d5b5),
	.w4(32'hb9ad3510),
	.w5(32'h3a835d8d),
	.w6(32'hba4fea09),
	.w7(32'h39085e96),
	.w8(32'h3a9639d8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39831ce9),
	.w1(32'hbb34ad5a),
	.w2(32'hba3d53de),
	.w3(32'h3a6a67b9),
	.w4(32'hba796a75),
	.w5(32'hb9ae8344),
	.w6(32'hbb84f479),
	.w7(32'hbafa6286),
	.w8(32'hba9be378),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d8feb),
	.w1(32'hb800e25a),
	.w2(32'hba9316cf),
	.w3(32'h3aca492d),
	.w4(32'h3a38e7bc),
	.w5(32'hbac83bae),
	.w6(32'hbadf72af),
	.w7(32'hbb285ef2),
	.w8(32'hba9e9604),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7db4e8),
	.w1(32'h396f8f6e),
	.w2(32'h39e57ea5),
	.w3(32'hba91732e),
	.w4(32'hb9f8d45b),
	.w5(32'hba1455c0),
	.w6(32'h3a135f6c),
	.w7(32'h3a603d23),
	.w8(32'h3a535f6d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f182de),
	.w1(32'hbb623f90),
	.w2(32'h3b732a51),
	.w3(32'hb92be77f),
	.w4(32'hbb15998d),
	.w5(32'hba2708cb),
	.w6(32'hbb587c2a),
	.w7(32'h3afc0bc9),
	.w8(32'hbaa2d411),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce4604),
	.w1(32'h3a57a01b),
	.w2(32'h3b1bd397),
	.w3(32'hbb28bf0e),
	.w4(32'hba052fca),
	.w5(32'h3ab07a63),
	.w6(32'h3a380f1d),
	.w7(32'h3abb968e),
	.w8(32'hb9c3322f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb489751),
	.w1(32'hba4da9ef),
	.w2(32'h3a3a40c1),
	.w3(32'hbb2018e9),
	.w4(32'hba250957),
	.w5(32'h38fec026),
	.w6(32'h392a98c3),
	.w7(32'h3a4f6896),
	.w8(32'hb9572328),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba901200),
	.w1(32'h394de0bb),
	.w2(32'h3a17191d),
	.w3(32'h3a1cda2e),
	.w4(32'h3a19dd3b),
	.w5(32'hba4c7d19),
	.w6(32'h3acc9f6b),
	.w7(32'h3a88ecfe),
	.w8(32'hbad2734d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bbd13),
	.w1(32'hba313409),
	.w2(32'hba976fce),
	.w3(32'h39facb0a),
	.w4(32'hbabfab26),
	.w5(32'hbac928c0),
	.w6(32'hbb3ec626),
	.w7(32'hba6c1516),
	.w8(32'hb93615d2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb168d8b),
	.w1(32'hbb0c6f30),
	.w2(32'h3ac634c2),
	.w3(32'h38bd69a2),
	.w4(32'hba0ed4bf),
	.w5(32'h3aeef60e),
	.w6(32'hb8ab14c9),
	.w7(32'hbb44cd6d),
	.w8(32'hbb42411b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09471d),
	.w1(32'h3b8ca5d5),
	.w2(32'h3b205c43),
	.w3(32'hbaeaa627),
	.w4(32'hba87c431),
	.w5(32'hbb8c7f4c),
	.w6(32'h3b9a7043),
	.w7(32'h3bbecf5c),
	.w8(32'h3b25abc8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf49c0a),
	.w1(32'hb7cb360c),
	.w2(32'h3a3ec88a),
	.w3(32'hbb0ae79b),
	.w4(32'h39a743e7),
	.w5(32'hb9e37995),
	.w6(32'hbab78f92),
	.w7(32'hb9f6d691),
	.w8(32'hba3637a5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9163a55),
	.w1(32'h373b3e74),
	.w2(32'hba94ed3c),
	.w3(32'h3a3d12f3),
	.w4(32'hbaa788da),
	.w5(32'hba7612e4),
	.w6(32'h3a5426b2),
	.w7(32'h3ae89629),
	.w8(32'h3a4a6122),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43e92e),
	.w1(32'hbb9cb9c0),
	.w2(32'hbb154df5),
	.w3(32'h39dcf396),
	.w4(32'hbab3e5ec),
	.w5(32'hbb44e3ef),
	.w6(32'hbbc09e5b),
	.w7(32'hbb02b307),
	.w8(32'hbb5d30a4),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb878c73),
	.w1(32'h3afff020),
	.w2(32'h3b017d7a),
	.w3(32'h37f6bfe2),
	.w4(32'h3b0104b3),
	.w5(32'h3a67f51f),
	.w6(32'h3ab5919f),
	.w7(32'h3a6625df),
	.w8(32'h3a8e55b5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0b04d),
	.w1(32'h39fbf3f7),
	.w2(32'hbb00e195),
	.w3(32'h3acf7fbd),
	.w4(32'h3aa5e800),
	.w5(32'hb8d72338),
	.w6(32'hba87f7a5),
	.w7(32'hba9bcd24),
	.w8(32'hba65f1e2),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e747f),
	.w1(32'hbbb23994),
	.w2(32'h3a6e2fa0),
	.w3(32'hba8ada88),
	.w4(32'hbbd9a96e),
	.w5(32'hb870cfd3),
	.w6(32'h394dbf3e),
	.w7(32'h3b65fded),
	.w8(32'h39e20756),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c38f3),
	.w1(32'hba584552),
	.w2(32'hbb2b0d54),
	.w3(32'hbb11101b),
	.w4(32'hba7151d0),
	.w5(32'hbba230ad),
	.w6(32'hbaaddda7),
	.w7(32'hbaaa511c),
	.w8(32'h3b0eb263),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66f145),
	.w1(32'h38fa3b4f),
	.w2(32'hb9b02163),
	.w3(32'h3a8ef0ff),
	.w4(32'hb99ee1d3),
	.w5(32'hb963e8ac),
	.w6(32'hb9ea3c59),
	.w7(32'hba0101b7),
	.w8(32'hb9bc65d6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9844fe3),
	.w1(32'h3ab7fe62),
	.w2(32'h3abab2cc),
	.w3(32'hb903e900),
	.w4(32'h3a10e2f2),
	.w5(32'h39ed9b5a),
	.w6(32'hba1fd654),
	.w7(32'h3a558be7),
	.w8(32'h3a20cd1c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396789de),
	.w1(32'h39804a5c),
	.w2(32'h3b8ffd09),
	.w3(32'h3a41a571),
	.w4(32'h3aaa9564),
	.w5(32'h3abf7dd5),
	.w6(32'h3a14b15f),
	.w7(32'h3b7f6a5e),
	.w8(32'h3783e6d8),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11340b),
	.w1(32'h3bbebea5),
	.w2(32'h3b5b9ac3),
	.w3(32'h3b02bf7d),
	.w4(32'h3c14828e),
	.w5(32'h39922f2f),
	.w6(32'h3bbcdb21),
	.w7(32'h3be19987),
	.w8(32'hba84d8f0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2b112),
	.w1(32'h39c1ea1e),
	.w2(32'hba883f15),
	.w3(32'hbae08bf8),
	.w4(32'hb94c7746),
	.w5(32'hba62af50),
	.w6(32'h3ad1db48),
	.w7(32'h3aa93d6a),
	.w8(32'hbad2a508),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb676561),
	.w1(32'h3afe0c6a),
	.w2(32'h3b1254f2),
	.w3(32'hbb0d5904),
	.w4(32'h3aaffaba),
	.w5(32'h3a00f9c8),
	.w6(32'h3aad7d3a),
	.w7(32'h3a931377),
	.w8(32'h3a36f39d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7426d5),
	.w1(32'hb9df9e34),
	.w2(32'hb96092bc),
	.w3(32'h3a4cd044),
	.w4(32'hb9bb0c7e),
	.w5(32'h39c6e39e),
	.w6(32'h398a8c58),
	.w7(32'hb8b85ab9),
	.w8(32'hba8548b9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb401466),
	.w1(32'h3a8e5583),
	.w2(32'h3b00db24),
	.w3(32'hbb14b59c),
	.w4(32'h3a03c46b),
	.w5(32'hb9b50abd),
	.w6(32'h3adea584),
	.w7(32'h3b014097),
	.w8(32'h3a44dbbd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51d15d),
	.w1(32'h3919f891),
	.w2(32'hb969167e),
	.w3(32'hba8ab510),
	.w4(32'hb6982ac9),
	.w5(32'hb9e454e2),
	.w6(32'hba328aaa),
	.w7(32'hba838d41),
	.w8(32'hba515388),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba524e84),
	.w1(32'hba4f25d7),
	.w2(32'hbafcf232),
	.w3(32'hb7fa25b9),
	.w4(32'h399826e5),
	.w5(32'hba596f73),
	.w6(32'h39784f50),
	.w7(32'h392c1f48),
	.w8(32'hb9999faf),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba888f5d),
	.w1(32'h3b93cac4),
	.w2(32'hbc0b5ebc),
	.w3(32'hb993091a),
	.w4(32'h3bc193a7),
	.w5(32'hbc73a74f),
	.w6(32'h3bd89376),
	.w7(32'hbad052f6),
	.w8(32'hb8db700f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdd307),
	.w1(32'hbacb2aa1),
	.w2(32'hba4f5630),
	.w3(32'hb9282ffd),
	.w4(32'hba22b768),
	.w5(32'hba09dce3),
	.w6(32'hb91ff009),
	.w7(32'hbb1a85a6),
	.w8(32'hba831bad),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b83856),
	.w1(32'h3a5f4e26),
	.w2(32'h3b2aa299),
	.w3(32'hba1f5734),
	.w4(32'h3a9e2368),
	.w5(32'h3a88b028),
	.w6(32'hb8ef2b2a),
	.w7(32'h3abb958e),
	.w8(32'h3a3ce743),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c23a6a),
	.w1(32'h3a010ff6),
	.w2(32'hb9a47f5d),
	.w3(32'h3a92d577),
	.w4(32'hbae14777),
	.w5(32'hbb7512d5),
	.w6(32'h3b339ae5),
	.w7(32'h3a622f44),
	.w8(32'hbac403e2),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f8816),
	.w1(32'hbafe8e0f),
	.w2(32'h37536530),
	.w3(32'hbb860937),
	.w4(32'hbb24e91c),
	.w5(32'hbb3c0938),
	.w6(32'hba83f0b1),
	.w7(32'h3b174930),
	.w8(32'hb97a21b3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ac568),
	.w1(32'hbb249648),
	.w2(32'hbb22c9e6),
	.w3(32'hbb8b7b74),
	.w4(32'hbb560546),
	.w5(32'hbb0ca392),
	.w6(32'h3951a0d2),
	.w7(32'hbac13f2d),
	.w8(32'hbaa9a51b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa5629),
	.w1(32'h3b373a55),
	.w2(32'h3b31cef9),
	.w3(32'hb92dcd6d),
	.w4(32'h3bb95daf),
	.w5(32'h3b59bd09),
	.w6(32'h3b0f5829),
	.w7(32'hbad32549),
	.w8(32'hbb1f6dbc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae77d41),
	.w1(32'h3ba070b7),
	.w2(32'h3c6648d5),
	.w3(32'hbaf5a592),
	.w4(32'h3b0ffa0f),
	.w5(32'h3c227931),
	.w6(32'h3b8dc33e),
	.w7(32'h3c705c94),
	.w8(32'h3ba27294),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb9cc5),
	.w1(32'h3a1855ee),
	.w2(32'h3b085235),
	.w3(32'hbb4a7ca7),
	.w4(32'h3735268f),
	.w5(32'hb9dfeb56),
	.w6(32'h39df416b),
	.w7(32'h3a81d2e6),
	.w8(32'h386884e7),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67d395),
	.w1(32'hba8535ab),
	.w2(32'hba774086),
	.w3(32'h3ab9bed3),
	.w4(32'hb9c7f4c2),
	.w5(32'hb95fb119),
	.w6(32'hbb224128),
	.w7(32'hbb0f194f),
	.w8(32'hba80837e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37636676),
	.w1(32'h3959d63a),
	.w2(32'hb98d4f61),
	.w3(32'h3a84d13c),
	.w4(32'hb8868fd6),
	.w5(32'hba6a6ae2),
	.w6(32'hb9ff9136),
	.w7(32'h399e0316),
	.w8(32'h3a89d81c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bd5e0),
	.w1(32'h3ab86712),
	.w2(32'hbb631b0f),
	.w3(32'h39c77f7a),
	.w4(32'h3b1f17c8),
	.w5(32'hbb4c1d39),
	.w6(32'hb999b8e2),
	.w7(32'h3aae5138),
	.w8(32'hbad66fc0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05054e),
	.w1(32'hba21775c),
	.w2(32'hba899273),
	.w3(32'h3b1859f0),
	.w4(32'hbac1292b),
	.w5(32'hbb6b1294),
	.w6(32'h3ae5cad3),
	.w7(32'h3a1d3720),
	.w8(32'h3a82ea83),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bb2e2),
	.w1(32'hbaaa6ba3),
	.w2(32'h3a989444),
	.w3(32'hbb09ac78),
	.w4(32'hbb017428),
	.w5(32'hbb201e9e),
	.w6(32'hb955e7e7),
	.w7(32'h3a9bfe7b),
	.w8(32'hba846a7d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a9b7d0),
	.w1(32'hbb147ce6),
	.w2(32'hb934caf5),
	.w3(32'hba6465ce),
	.w4(32'hbb130e8a),
	.w5(32'hbb6a07bd),
	.w6(32'hbaa7750c),
	.w7(32'h34823500),
	.w8(32'h38306ab4),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a60e9),
	.w1(32'hbb76b2ff),
	.w2(32'hbb99eae0),
	.w3(32'hba7c43c7),
	.w4(32'hbb5dbd5e),
	.w5(32'hbb82039b),
	.w6(32'hbaeb395a),
	.w7(32'hbb55cc28),
	.w8(32'hba4d4c0e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe5b94),
	.w1(32'hbb1f2f35),
	.w2(32'hbb5ba503),
	.w3(32'hbb0448ef),
	.w4(32'hbac99520),
	.w5(32'hbba85be0),
	.w6(32'h3a905949),
	.w7(32'h397a356f),
	.w8(32'h3b1b40cd),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4778fc),
	.w1(32'hba974305),
	.w2(32'hbb4e22d7),
	.w3(32'hbaf744c2),
	.w4(32'hbb64865f),
	.w5(32'hbb3d9a5d),
	.w6(32'hba8efcc9),
	.w7(32'hbb3ed839),
	.w8(32'hbb2583fa),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bedf1),
	.w1(32'h3a3511c4),
	.w2(32'h3a957ad9),
	.w3(32'h395ef0e9),
	.w4(32'h3a1ac982),
	.w5(32'h391e3903),
	.w6(32'h3a3820f3),
	.w7(32'h38fdbcf6),
	.w8(32'h39a7a705),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad76438),
	.w1(32'h3b171e9b),
	.w2(32'h3ad5c3b9),
	.w3(32'h3b5526c2),
	.w4(32'h3b3b079d),
	.w5(32'h3a10334c),
	.w6(32'h39f31ecf),
	.w7(32'hb9dba289),
	.w8(32'hba1c29e9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d797b),
	.w1(32'hbaf3aeab),
	.w2(32'hbb0f6412),
	.w3(32'hb88398bf),
	.w4(32'hba7479bf),
	.w5(32'hbb169990),
	.w6(32'hba01bc4d),
	.w7(32'h39ef99ed),
	.w8(32'hb9edb313),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94211a0),
	.w1(32'hbae996ef),
	.w2(32'hbaffe68c),
	.w3(32'hba015320),
	.w4(32'hb9a56222),
	.w5(32'hba571dac),
	.w6(32'hbb008377),
	.w7(32'hbb15bb4c),
	.w8(32'hba86204c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba215b7a),
	.w1(32'h3a4bb8e5),
	.w2(32'h39ca616d),
	.w3(32'hb9ce54a8),
	.w4(32'hbae638d5),
	.w5(32'hbb258035),
	.w6(32'h3a9e50d6),
	.w7(32'h3b4f83a5),
	.w8(32'h3a464b35),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7eed621),
	.w1(32'h3971d98f),
	.w2(32'hb8736671),
	.w3(32'hbb12344a),
	.w4(32'hbaac4627),
	.w5(32'hbb04adad),
	.w6(32'h3adad3ad),
	.w7(32'h3a5c8855),
	.w8(32'hb9fb75b6),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8b3a4),
	.w1(32'h38ac586f),
	.w2(32'h3ad9a8c7),
	.w3(32'hbb0d5079),
	.w4(32'hba4f25c9),
	.w5(32'h3a9b06b3),
	.w6(32'hb94b00b0),
	.w7(32'h39f5bcb7),
	.w8(32'h3a7605f3),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dfd89),
	.w1(32'hbab2290e),
	.w2(32'hba342289),
	.w3(32'hb91f0f59),
	.w4(32'hbb1efbfc),
	.w5(32'hba54a98d),
	.w6(32'hba09dff1),
	.w7(32'hb9575a57),
	.w8(32'hbafaa7ff),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d2205),
	.w1(32'h3a940c31),
	.w2(32'hbbbe86dd),
	.w3(32'hb92eee53),
	.w4(32'h3b44269e),
	.w5(32'hbc02ec82),
	.w6(32'h3b6ecfcb),
	.w7(32'hbb7b9248),
	.w8(32'hbb0d6f25),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba26390),
	.w1(32'h3c562dcb),
	.w2(32'h3b758fc5),
	.w3(32'hbad1a378),
	.w4(32'h3c086daa),
	.w5(32'hbbfd1d66),
	.w6(32'h3c2d932d),
	.w7(32'h3c654472),
	.w8(32'h3b870a06),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dc7d4),
	.w1(32'hbac9ca4b),
	.w2(32'hba1cffd4),
	.w3(32'hba7b465c),
	.w4(32'hba3ed4f2),
	.w5(32'hbb148ab6),
	.w6(32'hba23654c),
	.w7(32'hba72e7ef),
	.w8(32'hb926c49f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba816ed4),
	.w1(32'h390fe914),
	.w2(32'hbb2c056b),
	.w3(32'hba8833da),
	.w4(32'hba6a5df6),
	.w5(32'hbaa94694),
	.w6(32'hbad46fa0),
	.w7(32'hbb2a7e9a),
	.w8(32'hbb292aee),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3b836),
	.w1(32'h3a5d7ae8),
	.w2(32'h3a8da17b),
	.w3(32'h3a75c70c),
	.w4(32'hb95d1fb8),
	.w5(32'hb9a61840),
	.w6(32'h3abcd6e8),
	.w7(32'h3a3e1159),
	.w8(32'hba34ab54),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae4bab),
	.w1(32'h352d478f),
	.w2(32'h3a0bf014),
	.w3(32'hbaa70564),
	.w4(32'hb7b8a45d),
	.w5(32'h39a74039),
	.w6(32'hba29a3d7),
	.w7(32'hbaf8f435),
	.w8(32'hba24f47d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a414dcd),
	.w1(32'h3a24d95e),
	.w2(32'h3a31632b),
	.w3(32'h3a0fe227),
	.w4(32'h398cbbb0),
	.w5(32'h394fbf1b),
	.w6(32'hba239731),
	.w7(32'hba7c8b60),
	.w8(32'hb8b3d2fd),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a168646),
	.w1(32'h3b0a6d29),
	.w2(32'h3b0e9ba4),
	.w3(32'h3a16e8aa),
	.w4(32'h3ac00465),
	.w5(32'h3a01c391),
	.w6(32'hb9a2c594),
	.w7(32'h3a52caa9),
	.w8(32'h3a810e14),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b5e81),
	.w1(32'hba5b9c70),
	.w2(32'hbab76b4f),
	.w3(32'h3ae5b77b),
	.w4(32'h399881a8),
	.w5(32'hba7aca49),
	.w6(32'h39816ed0),
	.w7(32'h3aaab7d5),
	.w8(32'hba01ca60),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88ddf5),
	.w1(32'hb9800627),
	.w2(32'h3b5a39b1),
	.w3(32'hb9ad9816),
	.w4(32'h3a8356a7),
	.w5(32'h3a210a4a),
	.w6(32'hb9a9e9e2),
	.w7(32'hba780f5a),
	.w8(32'hbb4e2501),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f08629),
	.w1(32'hb9fb32e9),
	.w2(32'hba84b6b4),
	.w3(32'hbacab5f3),
	.w4(32'hba8b4aa3),
	.w5(32'hba9801f0),
	.w6(32'hba9675d5),
	.w7(32'hba6ff42f),
	.w8(32'hba9b9724),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aacdee),
	.w1(32'hba0e1c19),
	.w2(32'h3b528e66),
	.w3(32'h3a8a6673),
	.w4(32'hba46e93d),
	.w5(32'h398fb88a),
	.w6(32'hba67d779),
	.w7(32'h3a98f383),
	.w8(32'h3a281ad3),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7648f1),
	.w1(32'hbb9dc660),
	.w2(32'hbad87831),
	.w3(32'h3a7095ea),
	.w4(32'hbb7a182c),
	.w5(32'hbb97a9a9),
	.w6(32'hbb88b1ae),
	.w7(32'h3a06d6ff),
	.w8(32'hbb6faa73),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaecfd0),
	.w1(32'h3a8958b8),
	.w2(32'h39a5c6c4),
	.w3(32'hbab31330),
	.w4(32'hba1bc728),
	.w5(32'hb9bcf4ca),
	.w6(32'h39ba685a),
	.w7(32'h3a76e52a),
	.w8(32'hba3a3069),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5ae68),
	.w1(32'h3c50dc0d),
	.w2(32'hbac0a731),
	.w3(32'h3a288539),
	.w4(32'h3c2b0401),
	.w5(32'hbc11544b),
	.w6(32'h3c941d42),
	.w7(32'h3c33a63c),
	.w8(32'h3b9c2164),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedebe4),
	.w1(32'hbb228764),
	.w2(32'hb916677b),
	.w3(32'hbb6d94c0),
	.w4(32'hbb0f12b7),
	.w5(32'hba287c42),
	.w6(32'hb9d9440b),
	.w7(32'hba819268),
	.w8(32'hba02a438),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0a438),
	.w1(32'hba78fee9),
	.w2(32'hba84a78d),
	.w3(32'hba707bfc),
	.w4(32'hbad80b10),
	.w5(32'hbb084686),
	.w6(32'h39a3f34e),
	.w7(32'hba7a6384),
	.w8(32'h3a0f535e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf5a98),
	.w1(32'hba600b29),
	.w2(32'hba1337b8),
	.w3(32'hbaa1d6d8),
	.w4(32'hba11801a),
	.w5(32'hba8ebaca),
	.w6(32'h3a3922d9),
	.w7(32'h3aba3a1f),
	.w8(32'h39d57caf),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987f72f),
	.w1(32'h3c3723f1),
	.w2(32'h3c259d8d),
	.w3(32'hb73024f3),
	.w4(32'h3b72af90),
	.w5(32'h3afcc53d),
	.w6(32'h3cb0edb8),
	.w7(32'h3ce8c7b4),
	.w8(32'h3c5c88c0),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc99e2),
	.w1(32'hb9d5b924),
	.w2(32'h398eb5fb),
	.w3(32'hbbf18fe8),
	.w4(32'h38ca8309),
	.w5(32'hbb24abf9),
	.w6(32'h3a63e6c5),
	.w7(32'hb9313b39),
	.w8(32'hba588f2b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba682a64),
	.w1(32'hbb2d2283),
	.w2(32'h394f310c),
	.w3(32'hbab2ded8),
	.w4(32'hbb2c9c57),
	.w5(32'hbadde969),
	.w6(32'hbb8552ff),
	.w7(32'hbb5ae890),
	.w8(32'hbb21c909),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa9d89),
	.w1(32'hb98dcb12),
	.w2(32'hba16d314),
	.w3(32'hb9c32bcd),
	.w4(32'hb9db9b53),
	.w5(32'hba2f7636),
	.w6(32'hba920cae),
	.w7(32'hb9d095af),
	.w8(32'hb9303032),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba082b67),
	.w1(32'hbb03efa4),
	.w2(32'hb9be4c6c),
	.w3(32'hb91e3227),
	.w4(32'hbae7eb6d),
	.w5(32'hbb4b3465),
	.w6(32'hb948d4a9),
	.w7(32'hb90363fd),
	.w8(32'h3a4bef6e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e1e79),
	.w1(32'hba11d1d6),
	.w2(32'hbaf5c99a),
	.w3(32'hba4390a1),
	.w4(32'hbabcb107),
	.w5(32'hbb1033b0),
	.w6(32'hbb03aa49),
	.w7(32'hba0c5149),
	.w8(32'hba4b0593),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb058224),
	.w1(32'hbaa2a335),
	.w2(32'hba81aca9),
	.w3(32'h3915ff7d),
	.w4(32'hba729b3b),
	.w5(32'hba154063),
	.w6(32'hba81c23a),
	.w7(32'hb9f2ae67),
	.w8(32'h39f9b0d8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba331910),
	.w1(32'hb99e98f0),
	.w2(32'h3a3db8fc),
	.w3(32'hba23b6b6),
	.w4(32'hbb1c663f),
	.w5(32'hbb26015c),
	.w6(32'h3b4b1afc),
	.w7(32'h3b4594c1),
	.w8(32'h3a07c5eb),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e35e5),
	.w1(32'hba84c1d3),
	.w2(32'hbacc83e0),
	.w3(32'hbb5cd6d6),
	.w4(32'hbb111f25),
	.w5(32'hbb1daa25),
	.w6(32'h3a8cc62a),
	.w7(32'h39aec53e),
	.w8(32'h392b6e9d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24b33a),
	.w1(32'h3bdf4ffe),
	.w2(32'hbb83b17e),
	.w3(32'hbad97314),
	.w4(32'h3b4b9e77),
	.w5(32'hbc15e555),
	.w6(32'h3c5216f6),
	.w7(32'h3c03bdee),
	.w8(32'h3bb01234),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdaf4f8),
	.w1(32'hbabd1978),
	.w2(32'h3a835256),
	.w3(32'hbb2ebb2c),
	.w4(32'hba008caf),
	.w5(32'h3a224bc5),
	.w6(32'hbaa946f5),
	.w7(32'hbabb28ff),
	.w8(32'hba0228c1),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02e7ac),
	.w1(32'h3a5f2e27),
	.w2(32'h3b5896f2),
	.w3(32'h3a2587f9),
	.w4(32'hba70b80b),
	.w5(32'h3b034393),
	.w6(32'hba7096cc),
	.w7(32'hbb133bcd),
	.w8(32'hbb4915a3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eece7),
	.w1(32'h3c166cb5),
	.w2(32'h3abd7d98),
	.w3(32'hba70ff16),
	.w4(32'h3bcc83ec),
	.w5(32'hbb907791),
	.w6(32'h3b3dcbb7),
	.w7(32'h3a438c19),
	.w8(32'h384f7cee),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf5506),
	.w1(32'h3a38539c),
	.w2(32'hbacd289e),
	.w3(32'hba9fd30d),
	.w4(32'hbad06b80),
	.w5(32'hbb593cbb),
	.w6(32'hba03639f),
	.w7(32'hb9fe68f7),
	.w8(32'h39a98600),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07336e),
	.w1(32'hba835552),
	.w2(32'hba385f30),
	.w3(32'h3a496020),
	.w4(32'hbaac9cac),
	.w5(32'hba2e3643),
	.w6(32'h3a4a23b7),
	.w7(32'hba296e70),
	.w8(32'h3996e76d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b8cae),
	.w1(32'hb95b502e),
	.w2(32'hbaaf01f6),
	.w3(32'hbac50f53),
	.w4(32'hb9f7c943),
	.w5(32'hbaefe7f7),
	.w6(32'h3a0041f4),
	.w7(32'h3acf6ad4),
	.w8(32'hb98ea043),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1665b),
	.w1(32'h3a9bceee),
	.w2(32'hbb63880a),
	.w3(32'hbaf8b9e1),
	.w4(32'hbb3a9d45),
	.w5(32'hbbdfea8e),
	.w6(32'h3b34c8e4),
	.w7(32'hb97922b1),
	.w8(32'h3ada3478),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5d041),
	.w1(32'hba5a97e1),
	.w2(32'hba937ba6),
	.w3(32'h3a7fe71e),
	.w4(32'h38c98f4c),
	.w5(32'hbac729a0),
	.w6(32'h3b22e720),
	.w7(32'hbb44424d),
	.w8(32'hbb51e283),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc94e3),
	.w1(32'hbb2830c5),
	.w2(32'hba51cb37),
	.w3(32'hbaa3ed37),
	.w4(32'hbb451aa8),
	.w5(32'hbac85ec5),
	.w6(32'hbb584bd4),
	.w7(32'hbb263f82),
	.w8(32'hbae78d9b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52b4b0),
	.w1(32'h38eec773),
	.w2(32'hb886ed58),
	.w3(32'h3b1449fe),
	.w4(32'hb95b0036),
	.w5(32'hb9f40725),
	.w6(32'hb98a2224),
	.w7(32'hba975e12),
	.w8(32'hba37d693),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25dab2),
	.w1(32'hb8d55c70),
	.w2(32'h38e466bd),
	.w3(32'h3a92f150),
	.w4(32'hba7f056f),
	.w5(32'hb9a50033),
	.w6(32'hba9c1b92),
	.w7(32'hba81c8d2),
	.w8(32'hba2a2627),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389e1c18),
	.w1(32'h3acc2f1b),
	.w2(32'h3b2d270b),
	.w3(32'h3a758e3f),
	.w4(32'h3af34fb9),
	.w5(32'h3a95aaa0),
	.w6(32'h3a95011d),
	.w7(32'h3ac2d1b0),
	.w8(32'h38824aa7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c5719),
	.w1(32'hbae9f7ec),
	.w2(32'h393c3e95),
	.w3(32'h398fc973),
	.w4(32'hbb048a2b),
	.w5(32'hba9e8f63),
	.w6(32'hba076c18),
	.w7(32'hb9d777d1),
	.w8(32'hba3da308),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54b0be),
	.w1(32'hba80c0b1),
	.w2(32'hba95737e),
	.w3(32'hbac71f6a),
	.w4(32'hba9baeb9),
	.w5(32'hba66e9dc),
	.w6(32'hbb497fda),
	.w7(32'hba85c5d9),
	.w8(32'h38e71b71),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae4d9a),
	.w1(32'hb983a2ce),
	.w2(32'hb8a0ab8d),
	.w3(32'hba08e2de),
	.w4(32'hba52f258),
	.w5(32'hb990dcd8),
	.w6(32'hbaa5270c),
	.w7(32'hba94e385),
	.w8(32'hba3a6270),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b39cd2),
	.w1(32'hba16c032),
	.w2(32'h3ad5cc79),
	.w3(32'h3a8fff07),
	.w4(32'h38b02c07),
	.w5(32'hb8d9840e),
	.w6(32'hba9d1902),
	.w7(32'h3aaa5421),
	.w8(32'h3a39f865),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fd024),
	.w1(32'hb951630e),
	.w2(32'hbb0c9902),
	.w3(32'hba59f5b6),
	.w4(32'hb9b9cf34),
	.w5(32'hbb14a05f),
	.w6(32'hba953415),
	.w7(32'hb9735304),
	.w8(32'hba7596d9),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba246628),
	.w1(32'hbb8ef5fa),
	.w2(32'hbb5fe99f),
	.w3(32'h3aa2dcf4),
	.w4(32'hbb5cedce),
	.w5(32'hbbde6fc9),
	.w6(32'hbb6b582e),
	.w7(32'h3a780045),
	.w8(32'h3a21b215),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcc9fe),
	.w1(32'h3983a0b5),
	.w2(32'hb9f72b66),
	.w3(32'h3b37bb73),
	.w4(32'h3a017763),
	.w5(32'hbacb5c2f),
	.w6(32'h3a511a86),
	.w7(32'h3a227946),
	.w8(32'hba1ec224),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7716e),
	.w1(32'hba81c2df),
	.w2(32'hb85ac6e5),
	.w3(32'h3aa11c94),
	.w4(32'h3a33c677),
	.w5(32'h395eb815),
	.w6(32'hb9147fd8),
	.w7(32'hbabf674b),
	.w8(32'hbb06930d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e36dc),
	.w1(32'hbb00d9cd),
	.w2(32'hbae6cc5f),
	.w3(32'h3a2126b3),
	.w4(32'hba65336c),
	.w5(32'hbb41a41b),
	.w6(32'hbae07d7d),
	.w7(32'h397c6c48),
	.w8(32'hb93a0817),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fcf3e),
	.w1(32'hb9064f7c),
	.w2(32'h3861b8de),
	.w3(32'h38c632d1),
	.w4(32'hbaa20878),
	.w5(32'hb9dd7b12),
	.w6(32'hbad28f93),
	.w7(32'hbaa91cc9),
	.w8(32'hba658036),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e7ca8),
	.w1(32'h39c7b424),
	.w2(32'h3a390487),
	.w3(32'h3aca12bf),
	.w4(32'hba337a5a),
	.w5(32'hb8fe0a45),
	.w6(32'hb9213c52),
	.w7(32'hb971b6a8),
	.w8(32'hb92935f3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a250e9f),
	.w1(32'h3836049d),
	.w2(32'h3a0025e1),
	.w3(32'h39df4975),
	.w4(32'hba9b478a),
	.w5(32'hb99e2a80),
	.w6(32'hba2fad75),
	.w7(32'hba27bdc4),
	.w8(32'hba0cd2cc),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96763d9),
	.w1(32'h394e00d5),
	.w2(32'h3a9bf41d),
	.w3(32'hb9787d34),
	.w4(32'h3aa7e274),
	.w5(32'h3a79ff12),
	.w6(32'hba2acba0),
	.w7(32'hbadd84f7),
	.w8(32'hb7fd4cc1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66a704),
	.w1(32'h3b47f120),
	.w2(32'h3b880c73),
	.w3(32'h396888dc),
	.w4(32'hba01da17),
	.w5(32'h3a5203c5),
	.w6(32'h3ab156b6),
	.w7(32'h3b70a6fb),
	.w8(32'h3a4de24f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b9358),
	.w1(32'h3ac21141),
	.w2(32'h39bfa690),
	.w3(32'hba4bc134),
	.w4(32'hb92bc223),
	.w5(32'hba6a5056),
	.w6(32'h3ad11245),
	.w7(32'h379567cf),
	.w8(32'hb93a2a08),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9e671),
	.w1(32'h39df2d16),
	.w2(32'hba4a5ea8),
	.w3(32'hbaa8f3c6),
	.w4(32'hba31a9b9),
	.w5(32'hba9172a4),
	.w6(32'h37c8f067),
	.w7(32'hbaf79240),
	.w8(32'h38f707a4),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f6a61d),
	.w1(32'h39ee370d),
	.w2(32'h394cead5),
	.w3(32'hba8462bc),
	.w4(32'h39fd8bcf),
	.w5(32'h39b64c22),
	.w6(32'hbaa72060),
	.w7(32'hba9c1bcd),
	.w8(32'hb9959085),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a134887),
	.w1(32'h3a20f29d),
	.w2(32'h3b818f17),
	.w3(32'h3a9fabff),
	.w4(32'h3997e626),
	.w5(32'hb9a01a37),
	.w6(32'h3b85d075),
	.w7(32'h3a98b7dd),
	.w8(32'hb9ffbb88),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04f181),
	.w1(32'h395276f2),
	.w2(32'h3919094e),
	.w3(32'hbb2b30bf),
	.w4(32'hbb12046a),
	.w5(32'hbb5b8685),
	.w6(32'h3b298743),
	.w7(32'h3a16157c),
	.w8(32'hb961fd01),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb927b55),
	.w1(32'h3a352844),
	.w2(32'h3aa3a749),
	.w3(32'hbb95f02c),
	.w4(32'hba901d96),
	.w5(32'h38a5c3f7),
	.w6(32'hb9fec384),
	.w7(32'h399c1475),
	.w8(32'hb908f085),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b49c9b),
	.w1(32'h3aaa91b9),
	.w2(32'h3bbe3204),
	.w3(32'h3938b7a6),
	.w4(32'hbac36245),
	.w5(32'h3bae1161),
	.w6(32'hbb2147af),
	.w7(32'h3b3b5c02),
	.w8(32'hba25d32e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb452546),
	.w1(32'hb97b5135),
	.w2(32'hbb1675b1),
	.w3(32'hbb8be1b1),
	.w4(32'hbb56fe06),
	.w5(32'hbb579d53),
	.w6(32'hbb195c9a),
	.w7(32'hbadae1fb),
	.w8(32'hbb4af617),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule