module layer_10_featuremap_306(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc2e8c),
	.w1(32'h398b3ad5),
	.w2(32'hba323e7b),
	.w3(32'h3b9c035f),
	.w4(32'hb9927b89),
	.w5(32'h3b2a1040),
	.w6(32'h3bce3acc),
	.w7(32'hbad39088),
	.w8(32'h3bd6c553),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a467cac),
	.w1(32'hbbba2703),
	.w2(32'hbbdf2b24),
	.w3(32'hbbbea766),
	.w4(32'hbb69c342),
	.w5(32'hbbb8008f),
	.w6(32'hbb425af7),
	.w7(32'hbbd5c7b9),
	.w8(32'hbad1e708),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0c103),
	.w1(32'hbbed51f4),
	.w2(32'h3aabf237),
	.w3(32'hbbee2261),
	.w4(32'h39f26483),
	.w5(32'h3bab8169),
	.w6(32'h3b39a4c8),
	.w7(32'h39e5c5e3),
	.w8(32'h3b8fd855),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af715ec),
	.w1(32'hba9c8105),
	.w2(32'hb9945cfc),
	.w3(32'hbafac5f5),
	.w4(32'hbb43098d),
	.w5(32'hba2edb41),
	.w6(32'hbb813c6b),
	.w7(32'hbb180331),
	.w8(32'hbb43ea5a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9560d1),
	.w1(32'hbbc48f34),
	.w2(32'hba8371cd),
	.w3(32'hbc44500d),
	.w4(32'hbc272fa2),
	.w5(32'hbad91155),
	.w6(32'hbbd906b8),
	.w7(32'h3b60ad3a),
	.w8(32'hbb3b188f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fba3e),
	.w1(32'hbb55bc11),
	.w2(32'h3a9bad3f),
	.w3(32'h3a25e9ca),
	.w4(32'h3a8ecd1b),
	.w5(32'hbb128849),
	.w6(32'hbb357139),
	.w7(32'h3ab3e937),
	.w8(32'hbb7ec808),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb43b6e),
	.w1(32'hbb31af91),
	.w2(32'hba0e8fc5),
	.w3(32'hbb6ff67c),
	.w4(32'hb9f1f943),
	.w5(32'h3a50a27a),
	.w6(32'hbae134b0),
	.w7(32'hba943345),
	.w8(32'h3a807de2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70e368),
	.w1(32'hbb33797c),
	.w2(32'h3ae5aaf1),
	.w3(32'h3c1650ed),
	.w4(32'h3ba719a8),
	.w5(32'hba47e938),
	.w6(32'h3bdd42d0),
	.w7(32'h3a143328),
	.w8(32'hbb3409cd),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d0110),
	.w1(32'hbac7d078),
	.w2(32'h3a2adc97),
	.w3(32'h3b0ed0e1),
	.w4(32'h3b52f45a),
	.w5(32'hbac79604),
	.w6(32'hbb5862a4),
	.w7(32'hbac22ddc),
	.w8(32'hba84846a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5405be),
	.w1(32'h3a1a5ea6),
	.w2(32'h3b873c67),
	.w3(32'h3b1e2ae9),
	.w4(32'h3b3185c1),
	.w5(32'hb9b90493),
	.w6(32'hb8864b35),
	.w7(32'h3ab5c748),
	.w8(32'hbb8ce28c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb521e80),
	.w1(32'hbbf696af),
	.w2(32'h3abc77e6),
	.w3(32'hbb756e2f),
	.w4(32'hba8da6ff),
	.w5(32'hbb6db89f),
	.w6(32'hbc020763),
	.w7(32'hbaf6e262),
	.w8(32'hba5956d1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac60a0b),
	.w1(32'hbbe7f3f4),
	.w2(32'h3b7b7f4b),
	.w3(32'hbb1d9caf),
	.w4(32'hbac31857),
	.w5(32'hbc39eb1a),
	.w6(32'hbb3b7067),
	.w7(32'hbb6814a5),
	.w8(32'hbc04481a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b930a6d),
	.w1(32'h3c925eee),
	.w2(32'h3c7286be),
	.w3(32'h3c781ef6),
	.w4(32'h3bc6fa4e),
	.w5(32'h3aa63933),
	.w6(32'h3c620bd6),
	.w7(32'h3c420d77),
	.w8(32'h3c376368),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd46baf),
	.w1(32'hba66a0c0),
	.w2(32'hbb2778f4),
	.w3(32'h3c648852),
	.w4(32'h3a50321a),
	.w5(32'hbb63b64e),
	.w6(32'h3c404126),
	.w7(32'hbc18b97f),
	.w8(32'hbaa2b926),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b126433),
	.w1(32'hbb6818bc),
	.w2(32'h3bab7d50),
	.w3(32'h3a712f16),
	.w4(32'h3a47275a),
	.w5(32'h3b92756e),
	.w6(32'hbbcad535),
	.w7(32'hba3c93e2),
	.w8(32'h3bd1d188),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae9dd5),
	.w1(32'hbbdf36a2),
	.w2(32'hbaf2925b),
	.w3(32'hbb430897),
	.w4(32'hbb5571a5),
	.w5(32'h3983bc2d),
	.w6(32'hbb93718d),
	.w7(32'hbb725667),
	.w8(32'h399b9a84),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0c4bd),
	.w1(32'hbbde2a06),
	.w2(32'hba623783),
	.w3(32'h3a1fe25a),
	.w4(32'hba0c1226),
	.w5(32'hbbe88b9c),
	.w6(32'hbba27fb7),
	.w7(32'hbaac76dd),
	.w8(32'hbbdd5476),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a853bdd),
	.w1(32'h3bc45714),
	.w2(32'h3bfc2f19),
	.w3(32'hbb39353f),
	.w4(32'h3a73ee6e),
	.w5(32'h39b113ad),
	.w6(32'h3b988a43),
	.w7(32'h3bf0e7ba),
	.w8(32'hbb589e5a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc73f7d),
	.w1(32'hbbc8bf94),
	.w2(32'h3b3d2c58),
	.w3(32'hbb505bf0),
	.w4(32'h3b868d23),
	.w5(32'h3ba6058a),
	.w6(32'h3a6b86a4),
	.w7(32'h3b94f2a1),
	.w8(32'hba4dec00),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30b1c1),
	.w1(32'hbb319b01),
	.w2(32'h3baf697b),
	.w3(32'hbb8af462),
	.w4(32'hbc1e349b),
	.w5(32'hba75d542),
	.w6(32'hbbb7e19f),
	.w7(32'hbbf35566),
	.w8(32'h3b547c19),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba69ed7),
	.w1(32'h3a4687a1),
	.w2(32'hbb984524),
	.w3(32'hbb20ef12),
	.w4(32'hbb51fe37),
	.w5(32'hba2ac81a),
	.w6(32'h3b3f0ab0),
	.w7(32'hbbcb4c14),
	.w8(32'h39cf7a92),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ba011),
	.w1(32'hbb9310c2),
	.w2(32'hbbcd1e99),
	.w3(32'h3b43b993),
	.w4(32'hb9185e9f),
	.w5(32'hbb48c0c5),
	.w6(32'hb909b85f),
	.w7(32'hbb276e55),
	.w8(32'h3a9c954d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba779c39),
	.w1(32'h3ab4bda2),
	.w2(32'h3b98e3c3),
	.w3(32'h3b2aeed1),
	.w4(32'hbb52f3b1),
	.w5(32'h3bc33c6d),
	.w6(32'h3c6467ec),
	.w7(32'h3a9115f3),
	.w8(32'h3ba3728a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c045cee),
	.w1(32'h3b930f7f),
	.w2(32'h3c1509b2),
	.w3(32'h3ae564b2),
	.w4(32'h3bcfb3a7),
	.w5(32'h3bdb62c9),
	.w6(32'h3b81daf0),
	.w7(32'h3b7a21e6),
	.w8(32'h3a0f0afb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfae180),
	.w1(32'h3ab11c7e),
	.w2(32'h3b23d3e9),
	.w3(32'hbab3abb1),
	.w4(32'h3ad06edb),
	.w5(32'hbb81a277),
	.w6(32'hbb8f91da),
	.w7(32'h3c3e8251),
	.w8(32'hbbacf097),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac586fd),
	.w1(32'hbbd20dc3),
	.w2(32'h3b27c1a1),
	.w3(32'hbb4e9138),
	.w4(32'hbb8f47a0),
	.w5(32'h3b480bbe),
	.w6(32'hbbec3c89),
	.w7(32'h38091534),
	.w8(32'h3b9191c8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bb981),
	.w1(32'h3a1588bc),
	.w2(32'hb99f24ec),
	.w3(32'h3947baa6),
	.w4(32'hb9913edb),
	.w5(32'hba4ad6f3),
	.w6(32'h3a8c1aff),
	.w7(32'h39c947b2),
	.w8(32'h3ace2e3b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6f2d0),
	.w1(32'h3ba08d43),
	.w2(32'h3ac3565e),
	.w3(32'h3baa02cc),
	.w4(32'h3b8ceff4),
	.w5(32'h3b423d7e),
	.w6(32'h3b4adbb3),
	.w7(32'h3b46b302),
	.w8(32'h3b372a85),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae52d51),
	.w1(32'hbb8aefd6),
	.w2(32'hbb952f82),
	.w3(32'hba6ac10b),
	.w4(32'hbbb445ca),
	.w5(32'h3b7b4cba),
	.w6(32'hbbaab301),
	.w7(32'hbbe775db),
	.w8(32'h3b7de0c6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e4114),
	.w1(32'hba76e443),
	.w2(32'h390c1663),
	.w3(32'hbb91cc6f),
	.w4(32'hbb998dcb),
	.w5(32'hbbb41b39),
	.w6(32'h3ba244e8),
	.w7(32'hba769cd6),
	.w8(32'hb82c15a5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a9755),
	.w1(32'h3bc6e45e),
	.w2(32'h3c2e4a9b),
	.w3(32'h3c09568b),
	.w4(32'h3b0f773d),
	.w5(32'hbb6bf53b),
	.w6(32'h3c477f76),
	.w7(32'h3b380fd3),
	.w8(32'hbb08c31c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e268e),
	.w1(32'hbadb395a),
	.w2(32'h3a7f6a31),
	.w3(32'h39fb3360),
	.w4(32'h3af0377f),
	.w5(32'hbc5d6b5e),
	.w6(32'hbc2c6e88),
	.w7(32'h393c5c45),
	.w8(32'hbc80ab4e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ddd8f),
	.w1(32'hbafb517d),
	.w2(32'h3b0f066a),
	.w3(32'hbbc076f1),
	.w4(32'hb7ad0184),
	.w5(32'hbc445dc5),
	.w6(32'h3c5a579c),
	.w7(32'hb8e15bee),
	.w8(32'hbc5f7399),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2e58b),
	.w1(32'h3c55625c),
	.w2(32'h3c4fd43e),
	.w3(32'hbc1c3019),
	.w4(32'h3b49ff38),
	.w5(32'h3c297b6b),
	.w6(32'h3a21ca21),
	.w7(32'h3c6ae9e6),
	.w8(32'h3c13a34f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb12adc),
	.w1(32'hbb4fb44c),
	.w2(32'hbb8660a6),
	.w3(32'h3b368b25),
	.w4(32'hbb142102),
	.w5(32'hbbc316dc),
	.w6(32'hbbf469f6),
	.w7(32'h3adada5e),
	.w8(32'hbbc294b5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b706aba),
	.w1(32'h3c388fb8),
	.w2(32'h3b614851),
	.w3(32'h3b1c3ca0),
	.w4(32'h38e5f1d0),
	.w5(32'hbb70c5f9),
	.w6(32'h3c11b9c3),
	.w7(32'h3bd6e25f),
	.w8(32'h3a982d5d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba3a13),
	.w1(32'hbb5c13cf),
	.w2(32'h3c032dd7),
	.w3(32'hbbdea16c),
	.w4(32'hbbd189f9),
	.w5(32'hbad03cde),
	.w6(32'hbc2ef448),
	.w7(32'h3c14716d),
	.w8(32'hba71934d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a0d83),
	.w1(32'hba52534f),
	.w2(32'h3a0bc615),
	.w3(32'h3b082b91),
	.w4(32'hbb98ff79),
	.w5(32'h3935e7c5),
	.w6(32'h3b618747),
	.w7(32'hbad8d43d),
	.w8(32'hb71ccb76),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8687cb),
	.w1(32'hbb9f6192),
	.w2(32'hbaa05ac3),
	.w3(32'hbbe69a54),
	.w4(32'hbbadee6f),
	.w5(32'h3ba822dc),
	.w6(32'hbbe0156b),
	.w7(32'hbb7650bd),
	.w8(32'h3c1812a0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d64a5),
	.w1(32'hbadf912a),
	.w2(32'hbba8a82c),
	.w3(32'h3c4308c4),
	.w4(32'h371eeb6c),
	.w5(32'h3a4862bf),
	.w6(32'h3c0f189c),
	.w7(32'h3b7e2421),
	.w8(32'h3b9ec4b3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ce7ad),
	.w1(32'h3b80183c),
	.w2(32'h3ac884ea),
	.w3(32'h3c212109),
	.w4(32'h3bb07007),
	.w5(32'hbbc48df8),
	.w6(32'h3c978bde),
	.w7(32'hbb9e5017),
	.w8(32'hbb8fc775),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb411d),
	.w1(32'hbbc4baa6),
	.w2(32'h3a6c0a6f),
	.w3(32'hbba9f6b1),
	.w4(32'hbb209030),
	.w5(32'h3bde5a5d),
	.w6(32'hbbe94682),
	.w7(32'hbaf617ef),
	.w8(32'h3b3b651d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae21397),
	.w1(32'hbc2a96f9),
	.w2(32'hbbefd353),
	.w3(32'hbb9336c4),
	.w4(32'hbbb274d5),
	.w5(32'h3c0acbc0),
	.w6(32'hbc1b56a7),
	.w7(32'hbc100c20),
	.w8(32'h3b8ab58a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c118d9b),
	.w1(32'h3b10e39d),
	.w2(32'h3b0fd800),
	.w3(32'h39ef4b4f),
	.w4(32'h3b86c115),
	.w5(32'h39e48489),
	.w6(32'hbb2510ed),
	.w7(32'hbbd0a02f),
	.w8(32'hbb5466f0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19c4f5),
	.w1(32'hbbcafe8a),
	.w2(32'h3a9b1fe1),
	.w3(32'hbb9ff0f6),
	.w4(32'hbabe3af4),
	.w5(32'hbbc4f2d1),
	.w6(32'hbb8de57f),
	.w7(32'h3a970281),
	.w8(32'hbc00ea44),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81ce9e),
	.w1(32'h3c376954),
	.w2(32'h3c261435),
	.w3(32'h3afa8ca4),
	.w4(32'h3b9b2d6c),
	.w5(32'hbbacc7ef),
	.w6(32'hbb933e11),
	.w7(32'h3c262c3d),
	.w8(32'hbbbb7a28),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbacb8b),
	.w1(32'h3b84b0cc),
	.w2(32'h3bdb9d20),
	.w3(32'hba32055e),
	.w4(32'h3ae26acf),
	.w5(32'h3bb492e7),
	.w6(32'h3afd2c1d),
	.w7(32'h3c256b3a),
	.w8(32'h3bbaa323),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70ef75),
	.w1(32'hbc0791f7),
	.w2(32'hbbc07b3a),
	.w3(32'h3be4065f),
	.w4(32'h3a9e6ed9),
	.w5(32'hbc153e5f),
	.w6(32'h3b23f9ec),
	.w7(32'hbb58b5a1),
	.w8(32'hbc1bfa23),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaf1ae),
	.w1(32'h3ba6dc72),
	.w2(32'h3c1b8668),
	.w3(32'hba0dff44),
	.w4(32'h3a8fcc18),
	.w5(32'hba00d0bb),
	.w6(32'hbb189334),
	.w7(32'hb9b7556d),
	.w8(32'h3a31dc63),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3f16f),
	.w1(32'hbbed6454),
	.w2(32'hbbb76b7b),
	.w3(32'h39ad4937),
	.w4(32'hb9f790b7),
	.w5(32'hbb0ac4df),
	.w6(32'hba500721),
	.w7(32'hba5c4acc),
	.w8(32'hbc626fbc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a7b2e),
	.w1(32'h3b894347),
	.w2(32'hbc085197),
	.w3(32'hbb0c093b),
	.w4(32'hbb842cc2),
	.w5(32'h3beacf26),
	.w6(32'h3cc46fa6),
	.w7(32'hb9cfa640),
	.w8(32'h3b13568b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c5665),
	.w1(32'hb99d6787),
	.w2(32'h3b39feb5),
	.w3(32'h3a66496a),
	.w4(32'hbbcb154b),
	.w5(32'hbc403b15),
	.w6(32'hba32b948),
	.w7(32'hbaaaddb4),
	.w8(32'hbba801f6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c5698),
	.w1(32'hbacc8903),
	.w2(32'hbbb508de),
	.w3(32'h3b18062e),
	.w4(32'h3b27c707),
	.w5(32'hbb6c19d6),
	.w6(32'h3cb3d46d),
	.w7(32'hbb86ffbe),
	.w8(32'hbb5920f9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f774d),
	.w1(32'h3bc02299),
	.w2(32'h3b43672c),
	.w3(32'hbab65617),
	.w4(32'hbbbf5316),
	.w5(32'h3b616477),
	.w6(32'h3b061970),
	.w7(32'hbbb4fdc1),
	.w8(32'hbb556dfd),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb536864),
	.w1(32'hb927a028),
	.w2(32'h3c2e2c7f),
	.w3(32'hbba1884d),
	.w4(32'hbb8125bc),
	.w5(32'h3bce3dd5),
	.w6(32'hbb83a9cc),
	.w7(32'hba564869),
	.w8(32'h3b99746f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38fd32),
	.w1(32'h3a1712cc),
	.w2(32'hbba338ab),
	.w3(32'hbbaa94fd),
	.w4(32'hbb3a851f),
	.w5(32'h3b2b1247),
	.w6(32'hbbe80bb5),
	.w7(32'hbb6ad355),
	.w8(32'h3a94137a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b41be),
	.w1(32'h3a57e687),
	.w2(32'h3b2555cd),
	.w3(32'h3b71e859),
	.w4(32'h3b119be6),
	.w5(32'h39fe667d),
	.w6(32'hbabca068),
	.w7(32'hbb46b0c9),
	.w8(32'h3b5da936),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31c583),
	.w1(32'hbc84302a),
	.w2(32'hbb550c2f),
	.w3(32'hbbeaa07b),
	.w4(32'hbb22e2fa),
	.w5(32'hba8b0a19),
	.w6(32'hbc04f587),
	.w7(32'hbb23657d),
	.w8(32'hbaca1db4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc050c07),
	.w1(32'hbbd8a237),
	.w2(32'hbb963467),
	.w3(32'h38c0121c),
	.w4(32'hbad27728),
	.w5(32'hbbd9c370),
	.w6(32'hbab3c9e2),
	.w7(32'hbb3a4a79),
	.w8(32'hbc2980df),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74bdb9),
	.w1(32'h3bca242a),
	.w2(32'h3c0697f4),
	.w3(32'h3ad7b83a),
	.w4(32'h3bf54242),
	.w5(32'hb90b8528),
	.w6(32'h3b1e4d43),
	.w7(32'h3c8b1379),
	.w8(32'hba75ddf9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acccfdf),
	.w1(32'hbba151f9),
	.w2(32'h3af344a8),
	.w3(32'hbb3f03c6),
	.w4(32'hbb029a0c),
	.w5(32'hbafc3e7b),
	.w6(32'hbb907420),
	.w7(32'hba65e953),
	.w8(32'hba59bd89),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ec6897),
	.w1(32'hbb92da30),
	.w2(32'h3ba303d0),
	.w3(32'hbafe616a),
	.w4(32'hba879448),
	.w5(32'h3ad72885),
	.w6(32'hbb7f2004),
	.w7(32'h3b8889bb),
	.w8(32'hba63d947),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbe1c7),
	.w1(32'hbb99c40e),
	.w2(32'hbb323956),
	.w3(32'hbbb1e004),
	.w4(32'hbb932a81),
	.w5(32'h3bfb74e7),
	.w6(32'hbb053ac9),
	.w7(32'h3aa117fc),
	.w8(32'h3bd7947b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bdf12),
	.w1(32'h3bc7571d),
	.w2(32'hb884f9e6),
	.w3(32'h3c260516),
	.w4(32'h3a6d0ed7),
	.w5(32'h3c353bb3),
	.w6(32'h3bd81de0),
	.w7(32'hbaca8b9c),
	.w8(32'h3bf34f76),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22b77f),
	.w1(32'hbb216339),
	.w2(32'hbb00dfbd),
	.w3(32'hbb52d70b),
	.w4(32'hbc12344d),
	.w5(32'hbbbee2e0),
	.w6(32'hbc0b9f7d),
	.w7(32'hbb8bc0e4),
	.w8(32'hbbc81472),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4789bf),
	.w1(32'hbb71fa43),
	.w2(32'h3adc5b95),
	.w3(32'hbb0813f5),
	.w4(32'hb9b203a2),
	.w5(32'h3b7a8a0f),
	.w6(32'h39361003),
	.w7(32'h38dad68f),
	.w8(32'h3a3dc6e6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2efb49),
	.w1(32'hbb1560ea),
	.w2(32'h3b80a63e),
	.w3(32'hba05dc78),
	.w4(32'h3b3ba896),
	.w5(32'h3bc1361a),
	.w6(32'h39eb9acb),
	.w7(32'h3a6196e9),
	.w8(32'h3b6c8b35),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af54486),
	.w1(32'h3ab473fb),
	.w2(32'h3b9b4eec),
	.w3(32'h3b99b816),
	.w4(32'h3bbd0eda),
	.w5(32'h39274c94),
	.w6(32'hbbc37f4d),
	.w7(32'hbc08135c),
	.w8(32'hbc499a79),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7ccaa),
	.w1(32'h3abf6dbe),
	.w2(32'hbb7533bf),
	.w3(32'hbc0f9b73),
	.w4(32'hbb7f215c),
	.w5(32'hbbd7900e),
	.w6(32'h3bab542c),
	.w7(32'hbb7bc1ce),
	.w8(32'hbba3e801),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7909e),
	.w1(32'h3b161f4e),
	.w2(32'h3c0d9a21),
	.w3(32'hbb4a675c),
	.w4(32'h3b63dbf9),
	.w5(32'h3bf510f7),
	.w6(32'hbb901094),
	.w7(32'h3ab4ba60),
	.w8(32'h3c3e1907),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb78d1),
	.w1(32'hbb4d3247),
	.w2(32'hb7bfa8ee),
	.w3(32'h3b5bbe0e),
	.w4(32'hbb25295e),
	.w5(32'h3af8a1ed),
	.w6(32'hbad34582),
	.w7(32'hbbb1a2d7),
	.w8(32'h3a665d54),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdbc19),
	.w1(32'hb9e1173c),
	.w2(32'hba0b1dd1),
	.w3(32'h3ad70dea),
	.w4(32'h3aa3e669),
	.w5(32'hba525461),
	.w6(32'h3afa5994),
	.w7(32'hbb24a086),
	.w8(32'h3bdcfe57),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf52f1a),
	.w1(32'hbb474d6e),
	.w2(32'h3b5a56f3),
	.w3(32'hbb34bae5),
	.w4(32'hbb5e4c8d),
	.w5(32'hbc3cc35a),
	.w6(32'hbb53bb0f),
	.w7(32'hbbc4bb49),
	.w8(32'hbc5699b3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47bbca),
	.w1(32'h3b2f5111),
	.w2(32'h3c1c4284),
	.w3(32'hbc77f0d0),
	.w4(32'hbb0c6dab),
	.w5(32'h3ab11050),
	.w6(32'hbbc33281),
	.w7(32'h3c9346e6),
	.w8(32'hbb438a7b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcb38d),
	.w1(32'hbbd0c353),
	.w2(32'h3af064d8),
	.w3(32'hbb38d94c),
	.w4(32'h3ad5cf3e),
	.w5(32'hbc426408),
	.w6(32'hbb88dd64),
	.w7(32'hbbc178f9),
	.w8(32'hbc182b0c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3000bc),
	.w1(32'h3c43409a),
	.w2(32'h3c02d26a),
	.w3(32'hbaf7c5c5),
	.w4(32'h3b1ec7ee),
	.w5(32'hbbe55124),
	.w6(32'h3bcd3ef4),
	.w7(32'h3c08010b),
	.w8(32'hbb923602),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3cf3c),
	.w1(32'hbb0f5345),
	.w2(32'hba40fa16),
	.w3(32'h3ba0d54b),
	.w4(32'h38edd599),
	.w5(32'hb709a07a),
	.w6(32'h3c322480),
	.w7(32'hbb173b49),
	.w8(32'hb9c00c6e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84994f4),
	.w1(32'h3ac64173),
	.w2(32'h399db4f2),
	.w3(32'h3aaa8e35),
	.w4(32'hbb97b86c),
	.w5(32'hbc5a9759),
	.w6(32'h3c104393),
	.w7(32'h3972a190),
	.w8(32'hbc349e5b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab2462),
	.w1(32'h3b8543ae),
	.w2(32'h3ba836ae),
	.w3(32'hb8102412),
	.w4(32'h3b9c3253),
	.w5(32'h3b2bcf76),
	.w6(32'h3b9ea7b5),
	.w7(32'h3c0492dd),
	.w8(32'hb8210bf0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50f6c1),
	.w1(32'h3b7eadae),
	.w2(32'h3c1b41dd),
	.w3(32'h3b529034),
	.w4(32'h3aee8c71),
	.w5(32'h3c07d427),
	.w6(32'hb7ee362c),
	.w7(32'h3a981643),
	.w8(32'h3b00e49c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d2ebc),
	.w1(32'hbb826e39),
	.w2(32'hbbfa9f2e),
	.w3(32'h3b5a4efd),
	.w4(32'h3b51164f),
	.w5(32'hbc37e67b),
	.w6(32'hbac8c33f),
	.w7(32'hbc14b9a2),
	.w8(32'hbc363006),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba652eb),
	.w1(32'h3aa3a90f),
	.w2(32'h3c218397),
	.w3(32'hbba4b2aa),
	.w4(32'h3b94e5c7),
	.w5(32'hb895fab3),
	.w6(32'hba0d944d),
	.w7(32'h3bf08373),
	.w8(32'h3add9aed),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb24ba),
	.w1(32'h3b7d87f8),
	.w2(32'hbc1706d8),
	.w3(32'h3b14fd64),
	.w4(32'hbb13ed41),
	.w5(32'h3a1c32f2),
	.w6(32'h3c865624),
	.w7(32'hbaa93bfa),
	.w8(32'h3bb0623c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbcfe8),
	.w1(32'hb9d2321a),
	.w2(32'hbb86ee42),
	.w3(32'hba284980),
	.w4(32'hba81096a),
	.w5(32'h3be35512),
	.w6(32'h3ab9ad76),
	.w7(32'hba5bfe87),
	.w8(32'h3bd06e9b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920d732),
	.w1(32'h3b79533d),
	.w2(32'h3b03fcb1),
	.w3(32'h3b34b4ee),
	.w4(32'h3b087f9c),
	.w5(32'hbc07198f),
	.w6(32'h3c367340),
	.w7(32'h3bc16ccd),
	.w8(32'hbc5c6817),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5c125),
	.w1(32'h3b0a4e09),
	.w2(32'h3bbfb7ae),
	.w3(32'h396974cf),
	.w4(32'hbb176190),
	.w5(32'h3a987228),
	.w6(32'hbbe866e9),
	.w7(32'h3b8fec97),
	.w8(32'h3b26535a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07f450),
	.w1(32'hbc01173b),
	.w2(32'hbb3f72bc),
	.w3(32'hbb2eddae),
	.w4(32'h3a5f2869),
	.w5(32'h3a6b9efa),
	.w6(32'h3aec4e18),
	.w7(32'hbbdbb60e),
	.w8(32'hbb461f2b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb118f8b),
	.w1(32'hbb62f63e),
	.w2(32'hbb895bab),
	.w3(32'hbabde98c),
	.w4(32'hbb9cb855),
	.w5(32'hba9c192e),
	.w6(32'hbbc89003),
	.w7(32'hbae49468),
	.w8(32'hbb1c181d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cb1d0),
	.w1(32'hbb2392a7),
	.w2(32'h3b7b1b4f),
	.w3(32'h3b594949),
	.w4(32'h3b03be0e),
	.w5(32'h3c1e266c),
	.w6(32'hb92d373a),
	.w7(32'h3b085c75),
	.w8(32'h3c5c08ac),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c155747),
	.w1(32'h3b7e7ff8),
	.w2(32'h3bd8ce18),
	.w3(32'h3c2d17a3),
	.w4(32'h3c0c414f),
	.w5(32'h3b2611dc),
	.w6(32'h3c5ab6f2),
	.w7(32'h3bb5d8a0),
	.w8(32'h3b2d6c53),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cb0e1),
	.w1(32'h3bb96505),
	.w2(32'hba8fd623),
	.w3(32'h3c000a5f),
	.w4(32'h3b151aa2),
	.w5(32'h3c08ef07),
	.w6(32'h3bb57ab3),
	.w7(32'h3a5b5239),
	.w8(32'h3b5826cd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba766998),
	.w1(32'hbc2e6a4f),
	.w2(32'hbaa9ec9c),
	.w3(32'hbb833148),
	.w4(32'hbc12cbda),
	.w5(32'h3c12197a),
	.w6(32'hbb75a33f),
	.w7(32'hbb635ff7),
	.w8(32'h3b1028c9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb603134),
	.w1(32'hbbe19185),
	.w2(32'hbb48ee4d),
	.w3(32'hbc1965c0),
	.w4(32'hbb59856d),
	.w5(32'h3a7a7cc9),
	.w6(32'hbc77ac5a),
	.w7(32'hbb0e9676),
	.w8(32'h3b08fd72),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb16b02),
	.w1(32'hbbde3297),
	.w2(32'h3b773201),
	.w3(32'hbb95c8d4),
	.w4(32'h3b39081f),
	.w5(32'h3bcce354),
	.w6(32'hbbb9eed5),
	.w7(32'h3b51f150),
	.w8(32'h3b6bc65e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba394acf),
	.w1(32'hbb44dc19),
	.w2(32'h3b372f08),
	.w3(32'hbb099d5c),
	.w4(32'hbb20f44d),
	.w5(32'h3bad4c2a),
	.w6(32'h39c41caf),
	.w7(32'h3aa73155),
	.w8(32'h3bad070f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ddeb9),
	.w1(32'hbbc5c662),
	.w2(32'h3a866223),
	.w3(32'hbb68c94d),
	.w4(32'hbb400b80),
	.w5(32'hbbb610aa),
	.w6(32'hbb9d08ac),
	.w7(32'hbadf630c),
	.w8(32'hba0f8c77),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1917da),
	.w1(32'h3bb44425),
	.w2(32'h3a56f085),
	.w3(32'hbb1d3626),
	.w4(32'hba2cc9a7),
	.w5(32'hbbc1d3dd),
	.w6(32'h3bf74bd4),
	.w7(32'h3c12bf63),
	.w8(32'hbbbed631),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbf581),
	.w1(32'hbad67452),
	.w2(32'h3b1440bc),
	.w3(32'h39cdaf23),
	.w4(32'h3b89dba3),
	.w5(32'h3aceb3a8),
	.w6(32'h3c4d7e39),
	.w7(32'h3b760501),
	.w8(32'h3ab7388a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb3557),
	.w1(32'hbaab3013),
	.w2(32'hba4cc8b2),
	.w3(32'hba4411a2),
	.w4(32'hbb191fda),
	.w5(32'hbac086b7),
	.w6(32'hba0e6ea0),
	.w7(32'hba847d0b),
	.w8(32'hbacb5b64),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba284e4a),
	.w1(32'hba7fd6ce),
	.w2(32'hba6fd363),
	.w3(32'hb9257e02),
	.w4(32'hba48384e),
	.w5(32'hba061c03),
	.w6(32'h3a726a06),
	.w7(32'h3a867190),
	.w8(32'hb99c565b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11ad93),
	.w1(32'hbaf44017),
	.w2(32'h3b585b23),
	.w3(32'hbb01241b),
	.w4(32'hbb443dd2),
	.w5(32'h3b92d258),
	.w6(32'hba74e4fb),
	.w7(32'hba9339c2),
	.w8(32'h3bba6030),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b530f15),
	.w1(32'h3b800372),
	.w2(32'h3b8f4c33),
	.w3(32'h3b19087e),
	.w4(32'h3b2e5d96),
	.w5(32'h3b2796a6),
	.w6(32'h3bc36391),
	.w7(32'h3b0d9c97),
	.w8(32'h3ae9cdb6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7969f9f),
	.w1(32'h3a1c7196),
	.w2(32'h3b21bc3a),
	.w3(32'h398c30d9),
	.w4(32'h39eb5a7c),
	.w5(32'h3b7c2e6a),
	.w6(32'h39d2e42e),
	.w7(32'hb917f892),
	.w8(32'h3ba3353c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4a7f3),
	.w1(32'h3a5c413d),
	.w2(32'h3b34d013),
	.w3(32'h3b19ab3f),
	.w4(32'h3ac6fb30),
	.w5(32'hba0e6f16),
	.w6(32'h3aee410e),
	.w7(32'h3b0b3435),
	.w8(32'hba701fb3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b261005),
	.w1(32'h3a0b6c1a),
	.w2(32'h3ab263c3),
	.w3(32'hba8b86ba),
	.w4(32'hbac296ed),
	.w5(32'hb9b38605),
	.w6(32'h3a3ed7c5),
	.w7(32'h3999a255),
	.w8(32'hba026fc0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a964c45),
	.w1(32'hb904ff24),
	.w2(32'h3a81e245),
	.w3(32'h3a775743),
	.w4(32'h3a26be47),
	.w5(32'hba2cb27b),
	.w6(32'hb8256fc0),
	.w7(32'hb94db558),
	.w8(32'hbab2a3b2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1db906),
	.w1(32'hb9e65978),
	.w2(32'h3a89d1cf),
	.w3(32'hba0168a0),
	.w4(32'h3a0945c8),
	.w5(32'hba9dc28a),
	.w6(32'hbaf3abbe),
	.w7(32'hba0d08a2),
	.w8(32'hba3ba46c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f09fea),
	.w1(32'hb8af9ddc),
	.w2(32'h390553a0),
	.w3(32'hba521261),
	.w4(32'hba317641),
	.w5(32'h3a31a67e),
	.w6(32'h3a7ace0d),
	.w7(32'h3a311f6c),
	.w8(32'h39d7451e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66ab0b),
	.w1(32'h39896c0c),
	.w2(32'h3a832286),
	.w3(32'h3882e769),
	.w4(32'hb9fbb96e),
	.w5(32'hbb341ebb),
	.w6(32'h38878812),
	.w7(32'hb9e015df),
	.w8(32'hbaafed23),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38573a2d),
	.w1(32'hb72ebf87),
	.w2(32'h386a4c6f),
	.w3(32'hbad2cca0),
	.w4(32'hbb2e4d44),
	.w5(32'hba8f1706),
	.w6(32'hb861d108),
	.w7(32'hbad31cc7),
	.w8(32'hba28750f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4330d5),
	.w1(32'hb9af60e4),
	.w2(32'hb94db6a1),
	.w3(32'hbad55631),
	.w4(32'hb802a11c),
	.w5(32'h38be77dd),
	.w6(32'hbad107cd),
	.w7(32'h39d2736b),
	.w8(32'h3acd58b9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba805f7d),
	.w1(32'hb9958c19),
	.w2(32'h3970928e),
	.w3(32'hb8ee0c8b),
	.w4(32'hbadab33e),
	.w5(32'hb9bab91d),
	.w6(32'h3a622817),
	.w7(32'h3a82ecc7),
	.w8(32'h3ae4794f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35a7fd),
	.w1(32'h395e0e2b),
	.w2(32'hb8f92b8e),
	.w3(32'hba2f6a7e),
	.w4(32'hba8da2ae),
	.w5(32'hba2713be),
	.w6(32'hb9f3f2f4),
	.w7(32'hbabf4768),
	.w8(32'h39e792b4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf0803),
	.w1(32'h3a8f0b63),
	.w2(32'h3b0d0887),
	.w3(32'h39b22ac6),
	.w4(32'h3a932db1),
	.w5(32'h398588fc),
	.w6(32'h3b6ab9a6),
	.w7(32'h39c19334),
	.w8(32'h3ab38e14),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e32761),
	.w1(32'hba559e20),
	.w2(32'h39b35191),
	.w3(32'hbb17893b),
	.w4(32'hbb137248),
	.w5(32'h3a5a38da),
	.w6(32'hbac466e2),
	.w7(32'hba9e17c3),
	.w8(32'h3a09553a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c53f09),
	.w1(32'h3a126611),
	.w2(32'h3a5d38e8),
	.w3(32'hb99db0b9),
	.w4(32'hba5fa48c),
	.w5(32'h39d028da),
	.w6(32'h3aa65bf9),
	.w7(32'hb8da7a26),
	.w8(32'h39794d04),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14a2e3),
	.w1(32'hb9ca28ee),
	.w2(32'hba29afe1),
	.w3(32'hba1f8665),
	.w4(32'hb9f8f071),
	.w5(32'h3a9644ad),
	.w6(32'hba6dbd81),
	.w7(32'hb98e34ed),
	.w8(32'hb9ee1956),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace2f3b),
	.w1(32'hba81057e),
	.w2(32'h38b6400c),
	.w3(32'h3a3ad895),
	.w4(32'hb95f79b3),
	.w5(32'hbb118622),
	.w6(32'h3aae65b6),
	.w7(32'h39d801a8),
	.w8(32'hba80747a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f7ced),
	.w1(32'hbab1e4d8),
	.w2(32'hbab5b887),
	.w3(32'hbb1cdd1e),
	.w4(32'hbb07bef0),
	.w5(32'hbb01d3da),
	.w6(32'hba17c2c9),
	.w7(32'hb9d8f5ac),
	.w8(32'hb9ab6573),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86401b),
	.w1(32'hb9f86bd5),
	.w2(32'h3a6f3d5a),
	.w3(32'hbb00e0fb),
	.w4(32'hba26b871),
	.w5(32'h3aa7cdfa),
	.w6(32'hbabd7a6d),
	.w7(32'hb995152a),
	.w8(32'h3b023766),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfd2d7),
	.w1(32'hb91f03bf),
	.w2(32'hb94aee86),
	.w3(32'hb9a7591d),
	.w4(32'hbae8f945),
	.w5(32'hb99f2c18),
	.w6(32'h3af76e90),
	.w7(32'hb98be36b),
	.w8(32'h3a6130a6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af19b48),
	.w1(32'h39163633),
	.w2(32'hb93dad2c),
	.w3(32'h3a8e80d1),
	.w4(32'hba809681),
	.w5(32'h3ac21e23),
	.w6(32'h3a8f3add),
	.w7(32'h3925a7af),
	.w8(32'hbaccca11),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08d4a8),
	.w1(32'hbae4f732),
	.w2(32'hbb09fa04),
	.w3(32'h3b5fde55),
	.w4(32'h39983250),
	.w5(32'hbb34f04f),
	.w6(32'h3ac30bfc),
	.w7(32'hbaa87d19),
	.w8(32'hba04da7a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39230f7e),
	.w1(32'hb98cf211),
	.w2(32'hba6696d3),
	.w3(32'hb9e389fc),
	.w4(32'hb969e2f2),
	.w5(32'h3b00ce7d),
	.w6(32'hb9d9bf48),
	.w7(32'hbaa4c2b0),
	.w8(32'h3a8dc7de),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9520772),
	.w1(32'hb73136fb),
	.w2(32'hb97852e5),
	.w3(32'h3afec12e),
	.w4(32'h3aa904d9),
	.w5(32'hb9fd2098),
	.w6(32'h3ae790c7),
	.w7(32'h38a7a2ed),
	.w8(32'hb949a9eb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98480ab),
	.w1(32'hbab99e14),
	.w2(32'hbaa81790),
	.w3(32'hb9cbb466),
	.w4(32'hba806d99),
	.w5(32'hbb08db92),
	.w6(32'h3abb8978),
	.w7(32'h3a0978c4),
	.w8(32'hbacd9555),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9b490),
	.w1(32'hba400717),
	.w2(32'hba53a52a),
	.w3(32'hba9a7730),
	.w4(32'hbab6f5f6),
	.w5(32'h388785ec),
	.w6(32'hb817f4e3),
	.w7(32'hba6b5a6e),
	.w8(32'h39c59f2b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3429dc),
	.w1(32'h3ad928da),
	.w2(32'h3a45314f),
	.w3(32'h39b511ed),
	.w4(32'h376c59dc),
	.w5(32'hbad17aee),
	.w6(32'h3a539cff),
	.w7(32'hb98abb3f),
	.w8(32'hba75779d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba925138),
	.w1(32'hb9a63979),
	.w2(32'hba87a087),
	.w3(32'hbaf45195),
	.w4(32'hbb1064db),
	.w5(32'hb763ca22),
	.w6(32'h39ba2b81),
	.w7(32'hbadf4373),
	.w8(32'hba90a26b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39afd251),
	.w1(32'h38d35716),
	.w2(32'hb93482d9),
	.w3(32'h3a508be1),
	.w4(32'hb995f75a),
	.w5(32'hb8e0b010),
	.w6(32'h3a9b9b9a),
	.w7(32'hba9b9e6d),
	.w8(32'h39b71db3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39452b31),
	.w1(32'h3a18534a),
	.w2(32'h3ada5369),
	.w3(32'h397b883b),
	.w4(32'h38ea7f40),
	.w5(32'hba1317c7),
	.w6(32'h3aba194b),
	.w7(32'hb9f4ee78),
	.w8(32'h396d893a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39923e08),
	.w1(32'h3839333c),
	.w2(32'h3a0c1a5c),
	.w3(32'hb9134f6d),
	.w4(32'h39d0213c),
	.w5(32'hb95b688a),
	.w6(32'hb9693072),
	.w7(32'h37ae80d6),
	.w8(32'hbacdbbfa),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a981936),
	.w1(32'hb99425e6),
	.w2(32'h3a03c60b),
	.w3(32'hba88b9db),
	.w4(32'hbab877aa),
	.w5(32'hba243cc5),
	.w6(32'hbb226d3b),
	.w7(32'hbb1c2ace),
	.w8(32'h39c8ec4d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba579a8c),
	.w1(32'h398d57a2),
	.w2(32'h34ccc5d9),
	.w3(32'hbabe0f85),
	.w4(32'hba8244bc),
	.w5(32'h39675d39),
	.w6(32'hb9afb0c1),
	.w7(32'h38d17c0d),
	.w8(32'h39d08aab),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27c38e),
	.w1(32'h3a8f18a8),
	.w2(32'h3a66a8dd),
	.w3(32'h3a12c3ed),
	.w4(32'hb9bb5976),
	.w5(32'h39b8b78a),
	.w6(32'h3b0ec4a5),
	.w7(32'h38ce529b),
	.w8(32'hba367f32),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43724c),
	.w1(32'hb9ba3767),
	.w2(32'h39caa952),
	.w3(32'hbb04b0ce),
	.w4(32'hbae9cbf2),
	.w5(32'h3a19ef81),
	.w6(32'hba40e5c8),
	.w7(32'hba09b2d1),
	.w8(32'h3ad0f8f0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b211857),
	.w1(32'h39dc05ee),
	.w2(32'hb9550e6c),
	.w3(32'hb86e6744),
	.w4(32'hba492795),
	.w5(32'hbac945f8),
	.w6(32'h3a8c316b),
	.w7(32'hb9b6d290),
	.w8(32'hba407fad),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba999c01),
	.w1(32'hb9f91609),
	.w2(32'h39c289a1),
	.w3(32'hbab1b91a),
	.w4(32'hba917cdc),
	.w5(32'h39da6821),
	.w6(32'hba04b936),
	.w7(32'hb9a4aed3),
	.w8(32'h3a4ed69c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a7b6a),
	.w1(32'hba5a25ce),
	.w2(32'hb9b089c5),
	.w3(32'hba69d29f),
	.w4(32'hba24184c),
	.w5(32'hb90f5051),
	.w6(32'h39f38fb6),
	.w7(32'hb8b0b977),
	.w8(32'hb9f51ca6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0e47c),
	.w1(32'h3ad52b46),
	.w2(32'h3b8b1b70),
	.w3(32'hbabd082a),
	.w4(32'h39824b40),
	.w5(32'hba4606ab),
	.w6(32'h3990134c),
	.w7(32'h356a1f0b),
	.w8(32'h3977f9a6),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38da0807),
	.w1(32'hb98e95ca),
	.w2(32'h38345103),
	.w3(32'hbae4dcf2),
	.w4(32'hbaa90bfc),
	.w5(32'hb9d91a35),
	.w6(32'hba3aaac2),
	.w7(32'hbad6593e),
	.w8(32'hb9f77338),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72cb56),
	.w1(32'hbb7f5c5b),
	.w2(32'hbb24ae47),
	.w3(32'hbb4b7ce5),
	.w4(32'hbafc9532),
	.w5(32'hbaea4b30),
	.w6(32'hbb04f01d),
	.w7(32'hbae94774),
	.w8(32'hb9ef5b2d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ce37d),
	.w1(32'h38329c41),
	.w2(32'h39994a95),
	.w3(32'h383c07d9),
	.w4(32'h3a3eaf68),
	.w5(32'h39ef54d1),
	.w6(32'hba6548c4),
	.w7(32'h3900f7b2),
	.w8(32'h3a6140f4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83ba6b8),
	.w1(32'hba1ea9b4),
	.w2(32'h394b4319),
	.w3(32'hb960f97a),
	.w4(32'h3a4f1c63),
	.w5(32'hba8d99ef),
	.w6(32'hb6708a5f),
	.w7(32'h3a51b471),
	.w8(32'hba274668),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f06f0),
	.w1(32'h3ab0c818),
	.w2(32'h3a2501b9),
	.w3(32'hbaa14071),
	.w4(32'hba36bfe1),
	.w5(32'hba1558db),
	.w6(32'h3a952160),
	.w7(32'hb9b291fe),
	.w8(32'hba36233e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87b6e5),
	.w1(32'hba95c5f9),
	.w2(32'hba5a9b3a),
	.w3(32'h39442277),
	.w4(32'hba142367),
	.w5(32'hbb05f8bc),
	.w6(32'hb9b231d3),
	.w7(32'hb9fa73be),
	.w8(32'hbac4d954),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebed2f),
	.w1(32'h38229985),
	.w2(32'h37935896),
	.w3(32'hbb109883),
	.w4(32'hba55ba23),
	.w5(32'hb99b9e01),
	.w6(32'h3a9f5748),
	.w7(32'h3a79cd18),
	.w8(32'hba7280fa),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c2a7f),
	.w1(32'h396c79ce),
	.w2(32'hbab6cb05),
	.w3(32'h3b833134),
	.w4(32'hbaf21cb2),
	.w5(32'hbb76d4af),
	.w6(32'h3b3fadc5),
	.w7(32'hbae0b1aa),
	.w8(32'hbb8de8fb),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c6055),
	.w1(32'hb774fcdc),
	.w2(32'h3889d5c5),
	.w3(32'hba234419),
	.w4(32'h394b0f53),
	.w5(32'h39eed4e4),
	.w6(32'hb9659faf),
	.w7(32'h3a23bcfc),
	.w8(32'h39e3f23c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c151a),
	.w1(32'h3ac0bc1f),
	.w2(32'h3b1a3527),
	.w3(32'h3a7a0317),
	.w4(32'h39eaaa6a),
	.w5(32'h399d2030),
	.w6(32'h3a3ea6a2),
	.w7(32'h3a85faa8),
	.w8(32'h39ff9364),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49f493),
	.w1(32'h39f9b5f1),
	.w2(32'h3b0cc0c3),
	.w3(32'h381c8566),
	.w4(32'h3a5eb08e),
	.w5(32'h3944b040),
	.w6(32'h3ad537f1),
	.w7(32'h3a6c2e97),
	.w8(32'h388ecc5c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca8720),
	.w1(32'hb8f71de2),
	.w2(32'h37958779),
	.w3(32'hba8ea9dc),
	.w4(32'hbaf2b39a),
	.w5(32'hba0a144f),
	.w6(32'h399cc388),
	.w7(32'hba4803e6),
	.w8(32'hbb1098e6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939b37e),
	.w1(32'hb954f61f),
	.w2(32'h3aa03c61),
	.w3(32'hbabc78be),
	.w4(32'hbb21a949),
	.w5(32'h3900454d),
	.w6(32'h3aa7e29e),
	.w7(32'hbab9df41),
	.w8(32'h392957ca),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398de41d),
	.w1(32'hb9c46b00),
	.w2(32'h39df1b8c),
	.w3(32'h39aa7032),
	.w4(32'h3a08032a),
	.w5(32'h3a0c49fe),
	.w6(32'hb903b4a8),
	.w7(32'h3a20faf6),
	.w8(32'h3aa667c7),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944c101),
	.w1(32'hba8aabe8),
	.w2(32'h3a2a1d4d),
	.w3(32'hbaeba7cd),
	.w4(32'hb9853a61),
	.w5(32'hbb031889),
	.w6(32'hbaad9cc1),
	.w7(32'hba032270),
	.w8(32'hba95e28b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62c0c0),
	.w1(32'hb99fd4b8),
	.w2(32'hbac85a01),
	.w3(32'hbb1c1cec),
	.w4(32'hbb220197),
	.w5(32'hba7f71d9),
	.w6(32'hbac3ab9e),
	.w7(32'hbb0f0da2),
	.w8(32'hbaeccfdf),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe68a7),
	.w1(32'hbb0c8c45),
	.w2(32'hba10e396),
	.w3(32'h39689f39),
	.w4(32'h39673760),
	.w5(32'h3a2e5862),
	.w6(32'hba255565),
	.w7(32'h3ae37b32),
	.w8(32'h3ade0eca),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa648d7),
	.w1(32'hbae3d53a),
	.w2(32'hbabbc685),
	.w3(32'hbad32585),
	.w4(32'hbb265d9c),
	.w5(32'h3a69a474),
	.w6(32'hba7560b4),
	.w7(32'hba4a8e1d),
	.w8(32'h3a102fbd),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393129d2),
	.w1(32'h3a375881),
	.w2(32'hba816dc7),
	.w3(32'h3b1e6064),
	.w4(32'h3aa93fc2),
	.w5(32'h39a384d3),
	.w6(32'h3b5772fc),
	.w7(32'h39ae0602),
	.w8(32'h3aa74046),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77cd8a),
	.w1(32'h3b4ea7e8),
	.w2(32'h3b14af03),
	.w3(32'h3a5b729e),
	.w4(32'h38966134),
	.w5(32'h3a29b5ab),
	.w6(32'h3a07576c),
	.w7(32'hbabbf5ca),
	.w8(32'h3973bf72),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b133dc4),
	.w1(32'h3abbdc1f),
	.w2(32'hb88b84c8),
	.w3(32'h3a2b138b),
	.w4(32'hb9a38ebf),
	.w5(32'hba7bc6d9),
	.w6(32'h39ab6b44),
	.w7(32'hba401177),
	.w8(32'hbac292c8),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb191447),
	.w1(32'hbb0788ed),
	.w2(32'hba68cfb3),
	.w3(32'hba9cc7ab),
	.w4(32'hba74d10d),
	.w5(32'hba75a664),
	.w6(32'hba4e858d),
	.w7(32'hba1b5ad4),
	.w8(32'hbae75ebe),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9770c7b),
	.w1(32'hb8b4fd60),
	.w2(32'h39ee25c5),
	.w3(32'hbab9774b),
	.w4(32'hbafd28e1),
	.w5(32'hbb056afa),
	.w6(32'hbad27687),
	.w7(32'hba914554),
	.w8(32'hbae6c53d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c1323),
	.w1(32'hba94337f),
	.w2(32'hbac30714),
	.w3(32'hbb3223cf),
	.w4(32'hbb030f39),
	.w5(32'h39609bd1),
	.w6(32'hba449876),
	.w7(32'hba8e3fb6),
	.w8(32'hba54a756),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985f0d7),
	.w1(32'h39e3d09a),
	.w2(32'hbb0d233b),
	.w3(32'h35b92a83),
	.w4(32'hba2ad2b1),
	.w5(32'hbab3186e),
	.w6(32'h3a22183d),
	.w7(32'hba23f969),
	.w8(32'hba221fe8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da9948),
	.w1(32'hba96489d),
	.w2(32'hb939349f),
	.w3(32'hbae92f5d),
	.w4(32'hbaa34942),
	.w5(32'hba1af8e5),
	.w6(32'hbabb2cc7),
	.w7(32'hba0868bc),
	.w8(32'hb9aaa455),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9171733),
	.w1(32'h3a0ef18f),
	.w2(32'hb817421b),
	.w3(32'h3a167e91),
	.w4(32'hba14a42b),
	.w5(32'h39dc7b9f),
	.w6(32'h3a45d2bc),
	.w7(32'hba09a8c9),
	.w8(32'h3abb62b6),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a967cdb),
	.w1(32'h3a9de908),
	.w2(32'h3b2ae847),
	.w3(32'hb990da0b),
	.w4(32'hba05bcad),
	.w5(32'h378b22c8),
	.w6(32'h3966d25c),
	.w7(32'h3a808266),
	.w8(32'h39a1f454),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399cf649),
	.w1(32'h3a17a7e5),
	.w2(32'h3b2805fe),
	.w3(32'hba7336ca),
	.w4(32'h3af76a3b),
	.w5(32'h3a6c42c4),
	.w6(32'hba68a42c),
	.w7(32'h3aabdcff),
	.w8(32'h3ae4deb4),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f44b98),
	.w1(32'hba2ff286),
	.w2(32'h39ff48f6),
	.w3(32'hbab89d45),
	.w4(32'hba8714fb),
	.w5(32'hba1628ca),
	.w6(32'hba6571c1),
	.w7(32'hb8c24d7b),
	.w8(32'h3a4325d0),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a63e8),
	.w1(32'h3ace4c42),
	.w2(32'h3b51ef00),
	.w3(32'hba4e22f4),
	.w4(32'h3a42778f),
	.w5(32'h3a1d83cc),
	.w6(32'hb9bb7709),
	.w7(32'h3b1aee3e),
	.w8(32'hb9ea0d2d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad40085),
	.w1(32'hbb0dca2d),
	.w2(32'hbae14e95),
	.w3(32'hbb15df6e),
	.w4(32'hb9e88f3e),
	.w5(32'hbab19390),
	.w6(32'hb9c807ae),
	.w7(32'hbac073d8),
	.w8(32'hb9aec611),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90c62b),
	.w1(32'h3af5e13a),
	.w2(32'h3a781232),
	.w3(32'h3a2ee2c9),
	.w4(32'hbb462a27),
	.w5(32'hbb6acb96),
	.w6(32'h3a92f2a9),
	.w7(32'hbb265c05),
	.w8(32'hbb95c7a6),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8adaa),
	.w1(32'hbaa5198f),
	.w2(32'h3a9111a4),
	.w3(32'hba283ca3),
	.w4(32'hbaf8c0a0),
	.w5(32'hba8ea0d3),
	.w6(32'h3aabf666),
	.w7(32'hb9779ffa),
	.w8(32'hba868c0f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d42321),
	.w1(32'h39723e5d),
	.w2(32'h3ad8ed5b),
	.w3(32'hb91c4e0b),
	.w4(32'h3a009086),
	.w5(32'h3b247d85),
	.w6(32'h39bce134),
	.w7(32'hba21d76b),
	.w8(32'h3b0a6ac8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24a566),
	.w1(32'h3af793d4),
	.w2(32'h3a8f98ef),
	.w3(32'h3aa27f8a),
	.w4(32'h3a93c4e2),
	.w5(32'hbac6077f),
	.w6(32'h3a5ca53b),
	.w7(32'h39f3f60d),
	.w8(32'hba09cc45),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba223891),
	.w1(32'h3a8aeb08),
	.w2(32'h3a521ae5),
	.w3(32'hbad3faec),
	.w4(32'hb9a04508),
	.w5(32'h3af669e1),
	.w6(32'hba16c771),
	.w7(32'hb9f11c69),
	.w8(32'h3afe3b16),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab205a1),
	.w1(32'h3a072f71),
	.w2(32'h3ac471cd),
	.w3(32'h3a0d8507),
	.w4(32'h3ab758fc),
	.w5(32'h3a7c998c),
	.w6(32'hb89ce60c),
	.w7(32'h3a93885b),
	.w8(32'h37d75656),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a149b9),
	.w1(32'h392a2b55),
	.w2(32'h3921b973),
	.w3(32'hbae3c387),
	.w4(32'hbb1b99a5),
	.w5(32'hb99aeb51),
	.w6(32'hb9ecef54),
	.w7(32'hb9298bbe),
	.w8(32'hba7634d3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fcebb),
	.w1(32'hbac9b82a),
	.w2(32'hb938e299),
	.w3(32'hba9fe710),
	.w4(32'hbab074fd),
	.w5(32'h3abdd3a4),
	.w6(32'hba7a67aa),
	.w7(32'hba4584b5),
	.w8(32'h3a7c2869),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63ee44),
	.w1(32'hb9d10b36),
	.w2(32'h39e84d91),
	.w3(32'h3ae52ac7),
	.w4(32'h3a8feb29),
	.w5(32'hbabc8bed),
	.w6(32'h3b0bd827),
	.w7(32'h3a0c0222),
	.w8(32'hbaf388f3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d0b5f),
	.w1(32'hba983bbd),
	.w2(32'hb9072bfb),
	.w3(32'h3967202c),
	.w4(32'hba8d0996),
	.w5(32'hb797ed20),
	.w6(32'h3a824a9d),
	.w7(32'h395ef5ee),
	.w8(32'h39cf2390),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6c58a),
	.w1(32'h390b4dfc),
	.w2(32'hba4734c5),
	.w3(32'h3ab1a701),
	.w4(32'h3a8bfb60),
	.w5(32'hbb0070dd),
	.w6(32'h3a6cf4a3),
	.w7(32'h39e2345b),
	.w8(32'hbad20f40),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba663be1),
	.w1(32'hba848077),
	.w2(32'hba71fc1e),
	.w3(32'hbb0ada3f),
	.w4(32'hbaeb8250),
	.w5(32'hbaafad04),
	.w6(32'hba8ce876),
	.w7(32'hb91d60a6),
	.w8(32'hbaa3f219),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3257e),
	.w1(32'hba9676d4),
	.w2(32'hb8a7e91e),
	.w3(32'hbadaea29),
	.w4(32'hba2953e7),
	.w5(32'h39e3b6e2),
	.w6(32'hbaa57b59),
	.w7(32'hb9b5c427),
	.w8(32'h3a836587),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5585c7),
	.w1(32'h3a585c65),
	.w2(32'h39cbdec9),
	.w3(32'h3a7af5b1),
	.w4(32'h3a44f8e7),
	.w5(32'h3a9e7447),
	.w6(32'h3a3fb533),
	.w7(32'h3982d450),
	.w8(32'h3a92f4b5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade60c7),
	.w1(32'h3a10196a),
	.w2(32'h3ac89516),
	.w3(32'h39377458),
	.w4(32'h3a97be6e),
	.w5(32'h3a1914f9),
	.w6(32'hb9f4d66e),
	.w7(32'h3a40e18a),
	.w8(32'hb9e2fe6e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c234105),
	.w1(32'h3b442dd1),
	.w2(32'hba96b76a),
	.w3(32'h3b05d7ba),
	.w4(32'hbb4e8dd8),
	.w5(32'hbba17b98),
	.w6(32'h3a92574a),
	.w7(32'hbc092c34),
	.w8(32'hbbe4ffc4),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29b6e8),
	.w1(32'h3950ff4c),
	.w2(32'h38d7ac08),
	.w3(32'hba933add),
	.w4(32'hba590061),
	.w5(32'hba35cf09),
	.w6(32'hb985a145),
	.w7(32'hbaaee02f),
	.w8(32'hba3c5a06),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ea7cf),
	.w1(32'h3a1678b2),
	.w2(32'h3839c6cd),
	.w3(32'h390033ea),
	.w4(32'hb9a5b4c2),
	.w5(32'hba60af36),
	.w6(32'h3a38f578),
	.w7(32'hb9dc3275),
	.w8(32'hba42a166),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3710797d),
	.w1(32'hb9be8da5),
	.w2(32'hb991148a),
	.w3(32'hb9e22d74),
	.w4(32'hbb0e4d3a),
	.w5(32'hbaf9bbad),
	.w6(32'h3ade3c00),
	.w7(32'h39d95dba),
	.w8(32'hbaf421b6),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c9fe1),
	.w1(32'hba670b3d),
	.w2(32'h372666ee),
	.w3(32'hbad4d785),
	.w4(32'hba5e437f),
	.w5(32'hba9c2115),
	.w6(32'hbb1393d7),
	.w7(32'hba1213e8),
	.w8(32'hba03e3ec),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d787bb),
	.w1(32'hb8d71c9e),
	.w2(32'hbacb12d7),
	.w3(32'hba63daed),
	.w4(32'hba92ba1c),
	.w5(32'h3a9ec70e),
	.w6(32'hba3e3e49),
	.w7(32'hb9a238f5),
	.w8(32'h3aa73971),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ddb9d),
	.w1(32'h3820e136),
	.w2(32'h38d80a7f),
	.w3(32'h3b1648ee),
	.w4(32'h3a92d35d),
	.w5(32'hba1de14b),
	.w6(32'h3b5ee795),
	.w7(32'h3a00d09a),
	.w8(32'h3922dba3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4f1bc),
	.w1(32'h385d9e6f),
	.w2(32'h3ab231ba),
	.w3(32'hb959a63f),
	.w4(32'hb9f57caf),
	.w5(32'hbb04c270),
	.w6(32'h3abb5643),
	.w7(32'h3ab2249e),
	.w8(32'h3aa755e8),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a3317),
	.w1(32'h398b8b4a),
	.w2(32'hb8bf660a),
	.w3(32'hba8daf93),
	.w4(32'hbb166593),
	.w5(32'hbb2c3aaa),
	.w6(32'hba3686c4),
	.w7(32'hbb3008f4),
	.w8(32'hbb2b178b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a173adb),
	.w1(32'hba9803f9),
	.w2(32'hba7205de),
	.w3(32'hba8bf7bd),
	.w4(32'hba626f74),
	.w5(32'hbb763c86),
	.w6(32'hbb0b7501),
	.w7(32'hba07aa3e),
	.w8(32'hbb8349dd),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c29679),
	.w1(32'hbad9b87d),
	.w2(32'h3a36b56d),
	.w3(32'hbb8ff366),
	.w4(32'hbb3619e2),
	.w5(32'h3af5f658),
	.w6(32'hbb880471),
	.w7(32'hbaf4dea7),
	.w8(32'h3a0edf97),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee4c45),
	.w1(32'h39c6897c),
	.w2(32'h3a7ecc19),
	.w3(32'h3aa03b09),
	.w4(32'h3a9c2a07),
	.w5(32'hba2c8251),
	.w6(32'h3a055795),
	.w7(32'h3a5dad0f),
	.w8(32'h38a7e2e8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba825c0c),
	.w1(32'hba52fa29),
	.w2(32'h3adfc2ce),
	.w3(32'hba12c014),
	.w4(32'hba35e33a),
	.w5(32'h39e2f1d3),
	.w6(32'hb8e47687),
	.w7(32'h39006677),
	.w8(32'hbaba5717),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f13d2),
	.w1(32'h3a78cd76),
	.w2(32'h3a843378),
	.w3(32'h3a993c3e),
	.w4(32'h3a896523),
	.w5(32'hbab56f9d),
	.w6(32'hba66f8cc),
	.w7(32'hbaee2935),
	.w8(32'hba82614c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa90aea),
	.w1(32'hba1e0288),
	.w2(32'hb991104a),
	.w3(32'h378e2f1a),
	.w4(32'hb9d60043),
	.w5(32'h3921dde2),
	.w6(32'h3a14c0ec),
	.w7(32'hb9961303),
	.w8(32'h3959cf08),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac40588),
	.w1(32'hb9bf3d25),
	.w2(32'h39de683c),
	.w3(32'h3a3b67bb),
	.w4(32'hba9963f8),
	.w5(32'hbb24cf16),
	.w6(32'h3b024c76),
	.w7(32'h378f70c3),
	.w8(32'hbb059e8d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90fe23),
	.w1(32'hba45decd),
	.w2(32'hba27f5c0),
	.w3(32'hba9c0fdf),
	.w4(32'hba8a9302),
	.w5(32'hb90cab95),
	.w6(32'hba584b55),
	.w7(32'hba88f6d7),
	.w8(32'h3ac8a064),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d63ce),
	.w1(32'h388b7c2f),
	.w2(32'h3b1d7fc0),
	.w3(32'h39041a96),
	.w4(32'h3a455053),
	.w5(32'h3a87b5f3),
	.w6(32'h3b0729a2),
	.w7(32'h39f908fd),
	.w8(32'hb8b1c97a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad69382),
	.w1(32'hbad849e5),
	.w2(32'hba1535e5),
	.w3(32'hba6c8999),
	.w4(32'hba8de28a),
	.w5(32'h386048fa),
	.w6(32'hba9be4f9),
	.w7(32'hbac05aad),
	.w8(32'h3ad09f8b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1fde8),
	.w1(32'h3a5e644d),
	.w2(32'h3b1a7652),
	.w3(32'h3a4564c8),
	.w4(32'h38f1ef32),
	.w5(32'hb9c73d7d),
	.w6(32'h3b11d038),
	.w7(32'h39b8247b),
	.w8(32'h39d35450),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9651c2),
	.w1(32'h3ae0c339),
	.w2(32'h3ad17856),
	.w3(32'h3996128a),
	.w4(32'hb9a00b7a),
	.w5(32'h3b495fee),
	.w6(32'h3ab0737e),
	.w7(32'hb9e02e2a),
	.w8(32'h3ba0af5e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c483182),
	.w1(32'h3bdd1657),
	.w2(32'h3b9a7c94),
	.w3(32'h3bb85d94),
	.w4(32'h3b0d710a),
	.w5(32'hbb14e4de),
	.w6(32'h3bcce4f9),
	.w7(32'h3ab7720a),
	.w8(32'hbb6354a1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4063af),
	.w1(32'h3a302e28),
	.w2(32'h3902c099),
	.w3(32'hb9baa55c),
	.w4(32'hb7e9b9c2),
	.w5(32'h392e51fd),
	.w6(32'h3a02b563),
	.w7(32'h3a6e2f1b),
	.w8(32'hba69c55f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1fc29),
	.w1(32'hb8b20afa),
	.w2(32'hb9c38dd8),
	.w3(32'hba14bd1e),
	.w4(32'hba8a9e19),
	.w5(32'h3a2eea74),
	.w6(32'h3a0333df),
	.w7(32'hba6b21fa),
	.w8(32'h3a2decc6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae89253),
	.w1(32'h3a3613a6),
	.w2(32'h3aecb2eb),
	.w3(32'h3aa1aaff),
	.w4(32'h3a8ba7ec),
	.w5(32'hb896c635),
	.w6(32'h3a2da571),
	.w7(32'h3a16f706),
	.w8(32'h3a424afc),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ec6df),
	.w1(32'h3a4d5544),
	.w2(32'h3b1c3555),
	.w3(32'hbb23ce97),
	.w4(32'hba3fac48),
	.w5(32'h39f27ddf),
	.w6(32'h3a89a2ca),
	.w7(32'hba348346),
	.w8(32'h3a2f746d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a845b5f),
	.w1(32'h3a003f31),
	.w2(32'h3a76913c),
	.w3(32'h3a8f7dd7),
	.w4(32'hba290cfb),
	.w5(32'h39441a5d),
	.w6(32'h3af366c4),
	.w7(32'hb9c91241),
	.w8(32'hb9ba2319),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ecf29),
	.w1(32'h3a54f949),
	.w2(32'h3ab5f6ff),
	.w3(32'hba4faf80),
	.w4(32'hba504464),
	.w5(32'h39efdd11),
	.w6(32'hb9aea369),
	.w7(32'h3661901b),
	.w8(32'h3986f9ba),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1887a),
	.w1(32'hba7d7a81),
	.w2(32'hba7c140b),
	.w3(32'h3adb0a53),
	.w4(32'hb78869ec),
	.w5(32'hbaa64986),
	.w6(32'h3ac842d0),
	.w7(32'h3993abb0),
	.w8(32'hba8820e9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1282a),
	.w1(32'h39ab321b),
	.w2(32'hb9fba030),
	.w3(32'hbaa921a7),
	.w4(32'hba23fd9d),
	.w5(32'hb9f62e40),
	.w6(32'hb9cccc62),
	.w7(32'hba4652b9),
	.w8(32'h3aa78d63),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12e709),
	.w1(32'hb9820afa),
	.w2(32'hb8fd121c),
	.w3(32'hb8b18030),
	.w4(32'h38762635),
	.w5(32'hb9a504b9),
	.w6(32'hb9dd89f8),
	.w7(32'h3a44cbd3),
	.w8(32'h39284e9a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bceb60c),
	.w1(32'h3b2234ca),
	.w2(32'hb9a09084),
	.w3(32'h3af9c4ce),
	.w4(32'hbad665b6),
	.w5(32'hba594e72),
	.w6(32'h3afc2b31),
	.w7(32'hbb165c16),
	.w8(32'hbb06651b),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2e422),
	.w1(32'h38aa0f25),
	.w2(32'h3a0c3056),
	.w3(32'h3ab38813),
	.w4(32'h3929b06f),
	.w5(32'hbaf4bf18),
	.w6(32'h3a96bd1a),
	.w7(32'h3ab0b8ef),
	.w8(32'hb93953ac),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39afefc2),
	.w1(32'hba5718bd),
	.w2(32'hb8541c10),
	.w3(32'hbaa88184),
	.w4(32'hbaaeab28),
	.w5(32'hbace950f),
	.w6(32'h3a288c5b),
	.w7(32'hba5d6a1f),
	.w8(32'h3a1d1652),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc2b04),
	.w1(32'h3ad3f3cf),
	.w2(32'h3b0e6983),
	.w3(32'hba8cd67b),
	.w4(32'hba9df2e9),
	.w5(32'h3a7b2e8f),
	.w6(32'h386270c7),
	.w7(32'hb9a259d1),
	.w8(32'h3a031e56),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba525a11),
	.w1(32'hba7a2a1a),
	.w2(32'hb9692a08),
	.w3(32'hba57b7ac),
	.w4(32'hba106f1a),
	.w5(32'h3a1c2ffb),
	.w6(32'hbacf7463),
	.w7(32'hb93720c6),
	.w8(32'h3a122505),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1302b),
	.w1(32'h3b0482c1),
	.w2(32'h3b366374),
	.w3(32'hba67ae01),
	.w4(32'hb94aee10),
	.w5(32'h3b2019c0),
	.w6(32'hba8592c1),
	.w7(32'h3a5f0831),
	.w8(32'h3b49ef1d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad1684),
	.w1(32'h3a8e0a31),
	.w2(32'h3933b815),
	.w3(32'h3ae3a91e),
	.w4(32'h39e9aa27),
	.w5(32'h3a957e11),
	.w6(32'h3b299db0),
	.w7(32'h3a491d80),
	.w8(32'h3aa43f70),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67c725),
	.w1(32'h3a2940d6),
	.w2(32'hba568a23),
	.w3(32'h3a817bb1),
	.w4(32'h3abfb42b),
	.w5(32'h3bc3c2ab),
	.w6(32'h3a9e67ef),
	.w7(32'h39df971d),
	.w8(32'h3b1e636f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e45c61),
	.w1(32'hbb7876d8),
	.w2(32'hbb845965),
	.w3(32'h3b24c80b),
	.w4(32'hbacecb19),
	.w5(32'hbc057c84),
	.w6(32'hbbfc0464),
	.w7(32'hbac042e1),
	.w8(32'h3b08c9b8),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c229457),
	.w1(32'h3bf8c415),
	.w2(32'hbb83507f),
	.w3(32'h3b7028a8),
	.w4(32'h3c023d5e),
	.w5(32'h3c89899e),
	.w6(32'h3c68849b),
	.w7(32'h3bcd4f52),
	.w8(32'hba6fbf00),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39c0dd),
	.w1(32'hbc9fad67),
	.w2(32'hbc311dbf),
	.w3(32'h3ca386a4),
	.w4(32'h3c7cf551),
	.w5(32'h3bdc6a7d),
	.w6(32'hbb2bd0e9),
	.w7(32'hbb7daa50),
	.w8(32'hbba4a38e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5bec0),
	.w1(32'h3b5c1614),
	.w2(32'h3a77b8f3),
	.w3(32'h3b92632e),
	.w4(32'h3c18d0ec),
	.w5(32'h3a866b07),
	.w6(32'h3b6cde12),
	.w7(32'hbc40830c),
	.w8(32'h3b41c2df),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1d91f),
	.w1(32'h3b7c4b05),
	.w2(32'hbb0549c1),
	.w3(32'h39dced4c),
	.w4(32'h3993fac8),
	.w5(32'hbc857b07),
	.w6(32'h3bc89cb0),
	.w7(32'h36f6bb14),
	.w8(32'h3ba8edf2),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b5bbc),
	.w1(32'h3d03d33b),
	.w2(32'h3c6e6081),
	.w3(32'hbd0532d1),
	.w4(32'hbcb91183),
	.w5(32'h3c3c214a),
	.w6(32'hb9ae5867),
	.w7(32'hbb972f63),
	.w8(32'h3b38156d),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9afaa),
	.w1(32'hbcc82aba),
	.w2(32'hbc7a61a5),
	.w3(32'h3c2776b1),
	.w4(32'h3aeca0ed),
	.w5(32'hbb81f2ab),
	.w6(32'h3a9c5b22),
	.w7(32'h3bcc9001),
	.w8(32'h3b333c3e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80fc27),
	.w1(32'h3bcc05b7),
	.w2(32'hbaf4a322),
	.w3(32'hbae71daf),
	.w4(32'hbb9861b8),
	.w5(32'hbbc5a0aa),
	.w6(32'hbb9d1e72),
	.w7(32'hbbd048cd),
	.w8(32'hbbff868c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc928728),
	.w1(32'hbca28ebf),
	.w2(32'hbbc6a99b),
	.w3(32'hbb7d6d86),
	.w4(32'hbc556135),
	.w5(32'h3a7abbcc),
	.w6(32'hbbfb0e85),
	.w7(32'hbc808d33),
	.w8(32'h3b9c207f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b1688),
	.w1(32'hbb626340),
	.w2(32'hbba7c4ce),
	.w3(32'h3a1e0929),
	.w4(32'hba51d48b),
	.w5(32'h3bf3f15c),
	.w6(32'h3b792ca9),
	.w7(32'h39c3a777),
	.w8(32'hbb5557ec),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf80a81),
	.w1(32'hbc32937c),
	.w2(32'hbbc6813f),
	.w3(32'h3b901076),
	.w4(32'h3ac472c5),
	.w5(32'hbac0fec6),
	.w6(32'hbc49d5ea),
	.w7(32'hbb1f0827),
	.w8(32'hbb18f42f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8adc79),
	.w1(32'hbb8ea00f),
	.w2(32'hbbce5f02),
	.w3(32'hbb75d0e2),
	.w4(32'hba8f000f),
	.w5(32'h39ea3ed4),
	.w6(32'hbbd0b479),
	.w7(32'hbb75a125),
	.w8(32'h3c17f5ee),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04804e),
	.w1(32'hbc4c43ee),
	.w2(32'hbc32c19e),
	.w3(32'h3bb7b8f5),
	.w4(32'h3b321210),
	.w5(32'hbb66a752),
	.w6(32'h3ba77819),
	.w7(32'h3980dfb7),
	.w8(32'h3b0779bc),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dfaf3),
	.w1(32'h38949910),
	.w2(32'h3a7e12e7),
	.w3(32'hbac26e94),
	.w4(32'hbaf98079),
	.w5(32'h398026f6),
	.w6(32'h3bea315d),
	.w7(32'h3a8e47fb),
	.w8(32'h3adabb0a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3dad4),
	.w1(32'hbb857c03),
	.w2(32'hbbdfc893),
	.w3(32'hbab9adf6),
	.w4(32'hbaeecf64),
	.w5(32'h39b0d829),
	.w6(32'hbbac0091),
	.w7(32'hbb245923),
	.w8(32'hbaec6d60),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e4fca),
	.w1(32'h3b1dd53c),
	.w2(32'hb9ba6a87),
	.w3(32'hba98f92f),
	.w4(32'hba421e09),
	.w5(32'hb9aee6df),
	.w6(32'h3c37a90e),
	.w7(32'h3ab98492),
	.w8(32'hbc03608c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95fd46),
	.w1(32'hbc2f4067),
	.w2(32'hbc33ea3c),
	.w3(32'h3b6f5d27),
	.w4(32'hba5d240e),
	.w5(32'h39ac83d8),
	.w6(32'hbc3ef38a),
	.w7(32'hbc060333),
	.w8(32'h3b2337dc),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f0300),
	.w1(32'h3b8454f4),
	.w2(32'hbb7ec550),
	.w3(32'hbbbd4586),
	.w4(32'hba27def5),
	.w5(32'h3ae517dd),
	.w6(32'h3c16c4e4),
	.w7(32'h3b1bb375),
	.w8(32'hba146977),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb894388),
	.w1(32'hba8f6194),
	.w2(32'h3a8093cb),
	.w3(32'h3b58ef13),
	.w4(32'h3afc9a39),
	.w5(32'h3c89a872),
	.w6(32'hbb7ed456),
	.w7(32'hbae48a65),
	.w8(32'h3bf3c702),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe62c41),
	.w1(32'hbc207358),
	.w2(32'h3a5ef3ce),
	.w3(32'h3c453e7a),
	.w4(32'h3a8adb05),
	.w5(32'h3a907225),
	.w6(32'h3c555277),
	.w7(32'h3c8679dc),
	.w8(32'h3bada576),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5ecca),
	.w1(32'h3af9c6da),
	.w2(32'h3c078763),
	.w3(32'h3b69839f),
	.w4(32'hba2a3344),
	.w5(32'hbbdd4f2b),
	.w6(32'h3bb95f45),
	.w7(32'h3b1a0dfe),
	.w8(32'h3ab9fb69),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b688b3b),
	.w1(32'h3c0f9e48),
	.w2(32'h3bb99120),
	.w3(32'hbbc8b606),
	.w4(32'hbc10ff13),
	.w5(32'h3a82fbb3),
	.w6(32'hbaa0a34b),
	.w7(32'hbadfd391),
	.w8(32'h3a08f46b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996336f),
	.w1(32'hbb985d60),
	.w2(32'hbbea5cbd),
	.w3(32'hbc04e689),
	.w4(32'hbbd92ab8),
	.w5(32'hbc2e27b2),
	.w6(32'hbb7f8133),
	.w7(32'hbbac4cd3),
	.w8(32'hbba77e28),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b812455),
	.w1(32'h3be24cf2),
	.w2(32'h3b57d901),
	.w3(32'hbc5c61cf),
	.w4(32'hbc1c500f),
	.w5(32'hbb20d00c),
	.w6(32'hbb50c2f0),
	.w7(32'h3bba5a54),
	.w8(32'h39fe30e2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840a6b),
	.w1(32'h3c11c6fd),
	.w2(32'h3b4ef641),
	.w3(32'h3ba40c16),
	.w4(32'h3c1e49ce),
	.w5(32'hbbea9abb),
	.w6(32'h3bc92473),
	.w7(32'hbbda2122),
	.w8(32'hb9d10ec9),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed72e2),
	.w1(32'h3c0f2625),
	.w2(32'h3b8175b8),
	.w3(32'hbc097e99),
	.w4(32'hbafac8c9),
	.w5(32'hbab74e84),
	.w6(32'hbb3dd697),
	.w7(32'hbb2e36b0),
	.w8(32'h3bbe6c1f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14d5de),
	.w1(32'h3c94e2fa),
	.w2(32'h3b90deae),
	.w3(32'h3ae68efe),
	.w4(32'h391d3b0f),
	.w5(32'h3b3e76c1),
	.w6(32'h3c4827eb),
	.w7(32'h3af78430),
	.w8(32'h3a6fd095),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79fda8),
	.w1(32'h3bc13c37),
	.w2(32'h3b946c5d),
	.w3(32'hbac5cc1c),
	.w4(32'hbb8e8ec9),
	.w5(32'hbb089a6e),
	.w6(32'h3c875b1c),
	.w7(32'h3b4a15a6),
	.w8(32'hbb82a0f2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58e817),
	.w1(32'h38a64591),
	.w2(32'hbb3959e8),
	.w3(32'hbabfb4a9),
	.w4(32'hbb573abd),
	.w5(32'hbaffcbf7),
	.w6(32'hbba26476),
	.w7(32'hbbb39675),
	.w8(32'h38e2a802),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba28bf7),
	.w1(32'hbc2e5509),
	.w2(32'hbbec1f35),
	.w3(32'h3b390fc8),
	.w4(32'hbb54bf9e),
	.w5(32'hbbf7d6f2),
	.w6(32'hbb713542),
	.w7(32'hbc18d46a),
	.w8(32'hbbd66a6a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule