module layer_10_featuremap_188(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ad47c3),
	.w1(32'h391d2f66),
	.w2(32'hb91b794c),
	.w3(32'h38a5ee21),
	.w4(32'h399cad53),
	.w5(32'h393b959f),
	.w6(32'h39142e5f),
	.w7(32'h38eb62c3),
	.w8(32'h37f20788),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1792de),
	.w1(32'h3b8ba040),
	.w2(32'h3ad9cd88),
	.w3(32'h3b8de9c7),
	.w4(32'h3aa05077),
	.w5(32'hba11fc57),
	.w6(32'h3b56fc8f),
	.w7(32'hba24e3f7),
	.w8(32'hb7292939),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3894eb76),
	.w1(32'h3823fb89),
	.w2(32'h38fd9978),
	.w3(32'hb8183c88),
	.w4(32'hb91593cf),
	.w5(32'hb97b1d4c),
	.w6(32'h388cdeed),
	.w7(32'h38af54b5),
	.w8(32'h3912d8d3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da430a),
	.w1(32'h39bbb814),
	.w2(32'hba726d73),
	.w3(32'h38a3bd20),
	.w4(32'h39e78503),
	.w5(32'h3a05138d),
	.w6(32'hb8974d7c),
	.w7(32'h37f462a4),
	.w8(32'h39514cad),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a595149),
	.w1(32'h3a8f4bec),
	.w2(32'hb8ec6440),
	.w3(32'h3ab252f7),
	.w4(32'h3ac104d6),
	.w5(32'h399be7e7),
	.w6(32'h3afc6401),
	.w7(32'h3ad67c60),
	.w8(32'h3a7da07b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bd04a0),
	.w1(32'h392361c6),
	.w2(32'h37e6e503),
	.w3(32'h37d925e0),
	.w4(32'h39181082),
	.w5(32'h380e5a47),
	.w6(32'h398d6c4e),
	.w7(32'h38ac4e55),
	.w8(32'h38ac7ea6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef325b),
	.w1(32'h3ba82744),
	.w2(32'h3b5c6961),
	.w3(32'h3bd98af2),
	.w4(32'h3bab7877),
	.w5(32'h3a9f0a00),
	.w6(32'h3ae42c4d),
	.w7(32'h395ce919),
	.w8(32'hbadbb2ad),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc749dcb),
	.w1(32'hbc11704d),
	.w2(32'hbc2edee4),
	.w3(32'hbc9736f3),
	.w4(32'hbc0f1238),
	.w5(32'hbc25cf4e),
	.w6(32'hbc5b0547),
	.w7(32'hbc463154),
	.w8(32'hbae09bf8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bbfd90),
	.w1(32'hba90f6b2),
	.w2(32'hbae61512),
	.w3(32'h3a95d03a),
	.w4(32'hb936d669),
	.w5(32'hba96acde),
	.w6(32'h3a8c40d8),
	.w7(32'h39a474ac),
	.w8(32'hbaa3660d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad074d1),
	.w1(32'hba9fb0f1),
	.w2(32'h3b2f9107),
	.w3(32'h3abe6abc),
	.w4(32'h397248c5),
	.w5(32'hb9862ae8),
	.w6(32'hbb504f00),
	.w7(32'hbb65c9c9),
	.w8(32'hbb905d52),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc30bc),
	.w1(32'h3908c31e),
	.w2(32'hbb050eca),
	.w3(32'h3a1a025a),
	.w4(32'hba0aea2c),
	.w5(32'hbb20c6f7),
	.w6(32'h3a9ca8cf),
	.w7(32'h38f94f16),
	.w8(32'hbb021174),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc36904),
	.w1(32'h3bb48ce9),
	.w2(32'h3b92c4d2),
	.w3(32'h3bc09a7f),
	.w4(32'h3be8cf19),
	.w5(32'h3b8801b2),
	.w6(32'h3b8e9982),
	.w7(32'h3bce9d9a),
	.w8(32'hb8bf17fa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3157c),
	.w1(32'h3a1123f2),
	.w2(32'hba7011c3),
	.w3(32'h3b820952),
	.w4(32'h3a3cdbe2),
	.w5(32'hbb1f082d),
	.w6(32'h3b0f2cb2),
	.w7(32'hba1b049b),
	.w8(32'hbb60daca),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d855b),
	.w1(32'hba3db2b0),
	.w2(32'hba6fdf45),
	.w3(32'h3a3a71ec),
	.w4(32'hba266a41),
	.w5(32'hba39ffd5),
	.w6(32'h39d8825b),
	.w7(32'hb9e15f24),
	.w8(32'hba3a8229),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11d08e),
	.w1(32'h3ab5a26d),
	.w2(32'hbac0c29c),
	.w3(32'h3baa0895),
	.w4(32'h3a60547b),
	.w5(32'hba2ccf37),
	.w6(32'h3b0c9401),
	.w7(32'hba849c9f),
	.w8(32'h398cd0d1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb675fea),
	.w1(32'hbb0303cf),
	.w2(32'hbb44d7a5),
	.w3(32'hbbc1b3af),
	.w4(32'hbc0c4b17),
	.w5(32'hbb785d93),
	.w6(32'hbc0f4fbc),
	.w7(32'hbc426d9c),
	.w8(32'hbc4195fe),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a372c32),
	.w1(32'h391634ee),
	.w2(32'h39e3a736),
	.w3(32'h38e15afc),
	.w4(32'hba54db62),
	.w5(32'hb89d6be7),
	.w6(32'hb9197b82),
	.w7(32'hb9e35323),
	.w8(32'hb8a62939),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a49e4),
	.w1(32'hbc61c031),
	.w2(32'hbc96c9e6),
	.w3(32'hbcac5c89),
	.w4(32'hbc676b85),
	.w5(32'hbc57a87c),
	.w6(32'hbc59e683),
	.w7(32'hbc44684e),
	.w8(32'hbc365311),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48febd),
	.w1(32'hbb850372),
	.w2(32'hbb4ba644),
	.w3(32'hbbce7c6a),
	.w4(32'hbb8a3476),
	.w5(32'hbb4ee707),
	.w6(32'hbbdd42b2),
	.w7(32'hbb9a3a9d),
	.w8(32'hbb74d777),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81822aa),
	.w1(32'hb9102989),
	.w2(32'hb82cf148),
	.w3(32'hb9360f88),
	.w4(32'hb8fd1280),
	.w5(32'hb82f25bb),
	.w6(32'hb9219180),
	.w7(32'hb918b20a),
	.w8(32'hb8effbdb),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93dc5fa),
	.w1(32'hb98fe09d),
	.w2(32'h34ec0b57),
	.w3(32'hb91aa07b),
	.w4(32'hb9445123),
	.w5(32'hb9200988),
	.w6(32'h38af16fb),
	.w7(32'hb8a4aeb9),
	.w8(32'h38ae8282),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b334e6b),
	.w1(32'h3b51df7e),
	.w2(32'h3acb6e5f),
	.w3(32'h3b8210ed),
	.w4(32'h3b5ee2db),
	.w5(32'h3b1ce90a),
	.w6(32'h3b74e7fd),
	.w7(32'h3b096710),
	.w8(32'h3b04ecd1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc570528),
	.w1(32'hbcc77b06),
	.w2(32'hbc69c0c5),
	.w3(32'hbc856d3f),
	.w4(32'hbc30d61e),
	.w5(32'hbc67e182),
	.w6(32'hbcb1623e),
	.w7(32'hbc051fed),
	.w8(32'hbc98a671),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac1f32),
	.w1(32'hb7702434),
	.w2(32'h3b86a664),
	.w3(32'h3b34601d),
	.w4(32'h3aa5832b),
	.w5(32'h3b0ba9ea),
	.w6(32'h3975169e),
	.w7(32'hbab537ed),
	.w8(32'hba59e64e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c673ae),
	.w1(32'h3b3b8eca),
	.w2(32'hba351106),
	.w3(32'h3c243f22),
	.w4(32'h3bfab4c4),
	.w5(32'h3b24e043),
	.w6(32'h3be1ac5e),
	.w7(32'hbadaef2e),
	.w8(32'h381ab951),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63318f),
	.w1(32'h3a8b437f),
	.w2(32'h3a6606c1),
	.w3(32'h3a466eee),
	.w4(32'h3a1c95a3),
	.w5(32'h399c3095),
	.w6(32'h394f42e2),
	.w7(32'h3a63b224),
	.w8(32'h3a2dd314),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3850a954),
	.w1(32'h3838e004),
	.w2(32'h38d065f7),
	.w3(32'h385fc2fa),
	.w4(32'h3535c200),
	.w5(32'h388a49ff),
	.w6(32'h39288ec9),
	.w7(32'hb82c4fff),
	.w8(32'h381bc38a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a957247),
	.w1(32'h3be36bac),
	.w2(32'h3b2cf6f9),
	.w3(32'h3bb83405),
	.w4(32'h3c2511dc),
	.w5(32'h3ad13773),
	.w6(32'h3ba5c0ed),
	.w7(32'hb97071a8),
	.w8(32'hbbb7e185),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b8c9c),
	.w1(32'h3a8579e8),
	.w2(32'h39d53722),
	.w3(32'h3aa5abe7),
	.w4(32'h3adf43e8),
	.w5(32'h3af5af6e),
	.w6(32'h3a18502e),
	.w7(32'h3a505f15),
	.w8(32'h3afe5eac),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a720bff),
	.w1(32'h3b8f2240),
	.w2(32'h39b93a9c),
	.w3(32'h3c222b5b),
	.w4(32'h3bd3cd01),
	.w5(32'h3af4b656),
	.w6(32'h3c17661a),
	.w7(32'h3ae73ddb),
	.w8(32'hb9e5c914),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a6b388),
	.w1(32'hb802bb92),
	.w2(32'hb84eaecc),
	.w3(32'hb91ab900),
	.w4(32'h35034fe9),
	.w5(32'hb804e270),
	.w6(32'h39190337),
	.w7(32'hb801d621),
	.w8(32'h35a3eb3f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb945be0c),
	.w1(32'hb7d21b5c),
	.w2(32'h3959a971),
	.w3(32'hb8fc70ad),
	.w4(32'h382f47c7),
	.w5(32'h39a49080),
	.w6(32'hb7575494),
	.w7(32'h39004464),
	.w8(32'h39cc9d68),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60f23f),
	.w1(32'h39f8ebb1),
	.w2(32'h3aae8cc6),
	.w3(32'h39d0cdc7),
	.w4(32'h3a6f5abe),
	.w5(32'h3a3af43a),
	.w6(32'hbadede4f),
	.w7(32'hba1806fc),
	.w8(32'hba5e1e7e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba941188),
	.w1(32'hb8b9110d),
	.w2(32'hbaa7dc54),
	.w3(32'h3aa1e324),
	.w4(32'hb9a68459),
	.w5(32'hba8a4c9f),
	.w6(32'h399e0de8),
	.w7(32'hbac99a0f),
	.w8(32'hbaac330a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb811815a),
	.w1(32'h3a4401f2),
	.w2(32'h3a24d846),
	.w3(32'hb7a461a1),
	.w4(32'h3a2523d9),
	.w5(32'h3a7059f0),
	.w6(32'hb81a3bc0),
	.w7(32'hba032745),
	.w8(32'hb99a4660),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1aa528),
	.w1(32'h3b05be3f),
	.w2(32'h3b0c6606),
	.w3(32'hb9b56d5c),
	.w4(32'hb93026f8),
	.w5(32'h3ace3ecf),
	.w6(32'hbb0ed7ac),
	.w7(32'h39b1b453),
	.w8(32'h39a35982),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9018b),
	.w1(32'hbc656e90),
	.w2(32'hb6cf499c),
	.w3(32'h3a6fe12f),
	.w4(32'hbc2f4759),
	.w5(32'h3bc27982),
	.w6(32'hbc0c8d92),
	.w7(32'hbb6728fe),
	.w8(32'h3a69d8e3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27c608),
	.w1(32'h3c650b2d),
	.w2(32'h3bb550bd),
	.w3(32'h3c8d1786),
	.w4(32'h3c2c2185),
	.w5(32'h3b8f1efe),
	.w6(32'h3c292c03),
	.w7(32'h3b1eb5c0),
	.w8(32'h3b998f90),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a8a8f),
	.w1(32'h3cab920f),
	.w2(32'h3c0817b3),
	.w3(32'h3ca89789),
	.w4(32'h3c7d8274),
	.w5(32'h3b8f6d3a),
	.w6(32'h3ccd9803),
	.w7(32'h3c1c157f),
	.w8(32'h3ba76c6c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab78496),
	.w1(32'h3a53e890),
	.w2(32'h390b744c),
	.w3(32'h3b52c38f),
	.w4(32'h389459b4),
	.w5(32'hb7f62459),
	.w6(32'h3b05619d),
	.w7(32'hba0f1104),
	.w8(32'hb846327d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0fda7),
	.w1(32'hb9ce28cd),
	.w2(32'hb96876fe),
	.w3(32'hb9c2f64d),
	.w4(32'hb9da9066),
	.w5(32'hb9a03e2d),
	.w6(32'hb96029b0),
	.w7(32'h38168a06),
	.w8(32'h393b72b1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83ccdc3),
	.w1(32'h38531500),
	.w2(32'h39307cc5),
	.w3(32'hb88bb73a),
	.w4(32'h38a2ded6),
	.w5(32'h38bd2e09),
	.w6(32'h39a07a7b),
	.w7(32'hb5efde49),
	.w8(32'h38b9e4b6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44642b),
	.w1(32'hb91f635c),
	.w2(32'h3a741a15),
	.w3(32'hba6557ae),
	.w4(32'h38be2195),
	.w5(32'h39fa1e40),
	.w6(32'hba2feae2),
	.w7(32'h3932c3bc),
	.w8(32'h39c447e5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd87294),
	.w1(32'h3ae1d857),
	.w2(32'h3b183837),
	.w3(32'hbc0cc466),
	.w4(32'h3a592b80),
	.w5(32'hbac7b57d),
	.w6(32'hbbc72c72),
	.w7(32'hbb286950),
	.w8(32'hbb4a04ef),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a2518),
	.w1(32'hb9d040f6),
	.w2(32'hb9ddab4e),
	.w3(32'h3b47980f),
	.w4(32'h3b103222),
	.w5(32'h3aa479e2),
	.w6(32'h3aeb702d),
	.w7(32'hba6058e5),
	.w8(32'h3a0e69ef),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb836eb4),
	.w1(32'hba41cab1),
	.w2(32'h3b9d615f),
	.w3(32'h3b60c43a),
	.w4(32'h3aa69ba4),
	.w5(32'h3b1cf07f),
	.w6(32'h39c1c3b4),
	.w7(32'hb9ba6703),
	.w8(32'h3b5e0009),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8021e2),
	.w1(32'hbb314975),
	.w2(32'hba4988c7),
	.w3(32'hbb1c55ce),
	.w4(32'hba8a4505),
	.w5(32'h3b6bc2a6),
	.w6(32'hbbdbc506),
	.w7(32'hbb027e44),
	.w8(32'h3a529a7a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9a6f1),
	.w1(32'hbc7ffe2e),
	.w2(32'hbc7293c9),
	.w3(32'hbc76a29b),
	.w4(32'hbc2176d0),
	.w5(32'hbbd4f950),
	.w6(32'hbc78771e),
	.w7(32'hbbd3c089),
	.w8(32'hbbb29ae5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e52dac),
	.w1(32'h39acdebf),
	.w2(32'h3934576d),
	.w3(32'h3843aee0),
	.w4(32'h3a3cb33c),
	.w5(32'h3a10610e),
	.w6(32'h3978d043),
	.w7(32'h3a2d46cb),
	.w8(32'h39d569b3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad93b85),
	.w1(32'hba81e20f),
	.w2(32'hbaec757d),
	.w3(32'hbadfbec8),
	.w4(32'hbb0ba06f),
	.w5(32'hbb140c99),
	.w6(32'hbaea6df4),
	.w7(32'hbb221d4d),
	.w8(32'hbb4c4e6f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a380950),
	.w1(32'h3a744385),
	.w2(32'h37b0c059),
	.w3(32'h3a93ac2d),
	.w4(32'h3a871ccb),
	.w5(32'hb90bb852),
	.w6(32'h3a6db027),
	.w7(32'h3a5fe533),
	.w8(32'h394fd4f0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb518870),
	.w1(32'hbaa2bc02),
	.w2(32'hbb4687d3),
	.w3(32'hba57e0e3),
	.w4(32'h3b010f64),
	.w5(32'hbb48f86c),
	.w6(32'hba8b437a),
	.w7(32'hba356bd7),
	.w8(32'hbb927786),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a6155),
	.w1(32'hbb3252c4),
	.w2(32'hbb6e7c46),
	.w3(32'hbb0d5ca5),
	.w4(32'hbb144acf),
	.w5(32'hbb456e27),
	.w6(32'hbad5f571),
	.w7(32'hba90973e),
	.w8(32'hbb0d7e73),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea37be),
	.w1(32'hbbf6259a),
	.w2(32'hbbd58658),
	.w3(32'hbc75c834),
	.w4(32'hbc233755),
	.w5(32'hbbc51d5b),
	.w6(32'hbc4c98c7),
	.w7(32'hbba9f94e),
	.w8(32'hbc0e0508),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cf1ef),
	.w1(32'hbad7559e),
	.w2(32'hbb4e0acb),
	.w3(32'hb9efccc0),
	.w4(32'h39b83b65),
	.w5(32'hbb1acb55),
	.w6(32'h3ad722b5),
	.w7(32'h3a8fef74),
	.w8(32'hb9e76208),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39625406),
	.w1(32'hb9396fec),
	.w2(32'hb9e24db4),
	.w3(32'h3938ac6a),
	.w4(32'hb9b57cf3),
	.w5(32'hb9fd0bf9),
	.w6(32'hb91ff2f6),
	.w7(32'hb948e326),
	.w8(32'hb9180911),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9879248),
	.w1(32'hb855e7ee),
	.w2(32'hb48574e4),
	.w3(32'hb99b5cf6),
	.w4(32'hb941b874),
	.w5(32'hb938b041),
	.w6(32'h378ebabd),
	.w7(32'hb8ce84af),
	.w8(32'h3811af3d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb793397a),
	.w1(32'h398f6f80),
	.w2(32'hb966b51d),
	.w3(32'h39ccd623),
	.w4(32'h3a16de50),
	.w5(32'h38fc78eb),
	.w6(32'h3a44d15b),
	.w7(32'h38637d59),
	.w8(32'h399a8c7b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f8cd5),
	.w1(32'h3a266971),
	.w2(32'h39d5a7be),
	.w3(32'h3aab48fc),
	.w4(32'h3a86da6a),
	.w5(32'h3a13abe7),
	.w6(32'h3ab04ab6),
	.w7(32'h3a8c7a93),
	.w8(32'h3a41439d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996741c),
	.w1(32'h39ece175),
	.w2(32'h3a049531),
	.w3(32'h3a04e8ba),
	.w4(32'h39aa4f11),
	.w5(32'h3981aa43),
	.w6(32'h3a9ec9de),
	.w7(32'h39b3937d),
	.w8(32'h3985eded),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb616678),
	.w1(32'hbb7e8526),
	.w2(32'hbb48956f),
	.w3(32'hbba3ae5a),
	.w4(32'hbb5dbde1),
	.w5(32'hbb676d32),
	.w6(32'hbb726044),
	.w7(32'hbb618711),
	.w8(32'hbbb38483),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc295532),
	.w1(32'hbb357d15),
	.w2(32'hbb42b763),
	.w3(32'hbc531d2c),
	.w4(32'h3a8ed2c7),
	.w5(32'hbc1a4b3a),
	.w6(32'hbb8cf5ce),
	.w7(32'hbb07be97),
	.w8(32'hbc13c1f6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992e07d),
	.w1(32'hb98b7e0b),
	.w2(32'hb9fe28dc),
	.w3(32'hb828b8da),
	.w4(32'hb93424bc),
	.w5(32'hb9a68cb4),
	.w6(32'hba088a55),
	.w7(32'hba115f7e),
	.w8(32'hba06c580),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30e4cf),
	.w1(32'h391677d4),
	.w2(32'h382f5447),
	.w3(32'hba1a1454),
	.w4(32'h3934e5c2),
	.w5(32'h38d61cb9),
	.w6(32'h38db37d2),
	.w7(32'h35c3f947),
	.w8(32'h397cef02),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da6dfc),
	.w1(32'h38074d14),
	.w2(32'h38a44add),
	.w3(32'h39b8160e),
	.w4(32'hb8b1b90c),
	.w5(32'hb88e827b),
	.w6(32'h38ee1c00),
	.w7(32'h389d3d0a),
	.w8(32'h3973cd3e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386d7838),
	.w1(32'h35b71194),
	.w2(32'h38b41ceb),
	.w3(32'h379a0d5b),
	.w4(32'hb8598232),
	.w5(32'h392fed8f),
	.w6(32'h382d2c43),
	.w7(32'hb7733906),
	.w8(32'h390780a5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed09ab),
	.w1(32'h3b31b7ba),
	.w2(32'h3bb9a398),
	.w3(32'hbb562ee1),
	.w4(32'h3a0a1113),
	.w5(32'h39610535),
	.w6(32'hbbfde595),
	.w7(32'hbb8cb7d8),
	.w8(32'hbc129234),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0bb42),
	.w1(32'hbb12832f),
	.w2(32'hbb150b56),
	.w3(32'h3b048bcb),
	.w4(32'hbb827704),
	.w5(32'hbbe5b0ba),
	.w6(32'hbaf11a76),
	.w7(32'hbad48775),
	.w8(32'hbb79329d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23ae2a),
	.w1(32'hbc026f5c),
	.w2(32'hbc23f42d),
	.w3(32'hbbd92883),
	.w4(32'hbac0fec3),
	.w5(32'hbc2dd8e8),
	.w6(32'hbaf608f7),
	.w7(32'hbaa5e650),
	.w8(32'hbc141a94),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9425138),
	.w1(32'h3bb09dbf),
	.w2(32'h3b82e2b9),
	.w3(32'h3c367f57),
	.w4(32'h3bf8f801),
	.w5(32'h3b1bfa33),
	.w6(32'h3b7d3aec),
	.w7(32'hbad56039),
	.w8(32'h3b3e2a86),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397ecf85),
	.w1(32'h387fc759),
	.w2(32'h394182da),
	.w3(32'h399fc094),
	.w4(32'h390ddae5),
	.w5(32'h39391d22),
	.w6(32'h378a7209),
	.w7(32'h377a0cca),
	.w8(32'h390fbd93),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bc100d),
	.w1(32'hb8e1838a),
	.w2(32'hb88f815d),
	.w3(32'h386925c2),
	.w4(32'hb89a7294),
	.w5(32'hb88a4284),
	.w6(32'h38ae151a),
	.w7(32'hb84d4d88),
	.w8(32'h38862c7d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb897a1fb),
	.w1(32'hb7dd91cc),
	.w2(32'h38bef280),
	.w3(32'hb88dce7b),
	.w4(32'hb7648ad2),
	.w5(32'hb86f6197),
	.w6(32'h3937321b),
	.w7(32'hb66464c6),
	.w8(32'h38ecca28),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb916a39e),
	.w1(32'hbacdc7b2),
	.w2(32'hbae3fe0b),
	.w3(32'hba4e9db4),
	.w4(32'hbaa3a6b7),
	.w5(32'hbad488ee),
	.w6(32'hbac5ba6e),
	.w7(32'hbb17af17),
	.w8(32'hbb0bf1a3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380cc240),
	.w1(32'h38c768c1),
	.w2(32'h38f404c0),
	.w3(32'h390e5850),
	.w4(32'h386a2665),
	.w5(32'hb769b19b),
	.w6(32'h3967dc2f),
	.w7(32'h398ea37b),
	.w8(32'h39a2a249),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2876cb),
	.w1(32'hbc0d4838),
	.w2(32'hbb2c991d),
	.w3(32'hbc0cf017),
	.w4(32'hbc0aecbc),
	.w5(32'hba4b7d60),
	.w6(32'hbc21156d),
	.w7(32'hbb23d027),
	.w8(32'hbadf0335),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31cb48),
	.w1(32'hbc14057b),
	.w2(32'hbc069462),
	.w3(32'hbc2c0a8b),
	.w4(32'hbc948b1e),
	.w5(32'hbb8aa963),
	.w6(32'hbcade70c),
	.w7(32'hbc583b1d),
	.w8(32'hbc03456a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f3b8f),
	.w1(32'h3b6d3f49),
	.w2(32'hba3099c8),
	.w3(32'h3bb6476e),
	.w4(32'h3b50ec86),
	.w5(32'hb9bfbcab),
	.w6(32'h3b969504),
	.w7(32'h3a4c73ac),
	.w8(32'h3a62f062),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b60a3),
	.w1(32'hbb011ceb),
	.w2(32'hbb2f2cc6),
	.w3(32'hbb3c908b),
	.w4(32'hbaadef53),
	.w5(32'hbb3529f1),
	.w6(32'hbb12512f),
	.w7(32'hbad6c79a),
	.w8(32'hbb5ec4ee),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f8956),
	.w1(32'hbb5aab07),
	.w2(32'h3b1a7a01),
	.w3(32'hb7295f72),
	.w4(32'h39dfc0e8),
	.w5(32'h3b70fd5a),
	.w6(32'hbb45c745),
	.w7(32'hbafcc619),
	.w8(32'hbb1e7a25),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04baab),
	.w1(32'hba469b67),
	.w2(32'hbb36a3ca),
	.w3(32'h39f9619a),
	.w4(32'h3aae319b),
	.w5(32'hbb0ad185),
	.w6(32'hbafe44e6),
	.w7(32'hbb2fb370),
	.w8(32'hbb73cd55),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a97f4),
	.w1(32'hbbd1443d),
	.w2(32'hbb9912b5),
	.w3(32'hbbb6597f),
	.w4(32'hbb44638a),
	.w5(32'hba9c1970),
	.w6(32'hbb98e7e3),
	.w7(32'hbb2a71d4),
	.w8(32'hba85640f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374f6fd6),
	.w1(32'hb9801ca5),
	.w2(32'hb97cfdbd),
	.w3(32'hb89203da),
	.w4(32'hb93884cd),
	.w5(32'hb99806d3),
	.w6(32'hb9329437),
	.w7(32'hb944a311),
	.w8(32'hb8170c8d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d19e9),
	.w1(32'h38b6ba83),
	.w2(32'h3902fa33),
	.w3(32'hb966baec),
	.w4(32'hb85ca415),
	.w5(32'hb9216731),
	.w6(32'h38e1133c),
	.w7(32'h39338897),
	.w8(32'h39229e98),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f315d0),
	.w1(32'h38be7802),
	.w2(32'h3a15992e),
	.w3(32'h3a3cc36c),
	.w4(32'h3a21fbdf),
	.w5(32'h399a0346),
	.w6(32'h3a3f8a25),
	.w7(32'h399ff1b9),
	.w8(32'h399f1ed0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb99c4),
	.w1(32'h38a17b10),
	.w2(32'hb8c5c701),
	.w3(32'h3a176034),
	.w4(32'h392725d7),
	.w5(32'h394f948b),
	.w6(32'h3a216ea6),
	.w7(32'h38f22b7a),
	.w8(32'h39d2744b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb816fb49),
	.w1(32'h3b18c7f5),
	.w2(32'h3b5f7b66),
	.w3(32'h3bb4541c),
	.w4(32'h3add4963),
	.w5(32'h3b31ee06),
	.w6(32'h3b0b9036),
	.w7(32'hbb082e0a),
	.w8(32'h3aa4ced5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3785e342),
	.w1(32'hb92adb74),
	.w2(32'hba13f495),
	.w3(32'hb7ca24c5),
	.w4(32'h3886cf68),
	.w5(32'h3857bed2),
	.w6(32'hb9afd000),
	.w7(32'hb991be1a),
	.w8(32'h38d70142),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b9a09),
	.w1(32'hbb54c503),
	.w2(32'hbad2f87c),
	.w3(32'h38dd5756),
	.w4(32'hbabca988),
	.w5(32'h373ffdae),
	.w6(32'hbb20c056),
	.w7(32'hbb0ce243),
	.w8(32'h3a2e237d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27aaf3),
	.w1(32'hbc350392),
	.w2(32'hbbd1ab38),
	.w3(32'hbca8e858),
	.w4(32'hbc66abfc),
	.w5(32'hbb872470),
	.w6(32'hbcab9dfa),
	.w7(32'hbc1bfde3),
	.w8(32'hbbb38459),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1ad1e),
	.w1(32'h3b94f24b),
	.w2(32'hbac83b33),
	.w3(32'h3bdeafea),
	.w4(32'h3b98a6d4),
	.w5(32'h3b5d1dfb),
	.w6(32'h3bb6bd19),
	.w7(32'h3b26a275),
	.w8(32'h3b14d79c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0deffc),
	.w1(32'h3ab9b5fd),
	.w2(32'h3bc29e89),
	.w3(32'h3b7a39a4),
	.w4(32'h3ba67697),
	.w5(32'h3bdb2670),
	.w6(32'h3b32c825),
	.w7(32'h3c1ca177),
	.w8(32'h3a8738f5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11155a),
	.w1(32'h3bb4c4b2),
	.w2(32'h3b89a259),
	.w3(32'h3bb4cce9),
	.w4(32'h3bc06eab),
	.w5(32'h3b39b2fd),
	.w6(32'h3ba4b4e5),
	.w7(32'h3b911571),
	.w8(32'h3b727519),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9287f8),
	.w1(32'hbbb2a7fd),
	.w2(32'hbb87edd1),
	.w3(32'hbbe72dc8),
	.w4(32'hbbd5c20a),
	.w5(32'hbba129f2),
	.w6(32'hbbfae961),
	.w7(32'hbc0e5c57),
	.w8(32'hbc2faca3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8abd255),
	.w1(32'h3b35aac9),
	.w2(32'h3b8ff4d1),
	.w3(32'h3af6fc7e),
	.w4(32'h3af547ed),
	.w5(32'h3abad3a3),
	.w6(32'hba346ecb),
	.w7(32'hba2b0d83),
	.w8(32'hbb81a724),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac687f5),
	.w1(32'h3b392e2e),
	.w2(32'hbadf4862),
	.w3(32'h3bd6847b),
	.w4(32'h3b3b74a5),
	.w5(32'h3ac74b62),
	.w6(32'h3bb1042d),
	.w7(32'h39f2ca9a),
	.w8(32'h3a1f2a4d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af032ac),
	.w1(32'h3b02daff),
	.w2(32'h397f8ff7),
	.w3(32'h3b118164),
	.w4(32'h3ae34f77),
	.w5(32'h37c57f45),
	.w6(32'h3ac34643),
	.w7(32'h3a579684),
	.w8(32'hb9d1e832),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacabaa6),
	.w1(32'hb9ffb9de),
	.w2(32'hbae2239f),
	.w3(32'hbb49f906),
	.w4(32'hb9ec1356),
	.w5(32'hbb51a503),
	.w6(32'hbbaaeae5),
	.w7(32'hbb978d03),
	.w8(32'hbbc315f0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba551d6f),
	.w1(32'h3a2759a7),
	.w2(32'h3bbd4408),
	.w3(32'h3a758a8e),
	.w4(32'h3bc45dd6),
	.w5(32'h3b94f2a2),
	.w6(32'h3b53d38b),
	.w7(32'h3afc09f0),
	.w8(32'hbb1b1349),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12fbae),
	.w1(32'hbc92e295),
	.w2(32'hbbd30ca5),
	.w3(32'hbc88361d),
	.w4(32'hbc98df3e),
	.w5(32'h3b294354),
	.w6(32'hbcc16c8e),
	.w7(32'hbc0a98b0),
	.w8(32'h3b00dde7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5121c),
	.w1(32'h3c2e0570),
	.w2(32'hbb2a919f),
	.w3(32'h3ca4a382),
	.w4(32'h3c8baba8),
	.w5(32'h3b845b45),
	.w6(32'h3c87d457),
	.w7(32'h3c5344b6),
	.w8(32'h3ac39876),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb101035),
	.w1(32'h3b2cc23d),
	.w2(32'h3af2180d),
	.w3(32'h3be5b653),
	.w4(32'h3b83947c),
	.w5(32'h3b0cb00b),
	.w6(32'h3b17fd25),
	.w7(32'hbab3f560),
	.w8(32'h39f364c6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba131f03),
	.w1(32'hbbc55c75),
	.w2(32'h3aabf1e4),
	.w3(32'h3b3c5c29),
	.w4(32'h3b1709c6),
	.w5(32'h3b45015e),
	.w6(32'hbb2f851f),
	.w7(32'h3be2c32b),
	.w8(32'hba7a3981),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa41a38),
	.w1(32'h3aaeabf7),
	.w2(32'h3ad486f7),
	.w3(32'h3aeb0dc8),
	.w4(32'h3b29786a),
	.w5(32'h3b15b9c1),
	.w6(32'h3aaaca0a),
	.w7(32'h3b15d09e),
	.w8(32'h3af84114),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc190555),
	.w1(32'hbce0446a),
	.w2(32'hbcc75c64),
	.w3(32'hbc818da2),
	.w4(32'hbca69430),
	.w5(32'hbc0a6951),
	.w6(32'hbcba3f99),
	.w7(32'hbc5558b0),
	.w8(32'hbba19023),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba66304),
	.w1(32'h3a803f10),
	.w2(32'h3a9a3ff6),
	.w3(32'h3bce5d1d),
	.w4(32'h3b49913e),
	.w5(32'h38fcd8b6),
	.w6(32'h3b807d60),
	.w7(32'h3b2d84d0),
	.w8(32'h3ab6a7b7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de8c33),
	.w1(32'h398ef1d1),
	.w2(32'hb7c741de),
	.w3(32'h3a1039a3),
	.w4(32'h39e97762),
	.w5(32'hb842d655),
	.w6(32'h3a7c2232),
	.w7(32'h39e63cbf),
	.w8(32'h39989676),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4d577),
	.w1(32'hb783b778),
	.w2(32'hba36c303),
	.w3(32'hbad4d413),
	.w4(32'h3941d8e4),
	.w5(32'hbad49e64),
	.w6(32'hbb08fe75),
	.w7(32'hbb2c337e),
	.w8(32'hbab3f92c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d0675),
	.w1(32'h3b481f2c),
	.w2(32'h3b46fb28),
	.w3(32'h3afde2f7),
	.w4(32'h3b2b86c7),
	.w5(32'h3a7830cc),
	.w6(32'hba2d216a),
	.w7(32'hb9309508),
	.w8(32'hb8f1df0e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7d72a),
	.w1(32'h3b451cd2),
	.w2(32'h3af83eec),
	.w3(32'h3bcc18de),
	.w4(32'h3b8d9492),
	.w5(32'h3ae8e59e),
	.w6(32'h3b5a7839),
	.w7(32'h3a0507f4),
	.w8(32'h3b126cfe),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba994cb2),
	.w1(32'h3b95c10c),
	.w2(32'hbb6497d7),
	.w3(32'h3b83149d),
	.w4(32'h3b39e18f),
	.w5(32'hbaab4c16),
	.w6(32'h3b6c3137),
	.w7(32'h39ca13aa),
	.w8(32'hbaade8b6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba362f4a),
	.w1(32'hb929012f),
	.w2(32'hbb4a013c),
	.w3(32'h3ac2d776),
	.w4(32'h39806daa),
	.w5(32'hbb214a68),
	.w6(32'h38c48623),
	.w7(32'hbb1b7221),
	.w8(32'hbb7e9fc8),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8736a0),
	.w1(32'hb7aa2bfe),
	.w2(32'h3b8755cc),
	.w3(32'hbbd4cf8a),
	.w4(32'hbb51fc47),
	.w5(32'h3b7e1fc7),
	.w6(32'hbb042cf7),
	.w7(32'h3b33c02f),
	.w8(32'h3bc46c3b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ce0e1),
	.w1(32'hbbb6c161),
	.w2(32'hbb75c7a0),
	.w3(32'hbbc51e42),
	.w4(32'hbbda4d97),
	.w5(32'hbba104f1),
	.w6(32'hbbb6bc34),
	.w7(32'hbbfd169a),
	.w8(32'hbbef94d9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab40157),
	.w1(32'h39323331),
	.w2(32'h3a12ad3a),
	.w3(32'h3ae4f356),
	.w4(32'h3aba3228),
	.w5(32'h39c49e11),
	.w6(32'h3b3ae476),
	.w7(32'h3a264136),
	.w8(32'h386ec10e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9981c62),
	.w1(32'hb8d25db1),
	.w2(32'hb88dc62f),
	.w3(32'hb952e1ce),
	.w4(32'hb86798e9),
	.w5(32'hb84a6cb3),
	.w6(32'hb8e88e55),
	.w7(32'hb91f7f48),
	.w8(32'h386d4244),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a60b6f),
	.w1(32'hb9b727bb),
	.w2(32'hba03431f),
	.w3(32'h399e1739),
	.w4(32'hba630706),
	.w5(32'hba2629a9),
	.w6(32'h385a0716),
	.w7(32'hb9fa0b5a),
	.w8(32'hba4356b1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb705ef00),
	.w1(32'hb839f34b),
	.w2(32'hb876c796),
	.w3(32'hb7236755),
	.w4(32'hb7c439de),
	.w5(32'hb8c67ad8),
	.w6(32'h38ad7741),
	.w7(32'h362a262c),
	.w8(32'hb7b4f21c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398371cc),
	.w1(32'h3a29c707),
	.w2(32'h3abfca4d),
	.w3(32'h39f09bfb),
	.w4(32'h3a8de717),
	.w5(32'h3ad11d36),
	.w6(32'h3a2c1485),
	.w7(32'h39c104b6),
	.w8(32'hba14ac4b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cf190),
	.w1(32'h3b005066),
	.w2(32'h3b37d086),
	.w3(32'h3b9998e2),
	.w4(32'h3b4ac2ce),
	.w5(32'h3b2b117e),
	.w6(32'h3b1d35ae),
	.w7(32'hb9bafe66),
	.w8(32'h3aae3553),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa33cca),
	.w1(32'h39d9a9ae),
	.w2(32'hba1acf67),
	.w3(32'h3b027ac0),
	.w4(32'h3aedbf3a),
	.w5(32'h3932ad32),
	.w6(32'h3b271903),
	.w7(32'h3b102c79),
	.w8(32'h3a4a93d9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20ed98),
	.w1(32'hbb8290de),
	.w2(32'hbb0e86f2),
	.w3(32'hbb30eba2),
	.w4(32'hbb0d5fa3),
	.w5(32'hb89b4ab1),
	.w6(32'hbbad01bd),
	.w7(32'hbae68b15),
	.w8(32'hbadfd6b3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05d4da),
	.w1(32'h3bfecf47),
	.w2(32'h3afbd8bd),
	.w3(32'h3c0709a5),
	.w4(32'h3b90e84f),
	.w5(32'hb8ba2600),
	.w6(32'h3bf96530),
	.w7(32'h38ae5554),
	.w8(32'hbb18f21d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc4e25),
	.w1(32'h3a0758e3),
	.w2(32'h39d296ad),
	.w3(32'h39804386),
	.w4(32'h383520ff),
	.w5(32'h390da2cc),
	.w6(32'h39ab1f2c),
	.w7(32'h39532e84),
	.w8(32'h388f091e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae52c6),
	.w1(32'h37a2d8d9),
	.w2(32'hba511924),
	.w3(32'h3a10c3b4),
	.w4(32'h39c6c35e),
	.w5(32'hb9cbe0b0),
	.w6(32'h3a14f25f),
	.w7(32'h390a037b),
	.w8(32'hb97b1182),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e2f6d),
	.w1(32'hb90ae3c6),
	.w2(32'hb9303d33),
	.w3(32'hb9627108),
	.w4(32'hb88fa65e),
	.w5(32'hb89001b6),
	.w6(32'h38b1e3e7),
	.w7(32'hb9250a96),
	.w8(32'hb895767d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd036d),
	.w1(32'hbb41b754),
	.w2(32'hbb8a8a58),
	.w3(32'h3ae692b6),
	.w4(32'hba82d3df),
	.w5(32'hbc061782),
	.w6(32'hba8155aa),
	.w7(32'hbc1ad27d),
	.w8(32'h3892873e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23a9c7),
	.w1(32'h3c3fc648),
	.w2(32'h3c448cf6),
	.w3(32'hba978f3f),
	.w4(32'h3be57af3),
	.w5(32'h39c770ff),
	.w6(32'h3ad046ea),
	.w7(32'h3ac42595),
	.w8(32'hbc090448),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b7277),
	.w1(32'h3c64d39d),
	.w2(32'hbd1a31d6),
	.w3(32'hbc1556c3),
	.w4(32'h3c42c869),
	.w5(32'hbb6bc5cf),
	.w6(32'hbc81ce96),
	.w7(32'hbcb23582),
	.w8(32'hbc8386e8),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca7f096),
	.w1(32'h3bcb3b68),
	.w2(32'h3a6c50fb),
	.w3(32'hbca320e2),
	.w4(32'hbab69cc8),
	.w5(32'h3a027bcd),
	.w6(32'hba1eb5bb),
	.w7(32'hbb18a21a),
	.w8(32'hbc1d9c37),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ef571),
	.w1(32'hbbdabce0),
	.w2(32'hbb6519db),
	.w3(32'hbb543f72),
	.w4(32'hbbf2b349),
	.w5(32'hbaea92cc),
	.w6(32'hb99195b7),
	.w7(32'hbae488f1),
	.w8(32'h3a68bb22),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4b757),
	.w1(32'h3d2c4c82),
	.w2(32'h3b903754),
	.w3(32'h3c015e62),
	.w4(32'h3bc911de),
	.w5(32'hbb76b707),
	.w6(32'h3cec0fae),
	.w7(32'h3c8c2a61),
	.w8(32'hbb052788),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd6cd30),
	.w1(32'hbb2782c0),
	.w2(32'h3d35fd31),
	.w3(32'hb8db8e38),
	.w4(32'hba81c53c),
	.w5(32'hbc6a364c),
	.w6(32'hb9711c3c),
	.w7(32'hbc241c34),
	.w8(32'hbc4c9ff7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc976faa),
	.w1(32'h3cd2476e),
	.w2(32'h3c529f2d),
	.w3(32'hbc7f31e7),
	.w4(32'h3c4dd502),
	.w5(32'hba55c179),
	.w6(32'h3c56fd26),
	.w7(32'hbbdc4e7a),
	.w8(32'hbcc0b676),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1e5b47),
	.w1(32'hbc12313f),
	.w2(32'h3b038591),
	.w3(32'hbd02d62f),
	.w4(32'hbbf4c469),
	.w5(32'hbb890ad0),
	.w6(32'hbc678fd1),
	.w7(32'hbc410ad0),
	.w8(32'hbc578cc3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5f289),
	.w1(32'hbbef6e11),
	.w2(32'h3b93a5b4),
	.w3(32'h3bbcac61),
	.w4(32'hbaa5753b),
	.w5(32'hba9546bf),
	.w6(32'h3a74543d),
	.w7(32'hb866fc2f),
	.w8(32'h3b73abeb),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4a701),
	.w1(32'h3b265af0),
	.w2(32'hbb953074),
	.w3(32'hba75e948),
	.w4(32'h3b18e58b),
	.w5(32'h38a84885),
	.w6(32'hbba1469a),
	.w7(32'hbbb73e68),
	.w8(32'hbc1c94d3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a623f),
	.w1(32'h3be1d30c),
	.w2(32'hbc379e75),
	.w3(32'hbbf63ce1),
	.w4(32'hbb9f8b14),
	.w5(32'hbbb95e71),
	.w6(32'hba670ffc),
	.w7(32'hbc0d41e8),
	.w8(32'hbc437c0a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58527b),
	.w1(32'h3ca65fe4),
	.w2(32'h3bd17f1a),
	.w3(32'hbbb385e1),
	.w4(32'h3b83c57e),
	.w5(32'hba291841),
	.w6(32'h3ba25f10),
	.w7(32'h3c339b50),
	.w8(32'h3bb28ab3),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27f704),
	.w1(32'hbc5f8196),
	.w2(32'hbc3ee437),
	.w3(32'hbbb9efee),
	.w4(32'hbc8be0a1),
	.w5(32'hbc6e5107),
	.w6(32'hbc092f93),
	.w7(32'hbbb798e9),
	.w8(32'hbc5c7e09),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f6f74),
	.w1(32'hbb963bec),
	.w2(32'h3a28dcae),
	.w3(32'hbbf42dc3),
	.w4(32'hbb96cad3),
	.w5(32'hbb216b8f),
	.w6(32'hbb68d1ab),
	.w7(32'h3aa75b9b),
	.w8(32'h3bc83d96),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9576f),
	.w1(32'hbd3cf0ff),
	.w2(32'hbba1c5cd),
	.w3(32'h3c813866),
	.w4(32'hbccca955),
	.w5(32'hbc0e2584),
	.w6(32'hbc9096b0),
	.w7(32'h39a921a0),
	.w8(32'h3ca84e31),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4c97a8),
	.w1(32'hbbc992f3),
	.w2(32'h3c2bed95),
	.w3(32'h3c83d404),
	.w4(32'hbbe25236),
	.w5(32'hbc431731),
	.w6(32'h3b14b47c),
	.w7(32'h3c7ee522),
	.w8(32'hbbe8933e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd6f22b),
	.w1(32'h3c02f1e6),
	.w2(32'hba0fd0e8),
	.w3(32'hbc28c0de),
	.w4(32'h3b2f86a9),
	.w5(32'h3a94aa53),
	.w6(32'h3b451e21),
	.w7(32'hba025e44),
	.w8(32'hbbe1ee63),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf314df),
	.w1(32'h3bde2d35),
	.w2(32'h39ff7c09),
	.w3(32'hbbabcf01),
	.w4(32'h3bfbeffb),
	.w5(32'h3b1e4ee2),
	.w6(32'h3bb96259),
	.w7(32'h3aa2da42),
	.w8(32'hbbc7886f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc080b17),
	.w1(32'h3c03fa0a),
	.w2(32'h3b4bf7ff),
	.w3(32'hbb1edf6b),
	.w4(32'h3b594a70),
	.w5(32'h3b87db90),
	.w6(32'h3b6dfd03),
	.w7(32'hba29cd3f),
	.w8(32'h3b90032f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99b6c0),
	.w1(32'hb8112ab6),
	.w2(32'hbc133926),
	.w3(32'h3c8a9af9),
	.w4(32'hbb9e2130),
	.w5(32'hbb9107a9),
	.w6(32'hba7cb7ba),
	.w7(32'hbc26ad8e),
	.w8(32'hbbb3bacb),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba869581),
	.w1(32'h3b90215a),
	.w2(32'hbb858554),
	.w3(32'h3b42d882),
	.w4(32'h3b55c5eb),
	.w5(32'hbb365983),
	.w6(32'h3a961f7a),
	.w7(32'hbb862bd6),
	.w8(32'hbb84a220),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ef6a0),
	.w1(32'hbbc743ca),
	.w2(32'hbb94f081),
	.w3(32'hbb865ff2),
	.w4(32'hbb46df6d),
	.w5(32'hbb56023e),
	.w6(32'hbae1f2ba),
	.w7(32'hbbc91fb5),
	.w8(32'h3ac82520),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74b400),
	.w1(32'hbce7b044),
	.w2(32'h3bb11d5d),
	.w3(32'h3baa85d8),
	.w4(32'hbc869963),
	.w5(32'h3c1ef4b4),
	.w6(32'hbc2c6e93),
	.w7(32'h3b415479),
	.w8(32'h3bdcb3a1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdd20dd),
	.w1(32'h3ba88f3e),
	.w2(32'hba6577e1),
	.w3(32'h3ba89bad),
	.w4(32'h3b30bd97),
	.w5(32'hbbfa3fb3),
	.w6(32'h3b2dead3),
	.w7(32'hbc01ff08),
	.w8(32'hbb070810),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5efc9),
	.w1(32'hbc2127f6),
	.w2(32'hbbd56218),
	.w3(32'hbc134f87),
	.w4(32'hbb488d3c),
	.w5(32'hbb48c91d),
	.w6(32'hbc0004bb),
	.w7(32'hbb2deda0),
	.w8(32'hbbbd420c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb875524),
	.w1(32'h3c83717b),
	.w2(32'hbbb4ffab),
	.w3(32'h3b486c8a),
	.w4(32'h3b6ecdc8),
	.w5(32'hba4e3b4f),
	.w6(32'h3c735efb),
	.w7(32'h3b42f756),
	.w8(32'hbc571af5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc849f58),
	.w1(32'h3bcf3d17),
	.w2(32'hbb13d23e),
	.w3(32'hbb924d96),
	.w4(32'h3c45b6ff),
	.w5(32'h3b89ba1b),
	.w6(32'hba1f71a4),
	.w7(32'hbb5f8bce),
	.w8(32'h3b67bb4d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b6d805),
	.w1(32'h3b025f1b),
	.w2(32'hb9a0a1f3),
	.w3(32'h3b16c7cb),
	.w4(32'h3be2d82c),
	.w5(32'h3b77bbe0),
	.w6(32'h3ae9c5a6),
	.w7(32'h3b251e7d),
	.w8(32'h3b8c05f0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba1cbd),
	.w1(32'h3c892856),
	.w2(32'hbb5283f2),
	.w3(32'h3ba8f709),
	.w4(32'h3ba09db0),
	.w5(32'h3b6a7842),
	.w6(32'h3ba82262),
	.w7(32'hba8b9108),
	.w8(32'hbc16e51e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc944c8d),
	.w1(32'h3c8448d8),
	.w2(32'hbc74e22f),
	.w3(32'hbc072aed),
	.w4(32'h3c5f9d49),
	.w5(32'hbc6d96ff),
	.w6(32'h3ca694cb),
	.w7(32'hbc8792ae),
	.w8(32'hbbd1be5e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd28fdf),
	.w1(32'h3ba0fec6),
	.w2(32'h3bfe0d10),
	.w3(32'hbb444fb2),
	.w4(32'h3bb2e2f3),
	.w5(32'h3c08da4c),
	.w6(32'h3bc81e94),
	.w7(32'h3bc02b59),
	.w8(32'h3b64128a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39865a3d),
	.w1(32'hbb95b337),
	.w2(32'h3a91c298),
	.w3(32'hbb84d9a8),
	.w4(32'hb988b794),
	.w5(32'h3a35e48a),
	.w6(32'hbb092a16),
	.w7(32'hbabc8db9),
	.w8(32'h3b400da1),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8718bc),
	.w1(32'h3a2173c5),
	.w2(32'h3a4dadb2),
	.w3(32'h3b74272b),
	.w4(32'h3af2d65e),
	.w5(32'h3b4e0305),
	.w6(32'h3a563500),
	.w7(32'h3b4cec17),
	.w8(32'h3ba83a6f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a7ee1),
	.w1(32'hbb34c4f9),
	.w2(32'hbc8a4257),
	.w3(32'h39bab2e5),
	.w4(32'hbc0c0bd9),
	.w5(32'hbc1ccb86),
	.w6(32'hbc80a8b5),
	.w7(32'hbc99823e),
	.w8(32'hbcad31df),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8152f),
	.w1(32'h3be57554),
	.w2(32'hbc8fedb8),
	.w3(32'hbc3ad449),
	.w4(32'h3c029534),
	.w5(32'h3b5939f4),
	.w6(32'hba31c49c),
	.w7(32'h3bbd0b0a),
	.w8(32'h3ad47d1d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2caba0),
	.w1(32'h3ca0ae2d),
	.w2(32'hbbcfcc2f),
	.w3(32'hbb8a068c),
	.w4(32'h3bbf88d1),
	.w5(32'hbad7dec4),
	.w6(32'h3bdc312d),
	.w7(32'hbb904f18),
	.w8(32'hbc4ebec3),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce69d8),
	.w1(32'h3b541e1b),
	.w2(32'h3ad830d1),
	.w3(32'hbc1a480c),
	.w4(32'h3aa573b2),
	.w5(32'h3a228cbd),
	.w6(32'h3bd4c491),
	.w7(32'h3ac9536a),
	.w8(32'h3ac30ad0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd2409),
	.w1(32'h3ce08365),
	.w2(32'h3c9b77f6),
	.w3(32'h3bbcaa5b),
	.w4(32'h3c2c0948),
	.w5(32'h395edd3a),
	.w6(32'h3c934497),
	.w7(32'h3b94ea6c),
	.w8(32'hbbcc9c2c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc554003),
	.w1(32'hbb77a4c2),
	.w2(32'hbb5d40e0),
	.w3(32'hb8e9210e),
	.w4(32'hbb7eee83),
	.w5(32'hbaf5e52d),
	.w6(32'hbb8aa0ce),
	.w7(32'hbbafc55f),
	.w8(32'hbb3f3335),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb868acf),
	.w1(32'h3b0e3a2a),
	.w2(32'hbb5420eb),
	.w3(32'h39cbe628),
	.w4(32'h3b783174),
	.w5(32'hb9c2e7b1),
	.w6(32'h3b285d88),
	.w7(32'hba897a5d),
	.w8(32'hbb9534b2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9f2ea),
	.w1(32'hba66e256),
	.w2(32'hb98f7336),
	.w3(32'h3ad72153),
	.w4(32'h3a487a3b),
	.w5(32'hbb06be00),
	.w6(32'h3ad86f3d),
	.w7(32'h3a3fd04d),
	.w8(32'hbb1e96bc),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecd423),
	.w1(32'hbc84da01),
	.w2(32'h3b6ce941),
	.w3(32'hbbfa77fd),
	.w4(32'hbc6345f7),
	.w5(32'h3bb84150),
	.w6(32'hbc9b630a),
	.w7(32'hbaec2376),
	.w8(32'hba9d82a7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68c039),
	.w1(32'h3af5b00f),
	.w2(32'h3b4fcff8),
	.w3(32'h39925027),
	.w4(32'hbb08587a),
	.w5(32'h3b902296),
	.w6(32'h3b772942),
	.w7(32'h3bbe9578),
	.w8(32'hbb7dae49),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdffcc4),
	.w1(32'hbbb52339),
	.w2(32'hbc56e269),
	.w3(32'h3b33da9d),
	.w4(32'h39aa4a74),
	.w5(32'hbbb4a7b6),
	.w6(32'h3ae412b6),
	.w7(32'hbab9fbcc),
	.w8(32'h3ad2a5b3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b600fb3),
	.w1(32'h3c854887),
	.w2(32'h3be27c3c),
	.w3(32'h3b9d4d74),
	.w4(32'h3bd2220a),
	.w5(32'h3b40c160),
	.w6(32'h3c872e04),
	.w7(32'h3bf7c4ad),
	.w8(32'hb9a51e39),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7dc0c),
	.w1(32'hbd13d450),
	.w2(32'hbc957621),
	.w3(32'hbacd5ce1),
	.w4(32'hbca46d6f),
	.w5(32'hbc6b0c18),
	.w6(32'hbcbc60fe),
	.w7(32'hbb897bb4),
	.w8(32'h3c604dfa),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d261df1),
	.w1(32'hbcad6987),
	.w2(32'h3c13a077),
	.w3(32'h3b8124e8),
	.w4(32'hbc76aa35),
	.w5(32'hbba89aa2),
	.w6(32'hbc12c55b),
	.w7(32'hbc24d788),
	.w8(32'h3b49b0e9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbd0e3),
	.w1(32'hbbaa54f3),
	.w2(32'h3ae88a17),
	.w3(32'hbbad53ca),
	.w4(32'hbc5977e2),
	.w5(32'hbbc84514),
	.w6(32'hbbb20480),
	.w7(32'hb9b425ac),
	.w8(32'hbcb02bdc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6979bb),
	.w1(32'h3b3dc0da),
	.w2(32'h3b684e47),
	.w3(32'hbb6ff9bd),
	.w4(32'h3bbd26ce),
	.w5(32'h3bef70ba),
	.w6(32'h3c2c0f71),
	.w7(32'h3bccb53e),
	.w8(32'h3b921518),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9842e),
	.w1(32'h3a3da1f7),
	.w2(32'hbbebe171),
	.w3(32'hbad5916f),
	.w4(32'h3ad039f0),
	.w5(32'hbaec2cf9),
	.w6(32'hbb857fed),
	.w7(32'hbbc2865d),
	.w8(32'hbbba9273),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cfe78f),
	.w1(32'hbc5aca76),
	.w2(32'h3c232d49),
	.w3(32'h380d8a74),
	.w4(32'hbb81bb43),
	.w5(32'h3b80ef0c),
	.w6(32'hbbd34583),
	.w7(32'h3bac0968),
	.w8(32'h3c432ae1),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca821f3),
	.w1(32'hbcf5b1b7),
	.w2(32'h3c4e5686),
	.w3(32'h3c2941e8),
	.w4(32'hbc8ff0ef),
	.w5(32'hbaa87968),
	.w6(32'hbc8e1857),
	.w7(32'h3ae2944e),
	.w8(32'h3caa433e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0fe0b8),
	.w1(32'h3ca8ed84),
	.w2(32'hbd64fe7e),
	.w3(32'h3c8481a1),
	.w4(32'hbc5a0120),
	.w5(32'hbc6765ca),
	.w6(32'h3c44a1d9),
	.w7(32'hbc636c20),
	.w8(32'hbce84f8f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca18ee4),
	.w1(32'h3c916b30),
	.w2(32'h3b3a7ac9),
	.w3(32'hbcc92fc3),
	.w4(32'h3a73c6bf),
	.w5(32'hbae2e8db),
	.w6(32'h3c17e01e),
	.w7(32'hb9abfa94),
	.w8(32'hbcb3502d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdf56a4),
	.w1(32'h3bba0b84),
	.w2(32'h3c25221a),
	.w3(32'hbca003ba),
	.w4(32'hbb39bf1c),
	.w5(32'hbc845901),
	.w6(32'h3a9a6326),
	.w7(32'hbc3b28b6),
	.w8(32'hbc56cb26),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc901828),
	.w1(32'h3c418838),
	.w2(32'hbbe9321b),
	.w3(32'hbc79a35f),
	.w4(32'h3c0a0f02),
	.w5(32'hbadd5361),
	.w6(32'h3bd0fed0),
	.w7(32'hbb547249),
	.w8(32'hbbc27d96),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a97e4),
	.w1(32'hbc0bc97c),
	.w2(32'hbbd629a8),
	.w3(32'hbb9fe171),
	.w4(32'h3b3cf4c2),
	.w5(32'hbbbf563c),
	.w6(32'hbb1c46fa),
	.w7(32'hbba6945d),
	.w8(32'h3b99d07f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d729f),
	.w1(32'hbd0812ad),
	.w2(32'h3b88f5ce),
	.w3(32'h3b86dd25),
	.w4(32'hbc90b368),
	.w5(32'h3aab34c7),
	.w6(32'hbc86f5df),
	.w7(32'hbc0df620),
	.w8(32'h3c1fd62c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d047df9),
	.w1(32'hbc77de0f),
	.w2(32'h3cb08198),
	.w3(32'h3c012f00),
	.w4(32'hbc7e5093),
	.w5(32'hbd08a93b),
	.w6(32'hbcc7690b),
	.w7(32'hbcece8a2),
	.w8(32'hbc34c30d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2f78d),
	.w1(32'hbba0aa02),
	.w2(32'hbc20234d),
	.w3(32'hbcb68fb4),
	.w4(32'hbb9aa6b9),
	.w5(32'hbbab8f2e),
	.w6(32'hbb263851),
	.w7(32'hbb14d67e),
	.w8(32'hbb608abd),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc540e0b),
	.w1(32'hbbe5e3fd),
	.w2(32'hbc31f7c9),
	.w3(32'hbbd4c699),
	.w4(32'h39bd8cc5),
	.w5(32'hbbb30c35),
	.w6(32'hbc09e637),
	.w7(32'hbbef6d13),
	.w8(32'hbc12fee0),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e2180),
	.w1(32'h3bd476cb),
	.w2(32'h3b0ae26b),
	.w3(32'h3b5f6505),
	.w4(32'h3bd42bb0),
	.w5(32'h3acace3f),
	.w6(32'h3b1559c2),
	.w7(32'hbb76997f),
	.w8(32'hbc2d4f69),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa427c5),
	.w1(32'hbc361ae4),
	.w2(32'hbb969eec),
	.w3(32'h3a7beb85),
	.w4(32'hb92cac3f),
	.w5(32'hbb31e956),
	.w6(32'hbba1c204),
	.w7(32'hb714ad57),
	.w8(32'h3b97ad75),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c531c3f),
	.w1(32'hbb161f6c),
	.w2(32'hbb8ff775),
	.w3(32'h3b5f8dda),
	.w4(32'hbc1896e7),
	.w5(32'hbb0e57c4),
	.w6(32'hbbdad0e5),
	.w7(32'hbbd61506),
	.w8(32'hbcaa4af1),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34d052),
	.w1(32'h3c6a785f),
	.w2(32'h3b164aa2),
	.w3(32'hbc7a2e88),
	.w4(32'h3ba3983c),
	.w5(32'h3aae3c22),
	.w6(32'h3c4d1904),
	.w7(32'h3b9b8e0c),
	.w8(32'hbb5eeb75),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1848fa),
	.w1(32'h3bae5e19),
	.w2(32'hbbff96c9),
	.w3(32'hbb934f0f),
	.w4(32'hbae7546a),
	.w5(32'hbbefc5bc),
	.w6(32'hba8a3f8b),
	.w7(32'hbc278956),
	.w8(32'hbc0b92bc),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba25474),
	.w1(32'hbb80a882),
	.w2(32'h3c1a06ec),
	.w3(32'hbb9736b0),
	.w4(32'hbc50e9d0),
	.w5(32'hbce666f4),
	.w6(32'hbbb3ac74),
	.w7(32'hbcc7c4b6),
	.w8(32'hbc34943d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc128053),
	.w1(32'hbc36844c),
	.w2(32'hba995f62),
	.w3(32'hbb9132d0),
	.w4(32'hbc44d972),
	.w5(32'hbaae4c17),
	.w6(32'hbc52ebfc),
	.w7(32'hbaa582cc),
	.w8(32'hbbc443e8),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb443e4d),
	.w1(32'hbc28782d),
	.w2(32'h38c32ad7),
	.w3(32'hbb4cdcb6),
	.w4(32'hbb7d7179),
	.w5(32'h3ab3dfe8),
	.w6(32'h3b99a3a5),
	.w7(32'h3a4a7439),
	.w8(32'h3c3af663),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94fde9),
	.w1(32'h3b5d6b55),
	.w2(32'h3b87c759),
	.w3(32'h3ad93e11),
	.w4(32'h3a1e7026),
	.w5(32'h3b9fccc8),
	.w6(32'h3b5fc528),
	.w7(32'h3b6cc0e7),
	.w8(32'hbaf4ec5b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fbad6),
	.w1(32'hbd0068de),
	.w2(32'h3ceeefe2),
	.w3(32'h3ac15efa),
	.w4(32'hbca876bc),
	.w5(32'hbca1dbcc),
	.w6(32'hbcbd3957),
	.w7(32'hbc25dfbb),
	.w8(32'h3c8222c2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1dbcad),
	.w1(32'h3b2edbeb),
	.w2(32'hbb83d0f3),
	.w3(32'h3c86fdcb),
	.w4(32'h3a51c944),
	.w5(32'h3b3f1013),
	.w6(32'h3a347039),
	.w7(32'h3aca0c7f),
	.w8(32'h3aa18b1b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c0292),
	.w1(32'hbb1a342f),
	.w2(32'h3bfc19c5),
	.w3(32'h3bdb36fe),
	.w4(32'h3b275fd3),
	.w5(32'h3afc0f44),
	.w6(32'hbaa388f4),
	.w7(32'h3a50efb5),
	.w8(32'hb9d3e8f7),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9cfb4),
	.w1(32'hbb6f69ce),
	.w2(32'hbc0b43a0),
	.w3(32'hbb95d692),
	.w4(32'hbaccae98),
	.w5(32'hbb8416a9),
	.w6(32'h3a2b12ca),
	.w7(32'hbb326cc7),
	.w8(32'hbbad2854),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80b793),
	.w1(32'h39b2785c),
	.w2(32'hbaabf308),
	.w3(32'hbab5bc48),
	.w4(32'h3a6b114e),
	.w5(32'h3a93d236),
	.w6(32'h3b14e478),
	.w7(32'h3ad64794),
	.w8(32'h3bafd6d3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b065ee5),
	.w1(32'h3c2a116a),
	.w2(32'hbb8506a0),
	.w3(32'h3b0ce3c0),
	.w4(32'h3a4076fe),
	.w5(32'h3ad5e5ce),
	.w6(32'h3b8e99d2),
	.w7(32'h38541278),
	.w8(32'hbbf4d1d7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf04078),
	.w1(32'hbc85a157),
	.w2(32'h3a4f56c3),
	.w3(32'h3bf2c963),
	.w4(32'hbc892b9d),
	.w5(32'h3b4c8629),
	.w6(32'hbc95c8a0),
	.w7(32'hbb2b3dcb),
	.w8(32'hbb0c9ad4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe2691),
	.w1(32'hbc065a2f),
	.w2(32'h3b882aaa),
	.w3(32'h3bd023b3),
	.w4(32'h3aa8dad3),
	.w5(32'hbb85a623),
	.w6(32'h3b4b5ec4),
	.w7(32'h3a987165),
	.w8(32'h3beb6d17),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78a278),
	.w1(32'hbc442043),
	.w2(32'hbb8d2d5f),
	.w3(32'h3ba54548),
	.w4(32'hbbef6bf3),
	.w5(32'h39c5b206),
	.w6(32'hbc24da08),
	.w7(32'h3a1f8143),
	.w8(32'hbbd17c6a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cabf0),
	.w1(32'h3c3e8e06),
	.w2(32'hbcd6fcc4),
	.w3(32'h3b4940e2),
	.w4(32'h3c460a5d),
	.w5(32'hbc542d6a),
	.w6(32'h3c629b12),
	.w7(32'hbc6bd70d),
	.w8(32'hbc535aa8),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc285e53),
	.w1(32'hb988e845),
	.w2(32'h3aa69daa),
	.w3(32'hbc067d6e),
	.w4(32'hb89fdc81),
	.w5(32'hbb048317),
	.w6(32'hb8ffa266),
	.w7(32'hbbe3c179),
	.w8(32'h3a101a0a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c034869),
	.w1(32'hbc1aa8ef),
	.w2(32'hb9b59add),
	.w3(32'h3bdcbcbd),
	.w4(32'hbad910b3),
	.w5(32'h3aaa3c93),
	.w6(32'h3bc8b3ce),
	.w7(32'hba230e2d),
	.w8(32'h3b8c7738),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0db387),
	.w1(32'hb9bde6ae),
	.w2(32'h3c02567a),
	.w3(32'h3ac5f8a2),
	.w4(32'hbb9ff5de),
	.w5(32'h3bc74d78),
	.w6(32'hbb09668d),
	.w7(32'h3ba8b53d),
	.w8(32'hbb85dcfb),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfc303),
	.w1(32'h3be6b971),
	.w2(32'hbb2b3818),
	.w3(32'hbb12d331),
	.w4(32'hb986a8e5),
	.w5(32'h3b2cd260),
	.w6(32'h3c33b9c5),
	.w7(32'h3b96ac46),
	.w8(32'hbb9fb687),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6ea3f),
	.w1(32'h3bd542d8),
	.w2(32'h3abdfa65),
	.w3(32'h3a9bc35b),
	.w4(32'hbadc4eb6),
	.w5(32'h3b22451e),
	.w6(32'hba6f48b7),
	.w7(32'hba36fa2f),
	.w8(32'h3adbd1eb),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66f408),
	.w1(32'hbcc7b4b1),
	.w2(32'hbbb5fd53),
	.w3(32'hbc300942),
	.w4(32'hbc3f6492),
	.w5(32'hbb88a495),
	.w6(32'hbc58e0d6),
	.w7(32'hbb2e883a),
	.w8(32'hbc81c014),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc119828),
	.w1(32'hbbc29445),
	.w2(32'h3c6e783a),
	.w3(32'h3975a3ed),
	.w4(32'hbb88df1a),
	.w5(32'h3bdddb40),
	.w6(32'hbaeefe19),
	.w7(32'h3bbfdbb2),
	.w8(32'h3bc84cba),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12ad9b),
	.w1(32'hbd11d658),
	.w2(32'h3ba59b26),
	.w3(32'h3b8039f0),
	.w4(32'hbcb9ee59),
	.w5(32'h3ba4d6ec),
	.w6(32'hbcf6176d),
	.w7(32'hba9686de),
	.w8(32'h3b66321e),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d086cef),
	.w1(32'hbb0dc11b),
	.w2(32'hba8dbba7),
	.w3(32'h3c83989e),
	.w4(32'h39878d38),
	.w5(32'hb99bcbe5),
	.w6(32'hb8ff3655),
	.w7(32'hba76efb3),
	.w8(32'h3b5062c2),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae10223),
	.w1(32'h3c237299),
	.w2(32'hbada2796),
	.w3(32'h3b202cd0),
	.w4(32'h3b77421a),
	.w5(32'hb966b362),
	.w6(32'h3b783cbe),
	.w7(32'hbb36414a),
	.w8(32'hbc10e0e0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e392f),
	.w1(32'h3a495a72),
	.w2(32'h3b4fcbbc),
	.w3(32'hbb6d4f45),
	.w4(32'h3a0ece29),
	.w5(32'h3b90f406),
	.w6(32'hbc0bc1f8),
	.w7(32'h3ace3264),
	.w8(32'h3c10b64c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a364733),
	.w1(32'hbc3f8835),
	.w2(32'hbbdae512),
	.w3(32'hbb4aaac8),
	.w4(32'hbb922263),
	.w5(32'hba9c6d44),
	.w6(32'hbc06ca7a),
	.w7(32'hbb909161),
	.w8(32'hbb4f2297),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3847ea),
	.w1(32'hbc68e217),
	.w2(32'h3b7d9206),
	.w3(32'hbb9404a6),
	.w4(32'hbc8238d1),
	.w5(32'h3b61c5b2),
	.w6(32'hbcb2350a),
	.w7(32'hbbe2837e),
	.w8(32'h3bace7f1),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c412bc4),
	.w1(32'h3cef5cbc),
	.w2(32'h3b8b5779),
	.w3(32'h3c41844f),
	.w4(32'h3c8dbd75),
	.w5(32'h3c113eb8),
	.w6(32'h3c7de480),
	.w7(32'h3a9ae370),
	.w8(32'hbc4a352f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9fe580),
	.w1(32'hbada152a),
	.w2(32'hbc26a8d7),
	.w3(32'hb9b22b34),
	.w4(32'h3beac582),
	.w5(32'hbbb201b0),
	.w6(32'h3c5ec3a5),
	.w7(32'hbb604d90),
	.w8(32'h3b5be6b5),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba1808),
	.w1(32'h3ad2e9b5),
	.w2(32'h3b739af5),
	.w3(32'hbb01af49),
	.w4(32'h39df42fb),
	.w5(32'h3b34bddc),
	.w6(32'h3b5182e8),
	.w7(32'h3af896c7),
	.w8(32'h3936ea28),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa94ecf),
	.w1(32'h3b8488f9),
	.w2(32'h3c02cdc4),
	.w3(32'h3b42d35f),
	.w4(32'h3c3b6e95),
	.w5(32'h3ca7c794),
	.w6(32'h39229c42),
	.w7(32'hbc1a8515),
	.w8(32'hbc944718),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce31654),
	.w1(32'hbb9db1ff),
	.w2(32'h391c55aa),
	.w3(32'hbc0083d2),
	.w4(32'hba342ee8),
	.w5(32'hbbb2f9c1),
	.w6(32'hbb875d9b),
	.w7(32'h398ae1b4),
	.w8(32'h3ae63348),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9918f),
	.w1(32'h3c8def86),
	.w2(32'hbc4e1189),
	.w3(32'hbb60a5fb),
	.w4(32'h3bfe2e73),
	.w5(32'h3b93c6da),
	.w6(32'h3ab71a2b),
	.w7(32'h3a85ce40),
	.w8(32'hbbb70415),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a3790),
	.w1(32'h3bc1cb63),
	.w2(32'h3c0bf091),
	.w3(32'hbbe54ad4),
	.w4(32'h3ab7ba25),
	.w5(32'h3b96cd8a),
	.w6(32'h3b0d4d95),
	.w7(32'h3b913a91),
	.w8(32'hbaabd219),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f2b47),
	.w1(32'h3cc429a1),
	.w2(32'h398fff56),
	.w3(32'hbafca676),
	.w4(32'h3bbeb42a),
	.w5(32'hbb1d7a19),
	.w6(32'h3c2a36ae),
	.w7(32'h3b978dd9),
	.w8(32'hbca710a7),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc9a3ff),
	.w1(32'hbcbe7716),
	.w2(32'hbc541d02),
	.w3(32'hbbe72e71),
	.w4(32'hbc931997),
	.w5(32'hbd60f3a2),
	.w6(32'hbcab79d6),
	.w7(32'hbd3a2319),
	.w8(32'hbc4f0c51),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc905636),
	.w1(32'h3ba7e136),
	.w2(32'h3d0798a5),
	.w3(32'hbcbc80d2),
	.w4(32'h3b143289),
	.w5(32'hbbe0c1f5),
	.w6(32'h3b2f609b),
	.w7(32'hbaeed3f8),
	.w8(32'hbc2f8a50),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd23c9f4),
	.w1(32'hbcae2e32),
	.w2(32'h3b799f6d),
	.w3(32'hbcf1944b),
	.w4(32'hbbec465c),
	.w5(32'hbb43f902),
	.w6(32'hbc8f3ad0),
	.w7(32'hbbb4fdcb),
	.w8(32'h3c283640),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad637d),
	.w1(32'hbbc96475),
	.w2(32'h3c0d9ce3),
	.w3(32'h3baa180e),
	.w4(32'hb96a215a),
	.w5(32'h3a296bfa),
	.w6(32'hbbba5c8f),
	.w7(32'hbbe31c3a),
	.w8(32'hbbb31b73),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba41aa9),
	.w1(32'hbb8b3228),
	.w2(32'h3b1802ef),
	.w3(32'h39536ea9),
	.w4(32'h3a309b83),
	.w5(32'hbb485952),
	.w6(32'h39f82ff8),
	.w7(32'hb9c8a1a7),
	.w8(32'h3b77f691),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c3669),
	.w1(32'hbaf7240c),
	.w2(32'hbbba0bd5),
	.w3(32'hbb37cb57),
	.w4(32'h39ee0280),
	.w5(32'hbab6ddae),
	.w6(32'hbbbef303),
	.w7(32'hbbabf02d),
	.w8(32'hbac13532),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8773f9),
	.w1(32'h3984b81b),
	.w2(32'h3a241b93),
	.w3(32'h3b03425c),
	.w4(32'hbb1ec42e),
	.w5(32'hba99445f),
	.w6(32'hbaf8369f),
	.w7(32'hbab91d90),
	.w8(32'hba86ed24),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eadf24),
	.w1(32'hbbac9f86),
	.w2(32'hbb9a8edc),
	.w3(32'h39cfe97f),
	.w4(32'hba8221db),
	.w5(32'hba935a16),
	.w6(32'hba5198ef),
	.w7(32'hbb045811),
	.w8(32'h3b30e145),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad56fd7),
	.w1(32'hbc0df974),
	.w2(32'h3b9d6062),
	.w3(32'h3ac05f89),
	.w4(32'hba9489fc),
	.w5(32'hbb394f7d),
	.w6(32'hbafa1ccf),
	.w7(32'hb96eb333),
	.w8(32'h3bd6a439),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ef196),
	.w1(32'hbc92b667),
	.w2(32'hbc01db53),
	.w3(32'h3b845a9a),
	.w4(32'hbc86d658),
	.w5(32'hba15ab0f),
	.w6(32'hbc2f42ce),
	.w7(32'h3a7a9780),
	.w8(32'h3c5ee75f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0f794e),
	.w1(32'h3c40df97),
	.w2(32'hbc5c219c),
	.w3(32'h3c378cd5),
	.w4(32'h3b79f314),
	.w5(32'hbb0d36f0),
	.w6(32'h3c270551),
	.w7(32'hb7b61abb),
	.w8(32'hbbb98923),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc30bb3),
	.w1(32'hbcc74206),
	.w2(32'hbd1f305c),
	.w3(32'hbbd2f59c),
	.w4(32'hbcb208fb),
	.w5(32'hbc9bcb7b),
	.w6(32'hbcf28b46),
	.w7(32'hbcb965bb),
	.w8(32'hbd073fa5),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40f329),
	.w1(32'h3c3c2965),
	.w2(32'hbb8a68a8),
	.w3(32'hbd030c54),
	.w4(32'h3b2fb701),
	.w5(32'hb9ae9f76),
	.w6(32'h3c244a66),
	.w7(32'h3b266e24),
	.w8(32'hbc2e81ed),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c1b6d),
	.w1(32'hbbb0af75),
	.w2(32'hb9afc45c),
	.w3(32'hbc449aa4),
	.w4(32'hbb2f96d3),
	.w5(32'h3b22bf78),
	.w6(32'hbbb80f07),
	.w7(32'hbaa5824d),
	.w8(32'hbaeb699a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33f15d),
	.w1(32'hbccc2a4b),
	.w2(32'hba61f001),
	.w3(32'h3bf81433),
	.w4(32'hbc5f9857),
	.w5(32'hbad259e4),
	.w6(32'hbc9964f7),
	.w7(32'hbbc3244c),
	.w8(32'h3bcf77d3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf0b5f7),
	.w1(32'hbc1fa97a),
	.w2(32'h3b9bd97c),
	.w3(32'h3c1fbe05),
	.w4(32'hbaa33a1f),
	.w5(32'hbbb29b9e),
	.w6(32'hbaccefd7),
	.w7(32'hba829c1a),
	.w8(32'h3be88fc4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c812b4c),
	.w1(32'hba903fac),
	.w2(32'h3b420e3c),
	.w3(32'h3b9608aa),
	.w4(32'h3b4405b6),
	.w5(32'hbb257af1),
	.w6(32'hb8acc46b),
	.w7(32'hba740e1f),
	.w8(32'hbaa5b6a8),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb537f09),
	.w1(32'h3bb62f83),
	.w2(32'h3b847431),
	.w3(32'hbae6aaa6),
	.w4(32'h3be534ae),
	.w5(32'hbae43c87),
	.w6(32'h3bb281d0),
	.w7(32'hba3e3145),
	.w8(32'hbb66ff5d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e73fd),
	.w1(32'hbccea66e),
	.w2(32'hbc94e4b6),
	.w3(32'hbc10ed1d),
	.w4(32'hbc5d4bb0),
	.w5(32'hbc6cca04),
	.w6(32'hbc46070e),
	.w7(32'hbc1a9435),
	.w8(32'h3ae02a8c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7fd45),
	.w1(32'hbbb410e7),
	.w2(32'hbc215de9),
	.w3(32'hbc770cc4),
	.w4(32'hbbe19d92),
	.w5(32'hbc978f58),
	.w6(32'hb81e6a25),
	.w7(32'hbca7c5f4),
	.w8(32'hbb86e750),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1af718),
	.w1(32'h3bc4a053),
	.w2(32'h3c0d43c9),
	.w3(32'h3b509492),
	.w4(32'h3b99c10e),
	.w5(32'hbb1a35d8),
	.w6(32'h3bb3c70a),
	.w7(32'h3b066c54),
	.w8(32'hbb887fa4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ec221),
	.w1(32'h3c79a823),
	.w2(32'hbb9b2c80),
	.w3(32'hbc7cf1e1),
	.w4(32'h3ba248d9),
	.w5(32'hba1ba791),
	.w6(32'h3bad09eb),
	.w7(32'hbb622937),
	.w8(32'hbc4b45e9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ac7bf),
	.w1(32'hbb9e5c90),
	.w2(32'hbab6014a),
	.w3(32'hbc6d3edd),
	.w4(32'h3a1249f9),
	.w5(32'hbae1058c),
	.w6(32'hbabb3722),
	.w7(32'hba5de99b),
	.w8(32'hba8a8c3e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b261391),
	.w1(32'hbc3558bf),
	.w2(32'hbc4353c1),
	.w3(32'hba980b57),
	.w4(32'hbb866b19),
	.w5(32'h3b6ec553),
	.w6(32'hbb98d78e),
	.w7(32'hbc8d1a8f),
	.w8(32'hbb6677a1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72e471),
	.w1(32'h3cc74058),
	.w2(32'h3cad5583),
	.w3(32'hbc84a9a5),
	.w4(32'h3c3ffced),
	.w5(32'h3c465146),
	.w6(32'h3c5a2400),
	.w7(32'h3b8ff5c4),
	.w8(32'hbc90759c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd21a76b),
	.w1(32'h392a83d6),
	.w2(32'hbb3a3a72),
	.w3(32'hbcb2a9eb),
	.w4(32'h3a806c23),
	.w5(32'hbbd9af6e),
	.w6(32'hba838072),
	.w7(32'hbbc56d19),
	.w8(32'hbba2fd3e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a743791),
	.w1(32'h3905892a),
	.w2(32'hb7b9e8f2),
	.w3(32'h3b3ba89d),
	.w4(32'hb7c61f86),
	.w5(32'hb9003582),
	.w6(32'hb8f8427d),
	.w7(32'hb90c922a),
	.w8(32'hb9a00358),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf21264),
	.w1(32'hbb417fc0),
	.w2(32'hb9bcce5d),
	.w3(32'hbb0b3453),
	.w4(32'hbaea65e1),
	.w5(32'h3a92af49),
	.w6(32'hbb783999),
	.w7(32'h3a8efe08),
	.w8(32'hb9941a99),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule