module layer_8_featuremap_250(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d392d),
	.w1(32'h3c64cf94),
	.w2(32'h3c5fa10e),
	.w3(32'hbb1af8e5),
	.w4(32'h3adda091),
	.w5(32'h3c80e02a),
	.w6(32'h3b359bdb),
	.w7(32'h395b9029),
	.w8(32'h3ba5839b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f43ea),
	.w1(32'hbbf7a5f7),
	.w2(32'hbc4d72a9),
	.w3(32'h3b9b8ddf),
	.w4(32'hbb898d87),
	.w5(32'hbc09a40e),
	.w6(32'hbc04112b),
	.w7(32'hbc746b9a),
	.w8(32'hbc1f5515),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3fb12),
	.w1(32'hbb90f652),
	.w2(32'hbc3c0e74),
	.w3(32'hbb28610c),
	.w4(32'hbbc862a5),
	.w5(32'hbc6f231d),
	.w6(32'h3b41e40e),
	.w7(32'h3b889331),
	.w8(32'hb9d07f6d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc310615),
	.w1(32'h3b62bbef),
	.w2(32'h3c0d04c3),
	.w3(32'hbc08aeea),
	.w4(32'h3bd6562b),
	.w5(32'h3acbe5c2),
	.w6(32'h3b9f4fd3),
	.w7(32'h3c15bf3c),
	.w8(32'h3bec44aa),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20a847),
	.w1(32'hbaa64806),
	.w2(32'hbb007144),
	.w3(32'h3b96fb24),
	.w4(32'h3b34e110),
	.w5(32'h3b0a27de),
	.w6(32'hbb941ebc),
	.w7(32'hbb4afa03),
	.w8(32'hbb18a5c8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bc6b6),
	.w1(32'h3bacabeb),
	.w2(32'h3bba9167),
	.w3(32'h3b28c752),
	.w4(32'hb90a71ce),
	.w5(32'h3b868717),
	.w6(32'hbb1a09c0),
	.w7(32'hba482502),
	.w8(32'hba9b9803),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0dc488),
	.w1(32'h3c3ce83f),
	.w2(32'h3c6e99a4),
	.w3(32'hba094a5a),
	.w4(32'h3c2045f2),
	.w5(32'h3c6d4547),
	.w6(32'h3b18f637),
	.w7(32'h3c1fedb2),
	.w8(32'h3bf54f75),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3de687),
	.w1(32'h3b05bd2c),
	.w2(32'h3c43205f),
	.w3(32'h3c0d5cba),
	.w4(32'h3c26a55a),
	.w5(32'h3ced38f4),
	.w6(32'hbc8302c5),
	.w7(32'h3af932f4),
	.w8(32'hb9c22b8c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccbdba9),
	.w1(32'h3ac764e5),
	.w2(32'hbc5067df),
	.w3(32'h3ccca1c7),
	.w4(32'h3bf39607),
	.w5(32'hbc06952e),
	.w6(32'hbac95ad3),
	.w7(32'hbc546e2c),
	.w8(32'hbbc4806c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb538b54),
	.w1(32'h3c2aa664),
	.w2(32'h3c6bfdd2),
	.w3(32'hbb38ce50),
	.w4(32'h3bbb24d5),
	.w5(32'h3c3dd9bc),
	.w6(32'hbb143d6e),
	.w7(32'h3b1b6856),
	.w8(32'h3bcbe164),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77ed51),
	.w1(32'h3c1fc69c),
	.w2(32'h3cdfe6f5),
	.w3(32'h3c2b9fc8),
	.w4(32'h3af3dd91),
	.w5(32'h3c2b1f1a),
	.w6(32'h3b951bd9),
	.w7(32'h3b8f6a08),
	.w8(32'hbb802112),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e2b0e),
	.w1(32'h3a960984),
	.w2(32'h3ace7dfd),
	.w3(32'h3c81c13a),
	.w4(32'hba1e1deb),
	.w5(32'hbb102e88),
	.w6(32'hbba0d6a0),
	.w7(32'hb9ed1e24),
	.w8(32'hbbbba1f3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b1865),
	.w1(32'h3beafa6f),
	.w2(32'h3c65f5f7),
	.w3(32'hbc2c25b0),
	.w4(32'h39b5eabc),
	.w5(32'hbbc4173c),
	.w6(32'h3c387ef1),
	.w7(32'hbaccd4ed),
	.w8(32'h3ae9d774),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a1142),
	.w1(32'hbc81a5d0),
	.w2(32'hbd048423),
	.w3(32'h3b051c2e),
	.w4(32'hbc143261),
	.w5(32'hbc4eb164),
	.w6(32'h3ba0eb3d),
	.w7(32'hbc0178a3),
	.w8(32'hbbdc780b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb624c4),
	.w1(32'h3bb41bb2),
	.w2(32'h3b4cb119),
	.w3(32'hbbbc1041),
	.w4(32'h3ad219f9),
	.w5(32'h3a8eb5e1),
	.w6(32'h3b09ccba),
	.w7(32'h3b3c6e35),
	.w8(32'h3b4633b7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13f1a8),
	.w1(32'h3c9a9145),
	.w2(32'h3c991446),
	.w3(32'hbb8b4b36),
	.w4(32'h3c078214),
	.w5(32'h3c07cdd7),
	.w6(32'h3c45fcad),
	.w7(32'h3c816c0f),
	.w8(32'h3bdc9b54),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be48f6f),
	.w1(32'h3ce52318),
	.w2(32'h3c966f2d),
	.w3(32'h38c616fa),
	.w4(32'h3bc230e8),
	.w5(32'h3a182606),
	.w6(32'h3ca1a11e),
	.w7(32'h3c9a524e),
	.w8(32'h3a9d45da),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2be40),
	.w1(32'hbc11c8ce),
	.w2(32'hbcb36f65),
	.w3(32'hbaddb982),
	.w4(32'hbb47f8cf),
	.w5(32'hbc8ee5d3),
	.w6(32'hbb833e24),
	.w7(32'hbc48824b),
	.w8(32'h3bacdc7a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf11093),
	.w1(32'h3c6738e7),
	.w2(32'h3cb9ffae),
	.w3(32'hbb6b4fae),
	.w4(32'h3c65af24),
	.w5(32'h3cb33c9e),
	.w6(32'h3bfb76f5),
	.w7(32'h3ad57e04),
	.w8(32'h3af3099a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c176768),
	.w1(32'h3b007384),
	.w2(32'hba0de6f1),
	.w3(32'h3b9426fe),
	.w4(32'h3a2d7613),
	.w5(32'hbb51dfaa),
	.w6(32'h3abb5b17),
	.w7(32'hba4fa3f9),
	.w8(32'hbac42cb4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32b9d6),
	.w1(32'h3b30d9a0),
	.w2(32'h3bccba0f),
	.w3(32'hbb59bdff),
	.w4(32'h3c021c35),
	.w5(32'h3a3adbed),
	.w6(32'hbb32e3d6),
	.w7(32'h3bade416),
	.w8(32'h3916c0af),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccd48d),
	.w1(32'hbc0b48de),
	.w2(32'hbc82e00f),
	.w3(32'hba2f4248),
	.w4(32'hbc99db56),
	.w5(32'hbcadcf1c),
	.w6(32'hbc1ca5c9),
	.w7(32'hbca31de8),
	.w8(32'hbc75fc0f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f88c0),
	.w1(32'h37ab67c6),
	.w2(32'h3c5303bc),
	.w3(32'hbc550bbe),
	.w4(32'h3b8a6d6d),
	.w5(32'h3c090add),
	.w6(32'h3c327f95),
	.w7(32'h3bab94d7),
	.w8(32'h3b42098e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7154de),
	.w1(32'hbcdd587a),
	.w2(32'hbd171a31),
	.w3(32'h3c566d5c),
	.w4(32'hbcc7fbf5),
	.w5(32'hbce2c02c),
	.w6(32'hbc8e1d13),
	.w7(32'hbcce31f3),
	.w8(32'hbca0ac52),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce0a566),
	.w1(32'hbb602526),
	.w2(32'hbb1bb803),
	.w3(32'hbcc8cd4a),
	.w4(32'h3ab80d02),
	.w5(32'h3b345e02),
	.w6(32'hbb1e341d),
	.w7(32'hbc2d2039),
	.w8(32'hbc47eee0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc67ba),
	.w1(32'h3b9efc50),
	.w2(32'h3c7eed51),
	.w3(32'hbb786b2e),
	.w4(32'h3be6923e),
	.w5(32'h3cae4005),
	.w6(32'h3b91db1c),
	.w7(32'hba911a74),
	.w8(32'h3c4e108b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c696d52),
	.w1(32'h3bd1880a),
	.w2(32'h3c6cde7a),
	.w3(32'h3c7875da),
	.w4(32'h3c2c717a),
	.w5(32'h3c7f4347),
	.w6(32'hbbbc14b0),
	.w7(32'h3bd71942),
	.w8(32'h3b1433aa),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22f27a),
	.w1(32'h3c1459f8),
	.w2(32'h3c757051),
	.w3(32'h3b8c7b99),
	.w4(32'h3c9b216e),
	.w5(32'h3c42b2b4),
	.w6(32'h3c003ad3),
	.w7(32'h3c6528c0),
	.w8(32'h3bf3679c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c946bee),
	.w1(32'h3afe5a36),
	.w2(32'hbb433ad0),
	.w3(32'h3c7d4cb4),
	.w4(32'h3b9abb5d),
	.w5(32'h395ba480),
	.w6(32'hbb641fe2),
	.w7(32'hbc70c254),
	.w8(32'hbbfabbe5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65de17),
	.w1(32'hbb3ed0cd),
	.w2(32'hba97e29d),
	.w3(32'h39239266),
	.w4(32'h3bb042f2),
	.w5(32'h3c2b9db6),
	.w6(32'hbb6fcacb),
	.w7(32'hbacb0746),
	.w8(32'hbb8f5b9f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1a5fe),
	.w1(32'h3c1e8026),
	.w2(32'h3c851038),
	.w3(32'h3af2fb5d),
	.w4(32'h3a61529e),
	.w5(32'h3b555114),
	.w6(32'h3c0beaf6),
	.w7(32'h3c0d1c5f),
	.w8(32'h3b419dce),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82eb02),
	.w1(32'h3b1e6f2f),
	.w2(32'hbbb275f6),
	.w3(32'h3ba51267),
	.w4(32'h3a2238bb),
	.w5(32'hbc105316),
	.w6(32'h3b85f4d7),
	.w7(32'hbc1ba146),
	.w8(32'hbbe5af22),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e10ce),
	.w1(32'hbbdc86a8),
	.w2(32'hbc762531),
	.w3(32'hbbe8da4f),
	.w4(32'hbbc26891),
	.w5(32'hbc31c152),
	.w6(32'hbb98141a),
	.w7(32'hbbb33df1),
	.w8(32'h39ab08b8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9adeb4),
	.w1(32'h3c67f2f3),
	.w2(32'h3ca792b7),
	.w3(32'h3b2d9a7a),
	.w4(32'h3c20aa59),
	.w5(32'h3c6a45a5),
	.w6(32'h3c7f6dea),
	.w7(32'h3cbee978),
	.w8(32'h3c18a17c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d748d),
	.w1(32'hbaa7f74c),
	.w2(32'hbbc92fae),
	.w3(32'h3ca43ba0),
	.w4(32'h39d890be),
	.w5(32'hbb8e2d9c),
	.w6(32'h3ba03093),
	.w7(32'hbb9cd668),
	.w8(32'h3b03dfd2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ca4fb),
	.w1(32'h3cafd1e3),
	.w2(32'h3cebcb3f),
	.w3(32'h3b1b6163),
	.w4(32'h3c2de06e),
	.w5(32'h3c8672d0),
	.w6(32'h3c019b1f),
	.w7(32'h3c3990d1),
	.w8(32'h3c841878),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd7139e),
	.w1(32'h3a407a71),
	.w2(32'h3a8e868b),
	.w3(32'h3c4961de),
	.w4(32'h3b206849),
	.w5(32'h3afec1e0),
	.w6(32'hba999f21),
	.w7(32'hb9f406ef),
	.w8(32'h3a535dbc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba899a6b),
	.w1(32'h3b1a1ac1),
	.w2(32'hbbb97661),
	.w3(32'h3a6ce198),
	.w4(32'h3a5a019c),
	.w5(32'hbbab6a1e),
	.w6(32'h3b825a9f),
	.w7(32'hbaebc326),
	.w8(32'h3b6666ae),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9aaf48),
	.w1(32'h3b18f868),
	.w2(32'h3b6a0c70),
	.w3(32'h3adcb1b5),
	.w4(32'h3b276466),
	.w5(32'h3bc8fda7),
	.w6(32'hbb4243f3),
	.w7(32'hba0ecaf1),
	.w8(32'h3b2a3da9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8050fb),
	.w1(32'h3ce4d7e9),
	.w2(32'h3d68ce51),
	.w3(32'h3baf96f4),
	.w4(32'h3cdb30a7),
	.w5(32'h3d3139e2),
	.w6(32'h3c1df3be),
	.w7(32'h3cb11de6),
	.w8(32'h3cd35635),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2be4ca),
	.w1(32'hbbfd2930),
	.w2(32'hbcaf0ccc),
	.w3(32'h3cb03e70),
	.w4(32'hbb89f510),
	.w5(32'hbc9c1b54),
	.w6(32'h39d2b100),
	.w7(32'hbc4d0bd9),
	.w8(32'hba1d18d7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1554bf),
	.w1(32'h3bb12504),
	.w2(32'h3b80d66c),
	.w3(32'hbbfa8abb),
	.w4(32'h39e7551a),
	.w5(32'hbc065706),
	.w6(32'h3b9a0399),
	.w7(32'h3bc3103f),
	.w8(32'hbb46e9d8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe37dd),
	.w1(32'hb9b51737),
	.w2(32'hbb52dc59),
	.w3(32'h399ab15d),
	.w4(32'h3b6c11bc),
	.w5(32'h3c030e0c),
	.w6(32'hbbe859ee),
	.w7(32'hbb8c8b18),
	.w8(32'hbc14ec5a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde6dc6),
	.w1(32'h3b6935a4),
	.w2(32'hbc416a88),
	.w3(32'h352a5ad7),
	.w4(32'h3a1db074),
	.w5(32'h3a95708a),
	.w6(32'h3a865528),
	.w7(32'h3b8c00fe),
	.w8(32'h39accb53),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b072b),
	.w1(32'h3c0c72a5),
	.w2(32'hbbdfb22c),
	.w3(32'h3c0bd446),
	.w4(32'h3be436db),
	.w5(32'hbb43fdcf),
	.w6(32'h39ca85ab),
	.w7(32'hbcb99d3f),
	.w8(32'hbc13411f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40275b),
	.w1(32'hbbd605c4),
	.w2(32'hbbee3cb8),
	.w3(32'h3b99c23f),
	.w4(32'hbbf721bd),
	.w5(32'hbbe7f984),
	.w6(32'hbc467da8),
	.w7(32'hbc6accc7),
	.w8(32'hbbf1ac7b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3418bb),
	.w1(32'h3c8ece2a),
	.w2(32'h3ce39a5c),
	.w3(32'hbbad9062),
	.w4(32'h3c8424a8),
	.w5(32'h3cc1e59d),
	.w6(32'h39bf62fc),
	.w7(32'h3c2aba19),
	.w8(32'h3bc38301),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c913304),
	.w1(32'hbc6dbfb9),
	.w2(32'hbc85b977),
	.w3(32'h3bdbe53b),
	.w4(32'hbc7a58a2),
	.w5(32'hbc5fe156),
	.w6(32'hbc91bd72),
	.w7(32'hbc6b8648),
	.w8(32'hbc617d80),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc708ef6),
	.w1(32'hbcad9f40),
	.w2(32'hbcda4034),
	.w3(32'hbc264e2a),
	.w4(32'hbbd70cd5),
	.w5(32'hbc4c1a3a),
	.w6(32'hbbe853a1),
	.w7(32'hbc7f56f3),
	.w8(32'hbc3ccb15),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca05377),
	.w1(32'h3c05ee27),
	.w2(32'hba621c84),
	.w3(32'hbba7dee9),
	.w4(32'h3b6787a7),
	.w5(32'h39e85232),
	.w6(32'h3bdab38f),
	.w7(32'h3c1a7b38),
	.w8(32'h3c26ce2a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a246c),
	.w1(32'hbc00cf65),
	.w2(32'hbc1feede),
	.w3(32'h3b88d3d7),
	.w4(32'hbb0f9a00),
	.w5(32'hbc1effd2),
	.w6(32'hbb01ffe5),
	.w7(32'hbc014b58),
	.w8(32'hba18d195),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826974),
	.w1(32'h3ad36696),
	.w2(32'hbc1f5fcd),
	.w3(32'h3a92c4ae),
	.w4(32'h3b62a665),
	.w5(32'hbbe9d4b6),
	.w6(32'hbb200b0a),
	.w7(32'hbc536db1),
	.w8(32'hbb58e937),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8e654),
	.w1(32'hbaaee540),
	.w2(32'hbbd0757f),
	.w3(32'h3a049f22),
	.w4(32'hbb227cad),
	.w5(32'hbba464ed),
	.w6(32'hbbbb8514),
	.w7(32'hbc23129b),
	.w8(32'hbb05e892),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e58af),
	.w1(32'h3b860ecf),
	.w2(32'h3c8d9973),
	.w3(32'h3b8af95f),
	.w4(32'h3be7d18b),
	.w5(32'h3c48c0e1),
	.w6(32'h3b18be89),
	.w7(32'h3cb9f903),
	.w8(32'h3bde3bb6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09bdf2),
	.w1(32'h3c9da9a2),
	.w2(32'h3c2bc37e),
	.w3(32'h3c255da2),
	.w4(32'h3c43b8a5),
	.w5(32'h3c6bb023),
	.w6(32'h3c85505c),
	.w7(32'h3bc21fa3),
	.w8(32'h3c7f0ae8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3225d7),
	.w1(32'hbc8bfa6f),
	.w2(32'hbcfff265),
	.w3(32'h3c497156),
	.w4(32'hbc8deeb3),
	.w5(32'hbd0bf05c),
	.w6(32'hbc831749),
	.w7(32'hbc994e2d),
	.w8(32'hbc7e6dd7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92e92c),
	.w1(32'hba56f352),
	.w2(32'h3bc90dcd),
	.w3(32'hbc831ece),
	.w4(32'h3bcd156a),
	.w5(32'h3ba4832e),
	.w6(32'h3ba0359b),
	.w7(32'h3bb46e60),
	.w8(32'hbab90254),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b951e34),
	.w1(32'h3b9d9188),
	.w2(32'h3b296240),
	.w3(32'h3c835ea7),
	.w4(32'h3bb59420),
	.w5(32'h3b1d075f),
	.w6(32'h3b1431f5),
	.w7(32'hbb719f0b),
	.w8(32'hba2f3a75),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bc253),
	.w1(32'h3ab753a7),
	.w2(32'h3b6caa91),
	.w3(32'h394758f3),
	.w4(32'h3aee7fde),
	.w5(32'h3a9a669f),
	.w6(32'h3a73810b),
	.w7(32'h3b8f07b7),
	.w8(32'h3b15e9d8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8dd12),
	.w1(32'hbc9571be),
	.w2(32'hbc9286e9),
	.w3(32'hba9e4015),
	.w4(32'hbc46300e),
	.w5(32'hbc8ed439),
	.w6(32'hbc1ef48d),
	.w7(32'hbc952335),
	.w8(32'hbc9b575c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b04e0),
	.w1(32'h3c849dfd),
	.w2(32'h3bac832b),
	.w3(32'hbc0cb7ae),
	.w4(32'h3a504788),
	.w5(32'h3c367251),
	.w6(32'h3bbf0439),
	.w7(32'h3bba2771),
	.w8(32'h3b1542d9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6a627),
	.w1(32'hbb1558c0),
	.w2(32'h3a04b96e),
	.w3(32'h3c8553e4),
	.w4(32'hbbeefe03),
	.w5(32'h39f6e5b3),
	.w6(32'hbadffd30),
	.w7(32'hbbe7e5b0),
	.w8(32'hba2e98bb),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf5db6),
	.w1(32'hbabcabc4),
	.w2(32'hbc1c2cbb),
	.w3(32'hbbb9da4b),
	.w4(32'hbad0ae13),
	.w5(32'hbb7b6f70),
	.w6(32'hb8fc4b40),
	.w7(32'hbc5b31bb),
	.w8(32'hbc196f7b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd32155),
	.w1(32'hbb7fd259),
	.w2(32'hbc07ea3b),
	.w3(32'h39cb8740),
	.w4(32'hb9f58c15),
	.w5(32'hbbc3bd96),
	.w6(32'hb985e357),
	.w7(32'h3a2561fa),
	.w8(32'h3b3b720f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65af6a),
	.w1(32'h3b0ba9cb),
	.w2(32'h39370a1d),
	.w3(32'hbbc381a2),
	.w4(32'h3ba76535),
	.w5(32'h3ad711ee),
	.w6(32'h3ada7f11),
	.w7(32'h39e0bd01),
	.w8(32'h3a56b124),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba439c9f),
	.w1(32'h3c8dde32),
	.w2(32'h3d428d6c),
	.w3(32'hb97d58ce),
	.w4(32'h3caf02f4),
	.w5(32'h3d08e53e),
	.w6(32'h3ab43ae4),
	.w7(32'h3c5d6141),
	.w8(32'h3c703857),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd08277),
	.w1(32'h3c881857),
	.w2(32'h3c48a928),
	.w3(32'h3c66b8a5),
	.w4(32'h3c5e4c61),
	.w5(32'h3c211de0),
	.w6(32'hba216ad9),
	.w7(32'h3bfb428a),
	.w8(32'hbae34c80),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb45d92),
	.w1(32'h3c70b4f8),
	.w2(32'h3c991ed6),
	.w3(32'hbb8e0eda),
	.w4(32'h3bf53775),
	.w5(32'h3c1fceb3),
	.w6(32'h3b959cec),
	.w7(32'h3bc731f5),
	.w8(32'hbba118ac),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a3b31),
	.w1(32'hbc42acaf),
	.w2(32'hbd0f4a22),
	.w3(32'hbb5f5757),
	.w4(32'hbc683766),
	.w5(32'hbcc5f8fb),
	.w6(32'hbc112594),
	.w7(32'hbc8f216b),
	.w8(32'hbc277e1a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62ac5b),
	.w1(32'h3b5b935c),
	.w2(32'hbc5196e8),
	.w3(32'hbc36c50e),
	.w4(32'hbbf002ea),
	.w5(32'hbb007b4a),
	.w6(32'h3c36f7f3),
	.w7(32'hbadbcb07),
	.w8(32'h3b9a7e71),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7a211),
	.w1(32'hbb0709e1),
	.w2(32'hbba04c97),
	.w3(32'h3bd94445),
	.w4(32'h3c03d415),
	.w5(32'h3b8cc168),
	.w6(32'hbc26f8dd),
	.w7(32'hbc4e02c3),
	.w8(32'hbc61f2fe),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc84988),
	.w1(32'h3b08b374),
	.w2(32'hbb8e6d48),
	.w3(32'hbb167556),
	.w4(32'h3bb259e6),
	.w5(32'h3b3f4192),
	.w6(32'h3c10d0bb),
	.w7(32'h3bef2e08),
	.w8(32'h3bc0b965),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c83a5a),
	.w1(32'h3c17979b),
	.w2(32'h3a8cac71),
	.w3(32'h3b06e70b),
	.w4(32'h3b657de5),
	.w5(32'h3c1a64b0),
	.w6(32'h3bce2ebf),
	.w7(32'h3bd0e114),
	.w8(32'h3bd5ccdf),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb929c79),
	.w1(32'h3c40c3d8),
	.w2(32'h3bd0ebd9),
	.w3(32'h3c1c63bd),
	.w4(32'h3bbc1a06),
	.w5(32'h3bff99ca),
	.w6(32'h3c1933a3),
	.w7(32'h3b4c2a15),
	.w8(32'h3b2593c7),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7feac),
	.w1(32'h398def40),
	.w2(32'h3b2b4b2c),
	.w3(32'h3b96a50b),
	.w4(32'hbafbcd07),
	.w5(32'hba87e78e),
	.w6(32'h3b3ed2f3),
	.w7(32'h3b19ab02),
	.w8(32'h3a82c1bb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add4a99),
	.w1(32'h3c2c83e8),
	.w2(32'h3b0764c3),
	.w3(32'hba8a4702),
	.w4(32'h3bae949d),
	.w5(32'h3b88ad84),
	.w6(32'h3c482d24),
	.w7(32'h3c011e70),
	.w8(32'h3c434764),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44f92e),
	.w1(32'h3b7f850e),
	.w2(32'h3bf0b3dc),
	.w3(32'h3c2f3c2e),
	.w4(32'h3b41ddbe),
	.w5(32'h3bf401ec),
	.w6(32'hbb83145b),
	.w7(32'h3b174166),
	.w8(32'h3b01c9cf),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae82b0),
	.w1(32'hbb5b1b97),
	.w2(32'hbb148c3a),
	.w3(32'h3b04ee23),
	.w4(32'hbb2f2019),
	.w5(32'hbb573f93),
	.w6(32'hbbbefe14),
	.w7(32'hbaac70b6),
	.w8(32'h3b87bcbd),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94069fc),
	.w1(32'hba6a1ad1),
	.w2(32'h3bf7401a),
	.w3(32'hb926ae03),
	.w4(32'h3bbf899b),
	.w5(32'h3bc01df6),
	.w6(32'hbbb47970),
	.w7(32'h39987552),
	.w8(32'hbb0980d3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae90413),
	.w1(32'hbc82c300),
	.w2(32'hbc9a5f89),
	.w3(32'h3b0d285d),
	.w4(32'hbc5f206c),
	.w5(32'hbc68e3c6),
	.w6(32'hbb1662fd),
	.w7(32'hba954931),
	.w8(32'h3b1dfb73),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf80c5),
	.w1(32'h3ae8f6b8),
	.w2(32'hbb89ca87),
	.w3(32'h3bfc5123),
	.w4(32'h3ac99722),
	.w5(32'h3a8333bb),
	.w6(32'h3bca736e),
	.w7(32'h3b97bf06),
	.w8(32'h3c13c18f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc26f27),
	.w1(32'hbcca21e6),
	.w2(32'hbd1c9579),
	.w3(32'h3bd93419),
	.w4(32'hbca28a4d),
	.w5(32'hbce8473b),
	.w6(32'hbc85831c),
	.w7(32'hbcbf4e23),
	.w8(32'hbc97f6ae),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1ca30),
	.w1(32'hb81da890),
	.w2(32'hbbbb00fb),
	.w3(32'hbcb03c6e),
	.w4(32'h3afa1560),
	.w5(32'hbbe58581),
	.w6(32'h3bdb4691),
	.w7(32'hbb17e198),
	.w8(32'h3aebfae2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23f936),
	.w1(32'h3b0a78b1),
	.w2(32'h3c65454a),
	.w3(32'h3bd2ad8f),
	.w4(32'h3b911fb8),
	.w5(32'h3c846028),
	.w6(32'h3a144d5d),
	.w7(32'h3ba30c6a),
	.w8(32'h3c1eaff8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68cd3d),
	.w1(32'hbb8b7d6d),
	.w2(32'hbc560646),
	.w3(32'h3b7f27c5),
	.w4(32'hbc34969e),
	.w5(32'hbc47d31a),
	.w6(32'h3bd93b9c),
	.w7(32'h3b32874b),
	.w8(32'h3a32ca78),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc37260),
	.w1(32'hbb804d6d),
	.w2(32'hbadffd0a),
	.w3(32'hbbc6efe0),
	.w4(32'hbb57c137),
	.w5(32'hba2c9f03),
	.w6(32'h3b6da7d0),
	.w7(32'h3afc2801),
	.w8(32'h3bb3d34f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19640e),
	.w1(32'hba32a490),
	.w2(32'hbb90ffdb),
	.w3(32'h3be560f7),
	.w4(32'hbb3e940b),
	.w5(32'hbc022305),
	.w6(32'h3927ce23),
	.w7(32'hbb825b32),
	.w8(32'hbbcb3348),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81a31d),
	.w1(32'h3b289a04),
	.w2(32'hbc0d6038),
	.w3(32'hbc0a2697),
	.w4(32'h3c429956),
	.w5(32'h3bc0edf9),
	.w6(32'h3b720f15),
	.w7(32'hbbf13f4f),
	.w8(32'hbbd3e734),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc900d82),
	.w1(32'hbbaadc5d),
	.w2(32'hbba961dc),
	.w3(32'hbb8ee5da),
	.w4(32'hba9aa0c5),
	.w5(32'hbbae5bb1),
	.w6(32'h3ac719f0),
	.w7(32'h39e7ee11),
	.w8(32'h3a0e8d31),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8a6d2),
	.w1(32'h3b211e5b),
	.w2(32'hbc1d8cce),
	.w3(32'hbb05bfdb),
	.w4(32'hbc08482e),
	.w5(32'hbc23ab65),
	.w6(32'h3be4b231),
	.w7(32'h3b300b5a),
	.w8(32'h3bcd4d90),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1320f6),
	.w1(32'h3c2edd40),
	.w2(32'h3c3eed23),
	.w3(32'h3a6b2862),
	.w4(32'h3c54859a),
	.w5(32'h3bfb3864),
	.w6(32'h3c401e6d),
	.w7(32'h3c495aa7),
	.w8(32'h3c21a057),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5b8a1),
	.w1(32'h3c76f802),
	.w2(32'h3c878c7d),
	.w3(32'h3b67ae95),
	.w4(32'h3c12b504),
	.w5(32'h3c8c3d6c),
	.w6(32'h3c28ea94),
	.w7(32'h3c646b07),
	.w8(32'h3c31b8f1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb79886),
	.w1(32'hbba80ff2),
	.w2(32'hbb71a585),
	.w3(32'h3c8765a7),
	.w4(32'hbac7e5b3),
	.w5(32'hbaf6f344),
	.w6(32'hbb991e71),
	.w7(32'hbbe05874),
	.w8(32'hbbb21246),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a280c),
	.w1(32'h3b72c863),
	.w2(32'h3bce1cf2),
	.w3(32'h3ac226f1),
	.w4(32'h3bed8fc7),
	.w5(32'h3c0646ed),
	.w6(32'h3b318caa),
	.w7(32'h3b5e3d7a),
	.w8(32'h3b9f5f6b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f391d),
	.w1(32'h3cbecda0),
	.w2(32'h3c934d8c),
	.w3(32'h3beb196a),
	.w4(32'h3c23a3d5),
	.w5(32'h3c906b82),
	.w6(32'h3c500280),
	.w7(32'h3baaea6f),
	.w8(32'h3c65c1a2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca412c5),
	.w1(32'hba006948),
	.w2(32'hbb2ded43),
	.w3(32'h3c0936df),
	.w4(32'hbb3677a3),
	.w5(32'hbbc2dfd1),
	.w6(32'hba828fcc),
	.w7(32'hbb77bb2c),
	.w8(32'hbb0765f1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba889a62),
	.w1(32'h3b985ed2),
	.w2(32'h3be633bc),
	.w3(32'hbb06b78a),
	.w4(32'h3b05eece),
	.w5(32'h3b2f03ff),
	.w6(32'h3c5ac93b),
	.w7(32'h3bd006ff),
	.w8(32'h3c56fa7b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce535d),
	.w1(32'h3c323c58),
	.w2(32'hba6bc75a),
	.w3(32'h3b8012e4),
	.w4(32'h3bda0339),
	.w5(32'h3b5baed5),
	.w6(32'h3ba28d55),
	.w7(32'h3b7e443a),
	.w8(32'h3c1272f0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f2827),
	.w1(32'h3bfed7c0),
	.w2(32'hba349d65),
	.w3(32'h3c5c1a5a),
	.w4(32'h3bb9f182),
	.w5(32'h3b170e52),
	.w6(32'h3c0faeda),
	.w7(32'h3bedfbed),
	.w8(32'h3be2862a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc607cc),
	.w1(32'h3c38b6fc),
	.w2(32'h3ccf70b0),
	.w3(32'h3c573903),
	.w4(32'h3c0642eb),
	.w5(32'h3c81dc41),
	.w6(32'hb9243ff8),
	.w7(32'h3c1bea94),
	.w8(32'hbb1482ec),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96a9bc),
	.w1(32'h3c2c30ab),
	.w2(32'h3cb8e654),
	.w3(32'h3c7642f1),
	.w4(32'h3bcb7e37),
	.w5(32'h3be012fc),
	.w6(32'h3b192d83),
	.w7(32'h3c42814d),
	.w8(32'h3b2b3469),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be57a08),
	.w1(32'hbc0df94e),
	.w2(32'hbc1702c8),
	.w3(32'h3be2faea),
	.w4(32'hbb9e4307),
	.w5(32'h3662410b),
	.w6(32'hbc227c1f),
	.w7(32'hbc74c9c3),
	.w8(32'hbca2c144),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc172025),
	.w1(32'hbc3111ff),
	.w2(32'hbc8b1a80),
	.w3(32'hbbda33af),
	.w4(32'hbbfedb8a),
	.w5(32'hbc90ae08),
	.w6(32'hbac3ea3f),
	.w7(32'hbb64884c),
	.w8(32'hbc073d52),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3da830),
	.w1(32'h3c6d8b7a),
	.w2(32'h3c93f228),
	.w3(32'hbc55e151),
	.w4(32'h3bb34b4b),
	.w5(32'h3bef754a),
	.w6(32'h3c4b108e),
	.w7(32'h3c3b10f3),
	.w8(32'h3c2eb4ba),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf97dfe),
	.w1(32'h3ad57f0d),
	.w2(32'h3c1eb959),
	.w3(32'h3ca0e3ae),
	.w4(32'h3b506eab),
	.w5(32'h3b91b59a),
	.w6(32'h3bcfc06e),
	.w7(32'h3bd8a471),
	.w8(32'h3b8bf732),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb973a1d),
	.w1(32'h3b8d1641),
	.w2(32'hbb670dff),
	.w3(32'h3af14786),
	.w4(32'hb9c49166),
	.w5(32'hbbfbc25a),
	.w6(32'hba88f6f6),
	.w7(32'hbc09d0e2),
	.w8(32'hbb10c688),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26ba5f),
	.w1(32'h3bba5050),
	.w2(32'hb9cefeef),
	.w3(32'hb9fb0add),
	.w4(32'h3bd951e1),
	.w5(32'h3b698760),
	.w6(32'h3ba9a0ce),
	.w7(32'h3b84bcbb),
	.w8(32'h3b95540f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b991b02),
	.w1(32'h3b60a3f8),
	.w2(32'h3bee1851),
	.w3(32'h3ba5e9b3),
	.w4(32'h3bb53f4b),
	.w5(32'h3ba488dc),
	.w6(32'h3bb4f0d8),
	.w7(32'h3bc0c903),
	.w8(32'h3ba06d11),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a05b6),
	.w1(32'h3c95d47e),
	.w2(32'h3cec1515),
	.w3(32'h3bd45bed),
	.w4(32'h3c8be712),
	.w5(32'h3cc7c62a),
	.w6(32'h3a285e76),
	.w7(32'h3c2e01c3),
	.w8(32'h3c0df1e1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ce26d),
	.w1(32'h3c0bc26b),
	.w2(32'h3c0cfe00),
	.w3(32'h3c08048f),
	.w4(32'h3c11089c),
	.w5(32'h3c12b227),
	.w6(32'h3bf32ee8),
	.w7(32'h3bb07b05),
	.w8(32'h3bc66824),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28cdf1),
	.w1(32'hbc5e8d71),
	.w2(32'hbcc21fd4),
	.w3(32'h3c4046a6),
	.w4(32'hbc432b32),
	.w5(32'hbc7c9b0d),
	.w6(32'hbc1eb76d),
	.w7(32'hbb49d872),
	.w8(32'hbc1811e0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc851042),
	.w1(32'h3b5a8fe7),
	.w2(32'h3baa8b55),
	.w3(32'hbc267660),
	.w4(32'h3bff320f),
	.w5(32'h3b8daabd),
	.w6(32'h3ad07cc5),
	.w7(32'h3b5b9752),
	.w8(32'h3bb8c920),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf956a),
	.w1(32'h3d3e4695),
	.w2(32'h3dab0e18),
	.w3(32'h3a81c591),
	.w4(32'h3cf67709),
	.w5(32'h3d7942be),
	.w6(32'h3ce44de6),
	.w7(32'h3d5b7032),
	.w8(32'h3c212444),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2b7682),
	.w1(32'h3c1cb48e),
	.w2(32'h3c66a2d9),
	.w3(32'h3cadbf86),
	.w4(32'h3c87c6ec),
	.w5(32'h3c8fe62e),
	.w6(32'h3b9a501b),
	.w7(32'h3ad61159),
	.w8(32'hbabaa042),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20c0d7),
	.w1(32'hbc279a25),
	.w2(32'hbbfd16c8),
	.w3(32'h3c210b7b),
	.w4(32'hbc4d1dc3),
	.w5(32'hbc55d47b),
	.w6(32'hbb0245ba),
	.w7(32'hba3d9fb3),
	.w8(32'hbb6e9acd),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb857034),
	.w1(32'h3b024c16),
	.w2(32'hba1160b2),
	.w3(32'hbc0436d3),
	.w4(32'h3b6e1b6a),
	.w5(32'h3b3279aa),
	.w6(32'h3b142811),
	.w7(32'hbac728fc),
	.w8(32'h3ace281a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e49ec),
	.w1(32'h3a861eac),
	.w2(32'hbc250184),
	.w3(32'h3be939ef),
	.w4(32'h3ac72212),
	.w5(32'hbbc0d99b),
	.w6(32'h3aea4215),
	.w7(32'hbc445777),
	.w8(32'hbbbcd9bb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb918780),
	.w1(32'h3c9d2b32),
	.w2(32'h3d298ac4),
	.w3(32'h3b94e03d),
	.w4(32'h3c5f2003),
	.w5(32'h3cf88b8b),
	.w6(32'h3c6b2b01),
	.w7(32'h3d0247b3),
	.w8(32'h3c9b7d65),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce1b3a5),
	.w1(32'h3c55c00c),
	.w2(32'h3c8b74ce),
	.w3(32'h3cdde59e),
	.w4(32'h3c048975),
	.w5(32'h3ca71206),
	.w6(32'h3c6cea37),
	.w7(32'h3cb00914),
	.w8(32'h3c55d336),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c930960),
	.w1(32'hbad577af),
	.w2(32'h3b079130),
	.w3(32'h3ca0a63e),
	.w4(32'hbb4f5b9b),
	.w5(32'hbb94df7c),
	.w6(32'h391c839e),
	.w7(32'h3ae312a0),
	.w8(32'hbaa92083),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385375a4),
	.w1(32'hbcb66784),
	.w2(32'hbd16cc57),
	.w3(32'hbb8ebca3),
	.w4(32'hbcc82649),
	.w5(32'hbce2cde2),
	.w6(32'hbc8f8fa7),
	.w7(32'hbcbb5f36),
	.w8(32'hbc7982d5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86df79),
	.w1(32'hbaa86c27),
	.w2(32'hbb5fb1d9),
	.w3(32'hbc7338d5),
	.w4(32'hbb383018),
	.w5(32'hbb5a03ba),
	.w6(32'hba09d955),
	.w7(32'hbb06430b),
	.w8(32'hbc0e87c6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ae07a),
	.w1(32'h3b601f0e),
	.w2(32'h3bb69b33),
	.w3(32'hbb51c8ec),
	.w4(32'h3c0105c9),
	.w5(32'h3bb31dd1),
	.w6(32'h3b045dbf),
	.w7(32'h3b3bdb52),
	.w8(32'h3b7c716d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0079c1),
	.w1(32'h3d0c3839),
	.w2(32'h3d8111b6),
	.w3(32'h3bdf94f2),
	.w4(32'h3cb0b4d0),
	.w5(32'h3d20a962),
	.w6(32'h3c719abd),
	.w7(32'h3d27556f),
	.w8(32'h3c0ca8c1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf43289),
	.w1(32'h3c60a46f),
	.w2(32'h3c1e31de),
	.w3(32'h3c351e68),
	.w4(32'h3c6fcfe0),
	.w5(32'h3c5cc1e4),
	.w6(32'h3c3a5afd),
	.w7(32'h3ab587c2),
	.w8(32'h3c3c7e4c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38b779),
	.w1(32'hbc4c7ae0),
	.w2(32'hbbeef4f3),
	.w3(32'h3c595cea),
	.w4(32'hbc86ba0b),
	.w5(32'hbba7d7c4),
	.w6(32'hbc519b3e),
	.w7(32'hbc8bd4c4),
	.w8(32'hbc03582e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ef7d9),
	.w1(32'h3ab483a5),
	.w2(32'h3ad279dc),
	.w3(32'hba77e035),
	.w4(32'h3a18f0ce),
	.w5(32'hb9120460),
	.w6(32'h3a003e67),
	.w7(32'h3993fae2),
	.w8(32'h3a7b24a3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a876d7b),
	.w1(32'h3b5ab32a),
	.w2(32'hbc1e9767),
	.w3(32'h39be1cf0),
	.w4(32'hba3f140a),
	.w5(32'hbbc1c14c),
	.w6(32'h3b87fdec),
	.w7(32'hbbafb6c4),
	.w8(32'hbba349d5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule