module layer_8_featuremap_186(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b6bbf),
	.w1(32'hbbdbb8ee),
	.w2(32'h3badb9cc),
	.w3(32'hbb4a82ee),
	.w4(32'h3bc98a9a),
	.w5(32'h3b8263ba),
	.w6(32'hbb87b2fa),
	.w7(32'h3bfd94eb),
	.w8(32'h3bbdd4da),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3eae38),
	.w1(32'hbaf962b7),
	.w2(32'hbba8377e),
	.w3(32'hba439855),
	.w4(32'hbab62249),
	.w5(32'hba25c1f6),
	.w6(32'h396cae1b),
	.w7(32'hbb520dd0),
	.w8(32'hbbfe5b75),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37d0f7),
	.w1(32'hbb1f9115),
	.w2(32'hbbbbf4e3),
	.w3(32'hbbbb3cc1),
	.w4(32'hba6356de),
	.w5(32'h390c6362),
	.w6(32'hbb8665fc),
	.w7(32'hbb94691b),
	.w8(32'hbb142e81),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3dc08d),
	.w1(32'h3bb79f63),
	.w2(32'h3cc684f1),
	.w3(32'h3a89a9f5),
	.w4(32'hbb64d543),
	.w5(32'h3bc5cc69),
	.w6(32'h3b7b77f1),
	.w7(32'h3be18407),
	.w8(32'hbb733366),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad7c37),
	.w1(32'hbb0fd51e),
	.w2(32'h3b1ffab9),
	.w3(32'h3ba23d03),
	.w4(32'hbb735343),
	.w5(32'h3aa432e3),
	.w6(32'h39dc1aaf),
	.w7(32'hba0dbb1d),
	.w8(32'hbb967653),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b042d47),
	.w1(32'h3c3a461c),
	.w2(32'h3c8b15eb),
	.w3(32'h3b436edc),
	.w4(32'h3c42ce58),
	.w5(32'h3c8b18e8),
	.w6(32'h3c31b407),
	.w7(32'h3c5ee6de),
	.w8(32'h3b53348a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f1b43),
	.w1(32'hbbe2f0fd),
	.w2(32'hbb88b34d),
	.w3(32'h3c2a4283),
	.w4(32'hbba10b43),
	.w5(32'hbbd38008),
	.w6(32'hbb9394ae),
	.w7(32'hbb1ce1a6),
	.w8(32'h3a29787c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93aef0e),
	.w1(32'h3b9f1910),
	.w2(32'h3bf5058f),
	.w3(32'hb98f9038),
	.w4(32'h3bc822d0),
	.w5(32'h3be74d61),
	.w6(32'h3b6574ae),
	.w7(32'h3c13bbc4),
	.w8(32'h3b5b3c44),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c8c79),
	.w1(32'hbbf93695),
	.w2(32'h3a8eea7e),
	.w3(32'hbc085e22),
	.w4(32'hbbd35c8b),
	.w5(32'hb9bfc2c5),
	.w6(32'h3a8e10a6),
	.w7(32'h3be5d833),
	.w8(32'hbae3cc92),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba971e9c),
	.w1(32'h3bfd24f5),
	.w2(32'h3c87f916),
	.w3(32'h3af7c752),
	.w4(32'h3b3766d3),
	.w5(32'h3c587dea),
	.w6(32'h3bebf5da),
	.w7(32'h3c1d5c60),
	.w8(32'h3c0ea9b9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31fd1a),
	.w1(32'h3c33383c),
	.w2(32'hbc0c695c),
	.w3(32'h3c702a90),
	.w4(32'h3c9c5ecf),
	.w5(32'h3bc24f75),
	.w6(32'hbc06bd34),
	.w7(32'hbca7d405),
	.w8(32'hbc28c67a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca37492),
	.w1(32'h3926b3ce),
	.w2(32'h3a9064e5),
	.w3(32'hbc4ce1cd),
	.w4(32'hbaab1fad),
	.w5(32'h3b635f90),
	.w6(32'h3b328304),
	.w7(32'h3ae9f802),
	.w8(32'hbaa03ae9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f2985),
	.w1(32'h3ca7b532),
	.w2(32'h3ca55e69),
	.w3(32'h38aa0064),
	.w4(32'h3c249a43),
	.w5(32'h3c9679d6),
	.w6(32'h3c3ebc81),
	.w7(32'h3bf2135d),
	.w8(32'hbad3cf21),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cf621),
	.w1(32'hbb77ad81),
	.w2(32'hbc05ec73),
	.w3(32'h3c946dc5),
	.w4(32'hbc2a57d1),
	.w5(32'hbb426a14),
	.w6(32'hbc6d7fd7),
	.w7(32'hbbe43f31),
	.w8(32'hbb832461),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b9286),
	.w1(32'hbc5fd9bb),
	.w2(32'hbbdc5f4a),
	.w3(32'hbb5f24c8),
	.w4(32'hbc2ecca0),
	.w5(32'hbc37fe45),
	.w6(32'hbbf6fb6e),
	.w7(32'h3b256bfd),
	.w8(32'h3c0a766d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bdcd3),
	.w1(32'h3ba0ded6),
	.w2(32'h3b5798ff),
	.w3(32'hbb29f4f1),
	.w4(32'hbb40e196),
	.w5(32'h39f443ac),
	.w6(32'hbb98a3a9),
	.w7(32'hbbaa84ed),
	.w8(32'hbbc695a7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6dd921),
	.w1(32'hbb2a834b),
	.w2(32'h3bdb504a),
	.w3(32'h3bca8dc7),
	.w4(32'hbc0e8159),
	.w5(32'h3b749ac6),
	.w6(32'h3bf8af04),
	.w7(32'h3a54dc04),
	.w8(32'h3ad35da8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18601d),
	.w1(32'hbae7f941),
	.w2(32'hbc561551),
	.w3(32'h396e8974),
	.w4(32'hbc189a48),
	.w5(32'hbc0c475e),
	.w6(32'hbc0f7084),
	.w7(32'hbc553828),
	.w8(32'hbc346a6f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7fef71),
	.w1(32'h3d0bc022),
	.w2(32'h3cec679a),
	.w3(32'hbc7cdb24),
	.w4(32'h3be88b24),
	.w5(32'h3cf4d3f3),
	.w6(32'h3c88a026),
	.w7(32'h3aaf6818),
	.w8(32'hbc07e5e5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bf721f),
	.w1(32'hbb63a5f2),
	.w2(32'hbb9af559),
	.w3(32'h3c395dca),
	.w4(32'hbacc04ff),
	.w5(32'hbbc159a9),
	.w6(32'hbb8fc608),
	.w7(32'h390e4a1e),
	.w8(32'h3bad831f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f4972),
	.w1(32'hbc5ac361),
	.w2(32'hbbd94242),
	.w3(32'hb9bb9eea),
	.w4(32'hbc20e724),
	.w5(32'hbca3477a),
	.w6(32'hbbd9a809),
	.w7(32'hbbc05dd5),
	.w8(32'h3a9d9f2f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95cce4),
	.w1(32'h3a789d9f),
	.w2(32'hb9f91489),
	.w3(32'hbbf76047),
	.w4(32'h3b5c5793),
	.w5(32'h39416d19),
	.w6(32'h3b92e6bb),
	.w7(32'h3bc024cf),
	.w8(32'hba5f27b4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d0c00),
	.w1(32'h3a4a407b),
	.w2(32'hbb85c656),
	.w3(32'hbb42b582),
	.w4(32'hbb0be0b4),
	.w5(32'hbb996f39),
	.w6(32'h3b24054f),
	.w7(32'h3b807024),
	.w8(32'h3b6a9c58),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54d878),
	.w1(32'h3b9b7ab4),
	.w2(32'hbab399b3),
	.w3(32'h3af10bfd),
	.w4(32'hbb28fa65),
	.w5(32'hbbcc359b),
	.w6(32'h3ac142b6),
	.w7(32'hbba3149e),
	.w8(32'h3a3cef8a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cd712),
	.w1(32'hbc134645),
	.w2(32'hbc8d4304),
	.w3(32'hbaad305a),
	.w4(32'hba10d79c),
	.w5(32'hbb337f99),
	.w6(32'hbbf9a664),
	.w7(32'hbc31731f),
	.w8(32'hbc17ee24),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86425c),
	.w1(32'hbb31cf2f),
	.w2(32'hbc889551),
	.w3(32'hbbffa5d3),
	.w4(32'hbbd7475e),
	.w5(32'hbc1b55a6),
	.w6(32'hbbb07db7),
	.w7(32'hbc391ef2),
	.w8(32'hbb92e753),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc452fbc),
	.w1(32'hba2183f1),
	.w2(32'hbc162874),
	.w3(32'hba751b2d),
	.w4(32'h3c229f5b),
	.w5(32'hbba83976),
	.w6(32'h3b9e7fbd),
	.w7(32'hbb2eaf5b),
	.w8(32'h3b9adc5d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f5772),
	.w1(32'h3a2cc469),
	.w2(32'h3cc4322a),
	.w3(32'hbcb03223),
	.w4(32'hbcb3a1de),
	.w5(32'h3b5a70db),
	.w6(32'hbc3ad295),
	.w7(32'h3bc52129),
	.w8(32'hbc6359df),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b0e3d),
	.w1(32'hbc24c630),
	.w2(32'hbc98d9a3),
	.w3(32'h3c0801d4),
	.w4(32'hbbb26fb6),
	.w5(32'hbc51d4b4),
	.w6(32'hbb1d5825),
	.w7(32'hbc390f52),
	.w8(32'h3a31bc44),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00dad6),
	.w1(32'hbb10aa5c),
	.w2(32'hba457a60),
	.w3(32'hbc33218e),
	.w4(32'hbb203855),
	.w5(32'hbb727a7e),
	.w6(32'hba6cb360),
	.w7(32'h3b102da8),
	.w8(32'h3c4e5a66),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7dc3c5),
	.w1(32'h3b7e5717),
	.w2(32'h3c809354),
	.w3(32'h3c41546e),
	.w4(32'hbb53802d),
	.w5(32'h3c2b2e72),
	.w6(32'h3bf1817a),
	.w7(32'h3c4cf43f),
	.w8(32'h3b73395f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdada4f),
	.w1(32'h3c39176c),
	.w2(32'hbc459d66),
	.w3(32'h3c60b150),
	.w4(32'h3c8c4935),
	.w5(32'h3c429d56),
	.w6(32'hbbdd4f40),
	.w7(32'hbcc4287a),
	.w8(32'hbcc37a69),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd056df3),
	.w1(32'hbc386dec),
	.w2(32'hbc6db8a4),
	.w3(32'hbc5949e1),
	.w4(32'h3bc6a89d),
	.w5(32'hbc5aa386),
	.w6(32'hbb2649b0),
	.w7(32'h3a02aa22),
	.w8(32'h3ba6a9c4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dcf6c),
	.w1(32'h3c4f7802),
	.w2(32'h3c867317),
	.w3(32'hbc3c41b5),
	.w4(32'h3c3e824d),
	.w5(32'h3c0b423c),
	.w6(32'h3c47650f),
	.w7(32'h3c73fc04),
	.w8(32'h3bcf46fd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be27cd3),
	.w1(32'hbb8fb298),
	.w2(32'h3b1525b0),
	.w3(32'h3c3dbe38),
	.w4(32'h3b824070),
	.w5(32'h3b6250f0),
	.w6(32'hbb3005bc),
	.w7(32'h3b92df13),
	.w8(32'h3b9b61dc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade85bc),
	.w1(32'hbbc3cf00),
	.w2(32'hbbe4ee62),
	.w3(32'h3b27ed6d),
	.w4(32'hbbf7ef1f),
	.w5(32'hbc090c42),
	.w6(32'hbb96c1c8),
	.w7(32'hbc1b8bd8),
	.w8(32'h3a42bb5b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe127ea),
	.w1(32'hbc1b66bb),
	.w2(32'hbc8bfd26),
	.w3(32'hba4911dd),
	.w4(32'hbb761ab8),
	.w5(32'hbc19fbfb),
	.w6(32'hbbf9e8af),
	.w7(32'hbc3df654),
	.w8(32'hbbedf7d0),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc565987),
	.w1(32'hbc57b136),
	.w2(32'h3b66399f),
	.w3(32'hbc2b56a0),
	.w4(32'hbc6448b4),
	.w5(32'hbb9dbf05),
	.w6(32'hbbed2e20),
	.w7(32'h3c127ff8),
	.w8(32'h3bea0337),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c1daa),
	.w1(32'hbb4a67cf),
	.w2(32'hbc0914ab),
	.w3(32'h3b8221d9),
	.w4(32'hbbef762e),
	.w5(32'hbc208708),
	.w6(32'hbbe10ecd),
	.w7(32'hbc0dee4b),
	.w8(32'hbbb5af97),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e83f4),
	.w1(32'h3bb2dc4d),
	.w2(32'h3b6e0c0d),
	.w3(32'hbc246dfb),
	.w4(32'hba5a627a),
	.w5(32'h3ae6bda3),
	.w6(32'h3a654a3a),
	.w7(32'hbac9f402),
	.w8(32'h3ab3b9b9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9ea32),
	.w1(32'h3c064fba),
	.w2(32'h3c02ed99),
	.w3(32'h3baf4279),
	.w4(32'h3bf3099e),
	.w5(32'h3c0e00ac),
	.w6(32'h3b6d6ac4),
	.w7(32'h3aa0908a),
	.w8(32'hb9bc1884),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b259fc7),
	.w1(32'h3c625e1a),
	.w2(32'h3cd0c970),
	.w3(32'h3b2a5989),
	.w4(32'h3aba1116),
	.w5(32'h3c9c9f08),
	.w6(32'h3c70a651),
	.w7(32'h3c8edd9f),
	.w8(32'h3a8378a8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c092099),
	.w1(32'hbc6d12e3),
	.w2(32'hbca0386d),
	.w3(32'h3c3fa8fd),
	.w4(32'hbb0ec3d2),
	.w5(32'hbc499cd9),
	.w6(32'hbc48a240),
	.w7(32'hbc6dbb5a),
	.w8(32'hbb474543),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3816fc),
	.w1(32'hbb91633a),
	.w2(32'hbc6e29ed),
	.w3(32'hbc6b9404),
	.w4(32'hbba4fd11),
	.w5(32'hbc844495),
	.w6(32'hbc24b7f1),
	.w7(32'hbc447c93),
	.w8(32'hbb249415),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f1e86),
	.w1(32'hbc426bc8),
	.w2(32'hbbee8ab3),
	.w3(32'hbc7d3f47),
	.w4(32'hbc1ab657),
	.w5(32'hbc5d01f8),
	.w6(32'hbc15ce08),
	.w7(32'h3abeff1c),
	.w8(32'hbaf1d522),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8915ea),
	.w1(32'h3a5b4d8b),
	.w2(32'hbbfde16c),
	.w3(32'hbb85f226),
	.w4(32'h3b9d3dde),
	.w5(32'hbb582393),
	.w6(32'h3b9eafcf),
	.w7(32'h3a4d6c67),
	.w8(32'h3abf3765),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb714d82),
	.w1(32'hbc87a02e),
	.w2(32'hbc95b046),
	.w3(32'hbade29e9),
	.w4(32'hbc39b01b),
	.w5(32'hbca0f872),
	.w6(32'hbc7ea394),
	.w7(32'hbc457425),
	.w8(32'hbc35ba90),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3224ec),
	.w1(32'h3bd89249),
	.w2(32'h3b27d5fd),
	.w3(32'hbc85ec3a),
	.w4(32'hbb2c412f),
	.w5(32'hb9ce9907),
	.w6(32'h3ae062b2),
	.w7(32'h3bddb69c),
	.w8(32'h3b2e0956),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dd217),
	.w1(32'hbb5a9148),
	.w2(32'hbb716d89),
	.w3(32'h3ba04780),
	.w4(32'h3b19a052),
	.w5(32'hbb7fdc14),
	.w6(32'h3ba09c02),
	.w7(32'hba988861),
	.w8(32'h3baeb8f8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d255a),
	.w1(32'h3cdb8890),
	.w2(32'h3cbf5159),
	.w3(32'h3b6eaa49),
	.w4(32'h3b988e78),
	.w5(32'h3c8e0fc4),
	.w6(32'h3c799863),
	.w7(32'h3b12d9de),
	.w8(32'hba5460db),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f99d2),
	.w1(32'h3b4261ff),
	.w2(32'h393403f4),
	.w3(32'h3c9a04a6),
	.w4(32'h399f9038),
	.w5(32'h3a3118df),
	.w6(32'h3ac1dd86),
	.w7(32'hb97e69eb),
	.w8(32'h3a7ca8af),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e987b),
	.w1(32'h3c8359fb),
	.w2(32'h3c66534f),
	.w3(32'hbb3f7869),
	.w4(32'h3be7160f),
	.w5(32'h3c00176f),
	.w6(32'h3be9d960),
	.w7(32'h3bc37a74),
	.w8(32'h3b2700b7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20584f),
	.w1(32'hbba22a5b),
	.w2(32'hb90434be),
	.w3(32'h3c346064),
	.w4(32'hbb55a0dc),
	.w5(32'h3a618ac3),
	.w6(32'hbb43f0ec),
	.w7(32'h3919dea3),
	.w8(32'hbb9c1bc8),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52e870),
	.w1(32'h3b0a50ea),
	.w2(32'hbbd47291),
	.w3(32'hbaf820be),
	.w4(32'hbae5afa6),
	.w5(32'hbb93f4f5),
	.w6(32'hb9692ea9),
	.w7(32'hbb8c913a),
	.w8(32'h3abe6604),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbc6c5),
	.w1(32'hbcebb9db),
	.w2(32'hbcb5ecce),
	.w3(32'hb9d58498),
	.w4(32'hbc820456),
	.w5(32'hbcdb4386),
	.w6(32'hbccc50d7),
	.w7(32'hbc54a612),
	.w8(32'h3bc57990),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93d13b),
	.w1(32'hbc48f8d4),
	.w2(32'hbc85c7cb),
	.w3(32'hbcd54565),
	.w4(32'h3b02f567),
	.w5(32'hbc9bb78c),
	.w6(32'hbc924d3b),
	.w7(32'hbc888e4e),
	.w8(32'hbb1afce0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22ef9c),
	.w1(32'h3bef75a5),
	.w2(32'hba95f71d),
	.w3(32'hbc48a21a),
	.w4(32'h3ba68bee),
	.w5(32'h3ba19c18),
	.w6(32'h394ecd1a),
	.w7(32'hbbb1c63b),
	.w8(32'hbb4d0991),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f7e74),
	.w1(32'hbbeabc89),
	.w2(32'hbca6632f),
	.w3(32'h3b548896),
	.w4(32'hb9fd5949),
	.w5(32'hbc5e9e82),
	.w6(32'hbbeeba1b),
	.w7(32'hbc48a41c),
	.w8(32'hbb9d8e40),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc817537),
	.w1(32'hbb84f28e),
	.w2(32'hbb85bbbe),
	.w3(32'hbc6bf11b),
	.w4(32'hbbac1f81),
	.w5(32'hbb83dc14),
	.w6(32'hbaf68607),
	.w7(32'hbb61b99d),
	.w8(32'h3abc574f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a65ec),
	.w1(32'h3a88c2ce),
	.w2(32'hbbcaf2c9),
	.w3(32'h39f4321b),
	.w4(32'hbbd2e1eb),
	.w5(32'h3b24c79f),
	.w6(32'h3b81d4ae),
	.w7(32'hba108a98),
	.w8(32'hbbad352c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87f230),
	.w1(32'hbc813251),
	.w2(32'hbcd6682d),
	.w3(32'h3a99c3bf),
	.w4(32'h3b7be2fd),
	.w5(32'hbc4febda),
	.w6(32'hbc9428d6),
	.w7(32'hbbf8212f),
	.w8(32'h3adc2ea9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f9487),
	.w1(32'hbc88aae9),
	.w2(32'hbc319a7f),
	.w3(32'hbcb5c7db),
	.w4(32'hbc21971f),
	.w5(32'hbc127444),
	.w6(32'hbbe868bd),
	.w7(32'hbb4c4f8e),
	.w8(32'hbbca0cc3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc684a3b),
	.w1(32'hbbfb7920),
	.w2(32'h3b992842),
	.w3(32'hbc33d68c),
	.w4(32'hbc1fe366),
	.w5(32'h3ad781a6),
	.w6(32'hb8d208a5),
	.w7(32'h3b09df94),
	.w8(32'hba59bc2f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b2df1),
	.w1(32'h3bde0fc8),
	.w2(32'h3bcc8c42),
	.w3(32'h3b40977a),
	.w4(32'h3bb14de8),
	.w5(32'h3bbd64d0),
	.w6(32'h3c085391),
	.w7(32'h3bbe3548),
	.w8(32'h3ba43298),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf3ede),
	.w1(32'h3ba52afc),
	.w2(32'h3b8bca35),
	.w3(32'h3bd62583),
	.w4(32'h3ba1bc8e),
	.w5(32'h3bb72976),
	.w6(32'h3ba47846),
	.w7(32'h3b9752e1),
	.w8(32'h3b8f81e2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b3d07),
	.w1(32'h3a745c40),
	.w2(32'h3bfd42e1),
	.w3(32'h3b8727a7),
	.w4(32'h3ad7171b),
	.w5(32'h3b4d9854),
	.w6(32'h3bb26ef0),
	.w7(32'h3b2d0083),
	.w8(32'h3a6f466c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb13139),
	.w1(32'h3bdbe915),
	.w2(32'h3c24fc6e),
	.w3(32'hba339e4d),
	.w4(32'hbbc4ab96),
	.w5(32'h3c5d7e97),
	.w6(32'h3bee6ce0),
	.w7(32'h3c05e842),
	.w8(32'h3befbb9f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25c29c),
	.w1(32'hbc101d3a),
	.w2(32'hbc1fccd8),
	.w3(32'h3c60959e),
	.w4(32'hbb10b8f6),
	.w5(32'hbc682d0e),
	.w6(32'h3a84f4db),
	.w7(32'hbbb8e2df),
	.w8(32'h3b6ec972),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a271b),
	.w1(32'hbaba4f89),
	.w2(32'hbc5f8b0d),
	.w3(32'hbc2e756a),
	.w4(32'h3ac147cd),
	.w5(32'hbb4a5a19),
	.w6(32'hbbefb30b),
	.w7(32'hbbe0c32f),
	.w8(32'h3b2d3f7c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3b09f),
	.w1(32'h3bd6e2e3),
	.w2(32'hbbf738f4),
	.w3(32'hbc19d0f3),
	.w4(32'h3bd9605e),
	.w5(32'hba588ccb),
	.w6(32'hbbbbdf92),
	.w7(32'hbb8c540e),
	.w8(32'h3bb40e92),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09cd03),
	.w1(32'h3c20cf31),
	.w2(32'h3c92f932),
	.w3(32'hbc0c22c8),
	.w4(32'h3bdfda5c),
	.w5(32'h3c0cc37c),
	.w6(32'h3ad89507),
	.w7(32'h3c974dc1),
	.w8(32'h3c87d2e6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65eb17),
	.w1(32'hbc0f202f),
	.w2(32'hbc30e72c),
	.w3(32'h3c531cfe),
	.w4(32'hbb8a2af8),
	.w5(32'hbbed1541),
	.w6(32'hbba7e2e8),
	.w7(32'hbc05b9db),
	.w8(32'hbbe98281),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbacd6),
	.w1(32'hbb27c039),
	.w2(32'hbc3bead3),
	.w3(32'hbb9cb15a),
	.w4(32'hbb821ab5),
	.w5(32'hbac0bfec),
	.w6(32'hbc229ab4),
	.w7(32'hbc110af9),
	.w8(32'hbb554278),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc544797),
	.w1(32'h3b8fd0d8),
	.w2(32'h3aeec776),
	.w3(32'h37d6a21c),
	.w4(32'h3c2a05f1),
	.w5(32'h3bdafa8e),
	.w6(32'hbadca8a9),
	.w7(32'h3bd4fdfb),
	.w8(32'h3bb9eb94),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58fdd6),
	.w1(32'hbb30b5fa),
	.w2(32'hbbd293dd),
	.w3(32'h38a58cf6),
	.w4(32'h3bcb7533),
	.w5(32'hbbd1b98a),
	.w6(32'hba47e983),
	.w7(32'hbabbbf56),
	.w8(32'h3a50e53f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5c9f7),
	.w1(32'h3c833afc),
	.w2(32'h3ccd0347),
	.w3(32'hbc0b9422),
	.w4(32'hbaf077ba),
	.w5(32'h3c8bfbb2),
	.w6(32'h3c04c6cd),
	.w7(32'h3c5b0306),
	.w8(32'hbc3ff35a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2267c1),
	.w1(32'hbbe62486),
	.w2(32'hbbdd2be2),
	.w3(32'hbbc90faa),
	.w4(32'h39a69a53),
	.w5(32'hbc03a2c0),
	.w6(32'hba00520f),
	.w7(32'hbac0717c),
	.w8(32'h3bd1db53),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ba54c),
	.w1(32'hbc0b6ec4),
	.w2(32'hbc271738),
	.w3(32'hbb884d3e),
	.w4(32'hbba36760),
	.w5(32'hbc2384c0),
	.w6(32'hbbb7d9cd),
	.w7(32'hbc023eda),
	.w8(32'h3b2bffbf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48ad65),
	.w1(32'h3c30ab5c),
	.w2(32'h3c20ab3d),
	.w3(32'hb9e9d5c4),
	.w4(32'h3b3969fb),
	.w5(32'h3bc7e895),
	.w6(32'h3ba970a0),
	.w7(32'h3bd530b8),
	.w8(32'hbb3a4209),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4d542),
	.w1(32'hbbbc246f),
	.w2(32'h3b15703c),
	.w3(32'h3bb4d439),
	.w4(32'h3b6d2e9e),
	.w5(32'hbc034219),
	.w6(32'hbc0ca474),
	.w7(32'hb92f179d),
	.w8(32'hbb4a20ce),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc239f83),
	.w1(32'hbba56401),
	.w2(32'hbc36429f),
	.w3(32'hbb965374),
	.w4(32'h3b5e8e38),
	.w5(32'hba0511c0),
	.w6(32'hbc128f3f),
	.w7(32'hbb7d6cba),
	.w8(32'hbbd41c38),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1956a4),
	.w1(32'hbc92756b),
	.w2(32'hbc84b2e2),
	.w3(32'hbbe1159a),
	.w4(32'hbbbcabf9),
	.w5(32'hbbeb91cc),
	.w6(32'hbc66e7fc),
	.w7(32'h3b53555d),
	.w8(32'hbb0a18f7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4e2f1),
	.w1(32'h3c68a6af),
	.w2(32'h3c5ccc99),
	.w3(32'hbc47b637),
	.w4(32'h3b395cd0),
	.w5(32'h3a158aed),
	.w6(32'h3c589400),
	.w7(32'hbb5890b0),
	.w8(32'hbc2e083c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc440614),
	.w1(32'hbbe9be2a),
	.w2(32'hbbc28905),
	.w3(32'hbaede689),
	.w4(32'hbbbdfc1e),
	.w5(32'hbbf06a48),
	.w6(32'hbc58b624),
	.w7(32'hbc031d3c),
	.w8(32'hbbabade7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe50f38),
	.w1(32'hbb6ba1c0),
	.w2(32'h3c5e4152),
	.w3(32'hbbd3ec74),
	.w4(32'hbbc4b003),
	.w5(32'h3bf04891),
	.w6(32'hbc5d2d6f),
	.w7(32'hbc1f1bf4),
	.w8(32'hbc6e1aac),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb038d6b),
	.w1(32'hbbc729fc),
	.w2(32'hbbe2e38f),
	.w3(32'hbb5ade44),
	.w4(32'hbc41ff6b),
	.w5(32'hbbf290e0),
	.w6(32'hbc02c34d),
	.w7(32'hbad09c26),
	.w8(32'h3b5755ac),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf558d9),
	.w1(32'h3c4c3132),
	.w2(32'h3c4cc7f0),
	.w3(32'h3aecb1ce),
	.w4(32'h3bb8b66f),
	.w5(32'h3c3c4922),
	.w6(32'h3c0c36d6),
	.w7(32'h3bdac68b),
	.w8(32'h3b93098f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e56ed),
	.w1(32'hbc856e31),
	.w2(32'hbca1735c),
	.w3(32'h3c1ae4e1),
	.w4(32'hbb9da7bf),
	.w5(32'hbc33472a),
	.w6(32'hbc5c84bd),
	.w7(32'hbc249fd3),
	.w8(32'hbb53cbf2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc282ab9),
	.w1(32'h3c0bcc14),
	.w2(32'h3c0266ec),
	.w3(32'hbc42b471),
	.w4(32'h3bd77d58),
	.w5(32'h3c2ae6dd),
	.w6(32'h3ba31010),
	.w7(32'h3a74d0af),
	.w8(32'h3acb02ef),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16eab6),
	.w1(32'h3bf26321),
	.w2(32'h3b332648),
	.w3(32'h3bf44ad1),
	.w4(32'h3b914396),
	.w5(32'h3b0c9a28),
	.w6(32'hbb68fd0e),
	.w7(32'hbb8679aa),
	.w8(32'hbbc92d16),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21acb1),
	.w1(32'hbc82a4d6),
	.w2(32'hbc97dc5a),
	.w3(32'hbac54ca7),
	.w4(32'hbbb0b009),
	.w5(32'hbbad7f8c),
	.w6(32'hbb616f64),
	.w7(32'hbc031046),
	.w8(32'hbbf5e136),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cde6a),
	.w1(32'h3bb41947),
	.w2(32'h3a6f8733),
	.w3(32'h3ac08f6a),
	.w4(32'h3b02ca4c),
	.w5(32'h3c053d3a),
	.w6(32'h3c2dede8),
	.w7(32'h3bdd7c2b),
	.w8(32'h3bb1403d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91a721),
	.w1(32'h3b6e28ec),
	.w2(32'hbb072e54),
	.w3(32'h3b8ed739),
	.w4(32'h3be0f78f),
	.w5(32'h3b269e95),
	.w6(32'h3b4c6e24),
	.w7(32'hb9ab2cf2),
	.w8(32'hbb982b7e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcea2ed),
	.w1(32'hbb3323ec),
	.w2(32'hbc140821),
	.w3(32'hba5f1ec3),
	.w4(32'hbb385e47),
	.w5(32'hbb82aabd),
	.w6(32'hbb984077),
	.w7(32'hbc356825),
	.w8(32'hbc2c78ec),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1181dc),
	.w1(32'hbc79a309),
	.w2(32'hbcf83fe4),
	.w3(32'hbba30a02),
	.w4(32'hbbc3e458),
	.w5(32'hbcd7c9bd),
	.w6(32'hbbeaf9a5),
	.w7(32'hbc218a3b),
	.w8(32'h3bf16d47),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca51390),
	.w1(32'hbb86c9fa),
	.w2(32'hbba36771),
	.w3(32'hbcd2911c),
	.w4(32'hba2ff455),
	.w5(32'hbb8dba59),
	.w6(32'hba945d2a),
	.w7(32'hbb93696e),
	.w8(32'hba99c56f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdea49a),
	.w1(32'hba1e4ede),
	.w2(32'hbc878cef),
	.w3(32'hbbcbb9d4),
	.w4(32'h3b884f78),
	.w5(32'hbc5ed0c9),
	.w6(32'hbbf70601),
	.w7(32'hbc80f3f4),
	.w8(32'hbbe40372),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ee14f),
	.w1(32'hbb7ec27a),
	.w2(32'hbc887287),
	.w3(32'hbc6737ca),
	.w4(32'hbc1e0c20),
	.w5(32'hbcaeb255),
	.w6(32'hbc1e8ed8),
	.w7(32'hbc25043b),
	.w8(32'hbbea0540),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b01b4),
	.w1(32'hb8c0b84b),
	.w2(32'hbc45cd19),
	.w3(32'hbbd1f545),
	.w4(32'hbae987d9),
	.w5(32'hbc5bdf23),
	.w6(32'hbb04363d),
	.w7(32'hbbf08aa9),
	.w8(32'hbaadf0b8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e511b),
	.w1(32'h3c4693d3),
	.w2(32'hbc4ae6e4),
	.w3(32'hbc189166),
	.w4(32'h3c07d448),
	.w5(32'h3a4432c3),
	.w6(32'hbb8a1c09),
	.w7(32'hbc3e0318),
	.w8(32'h3a4631cc),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5444e7),
	.w1(32'h3c8d56d0),
	.w2(32'h3c50aac3),
	.w3(32'hbc68a3f4),
	.w4(32'h3c45904b),
	.w5(32'h3c942d5f),
	.w6(32'h3c3511c2),
	.w7(32'hbabebfd8),
	.w8(32'hbb77ee93),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d7667),
	.w1(32'h3c1f6f5f),
	.w2(32'h3b5b282d),
	.w3(32'h3b66aa74),
	.w4(32'h3c619eaa),
	.w5(32'h3c481105),
	.w6(32'h3bad7cdf),
	.w7(32'h3bbb278f),
	.w8(32'h3c096d73),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba1139),
	.w1(32'hbaafb947),
	.w2(32'h3b9cf9f2),
	.w3(32'h3c120c32),
	.w4(32'h39991f4a),
	.w5(32'h3ace0246),
	.w6(32'h3b80adab),
	.w7(32'hbbd2c2bd),
	.w8(32'h37faad8c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02ddcf),
	.w1(32'hbc0a8c98),
	.w2(32'hbc3be24a),
	.w3(32'hbb2b5618),
	.w4(32'h3b794cfb),
	.w5(32'hbb19aa0c),
	.w6(32'hba914c48),
	.w7(32'hbba369ce),
	.w8(32'hbc1f8148),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc486f23),
	.w1(32'hbb12967b),
	.w2(32'hbba8455e),
	.w3(32'hbc8b42d0),
	.w4(32'hbba3355c),
	.w5(32'hbc137991),
	.w6(32'hbb795ee6),
	.w7(32'h3b3d8a29),
	.w8(32'h3b66d558),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8755fe),
	.w1(32'hbbfae7d2),
	.w2(32'hbc3cf6b9),
	.w3(32'hbb9616ee),
	.w4(32'h391a6567),
	.w5(32'hbbc9ca1c),
	.w6(32'hbb181460),
	.w7(32'hbb4389d7),
	.w8(32'hba924562),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc078ee3),
	.w1(32'hbb2300b5),
	.w2(32'hba134907),
	.w3(32'hbbb0bbf0),
	.w4(32'h3b6a646b),
	.w5(32'h3bc77c5e),
	.w6(32'h3949c805),
	.w7(32'h3b8471fd),
	.w8(32'hba00302d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf30fa7),
	.w1(32'hbc6e887e),
	.w2(32'hbc95b4e6),
	.w3(32'h3aa60dd2),
	.w4(32'hbbd74df4),
	.w5(32'hbc073056),
	.w6(32'hbc51dfb9),
	.w7(32'hbc054492),
	.w8(32'hbb2b0282),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02f17b),
	.w1(32'h3a2da711),
	.w2(32'h3c08d334),
	.w3(32'hbc276b6b),
	.w4(32'hbb83e903),
	.w5(32'h3ac23865),
	.w6(32'h3bda0cbf),
	.w7(32'h3bc06304),
	.w8(32'h3c08c722),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ae819),
	.w1(32'hba4aaad7),
	.w2(32'hb9be1d0f),
	.w3(32'h3bb79165),
	.w4(32'hbb2774c1),
	.w5(32'h3b37e599),
	.w6(32'hbabf8716),
	.w7(32'hbb3ae0d9),
	.w8(32'hbbde5d38),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba603ae),
	.w1(32'hbb55d970),
	.w2(32'hbbb98327),
	.w3(32'hba73e766),
	.w4(32'hbaabc6ff),
	.w5(32'hbaea1acb),
	.w6(32'hbaef0e04),
	.w7(32'hbab31b18),
	.w8(32'hbb0b53e2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39a514),
	.w1(32'h3bef5579),
	.w2(32'h3a976b98),
	.w3(32'hbc541c36),
	.w4(32'h3c05419a),
	.w5(32'h3b995e08),
	.w6(32'h3b9d21ef),
	.w7(32'h38a83597),
	.w8(32'hbb273724),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27b774),
	.w1(32'hba8bf172),
	.w2(32'h3c4603b7),
	.w3(32'h3b4004d0),
	.w4(32'hbab1bad4),
	.w5(32'h3b50ecef),
	.w6(32'h39708c60),
	.w7(32'h3b825ec0),
	.w8(32'h3bec42e6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88a5ed),
	.w1(32'h3b945589),
	.w2(32'h3c30a681),
	.w3(32'hbafc7676),
	.w4(32'hbb5595a4),
	.w5(32'h3bc3b1e9),
	.w6(32'hbb028a07),
	.w7(32'h3afe63d7),
	.w8(32'hbb2f5ba3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedf350),
	.w1(32'h3c6ef201),
	.w2(32'h3c94c418),
	.w3(32'h3c0eb2b3),
	.w4(32'h3c0fc0dd),
	.w5(32'h3c954688),
	.w6(32'h3c1c335e),
	.w7(32'h3c09020c),
	.w8(32'h3bc48fcb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2301a1),
	.w1(32'h3b8de85e),
	.w2(32'h3b764407),
	.w3(32'h3c43bc17),
	.w4(32'h3b5c7c3d),
	.w5(32'h3bcae560),
	.w6(32'h3b3ad856),
	.w7(32'h3ad7219c),
	.w8(32'hbae97fc5),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa14e59),
	.w1(32'h3b99072b),
	.w2(32'h3b9264a8),
	.w3(32'h39cc5e71),
	.w4(32'h3ab3ea09),
	.w5(32'h3b52b1a8),
	.w6(32'h3afa1850),
	.w7(32'hb8509a93),
	.w8(32'h3be83611),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb37539),
	.w1(32'hb9538217),
	.w2(32'h3b775bd6),
	.w3(32'h3b768f8c),
	.w4(32'hbad4db3d),
	.w5(32'h3a4394ea),
	.w6(32'h394881c0),
	.w7(32'h3b9b5522),
	.w8(32'hb9a34c29),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8e549),
	.w1(32'h3c67b395),
	.w2(32'h3c73d082),
	.w3(32'h399c14f4),
	.w4(32'h3c31c40b),
	.w5(32'h3c983d05),
	.w6(32'hbb14cb3e),
	.w7(32'hbb719598),
	.w8(32'hbc0c9163),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e5bff),
	.w1(32'h3b32d51e),
	.w2(32'h3a895f45),
	.w3(32'h3c7f2cf6),
	.w4(32'h3b9a9a3f),
	.w5(32'h3a8e9fcd),
	.w6(32'h39ff1cbc),
	.w7(32'hbafd84a9),
	.w8(32'hbace08ca),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f0f45),
	.w1(32'hb8d2321c),
	.w2(32'hbb91c63f),
	.w3(32'h3a4f1aab),
	.w4(32'hbafdf714),
	.w5(32'hb99e604e),
	.w6(32'h3ac4fe0e),
	.w7(32'h3a8c3b94),
	.w8(32'hbb2b8ce7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ad6eb),
	.w1(32'h3b8e5652),
	.w2(32'hbb9dd48c),
	.w3(32'hba7e3bec),
	.w4(32'h3b98f3ad),
	.w5(32'h3a5167a3),
	.w6(32'hbbe18717),
	.w7(32'hbbd9e4df),
	.w8(32'h3b1d2c4d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa0169),
	.w1(32'h3b92178d),
	.w2(32'hbaeae8f6),
	.w3(32'hbc1ae082),
	.w4(32'h3ba684b0),
	.w5(32'h3b53b376),
	.w6(32'h3be26a56),
	.w7(32'hbad05305),
	.w8(32'hbba7fd80),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba87f07),
	.w1(32'hbb65e37f),
	.w2(32'h3bb3e59e),
	.w3(32'h39ee9e39),
	.w4(32'hbbbc0b18),
	.w5(32'hb94e0f1e),
	.w6(32'hbb98fdfa),
	.w7(32'h3b689e64),
	.w8(32'hbbe81bdc),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0e5d0),
	.w1(32'hbc40ba95),
	.w2(32'hbc56adcf),
	.w3(32'h3b63111d),
	.w4(32'hbbd4766d),
	.w5(32'hbc1d028d),
	.w6(32'hbc83d509),
	.w7(32'hbc53fc2f),
	.w8(32'hba8a3573),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fa938),
	.w1(32'h3c277e7d),
	.w2(32'h3bf2f5c3),
	.w3(32'hbbdb5a4e),
	.w4(32'h3b79bc54),
	.w5(32'h3b630489),
	.w6(32'h3b7d3ade),
	.w7(32'h3a6406d2),
	.w8(32'hb9d1acdf),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5152be),
	.w1(32'h3ae557b0),
	.w2(32'h3b1972cc),
	.w3(32'h3bea274c),
	.w4(32'h38c6eba9),
	.w5(32'h387e1a06),
	.w6(32'hb9910f61),
	.w7(32'hb8e120de),
	.w8(32'hb853cb82),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2347a3),
	.w1(32'h3b77485c),
	.w2(32'h39e18f28),
	.w3(32'h382037bd),
	.w4(32'h3aecd47e),
	.w5(32'hbb0a9151),
	.w6(32'h3bc7e8e7),
	.w7(32'h3bdd1784),
	.w8(32'h3bd46d81),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule