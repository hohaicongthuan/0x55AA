module layer_10_featuremap_195(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e0b05),
	.w1(32'h3ac387a3),
	.w2(32'hbbd30168),
	.w3(32'h3ab9df78),
	.w4(32'h3a86e6ab),
	.w5(32'h3bf75b12),
	.w6(32'h3a8f8714),
	.w7(32'h3b94444d),
	.w8(32'h3b666a30),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e91ff),
	.w1(32'hbac942c4),
	.w2(32'h39592b84),
	.w3(32'h3b28d322),
	.w4(32'h3a9caa0b),
	.w5(32'hb9d2a825),
	.w6(32'hbb05a886),
	.w7(32'hbb6a31f5),
	.w8(32'hba4b193f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3a8a4),
	.w1(32'hbb62a397),
	.w2(32'hbb36e2bb),
	.w3(32'hbb2dc11a),
	.w4(32'hbb529d01),
	.w5(32'hbb7f6a46),
	.w6(32'hbb16578b),
	.w7(32'hbb511162),
	.w8(32'h3943e7f1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ad14c),
	.w1(32'hbc2535fe),
	.w2(32'hbae74c22),
	.w3(32'hbb473e84),
	.w4(32'hba56040c),
	.w5(32'hb9e6b48e),
	.w6(32'hbacc2098),
	.w7(32'hbba4d25b),
	.w8(32'hbb22f9ef),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94693b),
	.w1(32'h3bcf2057),
	.w2(32'hbc03fffd),
	.w3(32'hba8e8650),
	.w4(32'h3b0e83f5),
	.w5(32'hb9ce5e58),
	.w6(32'h3b7746e4),
	.w7(32'hbb79a2c9),
	.w8(32'hbb7f6fd8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba840ac7),
	.w1(32'h3b70e22f),
	.w2(32'hbbae0f2c),
	.w3(32'hbab9e79e),
	.w4(32'h38fa700c),
	.w5(32'hbbe8fdbd),
	.w6(32'h3bc114c6),
	.w7(32'h3bf536d3),
	.w8(32'h3b705489),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e29c1),
	.w1(32'hbb1a128d),
	.w2(32'h37078ef4),
	.w3(32'hbbb98aa4),
	.w4(32'hb8cf45c6),
	.w5(32'h3a3e12e9),
	.w6(32'hbb3e6224),
	.w7(32'hbb636884),
	.w8(32'h3a257223),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc3734),
	.w1(32'h3ac9ceed),
	.w2(32'hbbe5e28b),
	.w3(32'hbc0398a8),
	.w4(32'hbb01a0b6),
	.w5(32'hbbbc8be7),
	.w6(32'h3b9ed5b0),
	.w7(32'h3c0969b6),
	.w8(32'h3bfd56bb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd827d5),
	.w1(32'hba499529),
	.w2(32'hbb9f6ffc),
	.w3(32'hbada9a8d),
	.w4(32'hb98bda0d),
	.w5(32'hbb9abc10),
	.w6(32'hba8f1207),
	.w7(32'h3b37a049),
	.w8(32'h3ae476a3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb360964),
	.w1(32'hbc27b0da),
	.w2(32'h3b069d65),
	.w3(32'hbae1c414),
	.w4(32'hbb41f370),
	.w5(32'h3c021c6b),
	.w6(32'hbbe0f28e),
	.w7(32'hbc134270),
	.w8(32'h38879f24),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcbf9b),
	.w1(32'hbb65a32e),
	.w2(32'h3b80a087),
	.w3(32'h3b4e53a4),
	.w4(32'hbb8e706a),
	.w5(32'hbbb0fe48),
	.w6(32'hbb82a0db),
	.w7(32'hbbd62d80),
	.w8(32'hbac45e13),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27c5c3),
	.w1(32'hbb2138ed),
	.w2(32'h3b1dd524),
	.w3(32'hbb1436a3),
	.w4(32'hbb4cb1a9),
	.w5(32'hba64983a),
	.w6(32'h3a9af2d5),
	.w7(32'h3b04f8fc),
	.w8(32'hbace722d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44f9ea),
	.w1(32'hb998a1e7),
	.w2(32'h3912fa12),
	.w3(32'hbb5c5014),
	.w4(32'h3abb7e24),
	.w5(32'h3aad0212),
	.w6(32'h3b065011),
	.w7(32'h3b0b4f1f),
	.w8(32'h3bddda86),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadefb7f),
	.w1(32'h3bdc948d),
	.w2(32'hbb83f47e),
	.w3(32'hb913c419),
	.w4(32'h39c3b2e4),
	.w5(32'hbc0d4c52),
	.w6(32'h3c047fb3),
	.w7(32'h3c106aad),
	.w8(32'h3afd0890),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc018202),
	.w1(32'hb9e89eb6),
	.w2(32'h3a8db38c),
	.w3(32'hbb4dbca7),
	.w4(32'hba5bb5dd),
	.w5(32'hbbbae8bd),
	.w6(32'hbacc2696),
	.w7(32'hb9ac128b),
	.w8(32'hbb516cf8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badfe46),
	.w1(32'h3b2df199),
	.w2(32'hbb2e4001),
	.w3(32'hbaf63f3f),
	.w4(32'h3a898ccf),
	.w5(32'hb8f4c7e0),
	.w6(32'h3bc587ea),
	.w7(32'h3be830d8),
	.w8(32'h3beffc0e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4a2d4),
	.w1(32'h3b25dc4a),
	.w2(32'h3b8c5009),
	.w3(32'h3b0a584b),
	.w4(32'h391d22f7),
	.w5(32'hbb8256ed),
	.w6(32'hba068012),
	.w7(32'h3b8673da),
	.w8(32'hbb83aaed),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13f4be),
	.w1(32'hbbe809a0),
	.w2(32'h3ace298b),
	.w3(32'hbbfb19db),
	.w4(32'h3a8293b0),
	.w5(32'h3bd3292e),
	.w6(32'hbb96a22d),
	.w7(32'hbb991847),
	.w8(32'h3b6fa606),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ba07b),
	.w1(32'hbb34bcfa),
	.w2(32'hba605dcb),
	.w3(32'hb93c0f20),
	.w4(32'hba87c927),
	.w5(32'h3ae4d395),
	.w6(32'hba50a0c7),
	.w7(32'h39ae383b),
	.w8(32'h3b095b5c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b26118),
	.w1(32'h38ce410e),
	.w2(32'hbb9cd377),
	.w3(32'hba212107),
	.w4(32'hb94b5aa5),
	.w5(32'hbb86222b),
	.w6(32'hba1234a7),
	.w7(32'h3b009b8d),
	.w8(32'h35ccbfc6),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ef082),
	.w1(32'hbb68fcbd),
	.w2(32'hbc217210),
	.w3(32'hb9e9a43d),
	.w4(32'h3a71df98),
	.w5(32'hbb2c73a7),
	.w6(32'hbba5face),
	.w7(32'hba03f81d),
	.w8(32'hb9d306ba),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9e879),
	.w1(32'hbbc81cdb),
	.w2(32'h3bd717d6),
	.w3(32'h3a91ac10),
	.w4(32'hbbcfe83d),
	.w5(32'hbc755ba0),
	.w6(32'hbb42c49a),
	.w7(32'hbc1385eb),
	.w8(32'hbba114b7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb63e31),
	.w1(32'hbb81b0c9),
	.w2(32'hba9c01bb),
	.w3(32'hbc33763d),
	.w4(32'hb9867159),
	.w5(32'h3aacf913),
	.w6(32'h3b30d9d6),
	.w7(32'hba03f825),
	.w8(32'hb6efc1fc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d0ed0),
	.w1(32'h3b8b8d16),
	.w2(32'hbb6d4c89),
	.w3(32'h39829bd0),
	.w4(32'h3b73671e),
	.w5(32'hbb515da2),
	.w6(32'h3bd49c03),
	.w7(32'h3c0927f3),
	.w8(32'h3ba7bf21),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82c15b),
	.w1(32'hbb2103cd),
	.w2(32'hbb146b3d),
	.w3(32'h3a0b5a7c),
	.w4(32'hba38d6c8),
	.w5(32'hbb3d06be),
	.w6(32'hbb45c2d2),
	.w7(32'hbb98110d),
	.w8(32'hba384115),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cf95e),
	.w1(32'hbc24e45a),
	.w2(32'hbc3eb99c),
	.w3(32'h397b423a),
	.w4(32'hbc3c0bef),
	.w5(32'hbc3d2c5e),
	.w6(32'hbb35a0b9),
	.w7(32'hbabe1aef),
	.w8(32'hbadf2598),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46807c),
	.w1(32'hbaf55953),
	.w2(32'hbbc2665b),
	.w3(32'hbb924d81),
	.w4(32'hbaac43ad),
	.w5(32'hbb986097),
	.w6(32'hba6229ac),
	.w7(32'h3b0ad673),
	.w8(32'h39cfef27),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba159b),
	.w1(32'hbb71bec1),
	.w2(32'h3b9e2806),
	.w3(32'hbb5048d9),
	.w4(32'h3b8ba49b),
	.w5(32'h3c0255c7),
	.w6(32'hbb99c442),
	.w7(32'hbb99fe97),
	.w8(32'h3b0f7f53),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03a32a),
	.w1(32'hbb867a15),
	.w2(32'hba757772),
	.w3(32'h3b8b5e09),
	.w4(32'hbb5ee10b),
	.w5(32'hbafa0995),
	.w6(32'hbba681ed),
	.w7(32'hba7b0ffc),
	.w8(32'h3b062adc),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968499b),
	.w1(32'h3ad91297),
	.w2(32'h3b8f944c),
	.w3(32'h3b1ada36),
	.w4(32'h3a9f75cc),
	.w5(32'hba9fccc4),
	.w6(32'h3b591162),
	.w7(32'h3b82e474),
	.w8(32'h39f852c6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31db80),
	.w1(32'hbb28d4ae),
	.w2(32'hbbd3ed2d),
	.w3(32'hbbbd5528),
	.w4(32'h38b0f644),
	.w5(32'hbacbbf8e),
	.w6(32'hbba494fd),
	.w7(32'hbb2ed507),
	.w8(32'hb8cc8356),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5696dc),
	.w1(32'hbaf9c29a),
	.w2(32'hbbd391a1),
	.w3(32'h3aebb75f),
	.w4(32'hb9c60f55),
	.w5(32'hbb0f2605),
	.w6(32'hbb061f58),
	.w7(32'h3a103827),
	.w8(32'h3a37f63d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fe415),
	.w1(32'hbb7862be),
	.w2(32'hbc10bf8d),
	.w3(32'h3a1bd21f),
	.w4(32'hbb2990ad),
	.w5(32'hbbf9c96d),
	.w6(32'hbb69edf8),
	.w7(32'hbb897df0),
	.w8(32'hbbe81cb6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ff177),
	.w1(32'h3bbe6ba0),
	.w2(32'h3b36438c),
	.w3(32'hbba5e961),
	.w4(32'h3b94e43e),
	.w5(32'h3b21cf1f),
	.w6(32'h3b39cdca),
	.w7(32'h3befb441),
	.w8(32'h3a65dba6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fdd8b),
	.w1(32'hbc083a31),
	.w2(32'h3ad13520),
	.w3(32'hbba68bcf),
	.w4(32'h3a17515d),
	.w5(32'h3c0f44d6),
	.w6(32'hbc0a28f6),
	.w7(32'hbbce558f),
	.w8(32'hb9dbe769),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b866c11),
	.w1(32'hbba17353),
	.w2(32'hbc0b582e),
	.w3(32'h3b698f08),
	.w4(32'hba49ce6a),
	.w5(32'hbafe992a),
	.w6(32'hbb06ceea),
	.w7(32'hbab0d8c2),
	.w8(32'h3b064f58),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafe656),
	.w1(32'hbbb34ad5),
	.w2(32'h3b58a999),
	.w3(32'hba833292),
	.w4(32'hb9a56c73),
	.w5(32'h3bff6b82),
	.w6(32'hba99eced),
	.w7(32'hbbb650b0),
	.w8(32'hbaa1e7f4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4de57),
	.w1(32'hb9f816fb),
	.w2(32'hba82a977),
	.w3(32'h3a704c5f),
	.w4(32'hba449def),
	.w5(32'hbb639b73),
	.w6(32'hbb2f2ee4),
	.w7(32'hbb04885f),
	.w8(32'hbb042bea),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bdbbd),
	.w1(32'h3b891e7b),
	.w2(32'hbb7c74ee),
	.w3(32'hbb814564),
	.w4(32'h3b9b1976),
	.w5(32'hbb7b9350),
	.w6(32'h3a1299a6),
	.w7(32'h3b8d2d76),
	.w8(32'h3b19f0dc),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42b477),
	.w1(32'hbabead0b),
	.w2(32'hb98f3a6f),
	.w3(32'h3aa80627),
	.w4(32'hba4de20b),
	.w5(32'h3a1cbff9),
	.w6(32'hbb0059e7),
	.w7(32'hbb204508),
	.w8(32'hbabaeea2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a964ad6),
	.w1(32'h3b6a7bad),
	.w2(32'h3b98c0c0),
	.w3(32'hbaa667e3),
	.w4(32'h3b47a445),
	.w5(32'h3b45d94b),
	.w6(32'h3b770f52),
	.w7(32'h3bab84de),
	.w8(32'h3a8ed5ab),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39401221),
	.w1(32'hb83b349a),
	.w2(32'h3a9d7b9b),
	.w3(32'hbac25d45),
	.w4(32'h3aac0202),
	.w5(32'hb940a297),
	.w6(32'hbb16b523),
	.w7(32'hbb73081a),
	.w8(32'hbafb4e89),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba430e84),
	.w1(32'h3acf34d4),
	.w2(32'hbb88daff),
	.w3(32'hbaf9137e),
	.w4(32'hb88b7cbd),
	.w5(32'hbb377a26),
	.w6(32'hbaa75ae8),
	.w7(32'h3b2a22b1),
	.w8(32'h3aa00df8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbedc88),
	.w1(32'hbb605eee),
	.w2(32'h3c206029),
	.w3(32'h3838dee0),
	.w4(32'h3baecf8d),
	.w5(32'h3c2e4d91),
	.w6(32'h39f85f82),
	.w7(32'hbb3e1d30),
	.w8(32'h3be73621),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6f18e),
	.w1(32'hbb9f2b5a),
	.w2(32'h39381125),
	.w3(32'hb90eec36),
	.w4(32'h3a063780),
	.w5(32'h3b90f9d3),
	.w6(32'hbbea6652),
	.w7(32'hbc0995fa),
	.w8(32'hbb870296),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bc137),
	.w1(32'hbb02bf95),
	.w2(32'h3bd6b923),
	.w3(32'h3b5c5e2c),
	.w4(32'h3b211b36),
	.w5(32'h3c058f3d),
	.w6(32'hb934e325),
	.w7(32'hb8a030df),
	.w8(32'h3bfa439d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfce2d2),
	.w1(32'hbb3a419e),
	.w2(32'h3c2084ed),
	.w3(32'h3bad3b19),
	.w4(32'h3a532ffe),
	.w5(32'h3af443fa),
	.w6(32'hbb9e23ce),
	.w7(32'hbc00966d),
	.w8(32'hbb98c30e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c168df8),
	.w1(32'hbb62b4bd),
	.w2(32'hba7bd4e5),
	.w3(32'hbb708688),
	.w4(32'hbb79af65),
	.w5(32'h39999668),
	.w6(32'hbadaae6c),
	.w7(32'h3b4b5520),
	.w8(32'h3bad9281),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53a2b1),
	.w1(32'h389c7bad),
	.w2(32'hbbc83032),
	.w3(32'hbb10c95b),
	.w4(32'hba55de40),
	.w5(32'hbb9bef45),
	.w6(32'hbab850b3),
	.w7(32'h3b0f741c),
	.w8(32'hb9d421a7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a18ab),
	.w1(32'h3ba949f8),
	.w2(32'hbb440f15),
	.w3(32'h392dae74),
	.w4(32'h3b50dfea),
	.w5(32'hbb8b4648),
	.w6(32'h3bb7b4e7),
	.w7(32'h3bcfbb07),
	.w8(32'h3b336d5c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d57df),
	.w1(32'hbbb8daaf),
	.w2(32'hba9a7ef7),
	.w3(32'hba7e2eea),
	.w4(32'hbb8b582a),
	.w5(32'h3aa35e39),
	.w6(32'hbbdfa27b),
	.w7(32'hbbdd3bc0),
	.w8(32'hba92210a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c8743),
	.w1(32'hbb2e3ac0),
	.w2(32'h3bdb2275),
	.w3(32'h3b0326ef),
	.w4(32'h38d99138),
	.w5(32'h3b1d8e1f),
	.w6(32'hbb76a55b),
	.w7(32'hbc0f0226),
	.w8(32'hbb4c8765),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc8c68),
	.w1(32'h387b24e6),
	.w2(32'hbbbf4004),
	.w3(32'hb950c8ac),
	.w4(32'hb8427766),
	.w5(32'hbb3424e4),
	.w6(32'h3a14485e),
	.w7(32'h3b3375e2),
	.w8(32'h3b8053d0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc40264),
	.w1(32'hbaef0c88),
	.w2(32'hbaaf2ff8),
	.w3(32'hbb94ba52),
	.w4(32'hbb1322f8),
	.w5(32'h3b9a956a),
	.w6(32'h3a8043c3),
	.w7(32'hba6ca6d9),
	.w8(32'hba84e3c8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961c112),
	.w1(32'h3ae90746),
	.w2(32'h3b1ac81a),
	.w3(32'h3b4cfb32),
	.w4(32'h3b43e001),
	.w5(32'h3b339f3b),
	.w6(32'h3aae31a0),
	.w7(32'h3ae1379a),
	.w8(32'h3b1a6e48),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51fab1),
	.w1(32'hba79f12f),
	.w2(32'hbb804a1c),
	.w3(32'h3a9d2e2d),
	.w4(32'h3b0940b0),
	.w5(32'hbad15ab4),
	.w6(32'h3b3e3ff8),
	.w7(32'hbabb683d),
	.w8(32'hba3b58bf),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab908f1),
	.w1(32'h3a9e11aa),
	.w2(32'h3ba78032),
	.w3(32'hba207897),
	.w4(32'h3b201ecc),
	.w5(32'h3b772b22),
	.w6(32'h3acfd6cf),
	.w7(32'h3b540274),
	.w8(32'h3b3fd94a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b5ffd),
	.w1(32'hbb29ffbc),
	.w2(32'hbb5d8eb7),
	.w3(32'hb98c5423),
	.w4(32'hbac95dca),
	.w5(32'h384846ca),
	.w6(32'hbb32832b),
	.w7(32'hbb6a2821),
	.w8(32'h3a3796c4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc058fad),
	.w1(32'hbab0a24e),
	.w2(32'h3a2726fe),
	.w3(32'hbb35505a),
	.w4(32'h3a36c116),
	.w5(32'hba92a545),
	.w6(32'hbb51f04d),
	.w7(32'hbb5ca40d),
	.w8(32'h39ac69cd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4296f9),
	.w1(32'h3b8f64c5),
	.w2(32'hbb6f3c93),
	.w3(32'hbbb71121),
	.w4(32'h3b4dd0c1),
	.w5(32'hbb69991b),
	.w6(32'h3b876a5e),
	.w7(32'h3bd9c856),
	.w8(32'h3b699b59),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3bdd6),
	.w1(32'hbb553f3b),
	.w2(32'hba0f4a00),
	.w3(32'hba95d6f6),
	.w4(32'hba500aa4),
	.w5(32'h3b151065),
	.w6(32'hba9632d2),
	.w7(32'hbb24333d),
	.w8(32'h3b2ca692),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b696cdb),
	.w1(32'h3a0b498f),
	.w2(32'hbb8f8138),
	.w3(32'hb9c539f3),
	.w4(32'h3a4fcbc7),
	.w5(32'hbb83a355),
	.w6(32'h3a82dfe3),
	.w7(32'h3b541cb5),
	.w8(32'h3b179b8d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d50af),
	.w1(32'h3b7cd920),
	.w2(32'hbc0c9057),
	.w3(32'hbab237ad),
	.w4(32'h3b11e968),
	.w5(32'hbb8a87f2),
	.w6(32'hb9038ad2),
	.w7(32'hbbcdf06e),
	.w8(32'hbc304411),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc637af),
	.w1(32'hbb2f3c0d),
	.w2(32'h3ba2bcae),
	.w3(32'hbb42b401),
	.w4(32'h3b0796ea),
	.w5(32'h3bbd5308),
	.w6(32'hbadaecf6),
	.w7(32'hbb99c5b8),
	.w8(32'h3a410b51),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb502ea),
	.w1(32'hbb54ec4a),
	.w2(32'hbb0581ce),
	.w3(32'hb87249d0),
	.w4(32'hb9e3751d),
	.w5(32'hba350eec),
	.w6(32'hbb50eaf4),
	.w7(32'hbb5ed315),
	.w8(32'h396e8255),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eb49a),
	.w1(32'hbb0be021),
	.w2(32'h3be4de16),
	.w3(32'h3b3f44a8),
	.w4(32'h3b09da42),
	.w5(32'h3b31ac66),
	.w6(32'hbba341cd),
	.w7(32'hbb33d94b),
	.w8(32'h3b7e2078),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d3ebe),
	.w1(32'h3b3e44af),
	.w2(32'h3bbbdff9),
	.w3(32'hbc375977),
	.w4(32'h39be36d2),
	.w5(32'h3b14a26d),
	.w6(32'h3b6f0459),
	.w7(32'h3ba2a99b),
	.w8(32'h3b4cd785),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f081e),
	.w1(32'hbac6acbb),
	.w2(32'hba0b4b5b),
	.w3(32'hbb7689bb),
	.w4(32'h3b1d9e3f),
	.w5(32'h3b15c8c4),
	.w6(32'h3a809f7d),
	.w7(32'hb9de610e),
	.w8(32'h3b9682bf),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47017a),
	.w1(32'h3b1a919b),
	.w2(32'hbb0a04ee),
	.w3(32'h3a99587b),
	.w4(32'h3b237779),
	.w5(32'hbab2f216),
	.w6(32'h3b4fb66a),
	.w7(32'h3beb6734),
	.w8(32'h3bcc822e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaefbe),
	.w1(32'hbbcbc688),
	.w2(32'h3a1bb444),
	.w3(32'h3b05d900),
	.w4(32'h39d3bf50),
	.w5(32'h3c14dab3),
	.w6(32'hbc0d06c9),
	.w7(32'hbc41164a),
	.w8(32'h395524b9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c207e8b),
	.w1(32'hbb3532a4),
	.w2(32'h3b144cd6),
	.w3(32'h3c1eb95d),
	.w4(32'h3a90fd99),
	.w5(32'h3a9780de),
	.w6(32'hbb44f677),
	.w7(32'hbb21e179),
	.w8(32'h3a42d66c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae05a52),
	.w1(32'h3a019620),
	.w2(32'hbb9f8eec),
	.w3(32'hbad0afe7),
	.w4(32'h3b23e97e),
	.w5(32'hbb51f5ae),
	.w6(32'h39f7d6a3),
	.w7(32'h3b352a13),
	.w8(32'h3afb46f5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dcdbf),
	.w1(32'h3b8ab281),
	.w2(32'hbb51cf3c),
	.w3(32'hba3a8fa4),
	.w4(32'h3b70226d),
	.w5(32'hbb2da47a),
	.w6(32'h3b7023f6),
	.w7(32'h3bb3c839),
	.w8(32'h3b5d0865),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb882068),
	.w1(32'hbb480abe),
	.w2(32'hbc1c6362),
	.w3(32'hb9f039bf),
	.w4(32'hb88dd1bb),
	.w5(32'hbb1b067e),
	.w6(32'hbb52aa7e),
	.w7(32'h3a37472f),
	.w8(32'h3a421e91),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc90f9b),
	.w1(32'hbaa052c5),
	.w2(32'h3b1eb269),
	.w3(32'h3b1914af),
	.w4(32'h3aa6e818),
	.w5(32'h3ace9fb9),
	.w6(32'hbb4a0f77),
	.w7(32'hbb203972),
	.w8(32'h3b038b39),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b2567),
	.w1(32'hbc218f8d),
	.w2(32'h3bedfbca),
	.w3(32'hbb27fd32),
	.w4(32'hbc010713),
	.w5(32'hbbff231d),
	.w6(32'hbba73c3e),
	.w7(32'hbc0410a7),
	.w8(32'hbbfc5ba6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac93904),
	.w1(32'h3b030d68),
	.w2(32'hbbd4a257),
	.w3(32'hbba59032),
	.w4(32'hba82c544),
	.w5(32'hbba533d3),
	.w6(32'h3bffd6df),
	.w7(32'h3bf98bc9),
	.w8(32'h3bc76411),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bb166),
	.w1(32'hbb0697a3),
	.w2(32'hbb2e51d0),
	.w3(32'h3ae0ebdd),
	.w4(32'h39b5c96d),
	.w5(32'hba8a0d34),
	.w6(32'hbaf82972),
	.w7(32'hbb769bab),
	.w8(32'hbb884cfc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3fa31),
	.w1(32'hbb068a65),
	.w2(32'h3b4c69a9),
	.w3(32'hbb972e1b),
	.w4(32'hbb1c222b),
	.w5(32'h3a848e9d),
	.w6(32'h3a1cde8d),
	.w7(32'h3b072ea6),
	.w8(32'h3a1c4d13),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b0c77),
	.w1(32'hbb3d96a0),
	.w2(32'hbbf5e207),
	.w3(32'h3a889ceb),
	.w4(32'hb9fa6c62),
	.w5(32'hbafbce32),
	.w6(32'hbbecfa67),
	.w7(32'hbb769d95),
	.w8(32'h3997b4e6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ee7f1),
	.w1(32'h3ac3f2a9),
	.w2(32'hb8e8da21),
	.w3(32'h3b3a54e2),
	.w4(32'h3b6983b0),
	.w5(32'h3ac6687b),
	.w6(32'hba351d0e),
	.w7(32'h397e868b),
	.w8(32'h392037b1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea0144),
	.w1(32'hba4b423a),
	.w2(32'h3abad3fc),
	.w3(32'hbac0a459),
	.w4(32'h3ac7c1ef),
	.w5(32'h3b8051f3),
	.w6(32'hba2b7ae9),
	.w7(32'hb88deb3e),
	.w8(32'h3a968dd4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a41c6),
	.w1(32'hbaa8f03e),
	.w2(32'hbb07e5aa),
	.w3(32'hbab99ecb),
	.w4(32'hba9abad8),
	.w5(32'hbb66699d),
	.w6(32'hbb26ebea),
	.w7(32'hbb1c48fb),
	.w8(32'hbaecd502),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa20fb),
	.w1(32'hba7ae26f),
	.w2(32'hb7de9ee7),
	.w3(32'hbb82367f),
	.w4(32'h3aff12aa),
	.w5(32'h3b0a5682),
	.w6(32'hbb157df2),
	.w7(32'hbadc90f2),
	.w8(32'hb8bdf6ac),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a003fe2),
	.w1(32'h3baeac82),
	.w2(32'h3ba0f84a),
	.w3(32'hbad8198e),
	.w4(32'hbb3fa99f),
	.w5(32'hba182b5b),
	.w6(32'h3b7eeb70),
	.w7(32'h3c072c39),
	.w8(32'h3b6358ed),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a015b),
	.w1(32'h38d275c0),
	.w2(32'h393b6cc8),
	.w3(32'hbb0f9da2),
	.w4(32'hbaf3a1c5),
	.w5(32'hbb4b1847),
	.w6(32'hb9e24720),
	.w7(32'h39230072),
	.w8(32'hbb3714d0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb148e30),
	.w1(32'hbb458a47),
	.w2(32'h3a943bee),
	.w3(32'hbbbcccb3),
	.w4(32'hbb870cf1),
	.w5(32'hbb8f61c4),
	.w6(32'hbb4ba9f6),
	.w7(32'hbb4d5f75),
	.w8(32'hbbbe5e36),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb575cff),
	.w1(32'hbaa03cf1),
	.w2(32'hbbb2f782),
	.w3(32'hbb9c3085),
	.w4(32'h3a906f72),
	.w5(32'hba9b84ac),
	.w6(32'hbb5a90ca),
	.w7(32'h36bd1314),
	.w8(32'h3a186293),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a461b),
	.w1(32'h3b31df8b),
	.w2(32'h3b0ec9f9),
	.w3(32'h3b183b07),
	.w4(32'h3b58061a),
	.w5(32'h3b2d6a5c),
	.w6(32'h3b081239),
	.w7(32'h3b0926b2),
	.w8(32'h3b034d88),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa4fce),
	.w1(32'hbb59ab16),
	.w2(32'hbbdcbc82),
	.w3(32'hbb229d38),
	.w4(32'h38a73c7f),
	.w5(32'hbafaacb3),
	.w6(32'hbb3e726b),
	.w7(32'h3a1e1178),
	.w8(32'h3b6be7e3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dc104),
	.w1(32'hbb4f0918),
	.w2(32'hbbd68a9f),
	.w3(32'h3af58ad4),
	.w4(32'h3ac0cfd6),
	.w5(32'hbaafd93f),
	.w6(32'hbbba7bfd),
	.w7(32'hbb343591),
	.w8(32'hbb298537),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ef82),
	.w1(32'hbbc29b8b),
	.w2(32'h3b29cac9),
	.w3(32'hb95757f4),
	.w4(32'hbaf12c74),
	.w5(32'h3ba4f085),
	.w6(32'hbbb29da0),
	.w7(32'hbb94dfbb),
	.w8(32'hbb1c060e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2d9a6),
	.w1(32'hbb3499cd),
	.w2(32'h3abf475d),
	.w3(32'hbb488e5a),
	.w4(32'h3b637a65),
	.w5(32'h3b96abba),
	.w6(32'hbb83362a),
	.w7(32'hbb08f5d4),
	.w8(32'h3a792d3b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d5172),
	.w1(32'h3add32c3),
	.w2(32'h3a6556b4),
	.w3(32'h3abc935d),
	.w4(32'h3b60760e),
	.w5(32'h3b3837a7),
	.w6(32'h3a86f341),
	.w7(32'hb77e1bd9),
	.w8(32'h3aa5b887),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ee09f),
	.w1(32'hbb867bb2),
	.w2(32'hbb6f1d55),
	.w3(32'h3a8a0487),
	.w4(32'hbad6dcd2),
	.w5(32'h39c1e977),
	.w6(32'hba55a1bb),
	.w7(32'hbb4fec9f),
	.w8(32'h390537bc),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc0a80),
	.w1(32'hbb05f3f6),
	.w2(32'hbb58463a),
	.w3(32'hb801d1a6),
	.w4(32'hbb5b1971),
	.w5(32'hbbb3a531),
	.w6(32'hbb411a81),
	.w7(32'hbbb03444),
	.w8(32'hbb84bdae),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95a058),
	.w1(32'hb9be5203),
	.w2(32'hbab21a9b),
	.w3(32'h3b211962),
	.w4(32'h3b6cf67b),
	.w5(32'h3b193f88),
	.w6(32'h3a7530ef),
	.w7(32'h3975fe04),
	.w8(32'hba8b7229),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f9c1d),
	.w1(32'hbba29f29),
	.w2(32'hba99273e),
	.w3(32'hbafd011e),
	.w4(32'hbab0f6c2),
	.w5(32'h3b154a7f),
	.w6(32'hbb62471a),
	.w7(32'hbbbb8c2c),
	.w8(32'h3b82e074),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63617b),
	.w1(32'hba775ee3),
	.w2(32'h3b9b043c),
	.w3(32'hbba48b15),
	.w4(32'h3b347ed3),
	.w5(32'h3bf88377),
	.w6(32'hbb44cc61),
	.w7(32'hbb09b824),
	.w8(32'h3a417f52),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae209a9),
	.w1(32'hbc0a5cfa),
	.w2(32'hbaa6bf15),
	.w3(32'hbb66c265),
	.w4(32'hbb67e6f2),
	.w5(32'h3aa72e9a),
	.w6(32'hbbc825f1),
	.w7(32'hbb8baf84),
	.w8(32'hb9c15a8a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bea5e),
	.w1(32'hbb5f68c1),
	.w2(32'hbc53172b),
	.w3(32'h3a3274d0),
	.w4(32'hbc17d8f2),
	.w5(32'hbb57068e),
	.w6(32'hbc319b2e),
	.w7(32'hbc7330ab),
	.w8(32'hbc0f9c5f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb917cb5),
	.w1(32'h3be8f4ea),
	.w2(32'h3c5c50a6),
	.w3(32'h3a076f81),
	.w4(32'h3a548a11),
	.w5(32'h3bb478e8),
	.w6(32'h3aa02e7f),
	.w7(32'h39383057),
	.w8(32'hbb836f63),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92b192),
	.w1(32'h3bc1321a),
	.w2(32'hbb8ec27a),
	.w3(32'hba796bc2),
	.w4(32'h3b3a48b9),
	.w5(32'hbb769a16),
	.w6(32'h3c0e517b),
	.w7(32'h3c044c22),
	.w8(32'h3b9800f7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc105e75),
	.w1(32'hba8dd7aa),
	.w2(32'hbbcd0b5f),
	.w3(32'h39221928),
	.w4(32'h3abce916),
	.w5(32'hbbaa125f),
	.w6(32'h39ea84bf),
	.w7(32'h3a812c8d),
	.w8(32'h3b2c3470),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97c60c),
	.w1(32'hba945d7b),
	.w2(32'hbbc98b3b),
	.w3(32'hbbab74a7),
	.w4(32'hbb83385d),
	.w5(32'hbbc1fc2b),
	.w6(32'h3b847feb),
	.w7(32'h3b8e2c3a),
	.w8(32'h3b1aa76a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb868375),
	.w1(32'hbb0da44a),
	.w2(32'hbbbfe2c2),
	.w3(32'hba267eae),
	.w4(32'hbb275c15),
	.w5(32'hbb507a37),
	.w6(32'hbab79339),
	.w7(32'h3b06cae8),
	.w8(32'hba522c8d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3214b),
	.w1(32'hbb56bad1),
	.w2(32'hbb14fa4d),
	.w3(32'hb9b4c9df),
	.w4(32'hb9a21b9d),
	.w5(32'hbacfebbb),
	.w6(32'hbb0f81e8),
	.w7(32'hbb2bf2f8),
	.w8(32'hba8b8a3c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba853cdc),
	.w1(32'hbb48c456),
	.w2(32'hbc031534),
	.w3(32'hbaa0da6f),
	.w4(32'h3a7af523),
	.w5(32'hbab86404),
	.w6(32'hbba53041),
	.w7(32'hbb31cbd0),
	.w8(32'hbb4760ab),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce661e),
	.w1(32'h3b5612ac),
	.w2(32'hbb44ae36),
	.w3(32'h3ae86502),
	.w4(32'h3b073af1),
	.w5(32'hbb4be74a),
	.w6(32'h3bcc073f),
	.w7(32'h3bd8404f),
	.w8(32'h3b9d9e3e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f6731),
	.w1(32'hbb1676b1),
	.w2(32'hbb331914),
	.w3(32'h3a9a544c),
	.w4(32'h3a828684),
	.w5(32'hbb0245f7),
	.w6(32'hbb90ab4b),
	.w7(32'hbba88a8d),
	.w8(32'hbbbdd2f8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae23777),
	.w1(32'h3bdadcda),
	.w2(32'hbb2a2f32),
	.w3(32'hbb1fd8bc),
	.w4(32'h3b6145cc),
	.w5(32'h3931dd98),
	.w6(32'h3be5dd04),
	.w7(32'h3c156222),
	.w8(32'h3baf5b43),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdb2cb),
	.w1(32'h3b33edd1),
	.w2(32'hbba89cda),
	.w3(32'h3b71d45d),
	.w4(32'h39e195ae),
	.w5(32'hb703237f),
	.w6(32'h3addb6b0),
	.w7(32'hbbbe1ff2),
	.w8(32'hbc08a90a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f4993),
	.w1(32'h3be072d9),
	.w2(32'hb9c19f81),
	.w3(32'h3b574c7f),
	.w4(32'h3b94e308),
	.w5(32'h3aaef3b7),
	.w6(32'h3c154861),
	.w7(32'h3c307948),
	.w8(32'h3c29e67c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cd0eb),
	.w1(32'hbb74e4a0),
	.w2(32'h3b0ac9c6),
	.w3(32'h3a9dee54),
	.w4(32'h38ece102),
	.w5(32'h3aa1bcd8),
	.w6(32'hbae2d1c9),
	.w7(32'hbb1b96de),
	.w8(32'h394f07ca),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9e269),
	.w1(32'h3b70835f),
	.w2(32'hbae5193c),
	.w3(32'hbaa9f0ab),
	.w4(32'h3b1373a1),
	.w5(32'hbb9e5816),
	.w6(32'h3b73354a),
	.w7(32'h3bcc1e34),
	.w8(32'h3b30d9c8),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48bc2f),
	.w1(32'h3b95c870),
	.w2(32'hbbc87352),
	.w3(32'h3b297ed5),
	.w4(32'h3b06c1e0),
	.w5(32'hbbc6d5b2),
	.w6(32'h3bcf1516),
	.w7(32'h3bdc7dd0),
	.w8(32'h3b5f384a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbbdb0),
	.w1(32'h3b0f364d),
	.w2(32'hbb5cf706),
	.w3(32'h38c8cffe),
	.w4(32'h3a07a96f),
	.w5(32'hbb9374c0),
	.w6(32'h3b270bd3),
	.w7(32'h3b85c5d4),
	.w8(32'h3aea3ecf),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e9e12),
	.w1(32'h3b079c47),
	.w2(32'hbb8202c8),
	.w3(32'hba39ce98),
	.w4(32'h3acf61c3),
	.w5(32'hbb6d2098),
	.w6(32'h3b45783d),
	.w7(32'h3bab740a),
	.w8(32'h3b077602),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafb4e7),
	.w1(32'h39ec0830),
	.w2(32'h3b7ae540),
	.w3(32'hb9715d84),
	.w4(32'h3ae073d6),
	.w5(32'hbaf0470f),
	.w6(32'h3b3745f9),
	.w7(32'hb67a029a),
	.w8(32'hba88d904),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafcd65),
	.w1(32'hbb820dfb),
	.w2(32'hb6e416ce),
	.w3(32'h3b9849ca),
	.w4(32'hbb3ab765),
	.w5(32'h3ac95f4b),
	.w6(32'hbb5af688),
	.w7(32'hbaaf6a46),
	.w8(32'h3af015a6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a417954),
	.w1(32'hbb90e094),
	.w2(32'hbbcc2bb1),
	.w3(32'hba0ab95e),
	.w4(32'hb99f70f6),
	.w5(32'h3a87e27b),
	.w6(32'hbb8303a9),
	.w7(32'hbaef00c8),
	.w8(32'hba255f62),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb546c9c),
	.w1(32'hbb17df7c),
	.w2(32'hbb27d00d),
	.w3(32'h3b5418d6),
	.w4(32'hba1fdb97),
	.w5(32'h3b31d51d),
	.w6(32'hbb918fdf),
	.w7(32'h39c4fea6),
	.w8(32'h36eaeb6e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f9082),
	.w1(32'h3bbba2da),
	.w2(32'hbbc0f59c),
	.w3(32'h39c12d55),
	.w4(32'h3b377783),
	.w5(32'hbbe999d6),
	.w6(32'h3b6cb28b),
	.w7(32'h3bb311f1),
	.w8(32'h3a24c0d1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdff39),
	.w1(32'hbb57c574),
	.w2(32'h3be1d338),
	.w3(32'hba6dd8d2),
	.w4(32'hbba53a76),
	.w5(32'hbb69d97c),
	.w6(32'hbad10ab7),
	.w7(32'hbba0c1e0),
	.w8(32'hbb924314),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7119c1),
	.w1(32'hba8c6e49),
	.w2(32'hbbaf3a62),
	.w3(32'h3a56b77b),
	.w4(32'hbadea0a2),
	.w5(32'hbbb99db3),
	.w6(32'hb914057c),
	.w7(32'h3b09418c),
	.w8(32'h3b7819f6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbff763),
	.w1(32'hbb8f251d),
	.w2(32'hbc0f3916),
	.w3(32'hbb0ebbbd),
	.w4(32'h3945351e),
	.w5(32'hbb230394),
	.w6(32'hbbfd5c55),
	.w7(32'hbb3f493f),
	.w8(32'h39053a3e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d7166),
	.w1(32'hbb09f630),
	.w2(32'hba37b5be),
	.w3(32'h3b19ca52),
	.w4(32'hba73b957),
	.w5(32'hba07029d),
	.w6(32'hbab2d938),
	.w7(32'hb9edaec7),
	.w8(32'h3af15e4a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb253e20),
	.w1(32'hbb7e4ede),
	.w2(32'hbb6fa1ea),
	.w3(32'h3a81605b),
	.w4(32'hbba0b26c),
	.w5(32'hbb547c6b),
	.w6(32'h3a33cfa7),
	.w7(32'hba4cec12),
	.w8(32'h3b4f2774),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b3623),
	.w1(32'hbaeb20a9),
	.w2(32'h3b867e34),
	.w3(32'hbb7fdb04),
	.w4(32'hbade0222),
	.w5(32'h3b04fef7),
	.w6(32'h3b2d1e5d),
	.w7(32'h3c1aae46),
	.w8(32'h3c05c7a1),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3baebc),
	.w1(32'hb7864c31),
	.w2(32'hba0e72a9),
	.w3(32'hbaf76e71),
	.w4(32'hbae7993a),
	.w5(32'hbad99a9a),
	.w6(32'hb902faed),
	.w7(32'hb9e6c3c3),
	.w8(32'hba494a50),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57377d),
	.w1(32'h3a8baddc),
	.w2(32'h3a73a06d),
	.w3(32'hba920aa4),
	.w4(32'hb99a9bd9),
	.w5(32'hb9ce7273),
	.w6(32'h3a157909),
	.w7(32'h3a0b1d27),
	.w8(32'h3a8f79b0),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2308d0),
	.w1(32'h3a040f73),
	.w2(32'hb9b9d02a),
	.w3(32'hb95d7fdd),
	.w4(32'hbb3182f7),
	.w5(32'hbb6a6948),
	.w6(32'h3bd0e3ff),
	.w7(32'h3b7dc20e),
	.w8(32'h3ba7ae96),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81e38d),
	.w1(32'h39a37c95),
	.w2(32'hbac46b39),
	.w3(32'hbafaf5f6),
	.w4(32'h39f96f08),
	.w5(32'hb99ce407),
	.w6(32'h3a28ee54),
	.w7(32'hbb34f89d),
	.w8(32'h39b2f6e6),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2113f),
	.w1(32'h3a42fe67),
	.w2(32'hb8b0a81f),
	.w3(32'h3b0ba14e),
	.w4(32'h392fe156),
	.w5(32'hbab3aad2),
	.w6(32'hbaab8af7),
	.w7(32'hbb2b2e6e),
	.w8(32'hb9abf640),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5b8cd),
	.w1(32'hba393f9b),
	.w2(32'hbab1d9b9),
	.w3(32'hbb43d2e7),
	.w4(32'hbb039129),
	.w5(32'hba66c99e),
	.w6(32'h3ab80159),
	.w7(32'hba1d1c46),
	.w8(32'h3ad4825b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78c0f0),
	.w1(32'hba87b961),
	.w2(32'hbb24848a),
	.w3(32'hba07de37),
	.w4(32'hb89e14e1),
	.w5(32'hbb13f53a),
	.w6(32'hba9b8c88),
	.w7(32'hbb395d03),
	.w8(32'hbb068f59),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae606c0),
	.w1(32'h3a0096c9),
	.w2(32'h3ac0667a),
	.w3(32'hbaf7ac84),
	.w4(32'h3abd4cf5),
	.w5(32'h3acf4a06),
	.w6(32'h3aa6e3d7),
	.w7(32'h3b07b8dd),
	.w8(32'h3ae189a1),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04465d),
	.w1(32'h3af0b541),
	.w2(32'h3b43c8de),
	.w3(32'hbb10487c),
	.w4(32'hb9f51cdc),
	.w5(32'h3abb81f7),
	.w6(32'h3b24bf9a),
	.w7(32'h3b13e9ed),
	.w8(32'h3b19f2df),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a671487),
	.w1(32'h3bd113c8),
	.w2(32'h3bec30f6),
	.w3(32'h3a413cb2),
	.w4(32'h3c0a3dee),
	.w5(32'h3c19dd36),
	.w6(32'h3c0765e0),
	.w7(32'h3bab2739),
	.w8(32'h3ba2fd88),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fa981),
	.w1(32'h3b05fb35),
	.w2(32'h3b7bb4e0),
	.w3(32'h3c04ce92),
	.w4(32'hba3b079c),
	.w5(32'h3a655154),
	.w6(32'h3b2f29eb),
	.w7(32'h3a31084d),
	.w8(32'h3b00da28),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4dc423),
	.w1(32'h38d44836),
	.w2(32'h39a619fa),
	.w3(32'hb964d765),
	.w4(32'h3ae2445d),
	.w5(32'h3adbffbb),
	.w6(32'h39f76067),
	.w7(32'h38bbb4e0),
	.w8(32'h3a4925c8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fa5e8),
	.w1(32'hbb3f778d),
	.w2(32'hbb8c73fb),
	.w3(32'h3b0297f7),
	.w4(32'hba13932a),
	.w5(32'hbb8714c8),
	.w6(32'hbb19d4fa),
	.w7(32'hbb8544cf),
	.w8(32'hbb5bb6e4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01fae6),
	.w1(32'h3b895e57),
	.w2(32'h3bace3ec),
	.w3(32'hbb1ae4aa),
	.w4(32'hba43417c),
	.w5(32'h39f9e0d7),
	.w6(32'h3b52acbe),
	.w7(32'hbb88e844),
	.w8(32'hbb7561ef),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17fa8c),
	.w1(32'hbaacaaac),
	.w2(32'hba2ea5a4),
	.w3(32'h3b1f5019),
	.w4(32'hb994bbdf),
	.w5(32'hb9ad1eb6),
	.w6(32'hbaa1565c),
	.w7(32'h3968c9dc),
	.w8(32'h3a3008bd),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38da29a9),
	.w1(32'h3b638b77),
	.w2(32'h3bfaaa23),
	.w3(32'hb792c1b8),
	.w4(32'h3a395d09),
	.w5(32'h3b2ef760),
	.w6(32'h39ec0381),
	.w7(32'h3b52b1b5),
	.w8(32'h3a5eda42),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8216e6),
	.w1(32'h33ac20b6),
	.w2(32'hbb06a13c),
	.w3(32'hbaab25b0),
	.w4(32'hbaf2b3b5),
	.w5(32'hbb24c6e9),
	.w6(32'h3a792b54),
	.w7(32'hb8e44a5e),
	.w8(32'h399d1052),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ce55ee),
	.w1(32'h3981732d),
	.w2(32'hba338b77),
	.w3(32'hb962f962),
	.w4(32'hb9dac3b8),
	.w5(32'hba5ca714),
	.w6(32'h3a99dc5d),
	.w7(32'h3a9ae4e1),
	.w8(32'h3a87fbbe),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf4d8e),
	.w1(32'h3abfd018),
	.w2(32'h3b7f16b0),
	.w3(32'h39de5564),
	.w4(32'h3af48ac3),
	.w5(32'h3b423c4f),
	.w6(32'h3b5edf4c),
	.w7(32'h3b90614a),
	.w8(32'h3b94a71f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a7f5f),
	.w1(32'hbafd1a18),
	.w2(32'hbaf340fc),
	.w3(32'h3ad73e63),
	.w4(32'hba88deea),
	.w5(32'hbad1a6b2),
	.w6(32'hbadc1b69),
	.w7(32'hbabc98ab),
	.w8(32'hba8f54fa),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb030372),
	.w1(32'h3b4743fa),
	.w2(32'h3baa5c97),
	.w3(32'hbb2a24a0),
	.w4(32'h3bcd396a),
	.w5(32'h3ba25717),
	.w6(32'h3b8e515e),
	.w7(32'h3be6dbc9),
	.w8(32'h3bdf794f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65cd45),
	.w1(32'h3b265c76),
	.w2(32'h3a8dfa27),
	.w3(32'h3a90320a),
	.w4(32'h3b5dca3f),
	.w5(32'h3aaf5210),
	.w6(32'h3a68416d),
	.w7(32'hb9f5d1f7),
	.w8(32'h3a77dd0a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af15345),
	.w1(32'hbb104975),
	.w2(32'hb9e83fa0),
	.w3(32'h3afc1198),
	.w4(32'hb944a484),
	.w5(32'h3a52fc5f),
	.w6(32'hb9fb4d91),
	.w7(32'hbb0066ba),
	.w8(32'h3984b771),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e5312),
	.w1(32'h3b8455b6),
	.w2(32'h3b8d38b9),
	.w3(32'hbaaa32b6),
	.w4(32'h3b555c61),
	.w5(32'h3ad8731f),
	.w6(32'h3b2c4880),
	.w7(32'h3b9793b0),
	.w8(32'h3b61b3c8),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e2c3d),
	.w1(32'h3c13e7fe),
	.w2(32'h3c91c4ec),
	.w3(32'h38e835b4),
	.w4(32'hb992d0bc),
	.w5(32'hb8c0a33a),
	.w6(32'h3bb3eda6),
	.w7(32'h3bf229a5),
	.w8(32'h3b8e7273),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c312f6b),
	.w1(32'h3b51cdbd),
	.w2(32'h3b63ed64),
	.w3(32'hb9e12304),
	.w4(32'h3b33b808),
	.w5(32'h3b0759e7),
	.w6(32'h3b2a5a77),
	.w7(32'h3b2bc078),
	.w8(32'h3b3bb60f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b0d45),
	.w1(32'h3b59abb0),
	.w2(32'h3b80186a),
	.w3(32'h3b35ad40),
	.w4(32'h3b844f53),
	.w5(32'h3b63b454),
	.w6(32'h3b502ac6),
	.w7(32'h3bb567cc),
	.w8(32'h3ba50a39),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f9ef1),
	.w1(32'h3b168b50),
	.w2(32'h3b030322),
	.w3(32'h3b17b115),
	.w4(32'h39b95948),
	.w5(32'hbac77188),
	.w6(32'h3b0aef67),
	.w7(32'h3a95a5cc),
	.w8(32'h3a88d6d5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e81a2),
	.w1(32'h3ba0e32b),
	.w2(32'h3bd0cde8),
	.w3(32'h38b8443c),
	.w4(32'h3a129b4b),
	.w5(32'h3aa8c02a),
	.w6(32'h3b7bb7bf),
	.w7(32'h3bad9d33),
	.w8(32'h3b3f9a25),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac95cf),
	.w1(32'hb9312d97),
	.w2(32'h397acb94),
	.w3(32'hba6f2739),
	.w4(32'h39eb83f8),
	.w5(32'h39de539c),
	.w6(32'hb8bd2a4e),
	.w7(32'h394540d3),
	.w8(32'h3a51cdf9),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d9591),
	.w1(32'h3afc5fce),
	.w2(32'h3afc14f8),
	.w3(32'h39444f85),
	.w4(32'h3b0f9efa),
	.w5(32'h3abfedc8),
	.w6(32'h3ae097e1),
	.w7(32'h3aab7520),
	.w8(32'h3aa73385),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77f818),
	.w1(32'h3c044640),
	.w2(32'h3c2d7540),
	.w3(32'hb8155332),
	.w4(32'h3c0308ba),
	.w5(32'h3c1fa55f),
	.w6(32'h3c12b4fa),
	.w7(32'h3c2f146d),
	.w8(32'h3b8ca82d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b97e52),
	.w1(32'h3b0a3999),
	.w2(32'h3c44b95c),
	.w3(32'h39218ea8),
	.w4(32'h3973f931),
	.w5(32'h3b80d0ba),
	.w6(32'h3b85a870),
	.w7(32'h3c2370ae),
	.w8(32'h3c10df83),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ffbde),
	.w1(32'h3a827f8f),
	.w2(32'h3a3ccb97),
	.w3(32'h3c286230),
	.w4(32'hba7c4da9),
	.w5(32'hbab13b58),
	.w6(32'h3b11ebc7),
	.w7(32'h3add2193),
	.w8(32'h3ac243cf),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b455eb),
	.w1(32'h3b52c64c),
	.w2(32'h3b3dadb7),
	.w3(32'hba8f34da),
	.w4(32'h3b443212),
	.w5(32'h3acee556),
	.w6(32'h3b2812f7),
	.w7(32'h3b0ef072),
	.w8(32'h3b50f586),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae297b8),
	.w1(32'h38c96937),
	.w2(32'hb9acb794),
	.w3(32'h3a647455),
	.w4(32'hbb4f90ee),
	.w5(32'hbb446947),
	.w6(32'h3ab518ad),
	.w7(32'hbb19fedb),
	.w8(32'hbab234e7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c6a70),
	.w1(32'h3a9d97b0),
	.w2(32'h3910a80f),
	.w3(32'hb90f8cb7),
	.w4(32'hb9b6429c),
	.w5(32'hba5230df),
	.w6(32'h3ace3d5f),
	.w7(32'h3a35a7c3),
	.w8(32'h3a43461f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33c9ef),
	.w1(32'hbae82549),
	.w2(32'hbb218c5d),
	.w3(32'h392d3880),
	.w4(32'hba2dfcde),
	.w5(32'hbb0398f0),
	.w6(32'hbaf4ef1e),
	.w7(32'hbb1b1a0e),
	.w8(32'hbaa13573),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b0d72),
	.w1(32'h3a78afc2),
	.w2(32'hb8b101ab),
	.w3(32'hba0112bc),
	.w4(32'h3903df82),
	.w5(32'hb9916f6c),
	.w6(32'h3a843ee5),
	.w7(32'hb9ede84f),
	.w8(32'hb7e3b324),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f632e),
	.w1(32'h3b549b59),
	.w2(32'h3c151e3e),
	.w3(32'hba46e2e0),
	.w4(32'h3a6b6dd2),
	.w5(32'h3bbebf74),
	.w6(32'h3bbce2d0),
	.w7(32'h3c3e0507),
	.w8(32'h3c385a90),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dd3d2),
	.w1(32'h3ad65e1c),
	.w2(32'h3b87d0fc),
	.w3(32'h3ba60a1b),
	.w4(32'hbb070bbd),
	.w5(32'hba28b680),
	.w6(32'h3ac60d7f),
	.w7(32'h3b7e4561),
	.w8(32'h3b541f46),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b020903),
	.w1(32'h3b615f47),
	.w2(32'h3ba32310),
	.w3(32'h3aa18854),
	.w4(32'h3b85bcd7),
	.w5(32'h3b867ddd),
	.w6(32'h3b7516d3),
	.w7(32'h3b3c89cb),
	.w8(32'h3b404923),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b349c9d),
	.w1(32'h3b3b5466),
	.w2(32'h3ac11b5c),
	.w3(32'h3b075a5a),
	.w4(32'h3b0f01dd),
	.w5(32'h3a374400),
	.w6(32'h3b1ec49c),
	.w7(32'h3aad2289),
	.w8(32'hb9846b5a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba870f4f),
	.w1(32'hbb674936),
	.w2(32'hbb850c71),
	.w3(32'h39d2b897),
	.w4(32'h39ecb893),
	.w5(32'hba9a4b32),
	.w6(32'hbaf7db28),
	.w7(32'hbb078cbf),
	.w8(32'h391f0557),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfa477),
	.w1(32'h3a36e083),
	.w2(32'h3a4cdbc6),
	.w3(32'hbba03559),
	.w4(32'h3a6f14b6),
	.w5(32'h3aa1d410),
	.w6(32'h3b3fd953),
	.w7(32'h3b01db58),
	.w8(32'h3b5aa868),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2a87d),
	.w1(32'hb9a83503),
	.w2(32'hba185174),
	.w3(32'h39a6108b),
	.w4(32'hbaed20b4),
	.w5(32'hb9cae7bd),
	.w6(32'h3b1af04d),
	.w7(32'hb9954942),
	.w8(32'h3b546791),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf2211),
	.w1(32'h3ab12f3b),
	.w2(32'h3b558284),
	.w3(32'h3907033e),
	.w4(32'h3a9ccb30),
	.w5(32'h3ab2d8d0),
	.w6(32'hb994a61f),
	.w7(32'h3ad7daf2),
	.w8(32'hba5b1111),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e8830),
	.w1(32'h3b8d1c71),
	.w2(32'h3bfbc348),
	.w3(32'hbaaf05d4),
	.w4(32'h3b7afa2a),
	.w5(32'h3b9ea5e3),
	.w6(32'h3b79e1ac),
	.w7(32'h3b86aa26),
	.w8(32'h3b81af58),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baad688),
	.w1(32'hbb0d6871),
	.w2(32'hbb53104e),
	.w3(32'h3b8c373a),
	.w4(32'hba5d7003),
	.w5(32'hbb35fae1),
	.w6(32'hbb01d032),
	.w7(32'hbb45e211),
	.w8(32'hbb0626e4),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2370cf),
	.w1(32'hbb4ed278),
	.w2(32'hbb167de2),
	.w3(32'hbb34050e),
	.w4(32'hbb8663fc),
	.w5(32'hbb88005f),
	.w6(32'hba124678),
	.w7(32'hbb033611),
	.w8(32'hb898e8bd),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89435b4),
	.w1(32'hbb478a4b),
	.w2(32'h3b85367b),
	.w3(32'hba6a8a50),
	.w4(32'h3af80fa3),
	.w5(32'h3bac2d11),
	.w6(32'hbb9c9db3),
	.w7(32'h3b57cb75),
	.w8(32'h3abf68f0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3745b6),
	.w1(32'h3b614a95),
	.w2(32'h3baf780f),
	.w3(32'h38757f3b),
	.w4(32'h3a736259),
	.w5(32'h3b3d961c),
	.w6(32'h3b3b18f1),
	.w7(32'h3b4e00f0),
	.w8(32'h3bac6ba4),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba89c15),
	.w1(32'h3b731ca8),
	.w2(32'h3930ce48),
	.w3(32'h3b2618f3),
	.w4(32'h3b22ace3),
	.w5(32'h3734f77c),
	.w6(32'h3b4be705),
	.w7(32'hbac5ec66),
	.w8(32'h39c412a4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b9812),
	.w1(32'h3bca0803),
	.w2(32'h3c0ac63f),
	.w3(32'h3b0b6793),
	.w4(32'h3b132200),
	.w5(32'h3bad9981),
	.w6(32'h3bbaf71e),
	.w7(32'h3bdda9ef),
	.w8(32'h3aadd2be),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac55a59),
	.w1(32'h3b724b3c),
	.w2(32'h3a721192),
	.w3(32'h3abea21d),
	.w4(32'h3b02fe2e),
	.w5(32'hb9ccef56),
	.w6(32'h3bad48c9),
	.w7(32'h3b89a892),
	.w8(32'h3c04c3ac),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3bcfe),
	.w1(32'hbb841a7b),
	.w2(32'h3aba2337),
	.w3(32'h3ba96511),
	.w4(32'hbb4b13f1),
	.w5(32'h3a7965dc),
	.w6(32'hba2b6306),
	.w7(32'h39b5d73d),
	.w8(32'h398d7a36),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa32199),
	.w1(32'hbb3124f6),
	.w2(32'hba973bbb),
	.w3(32'hbb5a8e1e),
	.w4(32'hbb24611c),
	.w5(32'hba8e8c21),
	.w6(32'h39383658),
	.w7(32'hbab8c2ec),
	.w8(32'h3b567343),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959362c),
	.w1(32'hb92857bf),
	.w2(32'hbaa73719),
	.w3(32'h3a802751),
	.w4(32'hb9f33d64),
	.w5(32'hbab2b325),
	.w6(32'hb9a0eaf7),
	.w7(32'hb8bade4c),
	.w8(32'hbabb2782),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba69c41),
	.w1(32'hbafb140e),
	.w2(32'h385db667),
	.w3(32'hbb75b4be),
	.w4(32'hb8b8863e),
	.w5(32'h3aeb9ebe),
	.w6(32'h3b88d4e2),
	.w7(32'h3b14e9b8),
	.w8(32'h3bc53369),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acf193),
	.w1(32'h39ca67b1),
	.w2(32'hbaac9fbe),
	.w3(32'hbacf14f0),
	.w4(32'h3b3861e3),
	.w5(32'hbad34967),
	.w6(32'hba69ffc0),
	.w7(32'h39cba1ac),
	.w8(32'hba830adb),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6d3a8),
	.w1(32'hba8884c0),
	.w2(32'hbaf06060),
	.w3(32'hbb1ef3cd),
	.w4(32'hb983c871),
	.w5(32'hba85da98),
	.w6(32'hbae5b45a),
	.w7(32'hbaa8e97a),
	.w8(32'hb9a3fcd5),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8921f),
	.w1(32'h3c23de07),
	.w2(32'h3bfaa803),
	.w3(32'hbaafa472),
	.w4(32'h3c3fe138),
	.w5(32'h3be0f99c),
	.w6(32'h3c0c8964),
	.w7(32'h3c1c3d2e),
	.w8(32'h3b8c3b36),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad634b4),
	.w1(32'h3b1d8347),
	.w2(32'h3a9afec9),
	.w3(32'h38f09afa),
	.w4(32'h3a956556),
	.w5(32'h3a062852),
	.w6(32'h3b0776e4),
	.w7(32'h3a844d94),
	.w8(32'hb914c5be),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39906a14),
	.w1(32'hb942f87f),
	.w2(32'hbaa5bf2e),
	.w3(32'h39e87e07),
	.w4(32'hb98d7f94),
	.w5(32'hba8273cf),
	.w6(32'h3979794a),
	.w7(32'hba874f71),
	.w8(32'hbaa154f2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb407c6b),
	.w1(32'hbaf0869b),
	.w2(32'h3a965f37),
	.w3(32'hbb0be124),
	.w4(32'hbae731f5),
	.w5(32'h3ae232a7),
	.w6(32'h3a8a7e0a),
	.w7(32'h3acd78b0),
	.w8(32'h3bc2b378),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba04245),
	.w1(32'h3b5af9cc),
	.w2(32'h3bed6906),
	.w3(32'h3b537ecd),
	.w4(32'hbb00e4d3),
	.w5(32'h3b188ce3),
	.w6(32'h3b4664d1),
	.w7(32'h3bd1a528),
	.w8(32'h3bc43962),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00ae6e),
	.w1(32'h3a35fd85),
	.w2(32'h3bb6435d),
	.w3(32'h3ba36b73),
	.w4(32'hba6a7f06),
	.w5(32'h3b31c2e0),
	.w6(32'hbb0d9a0e),
	.w7(32'h3a9e3593),
	.w8(32'h3b23cfea),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11ca01),
	.w1(32'h3a857d33),
	.w2(32'h3a7e6d0a),
	.w3(32'h3bc9ea45),
	.w4(32'h3a57ef6b),
	.w5(32'h3a1ee5e5),
	.w6(32'hb8c42a3b),
	.w7(32'h38da8896),
	.w8(32'h3a8460b1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b835a),
	.w1(32'hbbac2bb7),
	.w2(32'hbb7fb183),
	.w3(32'hba7e86f9),
	.w4(32'hbb735a98),
	.w5(32'hbb15616f),
	.w6(32'h3a98c21a),
	.w7(32'hba8e9256),
	.w8(32'h3b059059),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb119cb2),
	.w1(32'hb826fb47),
	.w2(32'hb9edb21b),
	.w3(32'hba81f4e6),
	.w4(32'hba6e4233),
	.w5(32'hb8942a9b),
	.w6(32'h3a4a14da),
	.w7(32'h39cf1c32),
	.w8(32'h3a85872f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc61c1),
	.w1(32'h3a508e13),
	.w2(32'hba6291c6),
	.w3(32'hb9a8714f),
	.w4(32'h3aa96fcb),
	.w5(32'hb92a60ac),
	.w6(32'h3a0f38d5),
	.w7(32'hb977fb8e),
	.w8(32'h3a85c8fc),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce3888),
	.w1(32'hbaf24144),
	.w2(32'hbad6c214),
	.w3(32'h3a242ebd),
	.w4(32'hba3a44ec),
	.w5(32'hba89f910),
	.w6(32'h3942bb04),
	.w7(32'hbabb68d1),
	.w8(32'hba0f06dc),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba744f7c),
	.w1(32'h3b476f14),
	.w2(32'h3b43f49e),
	.w3(32'hba6b5c07),
	.w4(32'h3b3f3735),
	.w5(32'h3b081d57),
	.w6(32'h3b1e8718),
	.w7(32'h3ac8991a),
	.w8(32'h3adca30b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27b3ba),
	.w1(32'hbabb44cf),
	.w2(32'hb9f26579),
	.w3(32'h3b012460),
	.w4(32'hbaf80901),
	.w5(32'hba81d6d5),
	.w6(32'hba3229f8),
	.w7(32'h396b30a0),
	.w8(32'hb92e7f1a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7155c0),
	.w1(32'h3bccbb81),
	.w2(32'h3c409f75),
	.w3(32'hba90a2ab),
	.w4(32'hbb8207f7),
	.w5(32'hbafba600),
	.w6(32'h3b641001),
	.w7(32'h3beb3711),
	.w8(32'h3b9c2102),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fa629),
	.w1(32'hba059b0c),
	.w2(32'hbb08d593),
	.w3(32'hba42eb07),
	.w4(32'h3a8b7d11),
	.w5(32'hbabdc467),
	.w6(32'h39c8e0c7),
	.w7(32'hbaeecb2b),
	.w8(32'hb919e346),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cb3fe),
	.w1(32'h398bb0b2),
	.w2(32'hb9938155),
	.w3(32'hbaa0d36a),
	.w4(32'hba1c5bcb),
	.w5(32'hbadc01ab),
	.w6(32'hb82c2c3a),
	.w7(32'h3aeb00fa),
	.w8(32'hbadeefdf),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ebd52),
	.w1(32'h3c2fbc80),
	.w2(32'h3c864bd1),
	.w3(32'hbb45db87),
	.w4(32'h3b7939fe),
	.w5(32'h3be6b4ff),
	.w6(32'h3bf520e5),
	.w7(32'h3c2dfcfa),
	.w8(32'h3b813919),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b986de6),
	.w1(32'hbaf5023f),
	.w2(32'hb9afc6d8),
	.w3(32'h39cb9f9b),
	.w4(32'hba7179d5),
	.w5(32'hb94147fe),
	.w6(32'hb9f357c7),
	.w7(32'h3985ddf7),
	.w8(32'h3ae921b2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba663ebd),
	.w1(32'hba2db200),
	.w2(32'h3ba45046),
	.w3(32'hb94fbbcb),
	.w4(32'hba9082d0),
	.w5(32'h3b8f7615),
	.w6(32'hbab7991e),
	.w7(32'h3b64dee1),
	.w8(32'h3bb1f37a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7ad63),
	.w1(32'hbb15aa74),
	.w2(32'h3996028a),
	.w3(32'h3ba7733c),
	.w4(32'hbb1bd3d9),
	.w5(32'h39c0e306),
	.w6(32'hbb330e27),
	.w7(32'hba0f927e),
	.w8(32'h3a67948a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940c011),
	.w1(32'h3bde418b),
	.w2(32'h3c1086c7),
	.w3(32'h39bdc197),
	.w4(32'h3b7ea46d),
	.w5(32'h3b994f75),
	.w6(32'h3baa92a1),
	.w7(32'h3bf3ebf4),
	.w8(32'h3ba0993f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b389362),
	.w1(32'hbaf67dde),
	.w2(32'hb9df37f5),
	.w3(32'h3ad02bda),
	.w4(32'hba4dd017),
	.w5(32'h39f57203),
	.w6(32'hb95da736),
	.w7(32'h3a289445),
	.w8(32'h3b263ffe),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49dce9),
	.w1(32'hbb3eb247),
	.w2(32'h3aa9bfec),
	.w3(32'hbb09beea),
	.w4(32'h3b7796da),
	.w5(32'h3bd4c261),
	.w6(32'hbb3db0a4),
	.w7(32'hbb238f0e),
	.w8(32'hbad3fe0a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba629c70),
	.w1(32'hba2c9eed),
	.w2(32'h3afd5c59),
	.w3(32'h3b9fcc56),
	.w4(32'hbacb7427),
	.w5(32'h3aaed807),
	.w6(32'h3a52a006),
	.w7(32'h3ab8c1db),
	.w8(32'h3b41b33f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61ba69),
	.w1(32'hba6b1495),
	.w2(32'h3ab63c0d),
	.w3(32'hbb5fb68a),
	.w4(32'hba9f33f7),
	.w5(32'h3a0edda9),
	.w6(32'hbacd22ff),
	.w7(32'h39b33fd9),
	.w8(32'hbb23eb9f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba512e3c),
	.w1(32'hb97b742e),
	.w2(32'hb987203e),
	.w3(32'hbb1e353b),
	.w4(32'h37ede091),
	.w5(32'hb9d99737),
	.w6(32'hb957e5a5),
	.w7(32'hb9fcbce8),
	.w8(32'hb96846a1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba275e18),
	.w1(32'h3b95d655),
	.w2(32'h3be73efc),
	.w3(32'hb9b5642b),
	.w4(32'h3ae6f30a),
	.w5(32'h3b98b608),
	.w6(32'h3bbf72c8),
	.w7(32'h3bd49a6e),
	.w8(32'h3b0975a9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b3272),
	.w1(32'hbb445f08),
	.w2(32'hbb2bf92a),
	.w3(32'hbb21b870),
	.w4(32'hbb3d0644),
	.w5(32'hba7df1d3),
	.w6(32'h394635ee),
	.w7(32'hbb0205db),
	.w8(32'h3ac08951),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a11f7),
	.w1(32'hba0fac3e),
	.w2(32'h3b0e6374),
	.w3(32'hbb134763),
	.w4(32'h3b08eca4),
	.w5(32'h3b76bf58),
	.w6(32'h3b828267),
	.w7(32'h3b72be3e),
	.w8(32'h3bb386e9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d37d1b),
	.w1(32'h3b4b949a),
	.w2(32'h3b7855dd),
	.w3(32'hba574d4d),
	.w4(32'h39cccb9f),
	.w5(32'h3b365256),
	.w6(32'h3b8a9203),
	.w7(32'h3b3b031f),
	.w8(32'h3b434f93),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48218e),
	.w1(32'h3a9a4c3c),
	.w2(32'h3b3fc9dd),
	.w3(32'h3b70bcab),
	.w4(32'h39300dc2),
	.w5(32'h3b14eb39),
	.w6(32'hba2d8821),
	.w7(32'h3a3006ee),
	.w8(32'hba6d9443),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac660c2),
	.w1(32'hbafeac4a),
	.w2(32'hb7768b80),
	.w3(32'h3a9f7a9f),
	.w4(32'hbb2bc3a6),
	.w5(32'hbb0aa19b),
	.w6(32'hbb936660),
	.w7(32'hbb37c280),
	.w8(32'h37796251),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb86787),
	.w1(32'h3a734caf),
	.w2(32'h3a9e4c70),
	.w3(32'h3b8db886),
	.w4(32'hba035a03),
	.w5(32'hbaa0c157),
	.w6(32'h3a9367a9),
	.w7(32'h3a44de22),
	.w8(32'h3a6f25a4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c1bfc),
	.w1(32'h3acb4f54),
	.w2(32'hbac60895),
	.w3(32'hba1d19ec),
	.w4(32'h392af7e2),
	.w5(32'hbb837b59),
	.w6(32'h3b2a020d),
	.w7(32'h3a64d3c0),
	.w8(32'h3aa953b8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaedbed),
	.w1(32'h3aeb9803),
	.w2(32'h3a1970a5),
	.w3(32'hbb87a68b),
	.w4(32'hb89efb1c),
	.w5(32'hba986d58),
	.w6(32'h3aa352de),
	.w7(32'h3b1b9a35),
	.w8(32'h3ad47792),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a856bbe),
	.w1(32'h3ac8576e),
	.w2(32'h3a9e5889),
	.w3(32'hb90ec81f),
	.w4(32'h3b267a7a),
	.w5(32'h3ac3f637),
	.w6(32'h3b453137),
	.w7(32'h3b4f6862),
	.w8(32'h3b0d4b57),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f27f0a),
	.w1(32'hba9ab44d),
	.w2(32'hbabb7204),
	.w3(32'hbaaa3e23),
	.w4(32'hbb1ed378),
	.w5(32'hb9b2ee64),
	.w6(32'hba7f40f9),
	.w7(32'hba8515a0),
	.w8(32'h3a98f8b7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab49688),
	.w1(32'h3aeed7af),
	.w2(32'h3bb18453),
	.w3(32'h3ad994f6),
	.w4(32'h392e123d),
	.w5(32'h3b750158),
	.w6(32'h3b918a7e),
	.w7(32'h3b8d281f),
	.w8(32'h3b98a280),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96e421),
	.w1(32'h3b82f7dd),
	.w2(32'h3bdda397),
	.w3(32'h3b491a1c),
	.w4(32'h3b126aef),
	.w5(32'h3b8465e3),
	.w6(32'h3bf72398),
	.w7(32'h3bbb5ea8),
	.w8(32'h3c4aa645),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f13e6),
	.w1(32'h3b06e375),
	.w2(32'h3ac5f2ef),
	.w3(32'h3c3cb122),
	.w4(32'h3acc8503),
	.w5(32'hbad1e53d),
	.w6(32'h37d6b9ef),
	.w7(32'hb933212b),
	.w8(32'h3aea759f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ac3e5),
	.w1(32'hbb7ef310),
	.w2(32'hbb9d1319),
	.w3(32'hbbe23e85),
	.w4(32'hbab43527),
	.w5(32'hbb06c155),
	.w6(32'h379284ac),
	.w7(32'hbb71a388),
	.w8(32'hb9eddf91),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb115e12),
	.w1(32'hb9100c88),
	.w2(32'hba7badfb),
	.w3(32'hbb12d3ef),
	.w4(32'h39bd7531),
	.w5(32'hb9c4ba6e),
	.w6(32'h3a8b9935),
	.w7(32'h39b01884),
	.w8(32'h3b25afe0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83c0b9),
	.w1(32'hba571e80),
	.w2(32'hbb0e812a),
	.w3(32'h3a0e2c2a),
	.w4(32'h3a2a5475),
	.w5(32'hbab270e7),
	.w6(32'hb9c776c3),
	.w7(32'hbaf94002),
	.w8(32'hba344dfc),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbb5e7),
	.w1(32'h3aeeaee9),
	.w2(32'h3b6821d2),
	.w3(32'hbb1efd8d),
	.w4(32'h3b11028e),
	.w5(32'h3b37b3f7),
	.w6(32'h3b134cf5),
	.w7(32'h3b8ea660),
	.w8(32'h3b849236),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1de51f),
	.w1(32'hb9773577),
	.w2(32'hba4e5c32),
	.w3(32'h3af48d04),
	.w4(32'hb9cceb1b),
	.w5(32'hb9c26ebf),
	.w6(32'hba4f62fb),
	.w7(32'hba11396a),
	.w8(32'hba79027f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7eb57d),
	.w1(32'hb8aa3443),
	.w2(32'h38457d22),
	.w3(32'hb698b621),
	.w4(32'h3aa41d43),
	.w5(32'h3a5ae81e),
	.w6(32'h36abc6ec),
	.w7(32'h393c3a6d),
	.w8(32'h36ae54da),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba417b95),
	.w1(32'hba4efe51),
	.w2(32'hbb1b9377),
	.w3(32'hb9caec1d),
	.w4(32'h39fd8c6d),
	.w5(32'hbaea1cde),
	.w6(32'hb9a9eb0d),
	.w7(32'hbb06cbf0),
	.w8(32'hba445d90),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e243f),
	.w1(32'hbb19ba4c),
	.w2(32'hbb61b349),
	.w3(32'hba473ea0),
	.w4(32'hbaff973e),
	.w5(32'hbb4d3d35),
	.w6(32'hbb25809f),
	.w7(32'hbae52948),
	.w8(32'hbad00e29),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f368d),
	.w1(32'hba84d4a8),
	.w2(32'hba5c2d58),
	.w3(32'hbb21470b),
	.w4(32'hb8ce30c0),
	.w5(32'hba8493b5),
	.w6(32'hba3f646b),
	.w7(32'hba4bc830),
	.w8(32'hba42ca4c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ada14),
	.w1(32'h3a7aade5),
	.w2(32'h3b8ceada),
	.w3(32'hbb28544c),
	.w4(32'h3b817b4d),
	.w5(32'h3b68a275),
	.w6(32'h39c0bc2b),
	.w7(32'h3bb2b1c6),
	.w8(32'h3a896fb6),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb766ae3),
	.w1(32'hbad364b2),
	.w2(32'hb8e50aec),
	.w3(32'hbb895971),
	.w4(32'hba14dbb8),
	.w5(32'h3a00f470),
	.w6(32'hba9393e1),
	.w7(32'hb956e079),
	.w8(32'h3afa1df6),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed2258),
	.w1(32'hbb25ea57),
	.w2(32'hba05b3b0),
	.w3(32'hbb3f1359),
	.w4(32'hbb3b8733),
	.w5(32'hbb1cce19),
	.w6(32'hb98241ce),
	.w7(32'h3a422ffe),
	.w8(32'h3a78c383),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ef15d),
	.w1(32'hbb811786),
	.w2(32'hbb887b99),
	.w3(32'hbb22f1d6),
	.w4(32'hbb428a3c),
	.w5(32'hbb80178d),
	.w6(32'hbb7d7c99),
	.w7(32'hbb9c43de),
	.w8(32'hbb916030),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba14d9a),
	.w1(32'hbaa0a937),
	.w2(32'hbb5a7ed0),
	.w3(32'hbb9c01a0),
	.w4(32'h39d7e35e),
	.w5(32'hbb25e2eb),
	.w6(32'hba0c7e46),
	.w7(32'hbb4cf69c),
	.w8(32'hba9db047),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bbc59),
	.w1(32'hbad07596),
	.w2(32'hbb42bb90),
	.w3(32'hba8ce071),
	.w4(32'hb9ff92ad),
	.w5(32'hbad33d02),
	.w6(32'hbad7ed6c),
	.w7(32'hbb3d2a89),
	.w8(32'hbaa391f2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca96c3),
	.w1(32'hbb15a0aa),
	.w2(32'hbb6944b3),
	.w3(32'hba53fe1a),
	.w4(32'hba8c0b98),
	.w5(32'hbb16da5d),
	.w6(32'hbb12da6f),
	.w7(32'hbb577339),
	.w8(32'hbacbb778),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5b394),
	.w1(32'hbaaf1b23),
	.w2(32'hbae4e855),
	.w3(32'hbae2fa8b),
	.w4(32'h3abca62d),
	.w5(32'h39284f10),
	.w6(32'hbaecb5eb),
	.w7(32'hbaf9be7a),
	.w8(32'hba90f3f1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b6b8d),
	.w1(32'h39fa0772),
	.w2(32'h3a828cf1),
	.w3(32'hbadc4b3d),
	.w4(32'hba634f52),
	.w5(32'hb9161209),
	.w6(32'h3b10a4da),
	.w7(32'h3adad448),
	.w8(32'h3bc78a2b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb39c2c),
	.w1(32'h3b15e325),
	.w2(32'h3b0fe564),
	.w3(32'h3bb0022c),
	.w4(32'h3b48bf30),
	.w5(32'h3adc377d),
	.w6(32'h3b48e35b),
	.w7(32'h3af66157),
	.w8(32'h3b997e74),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82e066),
	.w1(32'h3abf1fda),
	.w2(32'h3b5f63e9),
	.w3(32'h3b5c653c),
	.w4(32'h3b0dc89c),
	.w5(32'h3b64ddda),
	.w6(32'h3b156584),
	.w7(32'h3b9e7d55),
	.w8(32'h3ba89700),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96460a),
	.w1(32'hbaaf29ed),
	.w2(32'hbb1e15cc),
	.w3(32'h3b612024),
	.w4(32'hb91fb13c),
	.w5(32'hbaf08657),
	.w6(32'hbacbdd57),
	.w7(32'hbb2395f5),
	.w8(32'hbac82b9f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3b956),
	.w1(32'hbb09f3c7),
	.w2(32'hbb7db8e1),
	.w3(32'hbaf68c89),
	.w4(32'hbb792636),
	.w5(32'hbc05cac5),
	.w6(32'hbb00ff95),
	.w7(32'hbb0ac4d1),
	.w8(32'hbab236d8),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74b29b),
	.w1(32'h3b30c48f),
	.w2(32'h3b943c5d),
	.w3(32'hbc181b47),
	.w4(32'h3aa50eee),
	.w5(32'h3b59b80d),
	.w6(32'h3adacd60),
	.w7(32'h3af1574d),
	.w8(32'h3b912a97),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7c03a),
	.w1(32'h3998da1e),
	.w2(32'h3a588208),
	.w3(32'h3b078751),
	.w4(32'h3b13f8fd),
	.w5(32'h3a0222c1),
	.w6(32'hb8dedb06),
	.w7(32'h3ab7f3f5),
	.w8(32'h3b2b142d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a906260),
	.w1(32'hb955d3f7),
	.w2(32'hb8e19745),
	.w3(32'h3ac5dcb4),
	.w4(32'hb93f3518),
	.w5(32'hb842214e),
	.w6(32'hb963bec0),
	.w7(32'hb84f8bd0),
	.w8(32'hb73cbca1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2720b),
	.w1(32'h39c5a90d),
	.w2(32'h3a4c7fa4),
	.w3(32'h3a85a2b2),
	.w4(32'h3a310339),
	.w5(32'h3a4115e8),
	.w6(32'h3a0560c6),
	.w7(32'hb9618edc),
	.w8(32'h3b021cc4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule