module layer_10_featuremap_461(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381a6852),
	.w1(32'h3737a004),
	.w2(32'h3640da7b),
	.w3(32'h3802f8d4),
	.w4(32'h36aedaee),
	.w5(32'hb5d737a7),
	.w6(32'h382dff56),
	.w7(32'h37eb1b9f),
	.w8(32'h37a7c6fb),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8cb0c),
	.w1(32'h3a0d6d46),
	.w2(32'h3ab0fd6d),
	.w3(32'hba2abd2a),
	.w4(32'h3a7fa90d),
	.w5(32'h3a147013),
	.w6(32'hba4d0f6d),
	.w7(32'hb9f9104a),
	.w8(32'h3a0c9f59),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c791ce),
	.w1(32'h37cf8512),
	.w2(32'h37dbdd18),
	.w3(32'h3785b57b),
	.w4(32'h377727fc),
	.w5(32'h37a767c6),
	.w6(32'h378fdcd1),
	.w7(32'h3755e25b),
	.w8(32'h37d54323),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3780b6c7),
	.w1(32'h3a4c2755),
	.w2(32'h3984a1e8),
	.w3(32'h39fe5d40),
	.w4(32'h3a6c7b3b),
	.w5(32'h3946e7c0),
	.w6(32'h389db42c),
	.w7(32'h3a959440),
	.w8(32'h39a2af5a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3953e92e),
	.w1(32'h39688ac5),
	.w2(32'h3897e5c4),
	.w3(32'h3970f1cc),
	.w4(32'h397cfeaf),
	.w5(32'h390541b6),
	.w6(32'h3967e6ce),
	.w7(32'h398361fa),
	.w8(32'h393f1c83),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bca812),
	.w1(32'hb8249792),
	.w2(32'hb79824b9),
	.w3(32'h36e1b1c9),
	.w4(32'hb681bb04),
	.w5(32'h37bd1f15),
	.w6(32'h37e661ad),
	.w7(32'h37f7f0a9),
	.w8(32'h38735243),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b945c2a),
	.w1(32'h3af3d178),
	.w2(32'hba42bd11),
	.w3(32'h3b70cbb2),
	.w4(32'h3b020600),
	.w5(32'hbade000e),
	.w6(32'h3b8ab0aa),
	.w7(32'h39a74372),
	.w8(32'hbba2921d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19fa12),
	.w1(32'hbb84c9b6),
	.w2(32'hbbcd28a8),
	.w3(32'hbc03dd47),
	.w4(32'hbc171de9),
	.w5(32'hbbbe8e65),
	.w6(32'hbbe494d1),
	.w7(32'hbb8a02a2),
	.w8(32'hbb83fce1),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4c182),
	.w1(32'hba822c27),
	.w2(32'hbaa99a1c),
	.w3(32'hbb0df41b),
	.w4(32'hbab13db1),
	.w5(32'hbae6de28),
	.w6(32'hbb10e015),
	.w7(32'hbafc70af),
	.w8(32'hbb25d2bc),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa640fa),
	.w1(32'hba49e929),
	.w2(32'hbb26ae98),
	.w3(32'hbb34ba01),
	.w4(32'hba62ccc4),
	.w5(32'hbac77728),
	.w6(32'h3b00ae59),
	.w7(32'h3b7d4e31),
	.w8(32'hbad60029),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52ff9f),
	.w1(32'hba3b8510),
	.w2(32'hb90e33e2),
	.w3(32'hb9fb228a),
	.w4(32'hb7ee6f48),
	.w5(32'hb92f5252),
	.w6(32'h39e3f7e5),
	.w7(32'h3a30dc10),
	.w8(32'h3a5fcbf8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1a19a),
	.w1(32'h3bbf8931),
	.w2(32'hb90a40ee),
	.w3(32'h3bf3ee6d),
	.w4(32'h3bd1bce1),
	.w5(32'h3aecf6d7),
	.w6(32'h3be4f6e6),
	.w7(32'h3bd1ec12),
	.w8(32'h39efa230),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0130d2),
	.w1(32'h3b4df5d3),
	.w2(32'h397129c6),
	.w3(32'h3b2afec1),
	.w4(32'h3ac9c4b3),
	.w5(32'hbacdd612),
	.w6(32'h3b798791),
	.w7(32'h3aa50277),
	.w8(32'hbb976877),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92de304),
	.w1(32'h39b454ff),
	.w2(32'h3a5b6aa0),
	.w3(32'hba1adbda),
	.w4(32'hb95d49c7),
	.w5(32'h3ad7e0f7),
	.w6(32'h39eb05cc),
	.w7(32'h3a958cce),
	.w8(32'h3ac65f79),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa1cce),
	.w1(32'h39c66000),
	.w2(32'h39ab9687),
	.w3(32'hb9fd4496),
	.w4(32'h39aea6aa),
	.w5(32'h39b0b848),
	.w6(32'hba1fabef),
	.w7(32'hb988320d),
	.w8(32'hb9461958),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a96dd),
	.w1(32'hbb29c8ab),
	.w2(32'hbb242771),
	.w3(32'hbb335a46),
	.w4(32'hbb08bdf7),
	.w5(32'hbb1bb2cb),
	.w6(32'hbb2cd1ed),
	.w7(32'hbb1dc3a8),
	.w8(32'hbba0ee6a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c811c9),
	.w1(32'h398f5e50),
	.w2(32'h397a1719),
	.w3(32'h3583b259),
	.w4(32'h39ca203b),
	.w5(32'h3a89405b),
	.w6(32'hb8e96a89),
	.w7(32'h3a97525c),
	.w8(32'h3b0b6431),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad91923),
	.w1(32'hbbd483a8),
	.w2(32'hbc06c181),
	.w3(32'hbbccacbf),
	.w4(32'hbc121907),
	.w5(32'hbc0991b7),
	.w6(32'hba9427bc),
	.w7(32'hbbd736f8),
	.w8(32'hbc173643),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39585696),
	.w1(32'hbaa3e5d9),
	.w2(32'hbb47d55b),
	.w3(32'hbaaef9b9),
	.w4(32'hbb4f11f1),
	.w5(32'hbb83147a),
	.w6(32'h3a04e379),
	.w7(32'hbb2f1c75),
	.w8(32'hbbaf2a26),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb782b3be),
	.w1(32'h38a3bedd),
	.w2(32'h37d934d4),
	.w3(32'hb886e3eb),
	.w4(32'h38bd28ce),
	.w5(32'h384adb25),
	.w6(32'hb683f1f6),
	.w7(32'h38e0934e),
	.w8(32'hb7844ac6),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384228ab),
	.w1(32'hb88b75ab),
	.w2(32'hb6ff7538),
	.w3(32'h389986f4),
	.w4(32'hb5acce19),
	.w5(32'hb6564cab),
	.w6(32'h3807d3ae),
	.w7(32'hb76562cc),
	.w8(32'h39055210),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54fb04),
	.w1(32'h3a3c42b1),
	.w2(32'h3a344335),
	.w3(32'h3ac3c938),
	.w4(32'h3ac3d263),
	.w5(32'h3ad9bc70),
	.w6(32'h3a9d741a),
	.w7(32'h3aa1a586),
	.w8(32'h3aded1a8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e4688),
	.w1(32'hbb8fd84f),
	.w2(32'hbc609ce4),
	.w3(32'hbb704e6e),
	.w4(32'hbb96569d),
	.w5(32'hbc311af9),
	.w6(32'hbbb6702b),
	.w7(32'hbbf8d5fe),
	.w8(32'hbc6ceb71),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912ca92),
	.w1(32'h36a2feaa),
	.w2(32'h39f91cbe),
	.w3(32'hb93129fe),
	.w4(32'h3a974309),
	.w5(32'h3950ca12),
	.w6(32'h3b015141),
	.w7(32'h3b1fd587),
	.w8(32'h392c6454),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d42b07),
	.w1(32'h3a067c8f),
	.w2(32'h3a8d7108),
	.w3(32'h3a43e165),
	.w4(32'h3b51fc9c),
	.w5(32'h3b73b370),
	.w6(32'hbaa3a0ac),
	.w7(32'hbae66c24),
	.w8(32'h3aab4062),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41244a),
	.w1(32'h3a20c5df),
	.w2(32'h3a49d376),
	.w3(32'hba86df14),
	.w4(32'h3923f894),
	.w5(32'h38ff1bee),
	.w6(32'hba354111),
	.w7(32'h39e7a1e3),
	.w8(32'h398bc92b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974c3fd),
	.w1(32'h38717391),
	.w2(32'h39566698),
	.w3(32'h3932b760),
	.w4(32'h3851b164),
	.w5(32'h398206fa),
	.w6(32'h3978a1ac),
	.w7(32'h390b7b65),
	.w8(32'h39ab2949),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cc444),
	.w1(32'h3b4add08),
	.w2(32'h3a99dee8),
	.w3(32'h3b10c26d),
	.w4(32'h3b54e572),
	.w5(32'h3b11eb5f),
	.w6(32'h3b0646d0),
	.w7(32'hba394be9),
	.w8(32'h39562632),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b540e19),
	.w1(32'h3ab68ed9),
	.w2(32'h3a529b53),
	.w3(32'h3b4f4fd0),
	.w4(32'h3b2842b1),
	.w5(32'h3afc2e7c),
	.w6(32'h3b589b4c),
	.w7(32'h3b87683d),
	.w8(32'h3b98acce),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8270d3),
	.w1(32'h3b442cca),
	.w2(32'h3b99196a),
	.w3(32'hbb13920a),
	.w4(32'h3b1fb0fe),
	.w5(32'h3b262eac),
	.w6(32'hb9847de3),
	.w7(32'h3a2e114f),
	.w8(32'h3ae6cc52),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e01c2b),
	.w1(32'h38849d14),
	.w2(32'h3903cf80),
	.w3(32'h390bb32f),
	.w4(32'h3915fc39),
	.w5(32'h395c6d5c),
	.w6(32'h395e9d2c),
	.w7(32'h39781704),
	.w8(32'h399dc59b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6f464),
	.w1(32'hb980d585),
	.w2(32'h3a00607c),
	.w3(32'hb966dbd9),
	.w4(32'h3840406a),
	.w5(32'h3a774f09),
	.w6(32'hb8c98701),
	.w7(32'h3a02aff6),
	.w8(32'h3aa586ac),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e2831),
	.w1(32'h3a041279),
	.w2(32'hb8cfe466),
	.w3(32'hb9ddb7fc),
	.w4(32'h39d9cc97),
	.w5(32'hb89af6e3),
	.w6(32'h39e7247c),
	.w7(32'h3a8c1643),
	.w8(32'h38f38669),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb268835),
	.w1(32'hba03c523),
	.w2(32'hb78f5b15),
	.w3(32'hbaad29b3),
	.w4(32'h396008f7),
	.w5(32'hb9759054),
	.w6(32'hbad6fb96),
	.w7(32'hba92eae4),
	.w8(32'hba6ca222),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bb885),
	.w1(32'hb7610741),
	.w2(32'hb9d2f554),
	.w3(32'h395335f8),
	.w4(32'h39148cc1),
	.w5(32'h3833a4f4),
	.w6(32'h3a505f85),
	.w7(32'hb8dbab09),
	.w8(32'hb92266aa),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee3922),
	.w1(32'h3acddffa),
	.w2(32'h3793cb86),
	.w3(32'h3a5e1e3c),
	.w4(32'h3aca3fd3),
	.w5(32'hb9fc7a44),
	.w6(32'h3ac13962),
	.w7(32'h3b0b910a),
	.w8(32'hba9e3aae),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb87cd7),
	.w1(32'h3c053b94),
	.w2(32'hbbc6ef0b),
	.w3(32'hbb9c3811),
	.w4(32'h3b864b26),
	.w5(32'h3b4f618a),
	.w6(32'hba92839d),
	.w7(32'h3c25c764),
	.w8(32'h3ac09881),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f9ef),
	.w1(32'h3ba4ef63),
	.w2(32'h3c0192d8),
	.w3(32'h3ba2be22),
	.w4(32'h3c22fac6),
	.w5(32'h3c3e3554),
	.w6(32'hbad2d454),
	.w7(32'h3babf287),
	.w8(32'h3c27b8ee),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82c13f),
	.w1(32'h3bf14db1),
	.w2(32'h3bde1370),
	.w3(32'h3c1e10cf),
	.w4(32'h3c14a7f1),
	.w5(32'h3b82b78f),
	.w6(32'h3be36dbf),
	.w7(32'h3aa898c4),
	.w8(32'h3b65e265),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d9345),
	.w1(32'h3ac01dc6),
	.w2(32'h3af304b5),
	.w3(32'h39f0ee53),
	.w4(32'h3ae72e22),
	.w5(32'h3b18ca32),
	.w6(32'hb93125b8),
	.w7(32'h3a640936),
	.w8(32'h3abe61e3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89a47a),
	.w1(32'hba33b369),
	.w2(32'hba152f40),
	.w3(32'hba7a1e0c),
	.w4(32'hba46ba05),
	.w5(32'hb9df0156),
	.w6(32'hb9da72b3),
	.w7(32'hb99c6c45),
	.w8(32'hb71737cd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7db85),
	.w1(32'hb907d914),
	.w2(32'hb96f8085),
	.w3(32'h3a329eef),
	.w4(32'hb90a0381),
	.w5(32'hb9aaf7e2),
	.w6(32'h3a35e89e),
	.w7(32'h3889e965),
	.w8(32'hb7ed4468),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a942b64),
	.w1(32'h3b5552f6),
	.w2(32'h3b3f7df8),
	.w3(32'h3a2c664a),
	.w4(32'h3b258865),
	.w5(32'h3b311b10),
	.w6(32'h38c69226),
	.w7(32'h3b27d445),
	.w8(32'h3b0b5a78),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385bc682),
	.w1(32'h3aca5b3b),
	.w2(32'hbb1aabe9),
	.w3(32'hbaf33691),
	.w4(32'hb6dff0f8),
	.w5(32'hbbf3dc2c),
	.w6(32'h3924f962),
	.w7(32'hbae2a2e2),
	.w8(32'hbc05eee5),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f64b0),
	.w1(32'h3a123267),
	.w2(32'h3aa22e7c),
	.w3(32'hbb223d3e),
	.w4(32'h3ac9c24d),
	.w5(32'h3a4e84de),
	.w6(32'hba9a5f45),
	.w7(32'h3ac6d905),
	.w8(32'hb9a8c591),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25ba00),
	.w1(32'h3983ac8a),
	.w2(32'h3a818210),
	.w3(32'hb94ed877),
	.w4(32'h3b01e09c),
	.w5(32'hbabdd928),
	.w6(32'h3a235d49),
	.w7(32'h3aad64fb),
	.w8(32'hbb1562e4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce19b8),
	.w1(32'hbb0b7145),
	.w2(32'hbb292cd4),
	.w3(32'hbb9c2005),
	.w4(32'hbad7af3b),
	.w5(32'hbb5cf6f8),
	.w6(32'hbbac787b),
	.w7(32'hbb815447),
	.w8(32'hbbc06961),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e5f63),
	.w1(32'hbb383315),
	.w2(32'hbc2471c6),
	.w3(32'hba9f03b1),
	.w4(32'hbbefe47c),
	.w5(32'hbc25eb33),
	.w6(32'h39f3563f),
	.w7(32'hbb5b06ac),
	.w8(32'hbc46f381),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c83d2),
	.w1(32'h3a2b1d13),
	.w2(32'hb9e2dc28),
	.w3(32'h390b4d57),
	.w4(32'h3a881241),
	.w5(32'hb961e72e),
	.w6(32'h3984b2ae),
	.w7(32'h39af5383),
	.w8(32'hba947555),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9822894),
	.w1(32'hb91e9b15),
	.w2(32'hbb082c4a),
	.w3(32'hb9b5ac6c),
	.w4(32'hba9c45e8),
	.w5(32'hbb36bcfc),
	.w6(32'hba9aebd2),
	.w7(32'hbb2c471b),
	.w8(32'hbb96ad31),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b294cbc),
	.w1(32'h3b09f3d7),
	.w2(32'h3a1b0c54),
	.w3(32'h3b48e253),
	.w4(32'h3b1eea2d),
	.w5(32'h3a0865c4),
	.w6(32'h3b01eecf),
	.w7(32'h3ad4b861),
	.w8(32'h3a0548c4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabb3ad),
	.w1(32'hbaaeba17),
	.w2(32'hbb11bf21),
	.w3(32'hbaca4c12),
	.w4(32'h3a3c7cfa),
	.w5(32'h382bcff0),
	.w6(32'hba2a0536),
	.w7(32'h3919384f),
	.w8(32'hba45a6d6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c2d9d),
	.w1(32'hba63312d),
	.w2(32'hbac8355d),
	.w3(32'hb9bb7021),
	.w4(32'hba334f8f),
	.w5(32'hbac9a7cf),
	.w6(32'hba50a016),
	.w7(32'hba2ab443),
	.w8(32'hbaa6afb6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2880a8),
	.w1(32'hbb863b7f),
	.w2(32'hbbfe75ab),
	.w3(32'hbb39d5d7),
	.w4(32'hbbd57250),
	.w5(32'hbbc9f3e3),
	.w6(32'h39ed507f),
	.w7(32'hbb5e39a5),
	.w8(32'hbc0f5213),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6dd93),
	.w1(32'hba3d86a5),
	.w2(32'hba9242d7),
	.w3(32'h3a3d61c6),
	.w4(32'hb9977f44),
	.w5(32'hba64f62d),
	.w6(32'h3a8a1cc1),
	.w7(32'h39727743),
	.w8(32'hba20fdd8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3721a3e2),
	.w1(32'h39236c08),
	.w2(32'h3803f8a1),
	.w3(32'h36a04c7b),
	.w4(32'h39266db2),
	.w5(32'h37a5b043),
	.w6(32'hb8a54451),
	.w7(32'h3884f2f4),
	.w8(32'h371d0152),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6104b49),
	.w1(32'hb7bf96a8),
	.w2(32'hb6a3e4f8),
	.w3(32'h36e6e1e4),
	.w4(32'hb77c5908),
	.w5(32'hb61946fc),
	.w6(32'h377309ab),
	.w7(32'h37875391),
	.w8(32'h37d38f3e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396432c3),
	.w1(32'h36c3f969),
	.w2(32'h393f43e4),
	.w3(32'h399683c5),
	.w4(32'hb8c67f52),
	.w5(32'h394e5728),
	.w6(32'h39231bdb),
	.w7(32'hb981d7ad),
	.w8(32'h39660514),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f8389),
	.w1(32'h3a8a1759),
	.w2(32'h3aa3f2f3),
	.w3(32'h3a1f64bc),
	.w4(32'h3ab29f3a),
	.w5(32'h3a8b5ec1),
	.w6(32'h396c4de1),
	.w7(32'h3a852268),
	.w8(32'h3a0abd4f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a11ae8),
	.w1(32'h3a87673e),
	.w2(32'h3a297ca6),
	.w3(32'h38d95cda),
	.w4(32'h3989767e),
	.w5(32'h39bfb61d),
	.w6(32'h392b949e),
	.w7(32'h37b76d0e),
	.w8(32'h39319b67),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f38ef),
	.w1(32'hbafc8e3d),
	.w2(32'hbb53a276),
	.w3(32'hb99b098b),
	.w4(32'hbac37202),
	.w5(32'hbb56dbe2),
	.w6(32'h3aa08549),
	.w7(32'hbaaafcf3),
	.w8(32'hbb8dc854),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bedc9),
	.w1(32'hbb92ae7e),
	.w2(32'hbac0e930),
	.w3(32'hbb9d6c1a),
	.w4(32'hbb726061),
	.w5(32'hbb297122),
	.w6(32'hbb438cbe),
	.w7(32'hbb93fcfc),
	.w8(32'hbb660035),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb938c109),
	.w1(32'hb8444e4f),
	.w2(32'h386bac95),
	.w3(32'hb8432cb5),
	.w4(32'h38309e41),
	.w5(32'h3945e58f),
	.w6(32'h3870de50),
	.w7(32'h38b89d91),
	.w8(32'h3953fa7f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c7517c),
	.w1(32'hb7402433),
	.w2(32'h380e2161),
	.w3(32'hb8086cb6),
	.w4(32'hb7cf618b),
	.w5(32'h37e98250),
	.w6(32'hb7a4ae1d),
	.w7(32'hb726302e),
	.w8(32'h3828a9ec),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398de309),
	.w1(32'h38db1e48),
	.w2(32'h39a6eb13),
	.w3(32'h3987bf06),
	.w4(32'h39050856),
	.w5(32'h395a9c9a),
	.w6(32'h3930ff07),
	.w7(32'h3940bb1f),
	.w8(32'h399259eb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ef02fd),
	.w1(32'hb80dbe96),
	.w2(32'h38a4ff35),
	.w3(32'hb736c7d3),
	.w4(32'h3741fa14),
	.w5(32'h38f97bec),
	.w6(32'h381f58e3),
	.w7(32'h387c5435),
	.w8(32'h393f84a5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b853c5a),
	.w1(32'hbb26d829),
	.w2(32'hbb904f28),
	.w3(32'h3a496277),
	.w4(32'hba7d4220),
	.w5(32'h3ac44f4b),
	.w6(32'h3b348cce),
	.w7(32'hbb752ea3),
	.w8(32'hbba1de2f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93afd1d),
	.w1(32'hbb0ecb24),
	.w2(32'hbb4e78d1),
	.w3(32'h3b31dad1),
	.w4(32'h3ae0436e),
	.w5(32'hbbb311af),
	.w6(32'h3b2411da),
	.w7(32'h3a77577f),
	.w8(32'hbb7a1687),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba976bff),
	.w1(32'hbb9d5d3e),
	.w2(32'hbbadeb14),
	.w3(32'hbab9ca02),
	.w4(32'hbaef6fe4),
	.w5(32'hbba50ea0),
	.w6(32'hbb081f27),
	.w7(32'hbba18a9a),
	.w8(32'hbc004f9c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb793248),
	.w1(32'hbbac07b5),
	.w2(32'h3b2f28ae),
	.w3(32'h3b226fe5),
	.w4(32'h3b63726e),
	.w5(32'h3bfed312),
	.w6(32'hb9cba6c2),
	.w7(32'hbb366881),
	.w8(32'h3b466ab2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6f565),
	.w1(32'hbb1eeba1),
	.w2(32'hbaabff9b),
	.w3(32'hbaa69cb1),
	.w4(32'hbbc0be21),
	.w5(32'hbbb577c2),
	.w6(32'hbb31c77f),
	.w7(32'hbb7b1226),
	.w8(32'hbb7ed2e3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa3cc0),
	.w1(32'hbb34a75d),
	.w2(32'hbb4e3ba9),
	.w3(32'hbb83dbe8),
	.w4(32'hb9f2ae8b),
	.w5(32'h3b2635d6),
	.w6(32'hbba5ff64),
	.w7(32'hbae22998),
	.w8(32'hbbb0e191),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dadfe),
	.w1(32'hb8b1ee66),
	.w2(32'h3a8fbaea),
	.w3(32'hbb99e90f),
	.w4(32'hbad683b9),
	.w5(32'h3b2c85e1),
	.w6(32'hbb8617ae),
	.w7(32'h3a1712f3),
	.w8(32'h3bf9ff9b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdeb9eb),
	.w1(32'h3b03bc44),
	.w2(32'hbb7ad696),
	.w3(32'h3bcd7479),
	.w4(32'hbadbebf9),
	.w5(32'hbb6940ea),
	.w6(32'h3b2870d6),
	.w7(32'hbb124bfd),
	.w8(32'hbb5e9f25),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12aa1c),
	.w1(32'h3b99b7ac),
	.w2(32'h3baf5a6b),
	.w3(32'h3b5bce9c),
	.w4(32'h3a2f24df),
	.w5(32'hbb15bec1),
	.w6(32'h39a6bd53),
	.w7(32'h39899c8c),
	.w8(32'h3b40385b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d1cee),
	.w1(32'hbb39e081),
	.w2(32'hbbab37d4),
	.w3(32'hbba6b3e1),
	.w4(32'hbbab8e12),
	.w5(32'hbac93cbf),
	.w6(32'h3a80ba16),
	.w7(32'hb9fdbb38),
	.w8(32'hbb2a84a8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36548e),
	.w1(32'hbbb54c68),
	.w2(32'hbc4e8d8d),
	.w3(32'hbac4ff2d),
	.w4(32'hbb93798d),
	.w5(32'hbc0be6bd),
	.w6(32'hbb7bbd93),
	.w7(32'hbb8f6cc1),
	.w8(32'hbc3c3565),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb3eb3),
	.w1(32'h380e50df),
	.w2(32'h3bbe950e),
	.w3(32'hbb4d8a2b),
	.w4(32'hbb418cd4),
	.w5(32'hbb889f76),
	.w6(32'h3a9f2bd4),
	.w7(32'hbb2deb5f),
	.w8(32'hbb77f916),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cbeb7),
	.w1(32'hbb8a66cf),
	.w2(32'h3b050e2a),
	.w3(32'hbaef0aac),
	.w4(32'hbb6ef191),
	.w5(32'h3ab0a5e3),
	.w6(32'hbb80092d),
	.w7(32'hb8e967cc),
	.w8(32'hb91d8dd7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b546a93),
	.w1(32'hba1c42ef),
	.w2(32'hbb86f7b6),
	.w3(32'h39fdfa91),
	.w4(32'h37e2144b),
	.w5(32'hbaf02816),
	.w6(32'h3b882c40),
	.w7(32'h395f6199),
	.w8(32'hbb851e85),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad521f9),
	.w1(32'hba1a61f0),
	.w2(32'h3af71cd9),
	.w3(32'hbb9b1daf),
	.w4(32'h3b008bc4),
	.w5(32'h3b23aa86),
	.w6(32'hbb8d4e1a),
	.w7(32'h3af9cab8),
	.w8(32'h3b956257),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96d4ae),
	.w1(32'hbbbbbc0a),
	.w2(32'hbbec821b),
	.w3(32'h3bbd8295),
	.w4(32'hbbbd2aad),
	.w5(32'hbbec7a23),
	.w6(32'h3c04deb2),
	.w7(32'hbbb0f296),
	.w8(32'hbc169c35),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb409d89),
	.w1(32'h3aaf7fd6),
	.w2(32'h3ad6f02d),
	.w3(32'h3a371787),
	.w4(32'hba82bbb0),
	.w5(32'hb8ef5fc9),
	.w6(32'hba8e6cb7),
	.w7(32'h388b9f7b),
	.w8(32'h3948bf65),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcd0a3),
	.w1(32'hbaecaa96),
	.w2(32'h3b38ff1a),
	.w3(32'hba78775d),
	.w4(32'hbb2ed1c9),
	.w5(32'h39b5c8f3),
	.w6(32'h3ad449e7),
	.w7(32'hbb59613b),
	.w8(32'hbad6122d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3860f4d8),
	.w1(32'hbb43c993),
	.w2(32'hbb1aaedf),
	.w3(32'h3a3d4910),
	.w4(32'hbb1d5c3e),
	.w5(32'hbb82a9e9),
	.w6(32'h3a784daf),
	.w7(32'hbb9cec00),
	.w8(32'hbb564774),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea81b6),
	.w1(32'hbbf16cdc),
	.w2(32'hbb521b66),
	.w3(32'hba280164),
	.w4(32'h39e2c977),
	.w5(32'hbaf002bf),
	.w6(32'hbb440827),
	.w7(32'hbb2e89b1),
	.w8(32'hbbd3ef31),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f3f38),
	.w1(32'h394272a9),
	.w2(32'h3bd59f5a),
	.w3(32'hbb7e6281),
	.w4(32'hbaac5286),
	.w5(32'h3c0c6458),
	.w6(32'hbbcbc5eb),
	.w7(32'hbb8406b7),
	.w8(32'hbb23db92),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b4217),
	.w1(32'hb9f9c54c),
	.w2(32'hbb13dcf3),
	.w3(32'hbabfe7a8),
	.w4(32'h3a2726d5),
	.w5(32'h3a9d7819),
	.w6(32'hba8f9978),
	.w7(32'hba04f654),
	.w8(32'h3ba60220),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c0e57),
	.w1(32'hbbc9b741),
	.w2(32'hbb78e524),
	.w3(32'h3ab5a1b1),
	.w4(32'h395041ae),
	.w5(32'hbb1ab6bb),
	.w6(32'h3b7475fd),
	.w7(32'h3a4e8218),
	.w8(32'hba563a17),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c9192),
	.w1(32'hbb59fe5b),
	.w2(32'hbbae05c7),
	.w3(32'hbc175dd9),
	.w4(32'hbc26289f),
	.w5(32'hbb8358e2),
	.w6(32'hbbb907e9),
	.w7(32'hbb8fbc40),
	.w8(32'hbc152988),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a0ce3),
	.w1(32'hbadff46b),
	.w2(32'hbaebb081),
	.w3(32'h3af18792),
	.w4(32'hbad856a6),
	.w5(32'h3b64148e),
	.w6(32'h3a173df8),
	.w7(32'hbb3e89f1),
	.w8(32'h3a89ecb7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03a080),
	.w1(32'h3bb2fdac),
	.w2(32'hba6cfeda),
	.w3(32'hbb3f613d),
	.w4(32'h3c03e97f),
	.w5(32'h3a9d3d2b),
	.w6(32'hba91890b),
	.w7(32'h3c005560),
	.w8(32'h3ab9554d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b620896),
	.w1(32'h3af90f67),
	.w2(32'h3b1141de),
	.w3(32'h3b375222),
	.w4(32'h3b9bedeb),
	.w5(32'h3bdd7a26),
	.w6(32'h3b557829),
	.w7(32'h3bc4cdeb),
	.w8(32'h3b9fbdf3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50a7a3),
	.w1(32'hbbf1ae73),
	.w2(32'hbc118cdc),
	.w3(32'hb925e25f),
	.w4(32'hbb1020b9),
	.w5(32'hbaed0a40),
	.w6(32'h3ab86fc1),
	.w7(32'hbb9aad6e),
	.w8(32'hbbccb2d9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9e768),
	.w1(32'hba9d2237),
	.w2(32'hba5b4ed7),
	.w3(32'h39b20aa0),
	.w4(32'hbaeb44b1),
	.w5(32'hbb9c8085),
	.w6(32'hb9c5c4b3),
	.w7(32'h3b28c2ea),
	.w8(32'hb91a7098),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c941be),
	.w1(32'h3b325154),
	.w2(32'h3a9e0bb9),
	.w3(32'hbbb648bd),
	.w4(32'h3ab473de),
	.w5(32'h3ad79393),
	.w6(32'hbaf8164f),
	.w7(32'hbb6bdb99),
	.w8(32'hbb3e895e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a1344),
	.w1(32'h3acbdb45),
	.w2(32'h3a0967d1),
	.w3(32'hbabaf6a4),
	.w4(32'h39285390),
	.w5(32'hbb125fb6),
	.w6(32'hbb859b1f),
	.w7(32'hbb0c0bd0),
	.w8(32'hbbb7a42a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71d5e1),
	.w1(32'h3c026207),
	.w2(32'hbad97b3a),
	.w3(32'h3b21aa53),
	.w4(32'h3b994db3),
	.w5(32'hbb71a0d9),
	.w6(32'hbb1d989d),
	.w7(32'h3acbac7a),
	.w8(32'hbc18572c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a73db8),
	.w1(32'hbaf950ee),
	.w2(32'hbb80ba6e),
	.w3(32'h3a6be95a),
	.w4(32'hb9a880e0),
	.w5(32'hbaa34fd4),
	.w6(32'h3af557c1),
	.w7(32'hbb968f4b),
	.w8(32'hbc19be82),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad51aa8),
	.w1(32'h3c307c30),
	.w2(32'hbb4dbdff),
	.w3(32'hbc4ed684),
	.w4(32'h3ab56208),
	.w5(32'hbb33aed6),
	.w6(32'hbbbdbdda),
	.w7(32'h3c39ad42),
	.w8(32'h3c212589),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f4cfb),
	.w1(32'h3c20fd04),
	.w2(32'h3c1ea0d1),
	.w3(32'hbb1bc8bf),
	.w4(32'h3c363f57),
	.w5(32'h3c5a80a2),
	.w6(32'hbb8c0393),
	.w7(32'hbb409042),
	.w8(32'hba15ebb5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90fef96),
	.w1(32'hbab37528),
	.w2(32'h3778ef70),
	.w3(32'h3af5963b),
	.w4(32'hbb617ebe),
	.w5(32'hbb7d7f9b),
	.w6(32'hbb3e6ce1),
	.w7(32'hbb67cb4d),
	.w8(32'hbbad08ce),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba46d05),
	.w1(32'h3bca8e9b),
	.w2(32'hba8a6607),
	.w3(32'hbb9e04b4),
	.w4(32'h3b8408d0),
	.w5(32'h3a1712e2),
	.w6(32'hbb914741),
	.w7(32'h3bae5cf2),
	.w8(32'hbb2650b0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c182d2f),
	.w1(32'h3c0462b6),
	.w2(32'h3be162eb),
	.w3(32'h3af42187),
	.w4(32'h3a789518),
	.w5(32'hbae378a1),
	.w6(32'hba96709b),
	.w7(32'hbb82aae1),
	.w8(32'hbbc9e643),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ac8c0),
	.w1(32'hbbf378e9),
	.w2(32'hbc639485),
	.w3(32'hbc55d582),
	.w4(32'hbc0cf03c),
	.w5(32'hbb410076),
	.w6(32'hbc5732cc),
	.w7(32'hb9ca3a2e),
	.w8(32'hbb3d6c0d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52ee9c),
	.w1(32'hbaa0b59a),
	.w2(32'h39af5c9a),
	.w3(32'h3bde7182),
	.w4(32'h3aefe5e2),
	.w5(32'hbade4016),
	.w6(32'h3b60e0f5),
	.w7(32'h3b405494),
	.w8(32'hbb492678),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d2ea5),
	.w1(32'h3aa3699c),
	.w2(32'h3afcf31c),
	.w3(32'hba986fda),
	.w4(32'h380afd55),
	.w5(32'h3ad48506),
	.w6(32'hbadc8ae3),
	.w7(32'hba4dfda4),
	.w8(32'h3b16b7b5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c114fa),
	.w1(32'hbb884910),
	.w2(32'hbb739bce),
	.w3(32'h3b40cd87),
	.w4(32'hb9d73cf0),
	.w5(32'h3a403586),
	.w6(32'h3a3bc8e0),
	.w7(32'h3b28cd1f),
	.w8(32'h39dfe08b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba46156),
	.w1(32'h3bb76202),
	.w2(32'h3ac9d43d),
	.w3(32'h3b9517f0),
	.w4(32'hbac63464),
	.w5(32'hbbad91b2),
	.w6(32'h3a872f2e),
	.w7(32'hbbbe2836),
	.w8(32'hbbf71bf0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98d8d5),
	.w1(32'h3bc462ae),
	.w2(32'h3ac15f71),
	.w3(32'hba444ba2),
	.w4(32'h3b623a9d),
	.w5(32'h39a20ffe),
	.w6(32'h3a9e73f7),
	.w7(32'hbb364473),
	.w8(32'hbbadffe1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed3142),
	.w1(32'hbaaa533e),
	.w2(32'hbb2161fe),
	.w3(32'h3b6c8f55),
	.w4(32'h3b106117),
	.w5(32'h3a433093),
	.w6(32'hbaf9b6e9),
	.w7(32'hbb8261c6),
	.w8(32'hba47cd34),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1ed85),
	.w1(32'h393e3850),
	.w2(32'hb978e577),
	.w3(32'hbb7cec09),
	.w4(32'hbb883140),
	.w5(32'hbad811cb),
	.w6(32'hbbd01174),
	.w7(32'hbb621ee9),
	.w8(32'hbbcb38b8),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18a44c),
	.w1(32'h3bd0ae34),
	.w2(32'h395db34b),
	.w3(32'hbb8031a7),
	.w4(32'h3baebbd2),
	.w5(32'h3ac2d66a),
	.w6(32'hbb8227b6),
	.w7(32'h3c1cda01),
	.w8(32'h3bd11bbb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d287a),
	.w1(32'hbb84c1df),
	.w2(32'hbb8c77a4),
	.w3(32'hba600f89),
	.w4(32'hb9eb6910),
	.w5(32'h3b0fb8ee),
	.w6(32'hba83f6d1),
	.w7(32'hba253a36),
	.w8(32'hbb86ad16),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a948b),
	.w1(32'h3b81e5a0),
	.w2(32'h3bb77f7d),
	.w3(32'h3b8011b2),
	.w4(32'h3b8bc620),
	.w5(32'h3c1d0695),
	.w6(32'h3b2df6f3),
	.w7(32'h3bb7f6a1),
	.w8(32'h3b294a14),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00b557),
	.w1(32'hbbb1dfd5),
	.w2(32'hbb8dcbf5),
	.w3(32'hbabea2fb),
	.w4(32'hbb968027),
	.w5(32'hbb9459f7),
	.w6(32'h3b8461c5),
	.w7(32'hbb7f9ef8),
	.w8(32'hbb8874e0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d77a6),
	.w1(32'h3b45aa8d),
	.w2(32'hba6895a2),
	.w3(32'hbb27e483),
	.w4(32'h3b2b076e),
	.w5(32'h39bce09b),
	.w6(32'hbaf6e9a0),
	.w7(32'hbb9e54c3),
	.w8(32'hbb851295),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21c130),
	.w1(32'hbb60d72c),
	.w2(32'hbb86202f),
	.w3(32'h3b973ac8),
	.w4(32'h3b04eaad),
	.w5(32'h3ad1d8cf),
	.w6(32'h3ad7d388),
	.w7(32'h3a597bd7),
	.w8(32'hbb99b8a0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba657e7),
	.w1(32'h3ab3b5d3),
	.w2(32'h3abd36a3),
	.w3(32'hbb220aec),
	.w4(32'hba05d6a7),
	.w5(32'hb9b1ca74),
	.w6(32'hbb9dc640),
	.w7(32'hbb31f193),
	.w8(32'h39f109a1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27a69e),
	.w1(32'h38181bf8),
	.w2(32'h3aa290c9),
	.w3(32'h3ba8e901),
	.w4(32'hba844f10),
	.w5(32'hbb22b925),
	.w6(32'h3b1b5a99),
	.w7(32'h39f89355),
	.w8(32'hbb706575),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05d590),
	.w1(32'hbb979078),
	.w2(32'hb8e126cc),
	.w3(32'hbbad4b37),
	.w4(32'hba053abb),
	.w5(32'h39bedfe2),
	.w6(32'hbb9241b7),
	.w7(32'hbb1dbc22),
	.w8(32'h3b84b028),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f9c39),
	.w1(32'hbbc47248),
	.w2(32'hbbf86a39),
	.w3(32'h3b7cd30c),
	.w4(32'hbadc24cb),
	.w5(32'hbbe9208c),
	.w6(32'h3bcc132c),
	.w7(32'hbaadc3b1),
	.w8(32'hbb66466e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ed9fb),
	.w1(32'h3a0cca5c),
	.w2(32'h3a8666bc),
	.w3(32'hbbbb4758),
	.w4(32'hba94835f),
	.w5(32'hbb57935c),
	.w6(32'hbb9fed15),
	.w7(32'hbbc8c16f),
	.w8(32'hbb03fa60),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2317ca),
	.w1(32'h3a9c364d),
	.w2(32'hbb959cc5),
	.w3(32'hba639c4c),
	.w4(32'h3b48c5e6),
	.w5(32'hbb83b8c2),
	.w6(32'h3a4e6525),
	.w7(32'h3aaa74a0),
	.w8(32'hb905197e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6c5d6),
	.w1(32'h39226536),
	.w2(32'hbadcc96b),
	.w3(32'h3b41702c),
	.w4(32'h3ad0cbb3),
	.w5(32'hbb58ffeb),
	.w6(32'h3b2ed380),
	.w7(32'hbb6f2d4f),
	.w8(32'hbb5f8176),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b6552),
	.w1(32'hb93924d3),
	.w2(32'hb9d0be74),
	.w3(32'hbb7940d5),
	.w4(32'h3b8bf9f3),
	.w5(32'h3bb1027e),
	.w6(32'hbb6937e8),
	.w7(32'h3a29b7a6),
	.w8(32'hb9c68834),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c62f5),
	.w1(32'hba599032),
	.w2(32'hbb75e77c),
	.w3(32'h3b546ddf),
	.w4(32'h3abf19de),
	.w5(32'hba57b27e),
	.w6(32'h3aac9d09),
	.w7(32'h3afb12e5),
	.w8(32'hb9c429ad),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e7302),
	.w1(32'hbbde35d9),
	.w2(32'hbbae4fdb),
	.w3(32'hbb85f5e7),
	.w4(32'hbb206299),
	.w5(32'hbc1ec2be),
	.w6(32'hbb078ca6),
	.w7(32'hba99af7d),
	.w8(32'hbbb92b24),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd1dd5),
	.w1(32'hbacf92df),
	.w2(32'hbb8d132f),
	.w3(32'hbb58a05a),
	.w4(32'h3982248b),
	.w5(32'h39274423),
	.w6(32'h3a2d45f2),
	.w7(32'h3af7f9aa),
	.w8(32'hbb2b8ab8),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c73c8),
	.w1(32'hba472187),
	.w2(32'h39260d47),
	.w3(32'hbb4158c8),
	.w4(32'hba297ec5),
	.w5(32'h3a3cd5ef),
	.w6(32'h39fe2d81),
	.w7(32'hb9b2cd74),
	.w8(32'hbb3149bd),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dfb89),
	.w1(32'hbab3e202),
	.w2(32'hba903968),
	.w3(32'hbb830962),
	.w4(32'h3a9f6c1b),
	.w5(32'h3b526640),
	.w6(32'hbb54342c),
	.w7(32'hbb7a0fc6),
	.w8(32'hbb9215ba),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b82960),
	.w1(32'hbbb74051),
	.w2(32'h3aa05575),
	.w3(32'h3b96ffa3),
	.w4(32'hba918dbc),
	.w5(32'h3c0ac43b),
	.w6(32'h399533ec),
	.w7(32'hbb42983e),
	.w8(32'hbb87bbc7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8209b0),
	.w1(32'h3a4a139f),
	.w2(32'hbb6a43d3),
	.w3(32'hbbdb2188),
	.w4(32'h3b29919e),
	.w5(32'hbaf9a7d9),
	.w6(32'hbc0270bf),
	.w7(32'h3aa7b9a0),
	.w8(32'hbab11ea2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a901f),
	.w1(32'h3a84d885),
	.w2(32'hbb20b556),
	.w3(32'hbb272219),
	.w4(32'h3ae0fd79),
	.w5(32'hb88ca2c5),
	.w6(32'hba8de503),
	.w7(32'h3a6719bd),
	.w8(32'hb9a5d39c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7cdbe),
	.w1(32'hbb524ec6),
	.w2(32'hbbdc2033),
	.w3(32'hbb77668a),
	.w4(32'hbb5f34fb),
	.w5(32'hbbcd9971),
	.w6(32'h3b2a8fc4),
	.w7(32'hbb402bb7),
	.w8(32'hbc06cde8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba589c11),
	.w1(32'h3a2993b8),
	.w2(32'hbb90e37f),
	.w3(32'hb7eb05c0),
	.w4(32'h3b5682dd),
	.w5(32'h3bcbebec),
	.w6(32'hbad1d60a),
	.w7(32'hbb0e2420),
	.w8(32'hba2fd923),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb906650),
	.w1(32'hbb1ded06),
	.w2(32'hbb55195b),
	.w3(32'h3b5dfad7),
	.w4(32'hba94c1f1),
	.w5(32'hbb8c7a32),
	.w6(32'hbb785e3c),
	.w7(32'hbb5caba4),
	.w8(32'hbc32faf3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba747f6f),
	.w1(32'h3b9227fd),
	.w2(32'hbaf693b5),
	.w3(32'hbbe8af13),
	.w4(32'h3b02422d),
	.w5(32'hbace151e),
	.w6(32'hbc01e43c),
	.w7(32'hb79ca312),
	.w8(32'hba6118f2),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3cce3),
	.w1(32'h3ad9e467),
	.w2(32'hbb1166a5),
	.w3(32'hbb685bda),
	.w4(32'h3a91b6c9),
	.w5(32'hbb506c7d),
	.w6(32'hbaf877e9),
	.w7(32'h3ab6e719),
	.w8(32'hbabb17ad),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d4be3),
	.w1(32'hbb591f2f),
	.w2(32'hbb9e69ef),
	.w3(32'hbb1868f0),
	.w4(32'hbb9209a1),
	.w5(32'hbb5b7653),
	.w6(32'hbb0d4d94),
	.w7(32'hbb9c5510),
	.w8(32'hbb7a2f90),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf0f37),
	.w1(32'hbba81d7d),
	.w2(32'h3ab24aad),
	.w3(32'h3ab0bde5),
	.w4(32'hbbaffd7e),
	.w5(32'hba5b8568),
	.w6(32'h3b519b0b),
	.w7(32'hbbb495fc),
	.w8(32'hbbeedc55),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6ba28),
	.w1(32'h3a754fa7),
	.w2(32'h3ae3dd61),
	.w3(32'hba49b66c),
	.w4(32'hba2a2e64),
	.w5(32'hbb0cf919),
	.w6(32'hbba4fbfe),
	.w7(32'hbb15beca),
	.w8(32'hba72ad1e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9389f),
	.w1(32'hbb112c68),
	.w2(32'hbb477aaa),
	.w3(32'hbb375321),
	.w4(32'hbb695a79),
	.w5(32'hbba2f9c7),
	.w6(32'hbb7ba2a8),
	.w7(32'hbbd4d250),
	.w8(32'hbbc7ee12),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a521a72),
	.w1(32'hbb5f8b25),
	.w2(32'h3ab851d7),
	.w3(32'h3b0741f0),
	.w4(32'hbbad273d),
	.w5(32'hbb425210),
	.w6(32'hbaec6943),
	.w7(32'hbb8640a1),
	.w8(32'hbb1e9a9b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b863e0e),
	.w1(32'hbacc1971),
	.w2(32'hba1673f9),
	.w3(32'h3b3e7d28),
	.w4(32'hba993444),
	.w5(32'hb84fe55c),
	.w6(32'h3ab33583),
	.w7(32'hbb26d529),
	.w8(32'hbad24bed),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c4be86),
	.w1(32'h37818512),
	.w2(32'hbab4b29c),
	.w3(32'h3af66173),
	.w4(32'h3b037ba5),
	.w5(32'h3b93adc5),
	.w6(32'hb991f65b),
	.w7(32'h3ba40145),
	.w8(32'h3b5bd937),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba20706),
	.w1(32'hbb2ab362),
	.w2(32'hbb57f59a),
	.w3(32'hbb1b21ea),
	.w4(32'hbb4762ec),
	.w5(32'hba953529),
	.w6(32'hb9a3466a),
	.w7(32'hbb77672c),
	.w8(32'hbb6f2c0f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7bd00),
	.w1(32'hb993d820),
	.w2(32'h3aad26f4),
	.w3(32'h3b419479),
	.w4(32'h3b8ad99c),
	.w5(32'h3ab8ad7a),
	.w6(32'h3b56e229),
	.w7(32'hb912d296),
	.w8(32'h399f3b1b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d09e0),
	.w1(32'h3b816c20),
	.w2(32'h3b236aaa),
	.w3(32'hbaf0ea67),
	.w4(32'h3b813023),
	.w5(32'h3ac3e46a),
	.w6(32'hb9d2e289),
	.w7(32'h3abb8a13),
	.w8(32'hb985c57e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b141f40),
	.w1(32'hbac2eb26),
	.w2(32'h3a133cb7),
	.w3(32'h3b5a0c56),
	.w4(32'hbb4ded88),
	.w5(32'hba0e61b8),
	.w6(32'h3b952c62),
	.w7(32'hbb354777),
	.w8(32'hbbba4d3b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacebea4),
	.w1(32'h3ba5c7dd),
	.w2(32'hb95cda2b),
	.w3(32'hbb2f9f10),
	.w4(32'hba778bc5),
	.w5(32'hbbddced8),
	.w6(32'h3a8cb24a),
	.w7(32'hbb4d6c04),
	.w8(32'hbbc33284),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad94780),
	.w1(32'h3b1b9e74),
	.w2(32'hbb9cdeca),
	.w3(32'hbac1f362),
	.w4(32'hbac08ad8),
	.w5(32'hbbc70555),
	.w6(32'h3aa201ba),
	.w7(32'h3b2aa34f),
	.w8(32'hbb8aec96),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf4117),
	.w1(32'hbb886829),
	.w2(32'hb98c3c7a),
	.w3(32'h3b1926eb),
	.w4(32'hbb6cc4ed),
	.w5(32'h3b1bea88),
	.w6(32'h3bb8495a),
	.w7(32'hbbf7743d),
	.w8(32'h3b1541f0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92fe40e),
	.w1(32'h3b6112c8),
	.w2(32'hbb0c4c71),
	.w3(32'hba52eea1),
	.w4(32'h3b710716),
	.w5(32'hbb2e32b7),
	.w6(32'hbb94d211),
	.w7(32'h3b1458f4),
	.w8(32'h3c06723d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb556f),
	.w1(32'h3bfb4036),
	.w2(32'h3addc37b),
	.w3(32'h3b9baa15),
	.w4(32'h3c30d7e1),
	.w5(32'h3b80da77),
	.w6(32'h3bf08530),
	.w7(32'h3c03e50f),
	.w8(32'h3b16045f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf40c65),
	.w1(32'hba5aac91),
	.w2(32'hb9894198),
	.w3(32'hbb3aa8f7),
	.w4(32'hbb23558c),
	.w5(32'hbb83bf1b),
	.w6(32'hbb064009),
	.w7(32'h3992daed),
	.w8(32'hbac0b49b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d8d28),
	.w1(32'hba4fca2d),
	.w2(32'hbb25266b),
	.w3(32'h3b00fbca),
	.w4(32'h3aeef653),
	.w5(32'hb88a282c),
	.w6(32'hba2c5a45),
	.w7(32'hb9f047be),
	.w8(32'hbae3c78e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dcc53),
	.w1(32'h39013923),
	.w2(32'hba8f0b63),
	.w3(32'hbaa81dec),
	.w4(32'h3a955d30),
	.w5(32'h3b19328e),
	.w6(32'h399aa3c7),
	.w7(32'hb989fd0d),
	.w8(32'h3af5a752),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad62f98),
	.w1(32'h3a1abbb3),
	.w2(32'hb9d6cf1e),
	.w3(32'h3aa4dc51),
	.w4(32'h3c25d1b5),
	.w5(32'h3c19df71),
	.w6(32'h3b73cde4),
	.w7(32'h3b8907dd),
	.w8(32'h3a87d348),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f3e838),
	.w1(32'hb913b3ba),
	.w2(32'h3a8803a2),
	.w3(32'h3b8931fd),
	.w4(32'hbaa61186),
	.w5(32'h39fb8c58),
	.w6(32'h3b7a76a5),
	.w7(32'hbabff806),
	.w8(32'hbb148971),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeba726),
	.w1(32'h3b1389cc),
	.w2(32'h3bb7a2ba),
	.w3(32'h3a61c3a1),
	.w4(32'h397276ac),
	.w5(32'h399f4cc4),
	.w6(32'hb9c005f1),
	.w7(32'h39ab4221),
	.w8(32'hba9c93fa),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5cb74),
	.w1(32'h3b3d9365),
	.w2(32'h3a514439),
	.w3(32'h3a097804),
	.w4(32'h3aae534f),
	.w5(32'hbaf3f161),
	.w6(32'hbac4c513),
	.w7(32'h3aabd788),
	.w8(32'h3b95ec8d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913ad53),
	.w1(32'h3b4cca9e),
	.w2(32'h3b6e4bce),
	.w3(32'hbb4a74ee),
	.w4(32'hb9cb7dc4),
	.w5(32'h3ac41b8a),
	.w6(32'h3a86bf10),
	.w7(32'h3b57a8af),
	.w8(32'h3aeba650),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47f8df),
	.w1(32'h39b88049),
	.w2(32'h3bcc01b6),
	.w3(32'hbb35194a),
	.w4(32'h3af36d99),
	.w5(32'h3c0f4a97),
	.w6(32'h3a892059),
	.w7(32'h3bd53733),
	.w8(32'h3b8e2d0c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dc061),
	.w1(32'h3930498c),
	.w2(32'hb980c1b9),
	.w3(32'h3bb311ef),
	.w4(32'h3a868804),
	.w5(32'h3ad007bd),
	.w6(32'h3bd8ae36),
	.w7(32'h3ad46215),
	.w8(32'hba1204f3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c07d27),
	.w1(32'hba8e248d),
	.w2(32'h3ba90288),
	.w3(32'h3ae06dd1),
	.w4(32'hbae6be83),
	.w5(32'h3b478a50),
	.w6(32'h3a9b5a5a),
	.w7(32'hbb721cb0),
	.w8(32'hbb0c1be8),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79f469),
	.w1(32'h3bda8e5d),
	.w2(32'h3922109d),
	.w3(32'h3a9ede33),
	.w4(32'h3ba20967),
	.w5(32'h39c6ab7e),
	.w6(32'h3a71d56e),
	.w7(32'h3bac77bd),
	.w8(32'hba8c0d56),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27abe9),
	.w1(32'h3acc1e99),
	.w2(32'h3b72789b),
	.w3(32'hbb1c83a0),
	.w4(32'h3ac307b5),
	.w5(32'h3be53081),
	.w6(32'hb91b7277),
	.w7(32'h3b6430ca),
	.w8(32'h3b1205f9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae00cf),
	.w1(32'h3b3c9111),
	.w2(32'hbbaeaad5),
	.w3(32'hbaaf7e9a),
	.w4(32'hbaca48c6),
	.w5(32'hbc183cdf),
	.w6(32'hbb79586d),
	.w7(32'hb9ed76bb),
	.w8(32'hbc1474be),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb90e1),
	.w1(32'hb8e043f4),
	.w2(32'hbb159922),
	.w3(32'h3b830ea6),
	.w4(32'h3b5a78f2),
	.w5(32'hb9240225),
	.w6(32'h3b876478),
	.w7(32'hb9aa2668),
	.w8(32'hba730ed4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997259d),
	.w1(32'h3b38aeba),
	.w2(32'h3ba0423f),
	.w3(32'h3a40bbdb),
	.w4(32'h3b3459b1),
	.w5(32'h3c2f1b51),
	.w6(32'h3a570d19),
	.w7(32'h3be5f9ca),
	.w8(32'h3b80303c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b945c0a),
	.w1(32'hba06fc71),
	.w2(32'hba357175),
	.w3(32'h3ac88d14),
	.w4(32'hb9be4b61),
	.w5(32'h3b0c32b0),
	.w6(32'h3b3a6f42),
	.w7(32'hb91f9379),
	.w8(32'hbb89fea8),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55ef4c),
	.w1(32'hba395d30),
	.w2(32'hbb0385b0),
	.w3(32'hbbc3ea13),
	.w4(32'hba416fbf),
	.w5(32'hbb2267e3),
	.w6(32'hbb465e5b),
	.w7(32'hbb991316),
	.w8(32'hba8c1921),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab22298),
	.w1(32'hbbcf1014),
	.w2(32'hbbbff9b5),
	.w3(32'h3acee220),
	.w4(32'hbc0aa71b),
	.w5(32'hbba2c536),
	.w6(32'h3a203168),
	.w7(32'hbbc5ce7a),
	.w8(32'hbbe3edf8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b0d72),
	.w1(32'h3ade1be1),
	.w2(32'hbb8773d1),
	.w3(32'hbb673ef7),
	.w4(32'h39167f78),
	.w5(32'hbb42751f),
	.w6(32'hbb88957a),
	.w7(32'hbaae0671),
	.w8(32'hbbd56690),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff1a01),
	.w1(32'hbb041e34),
	.w2(32'h3b81af9a),
	.w3(32'h3b20591a),
	.w4(32'h3a74d06e),
	.w5(32'h3b791608),
	.w6(32'h3a4d1386),
	.w7(32'h3b3d7898),
	.w8(32'hb980b8c3),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a7441),
	.w1(32'hbb170c75),
	.w2(32'hbab282d7),
	.w3(32'hbbd40ef7),
	.w4(32'hba6bf1ba),
	.w5(32'hbb6a224d),
	.w6(32'hbb1c6755),
	.w7(32'hb75ff4d3),
	.w8(32'hbb3b566d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73d017),
	.w1(32'h3ae8df70),
	.w2(32'h3b23df4e),
	.w3(32'h3b305895),
	.w4(32'h39023dab),
	.w5(32'hb8c0e4cb),
	.w6(32'hba5b1e57),
	.w7(32'h3b0895c6),
	.w8(32'h3bd7d395),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f447f),
	.w1(32'h3b1cc9ae),
	.w2(32'hbabc42c0),
	.w3(32'h3b3101d7),
	.w4(32'h3a68587d),
	.w5(32'hba89b89b),
	.w6(32'h3bc58e6e),
	.w7(32'h3ada8799),
	.w8(32'hbae283f5),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9beaed),
	.w1(32'h3baf3ce1),
	.w2(32'h3af6cb71),
	.w3(32'hba36797b),
	.w4(32'h3b912734),
	.w5(32'h3a75feb1),
	.w6(32'hb95edac0),
	.w7(32'h3ae6edcf),
	.w8(32'hbab3e702),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba202116),
	.w1(32'hba5567ab),
	.w2(32'hba79cf8e),
	.w3(32'hb84b04b1),
	.w4(32'h3b91274d),
	.w5(32'h3be0a728),
	.w6(32'hba9c8b6f),
	.w7(32'h3bbfcc81),
	.w8(32'h3ba3792c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b353fd0),
	.w1(32'h3a111ab3),
	.w2(32'h3b4cc65f),
	.w3(32'h3be93f07),
	.w4(32'h3b92b920),
	.w5(32'h3bc9b6d5),
	.w6(32'h3bfc014b),
	.w7(32'hba2d1049),
	.w8(32'h3a8db7ff),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cf13c),
	.w1(32'hb9d37139),
	.w2(32'h3b8a32b9),
	.w3(32'h3bb692a0),
	.w4(32'hba1215fe),
	.w5(32'h3bae6a97),
	.w6(32'h3b9cbcf1),
	.w7(32'h3aaa5f63),
	.w8(32'h39c4009f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a940653),
	.w1(32'h3b906007),
	.w2(32'h3c1ceb37),
	.w3(32'h3acb64c7),
	.w4(32'hbb1216ff),
	.w5(32'h3aaed5da),
	.w6(32'hbaf90f0e),
	.w7(32'hbb1a5e8a),
	.w8(32'hba4452e3),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8045e),
	.w1(32'h3b2387a5),
	.w2(32'hbb55628a),
	.w3(32'h3a475386),
	.w4(32'h3bc8aac5),
	.w5(32'h3a990bbc),
	.w6(32'h3bb2aea8),
	.w7(32'h3bab4252),
	.w8(32'hb96b3d8c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba089347),
	.w1(32'h3a1a7778),
	.w2(32'hbbc4175e),
	.w3(32'hbaeb394a),
	.w4(32'hbb495667),
	.w5(32'hb9c94d2c),
	.w6(32'hba04629c),
	.w7(32'h3b8feff6),
	.w8(32'hb91c09ff),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e20a2),
	.w1(32'hba9c4150),
	.w2(32'hbadaeb2f),
	.w3(32'hbb61d06a),
	.w4(32'hbb12c2bd),
	.w5(32'h3a714e04),
	.w6(32'hbb9d77de),
	.w7(32'hbb2559c8),
	.w8(32'hbb2918e4),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6343dc),
	.w1(32'hba8a9a0a),
	.w2(32'hbbc4a5ee),
	.w3(32'h3b9cfb28),
	.w4(32'hbb68e7fe),
	.w5(32'hbbe94c0b),
	.w6(32'h3c1104ac),
	.w7(32'hbaf8d9fe),
	.w8(32'hbc89a4ad),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea74e2),
	.w1(32'h3bac2ee8),
	.w2(32'h3b419dc2),
	.w3(32'hbb72c178),
	.w4(32'h3c0d9d26),
	.w5(32'h3bbbee95),
	.w6(32'hbae2e819),
	.w7(32'h3b370557),
	.w8(32'h3a868019),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b4441),
	.w1(32'h3b0ce89c),
	.w2(32'hbaaba573),
	.w3(32'h3b4fe5fc),
	.w4(32'hb9bf7caa),
	.w5(32'hbb7ea662),
	.w6(32'h3b3b395e),
	.w7(32'hbaa8604b),
	.w8(32'hbb12f39a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dd50d),
	.w1(32'h39b3b432),
	.w2(32'h3bb200b7),
	.w3(32'h3bb50c7f),
	.w4(32'hbb93e146),
	.w5(32'h3b5ebb4c),
	.w6(32'h3b192044),
	.w7(32'hbb1e99be),
	.w8(32'hbad2f25d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e83fa),
	.w1(32'hbb91ffef),
	.w2(32'hbbf6c836),
	.w3(32'hbb9a5e6d),
	.w4(32'hbaebcd20),
	.w5(32'hbb786615),
	.w6(32'hbb27b93c),
	.w7(32'hbb4c57d3),
	.w8(32'hbb4da7dd),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb586f14),
	.w1(32'h3b539bfb),
	.w2(32'h3b9b45c8),
	.w3(32'hba6cf1df),
	.w4(32'h395b723b),
	.w5(32'h3b32b6aa),
	.w6(32'h3a500b31),
	.w7(32'h3aa82dd6),
	.w8(32'h3bafbbdf),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe791a),
	.w1(32'h3c0e24a0),
	.w2(32'hb98a049d),
	.w3(32'h3bb8b857),
	.w4(32'h3baf2e77),
	.w5(32'h3a41c217),
	.w6(32'h3c1284f8),
	.w7(32'h3c283d50),
	.w8(32'h3c10db7c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5555c),
	.w1(32'hbad5e4d2),
	.w2(32'hbb786f9c),
	.w3(32'h3bdfb149),
	.w4(32'hba9ace91),
	.w5(32'hbac27ab0),
	.w6(32'h3bea5d0e),
	.w7(32'hbb4ec3e6),
	.w8(32'hbb98b4df),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8df8),
	.w1(32'hba92ca2e),
	.w2(32'hbad1b01f),
	.w3(32'hbb21b69e),
	.w4(32'hba86f1f7),
	.w5(32'hbb5c9715),
	.w6(32'hbb06ea5e),
	.w7(32'h3a855e31),
	.w8(32'hbb48acdc),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f13b4c),
	.w1(32'hbab4fe39),
	.w2(32'h3bc2e9ca),
	.w3(32'hba5a28a5),
	.w4(32'hbb30ac6e),
	.w5(32'h3b9686f6),
	.w6(32'hbb1ab82a),
	.w7(32'hbb92b9f7),
	.w8(32'hbb3cc79c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3e0a3),
	.w1(32'h3b204255),
	.w2(32'hbb1c2690),
	.w3(32'hb9b2a288),
	.w4(32'h3a43f4ee),
	.w5(32'hbb6d310f),
	.w6(32'h39383860),
	.w7(32'h39519a26),
	.w8(32'hbba77e7e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad39044),
	.w1(32'h39b08377),
	.w2(32'hba296771),
	.w3(32'hb983165f),
	.w4(32'h3a3832e2),
	.w5(32'hb9520823),
	.w6(32'hb91ae086),
	.w7(32'h3b0fdb84),
	.w8(32'h3aa9dda3),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7f9fe),
	.w1(32'hb9c34cb6),
	.w2(32'hb71cced9),
	.w3(32'hb9f60188),
	.w4(32'hb9919eb4),
	.w5(32'hba2f99a5),
	.w6(32'h384e7e49),
	.w7(32'hba310b2a),
	.w8(32'hb9d19f82),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb416b0e),
	.w1(32'hba627160),
	.w2(32'hbb085a8a),
	.w3(32'hbb7b4608),
	.w4(32'hba29482e),
	.w5(32'hba91dcce),
	.w6(32'hbaf05a95),
	.w7(32'h3b1fe3f9),
	.w8(32'h3a9fa4c2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9a791),
	.w1(32'h3951b2f8),
	.w2(32'h394ae34d),
	.w3(32'hb9ec60e6),
	.w4(32'h39821468),
	.w5(32'h39b2ebec),
	.w6(32'hb9192d8a),
	.w7(32'h39dad75c),
	.w8(32'h39bd5a45),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace7435),
	.w1(32'h3aa858c0),
	.w2(32'hba8a1cef),
	.w3(32'h3a011d17),
	.w4(32'h3aa17a95),
	.w5(32'hba125eee),
	.w6(32'h3abe7b4c),
	.w7(32'h389bb7d8),
	.w8(32'hbb0874a3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59a742),
	.w1(32'hba012bff),
	.w2(32'h3a106547),
	.w3(32'h3a336f46),
	.w4(32'h3b31c1f3),
	.w5(32'h3b5d1a29),
	.w6(32'hbaed318d),
	.w7(32'hbae1bb42),
	.w8(32'h3a356dbe),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c20606),
	.w1(32'h3a53679b),
	.w2(32'hb8b41fbb),
	.w3(32'h3a9e8806),
	.w4(32'h3ae5b9dc),
	.w5(32'h3a581588),
	.w6(32'h3a85df65),
	.w7(32'h3ad3bd81),
	.w8(32'h3a6bbc7e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b6ddd),
	.w1(32'h39e4bfe8),
	.w2(32'hb7dc68b1),
	.w3(32'h3a04fad1),
	.w4(32'h399813de),
	.w5(32'hb96f956c),
	.w6(32'hb9294a35),
	.w7(32'hb97dcd30),
	.w8(32'h37fd2cec),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe563f),
	.w1(32'h3b1a978f),
	.w2(32'h3b47da77),
	.w3(32'hb81b1262),
	.w4(32'h3b02fdb0),
	.w5(32'h3b1bc041),
	.w6(32'h39f4cbbc),
	.w7(32'h3ae9924e),
	.w8(32'h3b514ecb),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba079a48),
	.w1(32'hba2e504e),
	.w2(32'hbae1900f),
	.w3(32'hbac9b069),
	.w4(32'hbaa891b9),
	.w5(32'hbb160a38),
	.w6(32'h3a84da4f),
	.w7(32'hba843d17),
	.w8(32'hbb51f6f4),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73a7ac),
	.w1(32'hba5c5a7b),
	.w2(32'hb976d273),
	.w3(32'h3a6c66e7),
	.w4(32'h38ad78f6),
	.w5(32'hb9761410),
	.w6(32'h3b1e97fc),
	.w7(32'h3a5e29b1),
	.w8(32'hbae5e730),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a406f7a),
	.w1(32'h39b14d47),
	.w2(32'h3915c208),
	.w3(32'h3a510f4d),
	.w4(32'h390b1a12),
	.w5(32'hb8b64b07),
	.w6(32'h3a7e76c3),
	.w7(32'h3993c56d),
	.w8(32'hb8c4d7a4),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3946c97f),
	.w1(32'h39b8a586),
	.w2(32'h39b24a51),
	.w3(32'h39127211),
	.w4(32'h39ba69a2),
	.w5(32'h395ec8ad),
	.w6(32'hb7b7f3ec),
	.w7(32'h39e8069d),
	.w8(32'h39f6c025),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aceef57),
	.w1(32'h3ae03c44),
	.w2(32'hb9e7bd75),
	.w3(32'h3ba107e2),
	.w4(32'h3b22de65),
	.w5(32'hbb0fbaec),
	.w6(32'h3b39a84a),
	.w7(32'h3b2339d6),
	.w8(32'hb9c125d7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba869fc7),
	.w1(32'hbb25355d),
	.w2(32'hbb8e75fc),
	.w3(32'hbac63685),
	.w4(32'hba9a833f),
	.w5(32'hbb8cc99b),
	.w6(32'hbae7872a),
	.w7(32'hbae4ff03),
	.w8(32'hbba34a5e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0e302),
	.w1(32'hbab238fa),
	.w2(32'hb98ddf1b),
	.w3(32'hbaa1d66d),
	.w4(32'hba1389f6),
	.w5(32'hba8ff825),
	.w6(32'h38e3ac1c),
	.w7(32'h3a535da5),
	.w8(32'h388e3874),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87ab8d),
	.w1(32'h3a7cec3e),
	.w2(32'hbacbf9df),
	.w3(32'h3a3bfb22),
	.w4(32'h3b59d935),
	.w5(32'h3b02750e),
	.w6(32'h3b59ed23),
	.w7(32'h3a82a025),
	.w8(32'hbac3f72d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6a50c),
	.w1(32'hba232083),
	.w2(32'hb984df06),
	.w3(32'hb9dbf600),
	.w4(32'hba1b0622),
	.w5(32'hba330182),
	.w6(32'hb9517625),
	.w7(32'hb9be0de9),
	.w8(32'h3819ca5d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c1c5a),
	.w1(32'hba5af703),
	.w2(32'hba1a50b5),
	.w3(32'hba7ac16a),
	.w4(32'hba13dd40),
	.w5(32'hb9449e45),
	.w6(32'hb86cafc2),
	.w7(32'hb9a5b4f0),
	.w8(32'hb93551ac),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8187be),
	.w1(32'h3c0ec729),
	.w2(32'hbb13b32f),
	.w3(32'h3b93ef33),
	.w4(32'h3beb3123),
	.w5(32'hbaea358e),
	.w6(32'h3b06ffd9),
	.w7(32'h3bc137eb),
	.w8(32'hb98d2155),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96bf22),
	.w1(32'hbb838934),
	.w2(32'hbb9df815),
	.w3(32'hba758bc8),
	.w4(32'hbba3f43e),
	.w5(32'hbbaaefff),
	.w6(32'h3afb3009),
	.w7(32'hbb1d869e),
	.w8(32'hbbe065f8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b494710),
	.w1(32'h3b2defe3),
	.w2(32'hbb08731a),
	.w3(32'h3a6db18c),
	.w4(32'hb9bc2d08),
	.w5(32'hbaa794d6),
	.w6(32'hbb09eaae),
	.w7(32'h3b22c4de),
	.w8(32'hbaa82c02),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16f832),
	.w1(32'h3ab4e77f),
	.w2(32'h3b459197),
	.w3(32'hba618912),
	.w4(32'h3b260537),
	.w5(32'h3b6a8fb9),
	.w6(32'hbace0163),
	.w7(32'h39f7fbf3),
	.w8(32'h3b2da0e9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8360a4),
	.w1(32'hba07ade5),
	.w2(32'h3a438b1a),
	.w3(32'hbaf630b1),
	.w4(32'h3a6d11f8),
	.w5(32'h3b007e84),
	.w6(32'hbb01530d),
	.w7(32'hbb01cc61),
	.w8(32'hb9af659e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d30395),
	.w1(32'hb7e2a6e4),
	.w2(32'h39c90d21),
	.w3(32'h39dc4cd9),
	.w4(32'hb9f30e35),
	.w5(32'hb9f516b4),
	.w6(32'h39e4918c),
	.w7(32'hb909a55c),
	.w8(32'hb841207d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b96b93),
	.w1(32'hb9487ed0),
	.w2(32'hb9e6c31b),
	.w3(32'hb98cf371),
	.w4(32'h3a684391),
	.w5(32'h377a513b),
	.w6(32'hb997c5af),
	.w7(32'h3a0c8346),
	.w8(32'hb9c55d37),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0870e5),
	.w1(32'hb9532a8c),
	.w2(32'hb9ad786c),
	.w3(32'h397055b1),
	.w4(32'hb97393e6),
	.w5(32'hba32c8ee),
	.w6(32'h38d30cd9),
	.w7(32'hb943b18c),
	.w8(32'hba2a76f5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384c87d6),
	.w1(32'h39579a3f),
	.w2(32'h3a589e4a),
	.w3(32'hb90678f7),
	.w4(32'h37c90940),
	.w5(32'h39df5a16),
	.w6(32'h386d33b5),
	.w7(32'hb9ba18d9),
	.w8(32'h3a6ba563),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1be177),
	.w1(32'h3a9c6768),
	.w2(32'hb953f55e),
	.w3(32'h3b1d6698),
	.w4(32'hb8d78587),
	.w5(32'hb9fc9851),
	.w6(32'h3afefb5c),
	.w7(32'h384b7ff4),
	.w8(32'hba0ad35f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf00f8),
	.w1(32'hbb916337),
	.w2(32'hbba46703),
	.w3(32'hbae0667a),
	.w4(32'hbb0b7dec),
	.w5(32'hbba367d6),
	.w6(32'hbabaa58c),
	.w7(32'hbb13d04a),
	.w8(32'hbbaa4789),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae75180),
	.w1(32'hb9145c6a),
	.w2(32'hb8d8c92c),
	.w3(32'hb9cb4b6c),
	.w4(32'h3a597717),
	.w5(32'h3a454c15),
	.w6(32'hbac57d22),
	.w7(32'h3a684b55),
	.w8(32'hba04cf24),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abf946),
	.w1(32'h39398da3),
	.w2(32'hb9c35918),
	.w3(32'h397282c8),
	.w4(32'h398b25ac),
	.w5(32'hb9294236),
	.w6(32'h395e1647),
	.w7(32'hb940a256),
	.w8(32'hb904a65f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a10e99),
	.w1(32'h3a7f0a2d),
	.w2(32'hbb8d6dda),
	.w3(32'hbb545c16),
	.w4(32'hb902a960),
	.w5(32'hbb2d9e81),
	.w6(32'hbb598ed9),
	.w7(32'h3ad6a614),
	.w8(32'hbb9bd078),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccc36a),
	.w1(32'hbadeef42),
	.w2(32'hbb22c133),
	.w3(32'hb9b6173e),
	.w4(32'hbad4fb5e),
	.w5(32'hbb46fc79),
	.w6(32'h38cb2a64),
	.w7(32'hba968615),
	.w8(32'hbb61b1d7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42276a),
	.w1(32'h3a18a40d),
	.w2(32'h3a187eb3),
	.w3(32'hba93f50c),
	.w4(32'h38c96af8),
	.w5(32'h3913387b),
	.w6(32'hba3f5f80),
	.w7(32'h3908a6ef),
	.w8(32'h3a18c6ee),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ee227),
	.w1(32'hba99d536),
	.w2(32'hbb28ec75),
	.w3(32'hb89c9f38),
	.w4(32'hbaa93fe0),
	.w5(32'hbad76b56),
	.w6(32'h3a0075e0),
	.w7(32'hb9bbb6ac),
	.w8(32'hbb57d70c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a152463),
	.w1(32'h3aa7939c),
	.w2(32'h3a2b39d2),
	.w3(32'h3a3e1b0a),
	.w4(32'h3a8c6f56),
	.w5(32'h39c54e8a),
	.w6(32'h3a05a859),
	.w7(32'h39e91c7f),
	.w8(32'hb793a3fb),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d92dd),
	.w1(32'h3a27a20a),
	.w2(32'hb9e61861),
	.w3(32'h39eff0d6),
	.w4(32'h39f4b130),
	.w5(32'hb9ffe7a7),
	.w6(32'h39537afb),
	.w7(32'h3a15beee),
	.w8(32'hb981f9b0),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943ceb3),
	.w1(32'h39de8666),
	.w2(32'h39a93931),
	.w3(32'hb8904431),
	.w4(32'h3a3f6c94),
	.w5(32'h3987ce33),
	.w6(32'h397fb9bc),
	.w7(32'h391ade9b),
	.w8(32'h39d7d13b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398addcf),
	.w1(32'h39ea3ca6),
	.w2(32'h390a637e),
	.w3(32'h39b1a36b),
	.w4(32'h39c698a9),
	.w5(32'hb92886f8),
	.w6(32'h398cff6d),
	.w7(32'h3a02f82e),
	.w8(32'h3a0dfb1d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba908e33),
	.w1(32'h3965b669),
	.w2(32'h3a9fb639),
	.w3(32'hba194804),
	.w4(32'h3a3d7c6f),
	.w5(32'h3aa0d5f8),
	.w6(32'hba3469a5),
	.w7(32'hb6f32592),
	.w8(32'h3adbd568),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0cd5f),
	.w1(32'hbb34ee0e),
	.w2(32'hbb7c6c25),
	.w3(32'hbb2d6474),
	.w4(32'hbb3f47bb),
	.w5(32'hbb448389),
	.w6(32'hb9cec6bf),
	.w7(32'hbb37c6d5),
	.w8(32'hbbbbc0a0),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba987828),
	.w1(32'hba1addaa),
	.w2(32'hbac7c87d),
	.w3(32'hba68a043),
	.w4(32'hba51aa8a),
	.w5(32'hbae27aa6),
	.w6(32'h3a916a5e),
	.w7(32'h3a1ecaac),
	.w8(32'hbb3694a5),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a52bfe),
	.w1(32'hba612944),
	.w2(32'hbafac225),
	.w3(32'hbaadb102),
	.w4(32'hba4514d2),
	.w5(32'hba8c794b),
	.w6(32'h3aa4d3d3),
	.w7(32'hba478a55),
	.w8(32'hbb543586),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15576e),
	.w1(32'h39eb95dd),
	.w2(32'h39dfb874),
	.w3(32'h39ad963e),
	.w4(32'h39659ed5),
	.w5(32'h39c4d870),
	.w6(32'h39a6f96f),
	.w7(32'h39841e2b),
	.w8(32'h391dc0d1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aeebce),
	.w1(32'hba41879d),
	.w2(32'hba1558d7),
	.w3(32'hb98f4f89),
	.w4(32'hb9710e2c),
	.w5(32'hb9daa2cb),
	.w6(32'h39825292),
	.w7(32'h3975a6b2),
	.w8(32'hb9c6674c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe2f10),
	.w1(32'h388fc3c4),
	.w2(32'h38d4f1e1),
	.w3(32'hb7cde06b),
	.w4(32'hb96f95b6),
	.w5(32'hb96567a1),
	.w6(32'h387dfc3a),
	.w7(32'h39734364),
	.w8(32'h38bf582a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399083cf),
	.w1(32'h39d8821a),
	.w2(32'hb89b71de),
	.w3(32'hb987f983),
	.w4(32'h390e7e95),
	.w5(32'h393bcd0b),
	.w6(32'hb923f2d3),
	.w7(32'hb91352d2),
	.w8(32'h3771eaf6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0193a9),
	.w1(32'hbb93ba87),
	.w2(32'hbb9bc656),
	.w3(32'hbad2fec3),
	.w4(32'hbb96ed8a),
	.w5(32'hbba1ea50),
	.w6(32'h3a32d061),
	.w7(32'hbb55c3f8),
	.w8(32'hbb9b7f43),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd03c3),
	.w1(32'hba885b95),
	.w2(32'hba842e5b),
	.w3(32'hbab92957),
	.w4(32'hbaa64f99),
	.w5(32'hbad69517),
	.w6(32'hbab2e080),
	.w7(32'hbae160d6),
	.w8(32'hbb081e2a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fc2e6),
	.w1(32'h3acae5b1),
	.w2(32'h3a49ae1c),
	.w3(32'h3a808659),
	.w4(32'h3af5391f),
	.w5(32'h3ac39881),
	.w6(32'h3a8d7b17),
	.w7(32'h3ada4e78),
	.w8(32'h3a9c2338),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9083553),
	.w1(32'h396ced71),
	.w2(32'h391abe21),
	.w3(32'h3a2abf9b),
	.w4(32'h3a2d6b00),
	.w5(32'h3ab7e790),
	.w6(32'h3a060003),
	.w7(32'h3a37b965),
	.w8(32'h3a8d95ed),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f30203),
	.w1(32'h38b9e5d3),
	.w2(32'hb99d0656),
	.w3(32'h3958783e),
	.w4(32'hb879f0af),
	.w5(32'hb9e23177),
	.w6(32'hb94ecf25),
	.w7(32'h3771ae53),
	.w8(32'hba20627b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eb225),
	.w1(32'h39f7da0c),
	.w2(32'hb9eee46d),
	.w3(32'h3a898a01),
	.w4(32'h3a28cfa8),
	.w5(32'hb8086bbd),
	.w6(32'h3ad21e5d),
	.w7(32'hb88c9405),
	.w8(32'hba8bd523),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4bff3),
	.w1(32'hb9836631),
	.w2(32'hb9e41432),
	.w3(32'hb948fa3c),
	.w4(32'hb96cf2d5),
	.w5(32'hba42c732),
	.w6(32'h39373930),
	.w7(32'hba1ac6d4),
	.w8(32'hba5bbbd3),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d26f1),
	.w1(32'hbb954aed),
	.w2(32'hbbad08d8),
	.w3(32'hbb0e562f),
	.w4(32'hbb384663),
	.w5(32'hbb0366a8),
	.w6(32'hbb449db0),
	.w7(32'hbbdd447a),
	.w8(32'hbbc073c9),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7f298),
	.w1(32'hb9caf50a),
	.w2(32'hba113f25),
	.w3(32'hb863a2ac),
	.w4(32'hba2cc3c8),
	.w5(32'hba7813ee),
	.w6(32'h3993efe1),
	.w7(32'hb9ccfcfb),
	.w8(32'hba6beb48),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72b656),
	.w1(32'h3a15cf0e),
	.w2(32'h3b3b06f9),
	.w3(32'hbb9d2a8c),
	.w4(32'hb9877e00),
	.w5(32'h3852a92e),
	.w6(32'hbb4a82d9),
	.w7(32'h3a296f2a),
	.w8(32'h3b0294f7),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule