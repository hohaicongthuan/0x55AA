module layer_8_featuremap_50(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60b7a78),
	.w1(32'h3896f6b1),
	.w2(32'h38b8fc66),
	.w3(32'hb986780c),
	.w4(32'hb89eb52b),
	.w5(32'hb6525d83),
	.w6(32'hb98f45e8),
	.w7(32'hb808bdea),
	.w8(32'h386d1680),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a21ed),
	.w1(32'h37819ac9),
	.w2(32'hb95ccdf6),
	.w3(32'h395186f7),
	.w4(32'h3908ce3c),
	.w5(32'hb850ae04),
	.w6(32'h37e80cf3),
	.w7(32'h3822149c),
	.w8(32'hb841600c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ae6874),
	.w1(32'h377d9d4f),
	.w2(32'hb7fbbf19),
	.w3(32'hb893a01d),
	.w4(32'hb76e3f16),
	.w5(32'h38e8fcc2),
	.w6(32'hb9775651),
	.w7(32'hb91122d7),
	.w8(32'hb8db23cc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81bcbad),
	.w1(32'hb8dde032),
	.w2(32'hb7c0d4c7),
	.w3(32'hb79f5fc5),
	.w4(32'hb8903450),
	.w5(32'hb8cb9cdd),
	.w6(32'hb8d8b1ea),
	.w7(32'hb89a4e5c),
	.w8(32'hb8235513),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c735b),
	.w1(32'hb97c311d),
	.w2(32'hb9054d5f),
	.w3(32'hb997f67d),
	.w4(32'hb9b1aad6),
	.w5(32'hb87b6698),
	.w6(32'hba1df9f0),
	.w7(32'h3492d62f),
	.w8(32'h39054f5a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ec8d7),
	.w1(32'hb950bf8d),
	.w2(32'hb9becc01),
	.w3(32'h37d0fa7b),
	.w4(32'hb8b18614),
	.w5(32'hb9b34664),
	.w6(32'h39082b07),
	.w7(32'h38afac24),
	.w8(32'hb92a7772),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89b8c47),
	.w1(32'hb90613e5),
	.w2(32'h385ad119),
	.w3(32'hb8dfd029),
	.w4(32'hb854eeda),
	.w5(32'h39285aa7),
	.w6(32'hb9a24b7c),
	.w7(32'hb9337b00),
	.w8(32'hb86b6488),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba471a80),
	.w1(32'hba27173e),
	.w2(32'hba4ede85),
	.w3(32'hba3c0bed),
	.w4(32'hb98e03b9),
	.w5(32'hba774df9),
	.w6(32'hba2cfa24),
	.w7(32'h39093edd),
	.w8(32'hba331f74),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a1126),
	.w1(32'hb9e1423f),
	.w2(32'hb95e4900),
	.w3(32'hba79e759),
	.w4(32'hba2834a5),
	.w5(32'hba174013),
	.w6(32'hba815867),
	.w7(32'hba0f8edb),
	.w8(32'hba0965e7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67905c),
	.w1(32'h3992e003),
	.w2(32'h39c23889),
	.w3(32'h39db34ad),
	.w4(32'h394ee768),
	.w5(32'hb8d20c12),
	.w6(32'h39baa03d),
	.w7(32'h38a2f6dd),
	.w8(32'hb9228b32),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa2cdd),
	.w1(32'hb9b66d38),
	.w2(32'hb92c5534),
	.w3(32'hba870873),
	.w4(32'hba62d803),
	.w5(32'hb9a6435f),
	.w6(32'hbaa25115),
	.w7(32'hba515486),
	.w8(32'hba23f335),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3836e8af),
	.w1(32'h385589e1),
	.w2(32'h38e2aae3),
	.w3(32'hb8bcb445),
	.w4(32'hb8c52343),
	.w5(32'hb9384bd0),
	.w6(32'hb89f4f2f),
	.w7(32'hb805f29c),
	.w8(32'hb91ebf2c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a1ddf),
	.w1(32'h3906319d),
	.w2(32'h38df16ff),
	.w3(32'h38685754),
	.w4(32'hb7daed14),
	.w5(32'hba524c69),
	.w6(32'hba8f5fba),
	.w7(32'hba442fc4),
	.w8(32'hb9e52c65),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09c546),
	.w1(32'hba1df3ec),
	.w2(32'hba57b991),
	.w3(32'hba643ec8),
	.w4(32'hba800316),
	.w5(32'hba7c688d),
	.w6(32'hbab46a9d),
	.w7(32'hba9b32b8),
	.w8(32'hba95e758),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b51a1a),
	.w1(32'h37df85b0),
	.w2(32'h382cf2a3),
	.w3(32'hb7efc91c),
	.w4(32'hb81c9947),
	.w5(32'hb74ec48d),
	.w6(32'hb9262746),
	.w7(32'hb87956f7),
	.w8(32'h37b0fb1f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8d554),
	.w1(32'hb8ce4b8d),
	.w2(32'hba07c861),
	.w3(32'hb9686622),
	.w4(32'h395f15fb),
	.w5(32'hb9022077),
	.w6(32'hba406c1a),
	.w7(32'h38d0e8f3),
	.w8(32'h3a3196ae),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ddad1),
	.w1(32'h39b5d46b),
	.w2(32'hb84c5e79),
	.w3(32'h3a366fb6),
	.w4(32'h39b24436),
	.w5(32'h38a2ddaa),
	.w6(32'h3abde2d8),
	.w7(32'h3a7d3d35),
	.w8(32'h3a2b5bae),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d01755),
	.w1(32'h3996bda2),
	.w2(32'h39af2d59),
	.w3(32'hb9c27996),
	.w4(32'h3a0f13dd),
	.w5(32'h38978d84),
	.w6(32'hbacc86f0),
	.w7(32'hba47f8c6),
	.w8(32'h39b590ff),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e503d7),
	.w1(32'hb962f737),
	.w2(32'h3a7d4c58),
	.w3(32'hba71848b),
	.w4(32'hba4512d3),
	.w5(32'hba3a2f18),
	.w6(32'hbb19b520),
	.w7(32'hbab6cf0f),
	.w8(32'hba7a65da),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad43c68),
	.w1(32'hbb377a8e),
	.w2(32'hbafb137c),
	.w3(32'hbb95f40a),
	.w4(32'hbb19b704),
	.w5(32'hb93d614a),
	.w6(32'hbba533f1),
	.w7(32'hbb139200),
	.w8(32'hba9cadbc),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba128aac),
	.w1(32'hb97df033),
	.w2(32'h3a1fddbc),
	.w3(32'h3a4762ac),
	.w4(32'h3965da7e),
	.w5(32'h3946b6a9),
	.w6(32'h39d28dfe),
	.w7(32'hb99cfff6),
	.w8(32'hba4355bf),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42d555),
	.w1(32'hbb531437),
	.w2(32'hb94eba54),
	.w3(32'hbb1f5fa0),
	.w4(32'hbb4975c8),
	.w5(32'hbb4ac101),
	.w6(32'hbbc33e93),
	.w7(32'hbbd7c65e),
	.w8(32'hbb97dec9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74f37cf),
	.w1(32'hb9e60552),
	.w2(32'hba544d9f),
	.w3(32'h3b0908a4),
	.w4(32'h3ae7ee56),
	.w5(32'hb93cef9a),
	.w6(32'h3a01858b),
	.w7(32'h3a82896c),
	.w8(32'h3a7d9295),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385c14ad),
	.w1(32'hb924a5ab),
	.w2(32'h399105a1),
	.w3(32'hbaae1fef),
	.w4(32'hba7b1f26),
	.w5(32'hb9d9faa3),
	.w6(32'hbb1fe599),
	.w7(32'hbaa64a3b),
	.w8(32'hb9e10b93),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1a4c9),
	.w1(32'h3b5af6d4),
	.w2(32'h3aad2e3e),
	.w3(32'h3b08110f),
	.w4(32'h3b3a452f),
	.w5(32'hb9ea85b3),
	.w6(32'h3b4df7f1),
	.w7(32'h3b8d62b6),
	.w8(32'h3b150db2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c6fdd9),
	.w1(32'hb98493f5),
	.w2(32'hb796640f),
	.w3(32'hb909ccbf),
	.w4(32'hb8b63a5a),
	.w5(32'h38c5121c),
	.w6(32'hba40c860),
	.w7(32'hba2354ad),
	.w8(32'h388a4915),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac80ef8),
	.w1(32'h3aa89daa),
	.w2(32'h3a6a7cc2),
	.w3(32'h3aeaf51e),
	.w4(32'h3aad6417),
	.w5(32'h3a84d13f),
	.w6(32'h3ae6c6de),
	.w7(32'h3ac665b1),
	.w8(32'h3a90dc83),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9526c9),
	.w1(32'h3a5c98dd),
	.w2(32'hba2ce8bf),
	.w3(32'hba852151),
	.w4(32'hb9a9415d),
	.w5(32'hb91141f7),
	.w6(32'hb9190afc),
	.w7(32'h3a69b9a8),
	.w8(32'hb88417ca),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3926f575),
	.w1(32'h3928b1cc),
	.w2(32'h399c8845),
	.w3(32'h390154fb),
	.w4(32'h3925bc1a),
	.w5(32'h39933975),
	.w6(32'h3969c3b8),
	.w7(32'h39bd37f7),
	.w8(32'h3a06a013),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba103f5b),
	.w1(32'hb9549152),
	.w2(32'h395878f1),
	.w3(32'hbb0d2474),
	.w4(32'hbad50ad0),
	.w5(32'hb95205eb),
	.w6(32'hbb394d66),
	.w7(32'hba9a6270),
	.w8(32'hba18d214),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba484f),
	.w1(32'h3abc296f),
	.w2(32'h3ad962b4),
	.w3(32'h3a979131),
	.w4(32'h3addd717),
	.w5(32'h3a9d8deb),
	.w6(32'h3b19b6fe),
	.w7(32'h3acf2dbe),
	.w8(32'h3a9c0aac),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968fb0b),
	.w1(32'hb9af9268),
	.w2(32'hb9ce6e36),
	.w3(32'h39d2b4a8),
	.w4(32'h39be798e),
	.w5(32'hb8046763),
	.w6(32'h3a6d2485),
	.w7(32'h3a0f9352),
	.w8(32'h3a146a3e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e68a9a),
	.w1(32'hb9371b32),
	.w2(32'hb90a672b),
	.w3(32'hb8a484cf),
	.w4(32'hb883332d),
	.w5(32'hb8937be0),
	.w6(32'hb876cb8b),
	.w7(32'hb7affe08),
	.w8(32'h36be7af3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dcbac5),
	.w1(32'hb717bc1d),
	.w2(32'hb65c0f03),
	.w3(32'h384b8b65),
	.w4(32'h359a3fce),
	.w5(32'hb6bd1d7e),
	.w6(32'h37be8a38),
	.w7(32'hb79ad21f),
	.w8(32'h35c24f1a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1107e5),
	.w1(32'h3a122b6c),
	.w2(32'h3a1c5997),
	.w3(32'hba0ec82e),
	.w4(32'hb9c58f4c),
	.w5(32'h39958a83),
	.w6(32'hba7f5535),
	.w7(32'hb9d87e72),
	.w8(32'hb93de74c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd7546),
	.w1(32'h38378ecd),
	.w2(32'h3921f31f),
	.w3(32'hb89b8512),
	.w4(32'h380115bb),
	.w5(32'h393ccedc),
	.w6(32'hb8dab220),
	.w7(32'hb7f5e643),
	.w8(32'h38c3dc5a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c158d6),
	.w1(32'hb76bcc40),
	.w2(32'hb9aa9b14),
	.w3(32'h39fd160e),
	.w4(32'h377d4625),
	.w5(32'hb8bad2e4),
	.w6(32'h39934a6b),
	.w7(32'h38020a83),
	.w8(32'hb99323cd),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998883e),
	.w1(32'hb8e04798),
	.w2(32'hb895eb11),
	.w3(32'hb9c7ff4a),
	.w4(32'hba404e1c),
	.w5(32'hba067cc5),
	.w6(32'hba97bcc5),
	.w7(32'hba423e3b),
	.w8(32'hb971049e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64dfc73),
	.w1(32'hb861a93d),
	.w2(32'hb8a68751),
	.w3(32'h385fafc5),
	.w4(32'h36d9cde6),
	.w5(32'h37acfa45),
	.w6(32'h38cb3c6e),
	.w7(32'h3876a0e8),
	.w8(32'h38947ae3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1b6bb),
	.w1(32'hb9c583d7),
	.w2(32'hb91517f4),
	.w3(32'hb9a3891f),
	.w4(32'hb97bb40a),
	.w5(32'hb95a1268),
	.w6(32'hb9c56b99),
	.w7(32'hb98995ac),
	.w8(32'hb9985238),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39072ac6),
	.w1(32'h394de2ef),
	.w2(32'h39b02796),
	.w3(32'h38d2ef45),
	.w4(32'h38bdec15),
	.w5(32'h3904bf07),
	.w6(32'hb945ac46),
	.w7(32'h373cf11a),
	.w8(32'h3a1a3b5c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c2e81),
	.w1(32'hba14446e),
	.w2(32'h3a77d42b),
	.w3(32'h39e3861c),
	.w4(32'h3abc883e),
	.w5(32'hb95be296),
	.w6(32'h3984d520),
	.w7(32'hb8f29352),
	.w8(32'h3a8715e9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae81be2),
	.w1(32'h3c305af4),
	.w2(32'hbbc225c2),
	.w3(32'hb9d11723),
	.w4(32'h3b5e8c86),
	.w5(32'hbb78855f),
	.w6(32'h3c04decb),
	.w7(32'hbb18f092),
	.w8(32'hb895ed75),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00f63d),
	.w1(32'hba8a020a),
	.w2(32'hbaad090a),
	.w3(32'hb96fb94c),
	.w4(32'h3aa9203f),
	.w5(32'hba84e1b1),
	.w6(32'hb9d801f5),
	.w7(32'hbaaca4c7),
	.w8(32'h3989e99a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a707acb),
	.w1(32'h3a8f25de),
	.w2(32'h3b172a44),
	.w3(32'h3aa13ee8),
	.w4(32'h3aa11529),
	.w5(32'h3af468e9),
	.w6(32'hba74687b),
	.w7(32'hb8871412),
	.w8(32'h3ab6c7ca),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39755f5e),
	.w1(32'hbb632a57),
	.w2(32'hbad09178),
	.w3(32'hba809c77),
	.w4(32'hba525e37),
	.w5(32'hbac9d095),
	.w6(32'h3a0ee94c),
	.w7(32'hbb7d3704),
	.w8(32'h3b39e2dd),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b7ed1),
	.w1(32'h399a3cd4),
	.w2(32'h3aeaeac8),
	.w3(32'hbb346c2d),
	.w4(32'hbb81b26e),
	.w5(32'h3aafdced),
	.w6(32'h3b775b0a),
	.w7(32'hbb9352bd),
	.w8(32'h3aa1c340),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26dd27),
	.w1(32'hbb3460fe),
	.w2(32'hb932b55b),
	.w3(32'hbaec9889),
	.w4(32'hb96956f1),
	.w5(32'hbb2968a9),
	.w6(32'hbb576e95),
	.w7(32'hb89f5dc6),
	.w8(32'h3b7eff43),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cef5e),
	.w1(32'h3aafd2ae),
	.w2(32'hbb117afa),
	.w3(32'h3b0ea99d),
	.w4(32'hbb01653f),
	.w5(32'hba09bea6),
	.w6(32'h3af6e45d),
	.w7(32'h388b6881),
	.w8(32'h3a87bd36),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad72ed4),
	.w1(32'h3a88b1e9),
	.w2(32'h3b2243c2),
	.w3(32'h3b10c4cd),
	.w4(32'h3b24d3c3),
	.w5(32'h3adc98ea),
	.w6(32'hb9576df5),
	.w7(32'hb985700c),
	.w8(32'hb84972d8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6448f9),
	.w1(32'hb8895e75),
	.w2(32'h39778060),
	.w3(32'hb96dcbe6),
	.w4(32'h3aadd6ba),
	.w5(32'h3a3d5e65),
	.w6(32'hb901a391),
	.w7(32'hb9ad3514),
	.w8(32'hba3f468d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d078e),
	.w1(32'hbb51cc22),
	.w2(32'hbb25f8e8),
	.w3(32'hbaf5838b),
	.w4(32'h3a06e06c),
	.w5(32'hbb019f6b),
	.w6(32'hbb9530b3),
	.w7(32'hbb688bac),
	.w8(32'hbbae41fd),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c750a),
	.w1(32'hbbdee2f7),
	.w2(32'hbbdf1286),
	.w3(32'hbbb657c3),
	.w4(32'hbc351e95),
	.w5(32'hbbe21768),
	.w6(32'hbba74e6a),
	.w7(32'hbbbdf50b),
	.w8(32'h3bd4d787),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8428d8),
	.w1(32'hbb5424fa),
	.w2(32'hbba8bf8c),
	.w3(32'h3a58e102),
	.w4(32'hbb97aa47),
	.w5(32'hbb6919e6),
	.w6(32'h3b019872),
	.w7(32'hbadf0bea),
	.w8(32'hbb3f66f2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921edbd),
	.w1(32'h3a12a5eb),
	.w2(32'hb98b5cb7),
	.w3(32'hbb5691b3),
	.w4(32'hbb27bf45),
	.w5(32'h3af9621d),
	.w6(32'hbba6841c),
	.w7(32'hbb03308f),
	.w8(32'h3847bd92),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fc92b),
	.w1(32'hbc0c104a),
	.w2(32'hbad75073),
	.w3(32'h3b73c63f),
	.w4(32'hba83d197),
	.w5(32'h3b2e5270),
	.w6(32'hbb940c5a),
	.w7(32'hbaac74af),
	.w8(32'h39ee8d60),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78f843),
	.w1(32'h3c4db069),
	.w2(32'h39601219),
	.w3(32'h3b2d0462),
	.w4(32'h3c05d7a3),
	.w5(32'hbb915ada),
	.w6(32'hbb68e7b0),
	.w7(32'h3a6fca0a),
	.w8(32'h3b6013d9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8daaf4),
	.w1(32'h3b802936),
	.w2(32'hbb691df7),
	.w3(32'hba3328db),
	.w4(32'h3b98417d),
	.w5(32'h3748199f),
	.w6(32'h3b0d38c3),
	.w7(32'h3a87d1ad),
	.w8(32'h3ae81ac5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b010926),
	.w1(32'h3a67d0ef),
	.w2(32'h3ac749b1),
	.w3(32'h3b228f56),
	.w4(32'h3a214ee3),
	.w5(32'h3b27cca3),
	.w6(32'hbae4189f),
	.w7(32'h3a6f6f0c),
	.w8(32'h3b8b127e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bf4cb),
	.w1(32'h3a90ca21),
	.w2(32'hbb397758),
	.w3(32'hbb16afd0),
	.w4(32'hbb6b736e),
	.w5(32'hbb8ef75c),
	.w6(32'h3c2c14c2),
	.w7(32'hbb0ccf47),
	.w8(32'hbb717e44),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87c628),
	.w1(32'h3be63322),
	.w2(32'hba1b64c7),
	.w3(32'hba50e7f8),
	.w4(32'h3ac44e42),
	.w5(32'hbb0ec301),
	.w6(32'h3b9de51c),
	.w7(32'h3b1a68c2),
	.w8(32'h3a0ec959),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb143b86),
	.w1(32'hbb0ed7c5),
	.w2(32'hbad401b9),
	.w3(32'h3aeb64d9),
	.w4(32'h3a71050c),
	.w5(32'hbb917575),
	.w6(32'hbb47da5e),
	.w7(32'hba5e13b4),
	.w8(32'h3a85b056),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afeb9ee),
	.w1(32'h3a59cab8),
	.w2(32'h3b4e1fcd),
	.w3(32'h3b252114),
	.w4(32'h3b4f24d0),
	.w5(32'h3bafc2ec),
	.w6(32'h3ae75a16),
	.w7(32'h3b6c1c68),
	.w8(32'h3bbe1426),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae2e8d),
	.w1(32'hb8453e7e),
	.w2(32'hbc264d07),
	.w3(32'hba971349),
	.w4(32'hb8ab2c78),
	.w5(32'hbb8ddf38),
	.w6(32'h3bd14036),
	.w7(32'hbac0f6fd),
	.w8(32'h39e5cd9c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba3eee),
	.w1(32'h3a99c25f),
	.w2(32'h395706f7),
	.w3(32'h3a9c0f55),
	.w4(32'h3b102b20),
	.w5(32'hb81b81be),
	.w6(32'h3adc4cf8),
	.w7(32'hb9a5ed73),
	.w8(32'hb9c359f3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c996d),
	.w1(32'hba71117c),
	.w2(32'hba90c543),
	.w3(32'h3a0dc4e3),
	.w4(32'h3a30893d),
	.w5(32'hb9f71988),
	.w6(32'hb970d2c0),
	.w7(32'hb99ff18a),
	.w8(32'hb83e956e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306eaa),
	.w1(32'hbb349cef),
	.w2(32'hbb27996d),
	.w3(32'hbb0589ee),
	.w4(32'hbab65a1a),
	.w5(32'hbab941be),
	.w6(32'hbb550aaa),
	.w7(32'hbae01c3e),
	.w8(32'hba23346e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fca33),
	.w1(32'hba737e14),
	.w2(32'h3abd4277),
	.w3(32'h3a3eebbe),
	.w4(32'hba2d7b1d),
	.w5(32'hbb25656e),
	.w6(32'h3aa42679),
	.w7(32'hba5ced33),
	.w8(32'h3a872be9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a354ca8),
	.w1(32'h3a1fa2c7),
	.w2(32'h3ae29d7a),
	.w3(32'h3b3a907b),
	.w4(32'h3b6119bb),
	.w5(32'h3b2edd9e),
	.w6(32'h3b495c45),
	.w7(32'h3b1c9873),
	.w8(32'hb7efdf9e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb127f79),
	.w1(32'hba86254b),
	.w2(32'h3b91b8c4),
	.w3(32'h3ab0e30f),
	.w4(32'h3b45dad1),
	.w5(32'h3ba6e322),
	.w6(32'hbbbd685a),
	.w7(32'h3a736895),
	.w8(32'hb9cc4409),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9098171),
	.w1(32'h3938e5ca),
	.w2(32'h3a3d7a9c),
	.w3(32'h3a9329ee),
	.w4(32'h3ae4baa0),
	.w5(32'h39e9b42a),
	.w6(32'h3a898196),
	.w7(32'h3a01b574),
	.w8(32'h3a5ca9aa),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1391a),
	.w1(32'hbaaf9676),
	.w2(32'h3a4a81da),
	.w3(32'hba661ff1),
	.w4(32'h3abfca6d),
	.w5(32'h3a0f9f0b),
	.w6(32'hbaa83142),
	.w7(32'hba981a16),
	.w8(32'hb9f43af0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c6a52),
	.w1(32'h39c94e61),
	.w2(32'h3a2a6f50),
	.w3(32'h3ad9e6f4),
	.w4(32'h3ac95fbd),
	.w5(32'h3992e80b),
	.w6(32'h3a420a70),
	.w7(32'hb8a758dc),
	.w8(32'h3b09d65e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be0340),
	.w1(32'hbb6a2700),
	.w2(32'hb89ea8d3),
	.w3(32'hbaa8c18f),
	.w4(32'hbba54fa5),
	.w5(32'hbbea4cb4),
	.w6(32'hbb441d83),
	.w7(32'hba44bc11),
	.w8(32'h39eb2a2c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904f6f5),
	.w1(32'hbaaf7594),
	.w2(32'hbaa7bbbf),
	.w3(32'h38b7cf39),
	.w4(32'h39abcf7c),
	.w5(32'hba50ddf3),
	.w6(32'h3a8f64f0),
	.w7(32'hbab6eda0),
	.w8(32'hb8e3903a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fdaeb),
	.w1(32'hba06f36a),
	.w2(32'hba97eb7e),
	.w3(32'h3aa5e95f),
	.w4(32'h3ad2ba6f),
	.w5(32'hb9c8fb6d),
	.w6(32'h3a86ead3),
	.w7(32'h3a741f3c),
	.w8(32'h3aab927b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c98b1b),
	.w1(32'hba931cbd),
	.w2(32'hba69ad43),
	.w3(32'h3a9da2e6),
	.w4(32'h3ab0f414),
	.w5(32'hba37cba4),
	.w6(32'hb8bab5c9),
	.w7(32'hba214755),
	.w8(32'hbb2bf0f9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0af3f3),
	.w1(32'hba87f7a4),
	.w2(32'h3bc1e4c1),
	.w3(32'h3af1c145),
	.w4(32'h3b5d4776),
	.w5(32'h3bc8eebb),
	.w6(32'hbbc33490),
	.w7(32'h3ada0619),
	.w8(32'hba8fb301),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43cda3),
	.w1(32'hbb001ffd),
	.w2(32'h3b9f5e14),
	.w3(32'h3ad21ba8),
	.w4(32'h3b56b26d),
	.w5(32'h3b2fb8f8),
	.w6(32'hbb3686e6),
	.w7(32'h3b2b2d07),
	.w8(32'h3afd4d4b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9e1b0),
	.w1(32'h3a1293d6),
	.w2(32'hbb336e22),
	.w3(32'hbac125a1),
	.w4(32'hba916ec8),
	.w5(32'hbaf8b43f),
	.w6(32'hba5357b8),
	.w7(32'hbae47760),
	.w8(32'h3b421d98),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bece8),
	.w1(32'hbb05c836),
	.w2(32'hba960dcb),
	.w3(32'h3bd11664),
	.w4(32'hbae38fd8),
	.w5(32'hbaadfce2),
	.w6(32'hba24f95a),
	.w7(32'hbb4dbbdd),
	.w8(32'h3a6f075f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba002ed7),
	.w1(32'hba546fe8),
	.w2(32'hbae36d53),
	.w3(32'h3ac66ddd),
	.w4(32'h3aa1cf04),
	.w5(32'hba96e3fe),
	.w6(32'hba714458),
	.w7(32'hbad84075),
	.w8(32'h3a757c6a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86d060),
	.w1(32'hbb04b9cc),
	.w2(32'hbad6cafa),
	.w3(32'hbb34a980),
	.w4(32'hb90ff5c2),
	.w5(32'hbb687133),
	.w6(32'hbbd6ecb1),
	.w7(32'hbbbd5972),
	.w8(32'hbb744869),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69824b),
	.w1(32'h3cc033c7),
	.w2(32'hbc2c90f9),
	.w3(32'h3c856fc6),
	.w4(32'hbbfac8de),
	.w5(32'hbbc48007),
	.w6(32'h3caed666),
	.w7(32'h3bef394e),
	.w8(32'h3bb454dc),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a169c77),
	.w1(32'hbad79efd),
	.w2(32'hbabb5b26),
	.w3(32'hbac6eae1),
	.w4(32'hbb121266),
	.w5(32'hbb3adbf0),
	.w6(32'h3a8d0b4b),
	.w7(32'h3a10f4b1),
	.w8(32'h3b688005),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63fc86),
	.w1(32'hb9eb6aac),
	.w2(32'h3905e15c),
	.w3(32'h3b2fbd60),
	.w4(32'h3b614974),
	.w5(32'h3ad5b09b),
	.w6(32'h3abaf89e),
	.w7(32'h3ad64510),
	.w8(32'h3bc54ef0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcccc12),
	.w1(32'h3ad1dde9),
	.w2(32'hbb4d2fe3),
	.w3(32'h3b38a132),
	.w4(32'hbb3a1b11),
	.w5(32'hba712762),
	.w6(32'h3b1b3e50),
	.w7(32'hb8dff280),
	.w8(32'h39c11699),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8452481),
	.w1(32'h3a63d511),
	.w2(32'h3b3571da),
	.w3(32'h3a498bcd),
	.w4(32'h3acd0c74),
	.w5(32'hb9752796),
	.w6(32'h3a08a1f9),
	.w7(32'hba662576),
	.w8(32'h3ba35c39),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c5516),
	.w1(32'h3c1f66dd),
	.w2(32'hbb85f41e),
	.w3(32'hba2149bc),
	.w4(32'hbb464198),
	.w5(32'hbb9d1eea),
	.w6(32'h3c144f59),
	.w7(32'h3b3660e5),
	.w8(32'h3bb8d588),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb86e79),
	.w1(32'h3acd105c),
	.w2(32'hbb3fa784),
	.w3(32'h3b28a7d1),
	.w4(32'hbb28b0a7),
	.w5(32'hba6cda5c),
	.w6(32'h3b0f7832),
	.w7(32'hb89ba5c9),
	.w8(32'h3b96a0df),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ea493),
	.w1(32'h3a80ff21),
	.w2(32'hbb4225db),
	.w3(32'h3b03ba45),
	.w4(32'hbb2738b3),
	.w5(32'hbaa63a71),
	.w6(32'h3ae82907),
	.w7(32'hba130a58),
	.w8(32'h3ba340d9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a656e),
	.w1(32'hb9a438e2),
	.w2(32'hbb2b8935),
	.w3(32'h39dbb6d8),
	.w4(32'hbb2226a4),
	.w5(32'hbb39ca8b),
	.w6(32'h3b4691bf),
	.w7(32'h39e02bea),
	.w8(32'h3b424e50),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69742d),
	.w1(32'h3c7665dd),
	.w2(32'hbb3bdfa8),
	.w3(32'hbb840c1c),
	.w4(32'h3bdfebff),
	.w5(32'hbb854a74),
	.w6(32'h3bdeea7a),
	.w7(32'hbb73242c),
	.w8(32'hba244bda),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14081a),
	.w1(32'h3982f2f7),
	.w2(32'h3973b71c),
	.w3(32'hba000d5e),
	.w4(32'h39b818ca),
	.w5(32'hba44e734),
	.w6(32'hbaff8c34),
	.w7(32'hba569b04),
	.w8(32'hba619c88),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb77ce),
	.w1(32'h3716c99e),
	.w2(32'hbbcc0cc0),
	.w3(32'hba723124),
	.w4(32'hbc166104),
	.w5(32'hbb30616b),
	.w6(32'hbc1a9103),
	.w7(32'h3af8b171),
	.w8(32'h3c3d0c0a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b194a8d),
	.w1(32'hbb5f4b0e),
	.w2(32'hbc12fe1a),
	.w3(32'hbb936139),
	.w4(32'hbc0d6eed),
	.w5(32'hbc1f3b56),
	.w6(32'h3bd27a12),
	.w7(32'h3a474789),
	.w8(32'h3ab6fff4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84fb1f),
	.w1(32'hbb7b5b11),
	.w2(32'h3bd540be),
	.w3(32'hbab273a8),
	.w4(32'hbb2fcd9c),
	.w5(32'hbb21102e),
	.w6(32'hbaf18978),
	.w7(32'h3afb019c),
	.w8(32'h3b115da5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc35638),
	.w1(32'hbbe8420f),
	.w2(32'hbbd09134),
	.w3(32'h3b405682),
	.w4(32'hbc37fb12),
	.w5(32'hbaf3d36e),
	.w6(32'h3bfc825a),
	.w7(32'h3ac3c608),
	.w8(32'hbb1f7371),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabadbd5),
	.w1(32'hb9fbd249),
	.w2(32'h3bae5f2c),
	.w3(32'h3b1622a5),
	.w4(32'h3b573814),
	.w5(32'h3bb4902f),
	.w6(32'hbb986871),
	.w7(32'h3ac4da78),
	.w8(32'h398a95b8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93734d),
	.w1(32'hb95cac05),
	.w2(32'hb89b2a75),
	.w3(32'h3aa1a354),
	.w4(32'h3ab64566),
	.w5(32'hbae8b2dd),
	.w6(32'hba78d870),
	.w7(32'hbb01f84d),
	.w8(32'h3c1a4809),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10cc19),
	.w1(32'hb85d6058),
	.w2(32'hbb5a595c),
	.w3(32'h3a87c766),
	.w4(32'hbb6b2ef3),
	.w5(32'hbb73ed95),
	.w6(32'h3c093029),
	.w7(32'h3988962a),
	.w8(32'h39d588ee),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0e639),
	.w1(32'hbb3ea52b),
	.w2(32'hbb27d687),
	.w3(32'hbb3712a1),
	.w4(32'hbad6a7f9),
	.w5(32'hbac0038f),
	.w6(32'hbb4def95),
	.w7(32'hbb350578),
	.w8(32'hbb16ec53),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9868d74),
	.w1(32'hb9fcd560),
	.w2(32'h3c2aa644),
	.w3(32'h3b94d4ca),
	.w4(32'h3bedcd34),
	.w5(32'h3bee1b6f),
	.w6(32'hbb4b3027),
	.w7(32'h3be44a8b),
	.w8(32'h3c071824),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b322c10),
	.w1(32'hbaa9cc42),
	.w2(32'hbba972f0),
	.w3(32'hba26a5a0),
	.w4(32'hbb8b40ef),
	.w5(32'hbbb19ac6),
	.w6(32'h3b20fdcf),
	.w7(32'hbab48d54),
	.w8(32'h3b062e7c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b3bd3),
	.w1(32'h3a664d5a),
	.w2(32'hba9290ed),
	.w3(32'h3aa0870e),
	.w4(32'hba8905e6),
	.w5(32'hb9b6616f),
	.w6(32'h3a73442d),
	.w7(32'hb7abdb8c),
	.w8(32'h3ba30b7c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed0173),
	.w1(32'hb9eb5470),
	.w2(32'hbc1afc8f),
	.w3(32'h3bfaf370),
	.w4(32'h3aa096e6),
	.w5(32'hbba18b74),
	.w6(32'h3a150121),
	.w7(32'hbb514f62),
	.w8(32'hbb546ac6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb29837),
	.w1(32'hbbf50091),
	.w2(32'hba7b054b),
	.w3(32'hbc638de3),
	.w4(32'hbc1c12ef),
	.w5(32'hbb4b1514),
	.w6(32'hbc414896),
	.w7(32'hbbb5c4dc),
	.w8(32'h3abf1b6b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d14b3),
	.w1(32'hbb6d8c26),
	.w2(32'hbc4a283e),
	.w3(32'h3bbbe786),
	.w4(32'hbabd035c),
	.w5(32'hbbdfd69c),
	.w6(32'hbbcb2e76),
	.w7(32'hbc26c15a),
	.w8(32'h3bdea17f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c397eea),
	.w1(32'h3a157606),
	.w2(32'hbc1d15f3),
	.w3(32'h3c25358c),
	.w4(32'h39579bc4),
	.w5(32'hbc192f15),
	.w6(32'hb8fecd52),
	.w7(32'hbc107f66),
	.w8(32'h3b5c37e3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77da2c),
	.w1(32'hbb9b6e73),
	.w2(32'hbc2ec4fc),
	.w3(32'h39045922),
	.w4(32'hbb005468),
	.w5(32'hbba0c8fd),
	.w6(32'hbbeea0d5),
	.w7(32'hbbfef9b7),
	.w8(32'h3be46c14),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab736d9),
	.w1(32'h3ba49e8a),
	.w2(32'h3abe1574),
	.w3(32'h3bed424e),
	.w4(32'h3c882848),
	.w5(32'h3c5818c6),
	.w6(32'hbb4e5c43),
	.w7(32'hbb194bac),
	.w8(32'hbc24928a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40bf9a),
	.w1(32'hbb9d2d60),
	.w2(32'h3a31d361),
	.w3(32'hbc40f4da),
	.w4(32'hbc171689),
	.w5(32'h39893abd),
	.w6(32'hbb8059fb),
	.w7(32'hbb12c978),
	.w8(32'hbca42b5b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdee0cd),
	.w1(32'h3824959d),
	.w2(32'h3d20f474),
	.w3(32'hbce8241a),
	.w4(32'hbc02a892),
	.w5(32'h3cd6e030),
	.w6(32'h3acca6ce),
	.w7(32'h3d096a43),
	.w8(32'h3c0133cd),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19c9c5),
	.w1(32'hbac0c89e),
	.w2(32'hbc4fd5c5),
	.w3(32'h3be7647b),
	.w4(32'hba3bcf8b),
	.w5(32'hbc256e59),
	.w6(32'hbac4b7ac),
	.w7(32'hbc2ff1b6),
	.w8(32'h3b9ccdc5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be348f3),
	.w1(32'hb87b83a2),
	.w2(32'hbc017c52),
	.w3(32'h3bd11e4f),
	.w4(32'h3a9e2665),
	.w5(32'hbba8d78f),
	.w6(32'hba619076),
	.w7(32'hbbcc7fba),
	.w8(32'h3c1a6640),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b1205),
	.w1(32'hbb0c96c4),
	.w2(32'hbc937404),
	.w3(32'h3c4bfb06),
	.w4(32'h3af0d345),
	.w5(32'hbc2d72f0),
	.w6(32'hbb9af908),
	.w7(32'hbc71ffe9),
	.w8(32'hbc716267),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23cb1e),
	.w1(32'hbc0309f0),
	.w2(32'hbd25c367),
	.w3(32'hbc0278c2),
	.w4(32'hbc5c60da),
	.w5(32'hbd12324a),
	.w6(32'hbc94ebdc),
	.w7(32'hbd0ba9d4),
	.w8(32'hbc4d34aa),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac680d),
	.w1(32'h396f4843),
	.w2(32'h3cbbdab9),
	.w3(32'hbc9b355d),
	.w4(32'hbb3bebe9),
	.w5(32'h3c81757f),
	.w6(32'h3ba9bdde),
	.w7(32'h3cc8ff5b),
	.w8(32'h3c0750ea),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31bfe8),
	.w1(32'hbba5b6ea),
	.w2(32'h3b59e084),
	.w3(32'h3bdefe99),
	.w4(32'h393d3989),
	.w5(32'h3bd3f1d2),
	.w6(32'hbb9c43d1),
	.w7(32'hbb7cf480),
	.w8(32'h3a6b13b0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09cb57),
	.w1(32'hbba39454),
	.w2(32'hbba0c5de),
	.w3(32'hbb6a7916),
	.w4(32'hbaefa9c6),
	.w5(32'h3abb81ad),
	.w6(32'hbc032b8d),
	.w7(32'hbb631c4b),
	.w8(32'hb9d0513f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91cd71),
	.w1(32'hbbc65b28),
	.w2(32'hbc024f0e),
	.w3(32'hbbf006e2),
	.w4(32'hbbde1a2d),
	.w5(32'hbb7de957),
	.w6(32'hbbedfe96),
	.w7(32'hbbfdcaef),
	.w8(32'h3c24c601),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca6e48),
	.w1(32'hb92d155b),
	.w2(32'hbaf7f872),
	.w3(32'h397facc5),
	.w4(32'h3bc62d9a),
	.w5(32'h3a678a57),
	.w6(32'h3bfeacb9),
	.w7(32'h38f8b081),
	.w8(32'h3c2d8468),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95d764),
	.w1(32'hb9c7874e),
	.w2(32'h3aa67dfc),
	.w3(32'h3c4b8748),
	.w4(32'hbba53df2),
	.w5(32'hbafa839e),
	.w6(32'hbbc5f076),
	.w7(32'hbb0c13ad),
	.w8(32'hbb04bea9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdac216),
	.w1(32'hbb4da6d4),
	.w2(32'hbc2ca139),
	.w3(32'hbb6028e3),
	.w4(32'hbb788d89),
	.w5(32'hbc305999),
	.w6(32'hbb1bdfdd),
	.w7(32'hbc25bd79),
	.w8(32'h3bf458aa),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a34290),
	.w1(32'h3bbb894a),
	.w2(32'h39dc1357),
	.w3(32'hbb57d809),
	.w4(32'h3bd19c5a),
	.w5(32'h3c2b7ca7),
	.w6(32'h3b36f0b6),
	.w7(32'h3b6cb3be),
	.w8(32'h3af67c30),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75c3bd),
	.w1(32'hbaee91a2),
	.w2(32'hbc29e8c1),
	.w3(32'h3b19657f),
	.w4(32'h3a91e363),
	.w5(32'hbb4a1461),
	.w6(32'hbb42f76e),
	.w7(32'hbc0e4d72),
	.w8(32'h3c22d677),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55fe60),
	.w1(32'h3a1b457f),
	.w2(32'hbc2fb699),
	.w3(32'h3c31f4e0),
	.w4(32'h3b5248f4),
	.w5(32'hbc2844e1),
	.w6(32'h3a994073),
	.w7(32'hbbe90909),
	.w8(32'h3b23884c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb982f60),
	.w1(32'h3b797f84),
	.w2(32'hbc32dd24),
	.w3(32'hbb5421ed),
	.w4(32'h3c0aafdb),
	.w5(32'hbc2b77c1),
	.w6(32'h3b862206),
	.w7(32'hbc33d417),
	.w8(32'h3b6552db),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule