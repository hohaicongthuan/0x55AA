module layer_10_featuremap_29(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91b4a5),
	.w1(32'hbc0a4dca),
	.w2(32'h3bfce5a9),
	.w3(32'h3c1f33c2),
	.w4(32'hbc9b5c5e),
	.w5(32'hbba8b144),
	.w6(32'h3bba5f38),
	.w7(32'hbb884aba),
	.w8(32'hbca0d3c9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f7dc7),
	.w1(32'hbc363cf5),
	.w2(32'hb87abc32),
	.w3(32'h3d068f55),
	.w4(32'hbbb4bc17),
	.w5(32'hbbd23c55),
	.w6(32'hbb7032ad),
	.w7(32'h3c5c9332),
	.w8(32'hbb059146),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24d9f7),
	.w1(32'hbc3e1c6f),
	.w2(32'hb7cf1111),
	.w3(32'hbcab3013),
	.w4(32'hbd1fa0c9),
	.w5(32'h3ac9d303),
	.w6(32'hbbf4fd66),
	.w7(32'hbcf3dabd),
	.w8(32'h3a856ba6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc232334),
	.w1(32'h3c229b0e),
	.w2(32'hbbc4263c),
	.w3(32'hbc3cbe36),
	.w4(32'h3c71b06e),
	.w5(32'hbc8ebfe3),
	.w6(32'hbb61001a),
	.w7(32'h3c03f6e3),
	.w8(32'hbb7a32dd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c3378),
	.w1(32'hbbf9110c),
	.w2(32'h3b0d139f),
	.w3(32'hba84fda0),
	.w4(32'hbc12da9c),
	.w5(32'h3cb86069),
	.w6(32'hbc2610c1),
	.w7(32'hbb98dfe6),
	.w8(32'h3c77d0d1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2a3a6),
	.w1(32'h3c10f475),
	.w2(32'h3b03ad18),
	.w3(32'h3add9d18),
	.w4(32'h3c646d0f),
	.w5(32'hbab49167),
	.w6(32'h3bc1e3d8),
	.w7(32'h3c769f68),
	.w8(32'h3acdd3af),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2622e6),
	.w1(32'h3bb93bb6),
	.w2(32'h3be78320),
	.w3(32'h3a2eabc6),
	.w4(32'h3b687163),
	.w5(32'h3c00a8da),
	.w6(32'h3b4e0013),
	.w7(32'h3becbdaa),
	.w8(32'h3b689b88),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba894335),
	.w1(32'hbc80c37e),
	.w2(32'hbb318dd7),
	.w3(32'hbb114e3a),
	.w4(32'hbc05e8da),
	.w5(32'h3c12ec8b),
	.w6(32'hbab91440),
	.w7(32'hba77855b),
	.w8(32'h3bcba231),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa15eaa),
	.w1(32'h3a718e07),
	.w2(32'h3ae15c03),
	.w3(32'hbc1e831b),
	.w4(32'hbb8ec40f),
	.w5(32'hbbde24f0),
	.w6(32'hbbecbad4),
	.w7(32'hbb9e507a),
	.w8(32'h3a81ddf3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0e96f),
	.w1(32'hbab53d7d),
	.w2(32'hbae2e4d1),
	.w3(32'hbbcaabfb),
	.w4(32'hb6d6ca85),
	.w5(32'hbb462dbc),
	.w6(32'hbbb5fb49),
	.w7(32'h3bf56f84),
	.w8(32'hbb8ac1b7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02fd0a),
	.w1(32'h3a1ac08f),
	.w2(32'hbb6f82d1),
	.w3(32'h3ad6a5b9),
	.w4(32'h3b38744f),
	.w5(32'hbbaa8701),
	.w6(32'hbb2d5c6e),
	.w7(32'h39331825),
	.w8(32'hbbd12109),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf78fb2),
	.w1(32'h3b53def9),
	.w2(32'h3b2a9a4d),
	.w3(32'hbc4bdb90),
	.w4(32'h3c487229),
	.w5(32'h3b6a533a),
	.w6(32'hbaef8cc4),
	.w7(32'h3c16e58a),
	.w8(32'h3b96a745),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb32b3d),
	.w1(32'hbad3a6c6),
	.w2(32'h3b4c7f8f),
	.w3(32'h3be27b08),
	.w4(32'hbba8bea2),
	.w5(32'h3ac75547),
	.w6(32'h3c11f8d2),
	.w7(32'hba94b2d3),
	.w8(32'h3b92341e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5076a1),
	.w1(32'hbb91f0dc),
	.w2(32'hbc17081f),
	.w3(32'hbb6ea0d6),
	.w4(32'hbb43bcb1),
	.w5(32'h3bb9671b),
	.w6(32'h3ae01e44),
	.w7(32'hbbe912c2),
	.w8(32'h3b8a7207),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae45d64),
	.w1(32'h3c05187d),
	.w2(32'hb9e026fa),
	.w3(32'hbc98a3a9),
	.w4(32'hbb814b18),
	.w5(32'hbb25518a),
	.w6(32'hbc4f68a8),
	.w7(32'h3b8a1cea),
	.w8(32'h3aae565c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2f3a8),
	.w1(32'h3b0e07b5),
	.w2(32'h39a55b85),
	.w3(32'h3b075106),
	.w4(32'h3b2580a8),
	.w5(32'hba5e6fdf),
	.w6(32'h3aeb136a),
	.w7(32'h3abbfe8a),
	.w8(32'hba291a5b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ad441),
	.w1(32'h3af6e5ee),
	.w2(32'h3b15c7dd),
	.w3(32'h3b57b4e0),
	.w4(32'h3a3f9fec),
	.w5(32'h3b1e4b3b),
	.w6(32'hb74841c2),
	.w7(32'h3a928cff),
	.w8(32'h3b1286a3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdedf11),
	.w1(32'hba15a285),
	.w2(32'h3a801671),
	.w3(32'hbc0cdf76),
	.w4(32'hbadde3e9),
	.w5(32'h3b76ad85),
	.w6(32'hbb3a4c3d),
	.w7(32'h385474d3),
	.w8(32'h3acae46a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb03238),
	.w1(32'h3b26fc9a),
	.w2(32'h3b17d92c),
	.w3(32'h3ad05335),
	.w4(32'hbbeabb33),
	.w5(32'h3c11150b),
	.w6(32'h3b3eab71),
	.w7(32'hbb0d137b),
	.w8(32'h389ad061),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc391ebb),
	.w1(32'h3b44fed5),
	.w2(32'hbb34df23),
	.w3(32'hbc5926a4),
	.w4(32'hba0fb51c),
	.w5(32'hbb4f259d),
	.w6(32'hbb7f6272),
	.w7(32'hbbbddb29),
	.w8(32'hbb608e9d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84f1f2),
	.w1(32'h3ad4e10b),
	.w2(32'h3a2d4c78),
	.w3(32'hbb5648b8),
	.w4(32'h37c2264d),
	.w5(32'hbaa58493),
	.w6(32'hbbac445b),
	.w7(32'h3b59f6cf),
	.w8(32'h3a37eabc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50e66d),
	.w1(32'h3ba15e08),
	.w2(32'h3b86c17b),
	.w3(32'hb9f6c883),
	.w4(32'h3c163248),
	.w5(32'h3b399cf6),
	.w6(32'h3c2a9996),
	.w7(32'h389c0908),
	.w8(32'hbb268188),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e442b),
	.w1(32'hbc219c76),
	.w2(32'hbb342168),
	.w3(32'hbbfe091c),
	.w4(32'hbc18db2c),
	.w5(32'h3a854767),
	.w6(32'hbbc6996b),
	.w7(32'hbb83998e),
	.w8(32'hba48aea3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0da52),
	.w1(32'h39f9f151),
	.w2(32'h3a656443),
	.w3(32'h3bb70ab3),
	.w4(32'h3ae93e1d),
	.w5(32'h3b1a16b8),
	.w6(32'h3b8107f6),
	.w7(32'h3b7672c4),
	.w8(32'h3b52869f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad31c2b),
	.w1(32'h3b16b820),
	.w2(32'hbbd7b3da),
	.w3(32'hb960790b),
	.w4(32'h3ab498e5),
	.w5(32'hbb255346),
	.w6(32'hb95be7e1),
	.w7(32'hbbaba94c),
	.w8(32'hbbd536ec),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd65d07),
	.w1(32'hbc33db9d),
	.w2(32'h3aa71684),
	.w3(32'h3c22ed3b),
	.w4(32'hbab21779),
	.w5(32'hbbb41282),
	.w6(32'h3b98b8ca),
	.w7(32'h3b1db360),
	.w8(32'h3af6f1ed),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c5378),
	.w1(32'h3a5870d9),
	.w2(32'h3a88e4b8),
	.w3(32'h3b3c6de9),
	.w4(32'h3bcc3ab0),
	.w5(32'hba326cbb),
	.w6(32'hbc86934e),
	.w7(32'h3c4b4273),
	.w8(32'h39c13698),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba95a6a),
	.w1(32'h3a142177),
	.w2(32'hbb6eab5b),
	.w3(32'h3b63ec06),
	.w4(32'hbaf0c3fa),
	.w5(32'h3a846a4c),
	.w6(32'h3b4d57e9),
	.w7(32'h3a180b2c),
	.w8(32'h3c526234),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00cc30),
	.w1(32'hbb495c4e),
	.w2(32'hb99bd8f9),
	.w3(32'h3aabd02d),
	.w4(32'hbb904264),
	.w5(32'hbc80114f),
	.w6(32'hbb939396),
	.w7(32'h3bbb07b7),
	.w8(32'hbc386d81),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8e85f),
	.w1(32'hbb689159),
	.w2(32'hbb2e9d79),
	.w3(32'hbc12d79d),
	.w4(32'hbc6f8918),
	.w5(32'hbb0acb96),
	.w6(32'hbc79fa74),
	.w7(32'hbc7d48c4),
	.w8(32'hbb3c2feb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96fd9b),
	.w1(32'hbba22a9f),
	.w2(32'h3b48ebff),
	.w3(32'hbb9a4597),
	.w4(32'hbb9d5c6b),
	.w5(32'h3c398d07),
	.w6(32'hbbe9c4d4),
	.w7(32'hbba04068),
	.w8(32'hbaf2fa0f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bf90a),
	.w1(32'hbbd0a1b3),
	.w2(32'h3a573845),
	.w3(32'hbb5d8b4b),
	.w4(32'hbbea3fe4),
	.w5(32'h3a5f9ed8),
	.w6(32'hbc1a22cb),
	.w7(32'h3a3c8b38),
	.w8(32'h3a4afc95),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05073e),
	.w1(32'hbc1e0095),
	.w2(32'hbba3750e),
	.w3(32'hbc970c1b),
	.w4(32'hbc9ea785),
	.w5(32'hbb975efd),
	.w6(32'hbc8976f3),
	.w7(32'hbc056938),
	.w8(32'hbb31076c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd67e61),
	.w1(32'h3b3c69f9),
	.w2(32'h3cd47548),
	.w3(32'h3b76917f),
	.w4(32'hbaf8a7cb),
	.w5(32'h3c9179d9),
	.w6(32'hbae384d7),
	.w7(32'hba9a1d08),
	.w8(32'hbb2bf025),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0925c0),
	.w1(32'h3ce97822),
	.w2(32'hbb10381d),
	.w3(32'h3a63513e),
	.w4(32'h3d6646a3),
	.w5(32'hb87a9159),
	.w6(32'h3d079aec),
	.w7(32'h3ca58d3e),
	.w8(32'h3a823cc2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b295783),
	.w1(32'hbb5b61b0),
	.w2(32'h3c8d812c),
	.w3(32'h3aa7749b),
	.w4(32'h39d7376e),
	.w5(32'h3c4fcc6e),
	.w6(32'hb8b36f6c),
	.w7(32'hba0d4b04),
	.w8(32'hbc24b2fe),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb98efc),
	.w1(32'h3b6092bb),
	.w2(32'hbba6607a),
	.w3(32'hbcfc3245),
	.w4(32'h3c5d7981),
	.w5(32'hbb0466a0),
	.w6(32'hb99227f4),
	.w7(32'h3c175cb4),
	.w8(32'hbb1f3de3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc86aa5),
	.w1(32'hbb35aa9a),
	.w2(32'hbc60281d),
	.w3(32'h3acdf2a8),
	.w4(32'hbaadc0de),
	.w5(32'h3b9e7abf),
	.w6(32'h3a54932d),
	.w7(32'h3ab507f7),
	.w8(32'h3b5b999b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7569e),
	.w1(32'hbc040569),
	.w2(32'hbc1f55b2),
	.w3(32'h3c330ff0),
	.w4(32'h3ab716ea),
	.w5(32'hbb78917d),
	.w6(32'h3c2d254e),
	.w7(32'h3b534d63),
	.w8(32'hba27de08),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4ac11),
	.w1(32'hbaaf1fc5),
	.w2(32'hba2a51f4),
	.w3(32'h3c3227de),
	.w4(32'hbba6e2f6),
	.w5(32'h3aac1a5e),
	.w6(32'h3b8c5e79),
	.w7(32'hbc880120),
	.w8(32'h3adb51c8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7dc17),
	.w1(32'h3a3bf32c),
	.w2(32'hbc5a8bf7),
	.w3(32'h3ab725a4),
	.w4(32'hbbcae8b7),
	.w5(32'hbbcfe535),
	.w6(32'h3bab266f),
	.w7(32'hbc017ff0),
	.w8(32'hbb9c3ab2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b942a85),
	.w1(32'h3bb06861),
	.w2(32'hbc28dc45),
	.w3(32'h3c166c80),
	.w4(32'hbbba46ff),
	.w5(32'hbb219e0b),
	.w6(32'hb94ed74c),
	.w7(32'hbc071156),
	.w8(32'hbb2a5a8d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18644b),
	.w1(32'hbc6045d4),
	.w2(32'hb9c81109),
	.w3(32'hbc1aba27),
	.w4(32'hbc429f4f),
	.w5(32'h3afffca9),
	.w6(32'hbcb4dbf5),
	.w7(32'hba75889b),
	.w8(32'h3a1156a4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7178d8),
	.w1(32'hbbfc58b3),
	.w2(32'hbbd51e78),
	.w3(32'hbae3a16f),
	.w4(32'hbb85b9b9),
	.w5(32'hbc58dd35),
	.w6(32'hbb15cd9c),
	.w7(32'hbaff7cc7),
	.w8(32'h3beefda3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95143e),
	.w1(32'hba8a2c77),
	.w2(32'h3b8dcecb),
	.w3(32'h3c96d648),
	.w4(32'hbce187cb),
	.w5(32'h3c87c22e),
	.w6(32'h3b3a59b4),
	.w7(32'hbc9d1aac),
	.w8(32'h3ce9dc29),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cce2587),
	.w1(32'hbca6ed6a),
	.w2(32'hbc20003a),
	.w3(32'h3c21d523),
	.w4(32'hbc1e43b6),
	.w5(32'hbc2fea3d),
	.w6(32'hbc852d6e),
	.w7(32'h3cb5e56c),
	.w8(32'hbc4546b7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09fb4c),
	.w1(32'hbc8ea078),
	.w2(32'h3c521ed8),
	.w3(32'hbcdc287b),
	.w4(32'hbd215989),
	.w5(32'h3bc844b8),
	.w6(32'hbcad2f19),
	.w7(32'hbce34d32),
	.w8(32'hbc6c6755),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf01780),
	.w1(32'h3c603e0d),
	.w2(32'hbb23963d),
	.w3(32'hbced191f),
	.w4(32'h3cc9f13f),
	.w5(32'hba76ef25),
	.w6(32'h3c0b0eef),
	.w7(32'h3ca3ad3b),
	.w8(32'hbb02312a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e59f9),
	.w1(32'hbbef839b),
	.w2(32'hbaeba5d7),
	.w3(32'hbb802c02),
	.w4(32'hbb6d3c3d),
	.w5(32'hbb53fb36),
	.w6(32'hbb7990fd),
	.w7(32'hb9bff412),
	.w8(32'h3a402585),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba54bc),
	.w1(32'hbb9d1905),
	.w2(32'hbb90c975),
	.w3(32'h3c0ff5da),
	.w4(32'h3a27d5bc),
	.w5(32'h3ac7b851),
	.w6(32'hbbc37d89),
	.w7(32'hbb1529cc),
	.w8(32'hbba6ff6e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc50df0),
	.w1(32'h3d1b4caa),
	.w2(32'hbc09a823),
	.w3(32'h3ce8f48e),
	.w4(32'h3d1a95f3),
	.w5(32'hbc3fc48f),
	.w6(32'h3cfba281),
	.w7(32'h3c3448cd),
	.w8(32'hbb5858b4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08708d),
	.w1(32'hba0f7c0a),
	.w2(32'h3a9d96a0),
	.w3(32'h3ce495b8),
	.w4(32'hbc2ee300),
	.w5(32'hbbbd82f9),
	.w6(32'h3c8a5f9a),
	.w7(32'hbc03b823),
	.w8(32'hbbc7ee7c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc133d50),
	.w1(32'h3c23426f),
	.w2(32'h3bee5b8f),
	.w3(32'h3c2e1b80),
	.w4(32'h3bcd3500),
	.w5(32'h39e06928),
	.w6(32'h3c877231),
	.w7(32'hbbabcd36),
	.w8(32'hbc00e344),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8cd90),
	.w1(32'h3c43d45d),
	.w2(32'h3bb660ff),
	.w3(32'hbc252346),
	.w4(32'h3b4c86ca),
	.w5(32'h3ab88776),
	.w6(32'hbac3d5b8),
	.w7(32'h3be15cb7),
	.w8(32'h3b3db1ac),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d3803),
	.w1(32'hbb39e143),
	.w2(32'h3c07f539),
	.w3(32'h3b080bb5),
	.w4(32'hbbadedc8),
	.w5(32'h3b79b54f),
	.w6(32'h3b67c6c4),
	.w7(32'hbbfe79c5),
	.w8(32'h3bb3dde0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e87e7),
	.w1(32'h3bcabe07),
	.w2(32'h3b42cc58),
	.w3(32'h3bc1fd64),
	.w4(32'h3baeccbc),
	.w5(32'h3bdcbf92),
	.w6(32'h3c6626b3),
	.w7(32'h3bcbbad3),
	.w8(32'h3b6a13a7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75019e),
	.w1(32'hbc9a3109),
	.w2(32'hbc29f9c8),
	.w3(32'hbc726ada),
	.w4(32'hbc95cd95),
	.w5(32'hbc2cd682),
	.w6(32'hbc56bc01),
	.w7(32'hbc2ecfbc),
	.w8(32'hbbb8e987),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0880da),
	.w1(32'h3b432c32),
	.w2(32'h3ad82853),
	.w3(32'h39ff6df6),
	.w4(32'hbb10c9a0),
	.w5(32'h3a1f51ea),
	.w6(32'hbbb6b378),
	.w7(32'hbabbdbc3),
	.w8(32'hbb4ccb9c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f50c9),
	.w1(32'hb9b59e73),
	.w2(32'hbb9678d4),
	.w3(32'h3bc76c7f),
	.w4(32'hbb44d499),
	.w5(32'hb97feb41),
	.w6(32'hbb4fc5d9),
	.w7(32'hbc0fc5b5),
	.w8(32'hb9fb311d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e8693),
	.w1(32'h3aed3b77),
	.w2(32'hb8d05e3a),
	.w3(32'h3bdc0a31),
	.w4(32'hbb5d4311),
	.w5(32'hbb91e470),
	.w6(32'hbb18da68),
	.w7(32'hba8e259e),
	.w8(32'hb9d39daf),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac370d2),
	.w1(32'h3a1a80c6),
	.w2(32'h3b69ab88),
	.w3(32'hba90809a),
	.w4(32'h3c0a8705),
	.w5(32'h3c86565c),
	.w6(32'hbb9749b6),
	.w7(32'hba8116fd),
	.w8(32'h3bd789a6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc90d11),
	.w1(32'hb8e1db2e),
	.w2(32'h3a9e9990),
	.w3(32'h3c45cf3f),
	.w4(32'hb98a3ca7),
	.w5(32'h3c12a4b2),
	.w6(32'h3c39688f),
	.w7(32'h3c05ff4e),
	.w8(32'h3b9e651e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe4bfa),
	.w1(32'hbb245ffc),
	.w2(32'hbb93b1a1),
	.w3(32'hbb413bae),
	.w4(32'h3b8619df),
	.w5(32'hbb8a2459),
	.w6(32'h3b2c176c),
	.w7(32'h3b933eb2),
	.w8(32'hb9a4eb77),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdde42),
	.w1(32'hba58e259),
	.w2(32'h3b3d681a),
	.w3(32'hb9cd3a91),
	.w4(32'hbc1037de),
	.w5(32'h3bee4e89),
	.w6(32'h3b0704f7),
	.w7(32'hbb4978cf),
	.w8(32'h3bd718bb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c266409),
	.w1(32'hbaf9ec51),
	.w2(32'h3b85cfd0),
	.w3(32'hbabdb2e8),
	.w4(32'h3a26a55f),
	.w5(32'h3ba52977),
	.w6(32'hbb0a57f6),
	.w7(32'h3aa7a97f),
	.w8(32'h3b8d7747),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b818cfb),
	.w1(32'h3b2241e9),
	.w2(32'hb9d7feda),
	.w3(32'h3aed5d81),
	.w4(32'hba383093),
	.w5(32'hba1b0570),
	.w6(32'hb9add2d0),
	.w7(32'h3a61c9e1),
	.w8(32'hb9da154f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc13826),
	.w1(32'hbbe45627),
	.w2(32'hbbfa8179),
	.w3(32'hbaaec2b3),
	.w4(32'hbc0661b0),
	.w5(32'hbba53a1e),
	.w6(32'hbaf1c165),
	.w7(32'hb95a90ce),
	.w8(32'hbc39a5e2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66d350),
	.w1(32'h3cae5dbc),
	.w2(32'hbbaf4ac6),
	.w3(32'h3cba0409),
	.w4(32'h3c03dced),
	.w5(32'hbb161bcf),
	.w6(32'h3cddc6ea),
	.w7(32'hbc0bac28),
	.w8(32'hbbfa78fe),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac309b),
	.w1(32'hbb5024fe),
	.w2(32'h3b21d990),
	.w3(32'hbb65d9d5),
	.w4(32'h3ac8a48a),
	.w5(32'h39743859),
	.w6(32'h3bc10821),
	.w7(32'hbb7da43c),
	.w8(32'h3a61106c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93e71b),
	.w1(32'h3ab2daea),
	.w2(32'h3c530334),
	.w3(32'hbbcdc6e4),
	.w4(32'h3a3c4818),
	.w5(32'h3c4fdacf),
	.w6(32'hbbb3217f),
	.w7(32'h38e31a91),
	.w8(32'h3b202057),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07ea28),
	.w1(32'hbb27d19e),
	.w2(32'hbb15c3b8),
	.w3(32'hbb2e8127),
	.w4(32'h3b837b8f),
	.w5(32'hbbae2424),
	.w6(32'h3b0ffaeb),
	.w7(32'hbaa23330),
	.w8(32'h3a0bb472),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b933f2c),
	.w1(32'hbb63f4b0),
	.w2(32'hbbc06241),
	.w3(32'h3c092e0f),
	.w4(32'hbc1c5345),
	.w5(32'hbbc1490c),
	.w6(32'h3b986cdf),
	.w7(32'hbbe5e83e),
	.w8(32'hbc58ad06),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ce844),
	.w1(32'hbae0e807),
	.w2(32'hbae227ba),
	.w3(32'hbc2ebfb3),
	.w4(32'hbc852c21),
	.w5(32'h3c6c30e8),
	.w6(32'hbc27d707),
	.w7(32'hbc3aa946),
	.w8(32'h3bfc9d8d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f2f4a),
	.w1(32'hbd09a14b),
	.w2(32'h3afb1476),
	.w3(32'hbbe1e5f0),
	.w4(32'hbcea549a),
	.w5(32'h3b23c968),
	.w6(32'hbca9df7b),
	.w7(32'h3952ed0e),
	.w8(32'h3a3afd63),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39adbd25),
	.w1(32'hbbd9dbd9),
	.w2(32'hbbe291db),
	.w3(32'hbb06e9ab),
	.w4(32'hbbc376c5),
	.w5(32'hbbf5b423),
	.w6(32'hbb5be810),
	.w7(32'hbabf5def),
	.w8(32'hbbb040bb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81ab6c),
	.w1(32'hba9bc06a),
	.w2(32'h3bacdf97),
	.w3(32'h3b98be69),
	.w4(32'hbbcbed3d),
	.w5(32'h3b9e4720),
	.w6(32'hbab8b297),
	.w7(32'hbb9b5ae3),
	.w8(32'h3bd2cb27),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6a740),
	.w1(32'hbbc47090),
	.w2(32'h3c37e4b8),
	.w3(32'hbc5126a7),
	.w4(32'hbb4e988c),
	.w5(32'h3be39eb9),
	.w6(32'hbc0c83dd),
	.w7(32'hbbe8a63e),
	.w8(32'h3afba921),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b755ab6),
	.w1(32'hbb20fb4a),
	.w2(32'hbb09bad2),
	.w3(32'h3aaad2b9),
	.w4(32'h3bb40c83),
	.w5(32'hbaf3a3bc),
	.w6(32'h3b98903b),
	.w7(32'h3b6bc0a9),
	.w8(32'h3bc1a7df),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0735e9),
	.w1(32'hbbc13140),
	.w2(32'h398b395e),
	.w3(32'hbbcad11b),
	.w4(32'hbc3eeb1a),
	.w5(32'hbac3fa36),
	.w6(32'hbb3f64ca),
	.w7(32'hbc1d2fa5),
	.w8(32'hba8115d6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05bbec),
	.w1(32'h39f156bb),
	.w2(32'h3bf964c4),
	.w3(32'hbb0fad8b),
	.w4(32'hb9d763cd),
	.w5(32'h3a035716),
	.w6(32'h37de13b5),
	.w7(32'h37d1aee5),
	.w8(32'hbaa29aac),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef0263),
	.w1(32'hb9f3e7f8),
	.w2(32'h3b71a6b8),
	.w3(32'hbbc29b5d),
	.w4(32'h3b96bcb4),
	.w5(32'h3b0330b0),
	.w6(32'h3bc65241),
	.w7(32'hbabcd5fd),
	.w8(32'h3aae7389),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a0965),
	.w1(32'hbb39b76f),
	.w2(32'h3cabc786),
	.w3(32'hbaa7c5c4),
	.w4(32'hbbdaa7b7),
	.w5(32'h3c637bd0),
	.w6(32'hbb69b71f),
	.w7(32'hbb6e43dd),
	.w8(32'hbc3a9f7d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc561158),
	.w1(32'h3cd13906),
	.w2(32'hb9f3f6f5),
	.w3(32'hbc5d07c5),
	.w4(32'h3cde9efa),
	.w5(32'hbab3fd09),
	.w6(32'h3c7c74db),
	.w7(32'h3beefbab),
	.w8(32'hbba3ab98),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eec07),
	.w1(32'hbc2cc2c6),
	.w2(32'h3b8b345c),
	.w3(32'hbc558134),
	.w4(32'hbc5d2899),
	.w5(32'h3abdaf73),
	.w6(32'hbc0e9720),
	.w7(32'hbaaeed63),
	.w8(32'h3c5fbf58),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64357f),
	.w1(32'hbbb3a200),
	.w2(32'hbc226445),
	.w3(32'hbbaf87ba),
	.w4(32'hbc828af7),
	.w5(32'h3c5632fc),
	.w6(32'hbc04f191),
	.w7(32'hbc16e03b),
	.w8(32'h3cc6ac23),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2c1f0b),
	.w1(32'hbc5bfd57),
	.w2(32'h3bd7f518),
	.w3(32'h3d36606e),
	.w4(32'hbce286e6),
	.w5(32'h3b931872),
	.w6(32'h3adce80b),
	.w7(32'hbc42bc54),
	.w8(32'h3bed2da8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb83fda),
	.w1(32'hbbaf61c5),
	.w2(32'hbb988c57),
	.w3(32'h3b900b18),
	.w4(32'hbc23c774),
	.w5(32'hbbaacba1),
	.w6(32'hbb387f7b),
	.w7(32'hbc28db6a),
	.w8(32'h3794e9a1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5baf6f),
	.w1(32'hbb743e2e),
	.w2(32'hba973413),
	.w3(32'hb7f313e6),
	.w4(32'hbb8ce251),
	.w5(32'hbc759a6d),
	.w6(32'hbaafaad3),
	.w7(32'hbb9a7b3f),
	.w8(32'hbc83d6be),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a9793),
	.w1(32'h3c658324),
	.w2(32'h3bfc5069),
	.w3(32'h3c10d1ef),
	.w4(32'h3c0768d8),
	.w5(32'h3bfc1c2a),
	.w6(32'h3c2a8e10),
	.w7(32'hbc4ee75a),
	.w8(32'hbc3093b3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e67ec),
	.w1(32'h3b7654fa),
	.w2(32'h3be7c496),
	.w3(32'hbc4e1cd9),
	.w4(32'h3bc86885),
	.w5(32'h3be4d308),
	.w6(32'h3b2afad2),
	.w7(32'hbae6ddfe),
	.w8(32'hba501043),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4de0ba),
	.w1(32'h3ba4398f),
	.w2(32'hba4780ea),
	.w3(32'hbbf19330),
	.w4(32'h3b90029d),
	.w5(32'h3a3f7aa0),
	.w6(32'hbc06ae1e),
	.w7(32'h3c2dfb64),
	.w8(32'h388a8f34),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aec2b),
	.w1(32'h3b852cf2),
	.w2(32'hb92f4a2d),
	.w3(32'h3a2cb84d),
	.w4(32'h3c2a1dcc),
	.w5(32'hb7bd67c9),
	.w6(32'h3b01cba0),
	.w7(32'h3bba8977),
	.w8(32'h3b24794f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6241ab),
	.w1(32'h3b77be6f),
	.w2(32'hba58e583),
	.w3(32'h3973561a),
	.w4(32'hb73c2126),
	.w5(32'hbae0a0e7),
	.w6(32'hb8a82bd1),
	.w7(32'hbacd9496),
	.w8(32'hbb79d80a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89a36e),
	.w1(32'hbb260934),
	.w2(32'h3ae81bfb),
	.w3(32'hbb0ae4d6),
	.w4(32'h39b55bde),
	.w5(32'hbc137421),
	.w6(32'hbb664038),
	.w7(32'hbb6b8fe6),
	.w8(32'hbc044cc0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7cd35c),
	.w1(32'hbac8c6c6),
	.w2(32'hbae0fdac),
	.w3(32'hbc221002),
	.w4(32'hbbb6bf16),
	.w5(32'hbc12d520),
	.w6(32'hbb4f8460),
	.w7(32'hbc07f666),
	.w8(32'hbc2a79e6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc90420),
	.w1(32'hbc15ebad),
	.w2(32'h3a8455f4),
	.w3(32'hbbb5d24e),
	.w4(32'hbc595b20),
	.w5(32'hb9d64f24),
	.w6(32'hbc165b57),
	.w7(32'h3b04758e),
	.w8(32'hbb95d4f0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c6c9a),
	.w1(32'h3c12f418),
	.w2(32'h3aeffaff),
	.w3(32'hbbc7a66b),
	.w4(32'hbb812556),
	.w5(32'h3bd21f94),
	.w6(32'hbb7e2e7f),
	.w7(32'h3a247e65),
	.w8(32'h3b61804f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee59d3),
	.w1(32'hbb8fab00),
	.w2(32'h3b5666b8),
	.w3(32'hbc40ca8f),
	.w4(32'hbbf12c3e),
	.w5(32'hbaa01311),
	.w6(32'h3a159474),
	.w7(32'h3c18653a),
	.w8(32'h3a81b458),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06da5a),
	.w1(32'hbb4cad56),
	.w2(32'h3c505087),
	.w3(32'h3bea4540),
	.w4(32'hbb95f82f),
	.w5(32'h3be3ad16),
	.w6(32'hbb7d829d),
	.w7(32'hbb077d87),
	.w8(32'h3b185d20),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a645c55),
	.w1(32'hbb28b51e),
	.w2(32'h3bc87d77),
	.w3(32'hbb9e5c9e),
	.w4(32'h3b5b7878),
	.w5(32'h3be8b20a),
	.w6(32'h3ab5830f),
	.w7(32'h3bd1cbec),
	.w8(32'h3c2ad29f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf83eb0),
	.w1(32'h3b0b4a64),
	.w2(32'h3c1d28bd),
	.w3(32'h3b5ef646),
	.w4(32'h3c12b853),
	.w5(32'h3c7658f5),
	.w6(32'h3aa3f7e0),
	.w7(32'h3c00b1a3),
	.w8(32'h3c88346e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ed4ba),
	.w1(32'hbb61b1f7),
	.w2(32'hbb6ce601),
	.w3(32'h3c139bef),
	.w4(32'h3bcd36d0),
	.w5(32'hba33f0b7),
	.w6(32'hbb8f2953),
	.w7(32'h3c6cc26e),
	.w8(32'h3bab2e26),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20e1f6),
	.w1(32'hbbad46d4),
	.w2(32'h3c10e7e0),
	.w3(32'h3bd1faf7),
	.w4(32'hbc880998),
	.w5(32'h3b97275e),
	.w6(32'hbbd0cb71),
	.w7(32'hbc3d2697),
	.w8(32'hbbb53a21),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cfc23),
	.w1(32'h3a95c72b),
	.w2(32'h3bb595f0),
	.w3(32'hbc3c1f33),
	.w4(32'hbb6f4b69),
	.w5(32'hbbc2ace0),
	.w6(32'hbba4146e),
	.w7(32'h3801fdcc),
	.w8(32'h3a85b08f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0329e),
	.w1(32'h3b81b159),
	.w2(32'h3a6d571f),
	.w3(32'h3c4d3938),
	.w4(32'h3c0b9123),
	.w5(32'h3a68cc2d),
	.w6(32'h3c1ad04b),
	.w7(32'hbba3beb7),
	.w8(32'h3bd9d96d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38b54b),
	.w1(32'h3b5fa914),
	.w2(32'hba8481ea),
	.w3(32'h3bcb2f17),
	.w4(32'hbbcab567),
	.w5(32'h38ecb9a6),
	.w6(32'h3bd6bb10),
	.w7(32'hbc2bca72),
	.w8(32'h3bbd841a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96c629),
	.w1(32'h3a82c70c),
	.w2(32'h3bd0b68d),
	.w3(32'h3b20d17a),
	.w4(32'hbacfd3da),
	.w5(32'hbb37dcc2),
	.w6(32'hb9699098),
	.w7(32'hbbc90ebf),
	.w8(32'hbbba6828),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc102d1f),
	.w1(32'hbb9fa4df),
	.w2(32'h3be17eec),
	.w3(32'hbbf8d57e),
	.w4(32'h3a56467c),
	.w5(32'h3b3e15b5),
	.w6(32'hbbdf565c),
	.w7(32'h3babee4b),
	.w8(32'h3a80f58a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6653bf),
	.w1(32'hbc10c7c1),
	.w2(32'hbb3b3701),
	.w3(32'hbc25ed5a),
	.w4(32'hbc7da7bd),
	.w5(32'h3c8f1a19),
	.w6(32'hbba697eb),
	.w7(32'hbc6715e6),
	.w8(32'h3c1b4f08),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9568e0),
	.w1(32'hbb9304b8),
	.w2(32'h3ba231f2),
	.w3(32'h3c312e31),
	.w4(32'hb99135d7),
	.w5(32'h3c18e3cc),
	.w6(32'hbadb23a2),
	.w7(32'h3c8ff1be),
	.w8(32'h3b406ea1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6bb2f),
	.w1(32'h3a86d2db),
	.w2(32'h3b3ad821),
	.w3(32'hbb0f10f7),
	.w4(32'h3bb35fbf),
	.w5(32'h3b8d425f),
	.w6(32'h3b83a54a),
	.w7(32'h3c2e7373),
	.w8(32'hbb7c2837),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fe054),
	.w1(32'h3c83f988),
	.w2(32'h3b8a86b7),
	.w3(32'hb928cdc5),
	.w4(32'h3c1c57ef),
	.w5(32'h3c6e5129),
	.w6(32'h3c3af58e),
	.w7(32'hbc3c727a),
	.w8(32'h3b4bf6c1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eea811),
	.w1(32'hbb76cccf),
	.w2(32'h3bfe452e),
	.w3(32'hbc5527b0),
	.w4(32'h3cc23ff6),
	.w5(32'h3c3886d8),
	.w6(32'h3a4297f9),
	.w7(32'h3d129504),
	.w8(32'hbb16ebbb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b47a8),
	.w1(32'hbc3fafa4),
	.w2(32'hbb5633a9),
	.w3(32'hbbe8419b),
	.w4(32'hbc2cbd80),
	.w5(32'hbc8a4184),
	.w6(32'hbc81a324),
	.w7(32'h3baca49f),
	.w8(32'hbbf181bb),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc39ec1),
	.w1(32'h3bc66a4e),
	.w2(32'hbaa3be11),
	.w3(32'h3c2e0436),
	.w4(32'hbc027032),
	.w5(32'hb9ddf228),
	.w6(32'h3b5e7686),
	.w7(32'hbcaa4177),
	.w8(32'h3b71b601),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e5051),
	.w1(32'h3ace10fd),
	.w2(32'hbb3dec62),
	.w3(32'h3a9681c0),
	.w4(32'h3b0f85db),
	.w5(32'hbbd38642),
	.w6(32'h3b5d217c),
	.w7(32'h3bc0d569),
	.w8(32'hbb70f896),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eb270),
	.w1(32'h3b0522c8),
	.w2(32'h3b4780cb),
	.w3(32'hbb2871a9),
	.w4(32'hbba8addb),
	.w5(32'h3b463a8f),
	.w6(32'h3a342b7f),
	.w7(32'hbb2025eb),
	.w8(32'h3b1aef45),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c2726),
	.w1(32'h3bbe8993),
	.w2(32'hbb9d2992),
	.w3(32'h3b28799c),
	.w4(32'hba2dd13d),
	.w5(32'hbc17a3d7),
	.w6(32'h3b08132a),
	.w7(32'h3b8b041b),
	.w8(32'hbba6f2f6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a9d8c),
	.w1(32'hbb591e23),
	.w2(32'h3c0db02c),
	.w3(32'hbad3d1be),
	.w4(32'hbc4d2a84),
	.w5(32'h3c82a938),
	.w6(32'hbc13f8fb),
	.w7(32'h3a5f26d6),
	.w8(32'h3c9d3d3d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90e136),
	.w1(32'h3b7ebd5b),
	.w2(32'hbba46e75),
	.w3(32'h3bf8f95f),
	.w4(32'h3b7c7814),
	.w5(32'hbb278ed3),
	.w6(32'h3a673d55),
	.w7(32'h3c617db8),
	.w8(32'h3b8c590e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f3369),
	.w1(32'hbadd12bc),
	.w2(32'hba514746),
	.w3(32'h3b3f9d54),
	.w4(32'hbb886ebb),
	.w5(32'hb9233748),
	.w6(32'hbaf8d6ed),
	.w7(32'h3bb9ba22),
	.w8(32'hb9b5ed06),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f890d2),
	.w1(32'hbae1040e),
	.w2(32'hbb6520fa),
	.w3(32'hba9da68e),
	.w4(32'hbb3e7662),
	.w5(32'hbb9aac08),
	.w6(32'hbad828b4),
	.w7(32'hbad7b6cb),
	.w8(32'hbb6affb7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b656e),
	.w1(32'h3ae0425e),
	.w2(32'hbc32a996),
	.w3(32'h3b0f5ff7),
	.w4(32'h3b036e5f),
	.w5(32'hbcc172c7),
	.w6(32'h3a4c679b),
	.w7(32'h382ca308),
	.w8(32'hbc881609),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87f26b),
	.w1(32'h39e31554),
	.w2(32'h3bd9783b),
	.w3(32'hbbe1e16a),
	.w4(32'hbc7ef111),
	.w5(32'h3c10fdcf),
	.w6(32'h3af576f9),
	.w7(32'hbc6f3485),
	.w8(32'h3ba0b215),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae2d6e),
	.w1(32'hbb6ba500),
	.w2(32'h3b1841bd),
	.w3(32'hbb3a3471),
	.w4(32'hbb5910d0),
	.w5(32'hbc31155f),
	.w6(32'hbba3f491),
	.w7(32'h3a3007cc),
	.w8(32'h3b51a245),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b89e4),
	.w1(32'h3c041672),
	.w2(32'h3bcb73e9),
	.w3(32'hb94087a7),
	.w4(32'h3c5f4a6b),
	.w5(32'hbc085074),
	.w6(32'hbb0ece67),
	.w7(32'h3bdaa308),
	.w8(32'hbcafe2f7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc731f3b),
	.w1(32'h3caf8241),
	.w2(32'hbbc779cc),
	.w3(32'h3c257756),
	.w4(32'h3ccbf368),
	.w5(32'hbc2884ac),
	.w6(32'h3c83cf80),
	.w7(32'h3ac38350),
	.w8(32'hbc19da17),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41b087),
	.w1(32'h3c12a6a1),
	.w2(32'hbc298cbe),
	.w3(32'h3cc141d0),
	.w4(32'h3bf893f7),
	.w5(32'hbc484f9b),
	.w6(32'h3c83f837),
	.w7(32'hbafec342),
	.w8(32'hbbb33079),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b948c50),
	.w1(32'h3b9ca4ae),
	.w2(32'hbb9245d6),
	.w3(32'h3ba58f8b),
	.w4(32'h3af43fc1),
	.w5(32'hbb9f7e8f),
	.w6(32'h3be1da10),
	.w7(32'h3bd42ea5),
	.w8(32'hbbf540f4),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f47d7),
	.w1(32'hbab662e5),
	.w2(32'h3a4565ef),
	.w3(32'h3a083a45),
	.w4(32'hbc357f40),
	.w5(32'h3c99ac63),
	.w6(32'h3b353880),
	.w7(32'hbc43ef36),
	.w8(32'h3b5564d5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bbec7),
	.w1(32'hbcd77308),
	.w2(32'hbb58c0db),
	.w3(32'hbcaf887e),
	.w4(32'hba0778b6),
	.w5(32'h3ad69b31),
	.w6(32'hbcb844b6),
	.w7(32'h3c419385),
	.w8(32'h3bc6198a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b560d4c),
	.w1(32'hbbb4fa35),
	.w2(32'hbb2a0970),
	.w3(32'h3bc7961e),
	.w4(32'hbb888ba3),
	.w5(32'hbb85748f),
	.w6(32'hbc08ff62),
	.w7(32'h3bd0307a),
	.w8(32'h3bc1dbc6),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfad0ec),
	.w1(32'hbc023795),
	.w2(32'hbc2a1110),
	.w3(32'hbc011818),
	.w4(32'hbc645272),
	.w5(32'hbc2fe830),
	.w6(32'hbcbedf3a),
	.w7(32'hbbd8e327),
	.w8(32'hbb635588),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4aff21),
	.w1(32'hbcaba08a),
	.w2(32'h3b562b25),
	.w3(32'h3b5d682a),
	.w4(32'hbce334be),
	.w5(32'h3af4845d),
	.w6(32'hbc5968ee),
	.w7(32'hbbc5a425),
	.w8(32'h3aea9d09),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bc767),
	.w1(32'hbb1a7984),
	.w2(32'hb9a5c1b9),
	.w3(32'hba25ce8e),
	.w4(32'hbb467624),
	.w5(32'h3a980e9b),
	.w6(32'hba973934),
	.w7(32'h39a924e5),
	.w8(32'hbaa1ebda),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c294285),
	.w1(32'h3bb8751c),
	.w2(32'h3b57c0c4),
	.w3(32'h3b9187e7),
	.w4(32'hbb99519a),
	.w5(32'h39a4ee41),
	.w6(32'h39919a64),
	.w7(32'hbbf4856a),
	.w8(32'h3bc106d6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2b2cb),
	.w1(32'hbb51d505),
	.w2(32'hba5775e6),
	.w3(32'h3aef58e4),
	.w4(32'hbc0b693d),
	.w5(32'hbad39b02),
	.w6(32'hbc03004f),
	.w7(32'hb7b5b681),
	.w8(32'h3ae7cc08),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ad11e),
	.w1(32'h3c5eb76f),
	.w2(32'h3adf39c3),
	.w3(32'h3b08575f),
	.w4(32'h3c3eb174),
	.w5(32'h3a4f559d),
	.w6(32'h3bf89560),
	.w7(32'h3bfa6072),
	.w8(32'h3a39fa29),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb013d79),
	.w1(32'h3b387592),
	.w2(32'hb9bb2618),
	.w3(32'h38f2202f),
	.w4(32'h3b4d39b7),
	.w5(32'hbbb8fe36),
	.w6(32'h3a3e771c),
	.w7(32'h3b02694a),
	.w8(32'hbbb892a2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4be4a),
	.w1(32'hbc0ce381),
	.w2(32'h3ac2fc7d),
	.w3(32'hbb00e046),
	.w4(32'hbc11da5a),
	.w5(32'hba1f3a69),
	.w6(32'hbc56be31),
	.w7(32'hbafa13b4),
	.w8(32'h3a1a049c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06b066),
	.w1(32'hb9bed7a0),
	.w2(32'h3b0a066d),
	.w3(32'hbaf01bd3),
	.w4(32'h3ab03cc2),
	.w5(32'hba7ebb28),
	.w6(32'hba1f6c8d),
	.w7(32'h3a928c82),
	.w8(32'hba8f79cf),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab26266),
	.w1(32'hb9a55007),
	.w2(32'h3c7e4035),
	.w3(32'hba7f55fe),
	.w4(32'h3b94f866),
	.w5(32'h3bd0d9f2),
	.w6(32'hbb0f0c7b),
	.w7(32'hbb66273d),
	.w8(32'h3b44b845),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd08b61),
	.w1(32'h3bdff1d9),
	.w2(32'h3b9772d5),
	.w3(32'hbc084ee9),
	.w4(32'h3b8d8f36),
	.w5(32'hbb07d22a),
	.w6(32'hbbc96738),
	.w7(32'h3c0174e4),
	.w8(32'h39efbaf1),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3719d),
	.w1(32'hb934e806),
	.w2(32'h3ab4c6f4),
	.w3(32'hbb98aa20),
	.w4(32'h3a247120),
	.w5(32'h3a251a3a),
	.w6(32'hbb4e57a3),
	.w7(32'h3af235f6),
	.w8(32'h3994b4b7),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf978a7),
	.w1(32'h3a1e84f7),
	.w2(32'h3bee459d),
	.w3(32'hb740b20b),
	.w4(32'h3a7d8ce2),
	.w5(32'h3afb1d97),
	.w6(32'h39cca3cf),
	.w7(32'hba9c1659),
	.w8(32'hbab4904f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bfd27),
	.w1(32'h3b84a810),
	.w2(32'hbb0f95d2),
	.w3(32'hbc17d40f),
	.w4(32'h3bcc1746),
	.w5(32'h3a3eb93c),
	.w6(32'hbc1fd925),
	.w7(32'h3c48ccec),
	.w8(32'hbad8b9d3),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31918b),
	.w1(32'hbb9c2aaa),
	.w2(32'h3bddc507),
	.w3(32'h3b1a3c0a),
	.w4(32'hbb138b41),
	.w5(32'h3c21a420),
	.w6(32'h39bd2603),
	.w7(32'hbb223912),
	.w8(32'h3c1a5c60),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb51dcf),
	.w1(32'hbbba8b10),
	.w2(32'h3c0bfc2a),
	.w3(32'h3bbca799),
	.w4(32'h3b4ba74f),
	.w5(32'h3ba916d3),
	.w6(32'h3b308cc4),
	.w7(32'h3c7a8620),
	.w8(32'hb9c8f285),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f42e6),
	.w1(32'hba13abae),
	.w2(32'h3c5dffb6),
	.w3(32'hbbd469d0),
	.w4(32'hbb4a86be),
	.w5(32'h3c8e1e8e),
	.w6(32'hbb1e2e83),
	.w7(32'hbb7e2125),
	.w8(32'h3c9a4d8f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7594c6),
	.w1(32'h3bb2380c),
	.w2(32'hba821407),
	.w3(32'h3c860968),
	.w4(32'h3be1d17f),
	.w5(32'h37e6e3c7),
	.w6(32'h3c3eedf6),
	.w7(32'h3c5b9ef5),
	.w8(32'hbb385914),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95ad81),
	.w1(32'hbaabaf46),
	.w2(32'hbbc14e24),
	.w3(32'hbc0aa5ef),
	.w4(32'h3b301491),
	.w5(32'hbbfd6aa0),
	.w6(32'hbbd83440),
	.w7(32'h3b6f26aa),
	.w8(32'hbbaadaae),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed2d4e),
	.w1(32'h3b7e7e8d),
	.w2(32'hbb0d0c06),
	.w3(32'h3a20f4bf),
	.w4(32'hba929263),
	.w5(32'hbb0a278c),
	.w6(32'hbaee1196),
	.w7(32'hbb6da754),
	.w8(32'hbacb233c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb806e20),
	.w1(32'h3b123e8a),
	.w2(32'hbc329c00),
	.w3(32'h3bf1ab82),
	.w4(32'h3a914e81),
	.w5(32'hbbe4efc2),
	.w6(32'h3b5f53d1),
	.w7(32'h39637c0e),
	.w8(32'hbc026fbd),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc422cd2),
	.w1(32'hbc8fd3f5),
	.w2(32'h3ba5b0d1),
	.w3(32'hbcf73fc7),
	.w4(32'hbc9cda95),
	.w5(32'h3a27203f),
	.w6(32'hbc990e99),
	.w7(32'hbbcd99c1),
	.w8(32'h3af0ddae),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff63ba),
	.w1(32'hbb0511bf),
	.w2(32'hbc422061),
	.w3(32'hbc446f78),
	.w4(32'h39f5e662),
	.w5(32'hbc2e63cd),
	.w6(32'h3b5a540d),
	.w7(32'hbb238aaa),
	.w8(32'hbc058757),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4b0e0),
	.w1(32'h3be7d736),
	.w2(32'h3b6a757b),
	.w3(32'h3d1d8843),
	.w4(32'h3c9e5f18),
	.w5(32'hbb09332e),
	.w6(32'h3c91dd7f),
	.w7(32'h3c38eb78),
	.w8(32'hbb3da1c8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfac4fe),
	.w1(32'h3c456a05),
	.w2(32'hbb15d1d6),
	.w3(32'h3bb21ad3),
	.w4(32'h3c7e8e35),
	.w5(32'h3b75575b),
	.w6(32'hba697652),
	.w7(32'h3be108ab),
	.w8(32'h3c415084),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba608055),
	.w1(32'hba49dc47),
	.w2(32'hbb9242d9),
	.w3(32'hbc037c42),
	.w4(32'hbbd58594),
	.w5(32'hbc274582),
	.w6(32'h3bd03df8),
	.w7(32'hbb10fe5e),
	.w8(32'hb995926a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a8799),
	.w1(32'h3b0f4727),
	.w2(32'h3b5b0e31),
	.w3(32'hbaf61d1f),
	.w4(32'h3bf42562),
	.w5(32'hbb05b1a6),
	.w6(32'h3bdeb1ca),
	.w7(32'h3c6836aa),
	.w8(32'hbb410a06),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a746277),
	.w1(32'hb8b792d5),
	.w2(32'hbc02f5ac),
	.w3(32'h39ed90f4),
	.w4(32'h3b01f20e),
	.w5(32'h39b7f4a4),
	.w6(32'hba9331fe),
	.w7(32'hb9dab82d),
	.w8(32'hba8771d0),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1beda),
	.w1(32'h3899b79a),
	.w2(32'h3d251c05),
	.w3(32'h3c023f54),
	.w4(32'h3bf4ed73),
	.w5(32'h3d05f033),
	.w6(32'h3b0d744d),
	.w7(32'h3b5119d9),
	.w8(32'h3ceda6cb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c079004),
	.w1(32'hbbe9066c),
	.w2(32'h3be8f24c),
	.w3(32'hbcb63618),
	.w4(32'hbd25ec09),
	.w5(32'h3b872bf2),
	.w6(32'hbc743462),
	.w7(32'hbcc698a7),
	.w8(32'h3bd1ba25),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc32470),
	.w1(32'h3baad98a),
	.w2(32'h3c05cef1),
	.w3(32'h3aec2a8d),
	.w4(32'h3a6e76a6),
	.w5(32'h3c099260),
	.w6(32'h3b34934f),
	.w7(32'h3b6dad39),
	.w8(32'h3b281e61),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc024eec),
	.w1(32'hbc92f5f4),
	.w2(32'hbb447516),
	.w3(32'hbc8c4318),
	.w4(32'hbcf3fd0b),
	.w5(32'h3b898f6f),
	.w6(32'hbc92fdf1),
	.w7(32'hbce225f1),
	.w8(32'h3af86f41),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bcb05),
	.w1(32'hbbdafa02),
	.w2(32'h3d572873),
	.w3(32'h3b0e84d3),
	.w4(32'hbb055e6c),
	.w5(32'h3d11c29f),
	.w6(32'h3a499638),
	.w7(32'hbab83ae2),
	.w8(32'h3d0badf8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b332719),
	.w1(32'hbca3148f),
	.w2(32'hba3b45d9),
	.w3(32'hbcf887ef),
	.w4(32'hbd658094),
	.w5(32'hbb7be687),
	.w6(32'hbc9c7b9f),
	.w7(32'hbd09a0be),
	.w8(32'hbc16b970),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e3910),
	.w1(32'hbb6049f0),
	.w2(32'h3a96e7cb),
	.w3(32'hba95396a),
	.w4(32'hbb0bd0ee),
	.w5(32'hb9f217c7),
	.w6(32'hbb27c2cb),
	.w7(32'h3ba1f306),
	.w8(32'h3bc7b521),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14e53c),
	.w1(32'h3b877c68),
	.w2(32'h3afeef42),
	.w3(32'h3bad1bae),
	.w4(32'h3baa9999),
	.w5(32'h3aff4b0e),
	.w6(32'h3c04af59),
	.w7(32'h3c0b2db1),
	.w8(32'hbbadb45e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3798ca6e),
	.w1(32'hb9b9cd3f),
	.w2(32'hbbd2e2f3),
	.w3(32'hba964d0e),
	.w4(32'hb8aaa96c),
	.w5(32'hbb89846e),
	.w6(32'h3b117f84),
	.w7(32'hbb0c9992),
	.w8(32'hbb2760ce),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927567f),
	.w1(32'h3a6ba5f8),
	.w2(32'h3b06d633),
	.w3(32'hbb7ef2f4),
	.w4(32'hb9612230),
	.w5(32'h3b13137b),
	.w6(32'h3b4ce60e),
	.w7(32'h3b156177),
	.w8(32'h396b28f4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b671bba),
	.w1(32'h3b1e58f6),
	.w2(32'hbd19c1b2),
	.w3(32'h3b175595),
	.w4(32'h3b802cc9),
	.w5(32'hbd0b6df9),
	.w6(32'hbab3ba88),
	.w7(32'h3b41eb26),
	.w8(32'hbd143bfa),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1395f),
	.w1(32'h3d0167cb),
	.w2(32'hbb15bb07),
	.w3(32'h3d507ca5),
	.w4(32'h3d9cf505),
	.w5(32'hbae000ff),
	.w6(32'h3d04821c),
	.w7(32'h3d5006e7),
	.w8(32'hbb55b02d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa773c7),
	.w1(32'h3bad9e1b),
	.w2(32'hbb54f397),
	.w3(32'hbb836d3c),
	.w4(32'h3c12fc0b),
	.w5(32'hbad21fe3),
	.w6(32'hb9b09efd),
	.w7(32'h3c06e74f),
	.w8(32'hba39e5e9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60a40a),
	.w1(32'h3b2f6516),
	.w2(32'hba7a0095),
	.w3(32'h3b4c1c1e),
	.w4(32'h3aa74636),
	.w5(32'hbbcae059),
	.w6(32'h3a06c503),
	.w7(32'hbabdd72e),
	.w8(32'hba33f7cd),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4b0b7),
	.w1(32'h3bfe8461),
	.w2(32'hbb106d6c),
	.w3(32'hbb20a7e9),
	.w4(32'h3bb4e523),
	.w5(32'h3a106b15),
	.w6(32'hbb7dad7d),
	.w7(32'h3adf3df9),
	.w8(32'hba24adae),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21f39a),
	.w1(32'h3bcf2cb5),
	.w2(32'h3c1c8c9b),
	.w3(32'hbb1933ce),
	.w4(32'h3a2a7022),
	.w5(32'h3c33d2af),
	.w6(32'h3b64bfc5),
	.w7(32'hba58d2d0),
	.w8(32'h3be4e584),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba504d56),
	.w1(32'hbc370f21),
	.w2(32'hbb8de522),
	.w3(32'hbc2b1e07),
	.w4(32'hbcb8421d),
	.w5(32'hbbf9c9f2),
	.w6(32'hbc4e5203),
	.w7(32'hbcbb2630),
	.w8(32'hbc0de2a0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba60695),
	.w1(32'hba218690),
	.w2(32'h3add6e97),
	.w3(32'h3a94411e),
	.w4(32'h3a572269),
	.w5(32'h3aed83c5),
	.w6(32'hbb6303b9),
	.w7(32'h3b4326a7),
	.w8(32'h3b39aa97),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa6352),
	.w1(32'hbb4a0236),
	.w2(32'hbb4d6d7d),
	.w3(32'h3b4cf82f),
	.w4(32'h39b22d3f),
	.w5(32'hbc0aa618),
	.w6(32'hbae5b12d),
	.w7(32'hb9a6b34c),
	.w8(32'hbba13a72),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f0cbe),
	.w1(32'h3b5af888),
	.w2(32'hba80ee2c),
	.w3(32'hbb667342),
	.w4(32'h3b5dc6ca),
	.w5(32'h389d5e3c),
	.w6(32'hbb7e4e09),
	.w7(32'h3b22f885),
	.w8(32'h3ae4f9b7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86af7e),
	.w1(32'hbbf967eb),
	.w2(32'hba71bb97),
	.w3(32'hbb66fc62),
	.w4(32'hba91eb69),
	.w5(32'hbbb34b05),
	.w6(32'hba699e7c),
	.w7(32'hbae9efc5),
	.w8(32'hbb121f72),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fbf27),
	.w1(32'h3aca8e56),
	.w2(32'hbbab2bf7),
	.w3(32'hbb7d743a),
	.w4(32'h3b72a80f),
	.w5(32'h3b10f1f4),
	.w6(32'h3afaf9fa),
	.w7(32'h3adc0d52),
	.w8(32'h3b9eecc1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a6acb),
	.w1(32'h37363241),
	.w2(32'hbb09371f),
	.w3(32'hbbe3666f),
	.w4(32'hbb61c610),
	.w5(32'hbb220c35),
	.w6(32'h3a5f10fd),
	.w7(32'hbc004b80),
	.w8(32'hbaaee133),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3206b2),
	.w1(32'h37d70a69),
	.w2(32'h392c0ec2),
	.w3(32'h3a240a22),
	.w4(32'h3bf62601),
	.w5(32'h3b065554),
	.w6(32'hb9e1010d),
	.w7(32'h395fc987),
	.w8(32'hbab42176),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eff9f),
	.w1(32'h3c06b22f),
	.w2(32'hbaf6032a),
	.w3(32'h3bb1c5ca),
	.w4(32'h3bc4e097),
	.w5(32'hbc1b55c8),
	.w6(32'h3b13a76d),
	.w7(32'h3baf3733),
	.w8(32'hbbe44f9d),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf375c5),
	.w1(32'hbbc17dff),
	.w2(32'hbb93fb36),
	.w3(32'hbac9bbef),
	.w4(32'hbb90da5f),
	.w5(32'hbc236490),
	.w6(32'hba48ce68),
	.w7(32'hbb66a3b1),
	.w8(32'hbc37b1d2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a2cec),
	.w1(32'h3c3b6de5),
	.w2(32'hbb208957),
	.w3(32'h3bb39660),
	.w4(32'h3c8a42a5),
	.w5(32'hbc339a69),
	.w6(32'h3ba47005),
	.w7(32'h3cc7dd77),
	.w8(32'hbbc643e5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa49ba5),
	.w1(32'h3bab1d25),
	.w2(32'h3b7c1d63),
	.w3(32'hbba00191),
	.w4(32'hba854639),
	.w5(32'h378aacb3),
	.w6(32'hbb72b2be),
	.w7(32'hbb34581a),
	.w8(32'h3ba5af4f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dcc86),
	.w1(32'hbc0b0d2a),
	.w2(32'hbab215ce),
	.w3(32'hbb4c5c70),
	.w4(32'hbbcf75d5),
	.w5(32'hbb1c63cf),
	.w6(32'h3b95a6e9),
	.w7(32'hba616fec),
	.w8(32'hbb56d584),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a299089),
	.w1(32'h3b3bdcb1),
	.w2(32'h3b16ed68),
	.w3(32'hb924a1a4),
	.w4(32'h3b040e89),
	.w5(32'hbae1351b),
	.w6(32'hbad07bb0),
	.w7(32'h3aadaf7f),
	.w8(32'hbb8e563c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b789057),
	.w1(32'hbb7b2e4e),
	.w2(32'hbafeb5c9),
	.w3(32'h3af08ca1),
	.w4(32'hbb624bfa),
	.w5(32'hbb92351d),
	.w6(32'h3bcd9690),
	.w7(32'hbbb3686f),
	.w8(32'hbb58af78),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c953b),
	.w1(32'h3b998722),
	.w2(32'hbb4ccc78),
	.w3(32'hbaefafb6),
	.w4(32'h3b0e2a92),
	.w5(32'h399e9d96),
	.w6(32'hbae3256c),
	.w7(32'h3ba30258),
	.w8(32'hbab4124b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2aea98),
	.w1(32'hbb81d114),
	.w2(32'h3af717d7),
	.w3(32'h39040ac7),
	.w4(32'hbb31f695),
	.w5(32'h3b86cca5),
	.w6(32'hbb820ba5),
	.w7(32'hbbe22fef),
	.w8(32'h3b89cba7),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b952cb1),
	.w1(32'h3c07381a),
	.w2(32'hbd58e545),
	.w3(32'h3b83963d),
	.w4(32'h3c1041cb),
	.w5(32'hbd5c5d22),
	.w6(32'h3bd1920a),
	.w7(32'h3c0e6710),
	.w8(32'hbd434abb),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95aca8),
	.w1(32'h3d35c80b),
	.w2(32'hbb7b5bc1),
	.w3(32'h3d746879),
	.w4(32'h3dcbaae0),
	.w5(32'hbb3200df),
	.w6(32'h3d26acf1),
	.w7(32'h3d9484d4),
	.w8(32'hbaef2b68),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25f2b9),
	.w1(32'h3bcbdb42),
	.w2(32'hba522851),
	.w3(32'hbacc3f68),
	.w4(32'h3b7a59e2),
	.w5(32'hbb866dc6),
	.w6(32'h3ad0e565),
	.w7(32'h3b5f7a90),
	.w8(32'hbadd87b8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53df9e),
	.w1(32'hbae53054),
	.w2(32'hbb8eebd9),
	.w3(32'hbb170559),
	.w4(32'hbb43e73a),
	.w5(32'h3a08d9c0),
	.w6(32'h3af4e5f8),
	.w7(32'hbaa18158),
	.w8(32'h3a329ab7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf41c82),
	.w1(32'hbb391876),
	.w2(32'h3b8ef378),
	.w3(32'h3c209153),
	.w4(32'h3bb79624),
	.w5(32'hbbb557fc),
	.w6(32'h3c36e916),
	.w7(32'h3b788625),
	.w8(32'hbb01faad),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf24fcd),
	.w1(32'h3c2077c5),
	.w2(32'hb90f5f16),
	.w3(32'h3b60724b),
	.w4(32'h3c660891),
	.w5(32'hbb261199),
	.w6(32'h3bbe4447),
	.w7(32'h3c75a02e),
	.w8(32'h39bd7ad1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368e8aa2),
	.w1(32'h3baabdbf),
	.w2(32'h39b5630d),
	.w3(32'hb9675918),
	.w4(32'h3b309709),
	.w5(32'hbbb853f4),
	.w6(32'h3b88e1e5),
	.w7(32'h3bc965eb),
	.w8(32'hbb547f87),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4be688),
	.w1(32'h3b153bea),
	.w2(32'h3b71be3d),
	.w3(32'h3b638002),
	.w4(32'hba1d0ad8),
	.w5(32'hba80bddf),
	.w6(32'h398e85ff),
	.w7(32'hbb03830c),
	.w8(32'hbb68b8ab),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4906bc),
	.w1(32'hbb7752eb),
	.w2(32'hbc418c1b),
	.w3(32'h3a26899b),
	.w4(32'h39a249c4),
	.w5(32'hbc096817),
	.w6(32'hbaefab25),
	.w7(32'hbab0f474),
	.w8(32'hbc298a1e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2de240),
	.w1(32'hbc55a4da),
	.w2(32'h3b4ed56f),
	.w3(32'hba845212),
	.w4(32'hbc0a984b),
	.w5(32'hbb7e3a48),
	.w6(32'hba8fdc4d),
	.w7(32'hbc4a7bb6),
	.w8(32'hbb18544d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ca053),
	.w1(32'hb92c6437),
	.w2(32'hb9e2b1cb),
	.w3(32'hbbe52590),
	.w4(32'hbb9c17c0),
	.w5(32'hbac776b8),
	.w6(32'hbbb876ab),
	.w7(32'hba9565d6),
	.w8(32'h3b8d73a5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92c9fd),
	.w1(32'h38c40140),
	.w2(32'h3b31989c),
	.w3(32'hbb9254ba),
	.w4(32'hb9c2b4b9),
	.w5(32'hba306820),
	.w6(32'hbb987594),
	.w7(32'hbad32cf9),
	.w8(32'h3b88f09b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af18b58),
	.w1(32'h3a99bf11),
	.w2(32'hbbe9bd5b),
	.w3(32'hbbdb3897),
	.w4(32'hbb92b22c),
	.w5(32'hbb861ea3),
	.w6(32'hbb18a0fe),
	.w7(32'h3b6d4ee6),
	.w8(32'hbadcf5d9),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8103b6),
	.w1(32'h3bc72f5e),
	.w2(32'hbc91ae49),
	.w3(32'h3aad6692),
	.w4(32'h3c33e47b),
	.w5(32'hbc895bd5),
	.w6(32'h3a8e5688),
	.w7(32'h3b9493ba),
	.w8(32'hbc45f88b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd93f0e),
	.w1(32'h3c0ca156),
	.w2(32'hba71ee47),
	.w3(32'h3d5a5665),
	.w4(32'h3cf1e2a5),
	.w5(32'hbb60b5fe),
	.w6(32'h3ceb0ee4),
	.w7(32'h3c855b60),
	.w8(32'hbb38f6fb),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf64881),
	.w1(32'h3a504b1e),
	.w2(32'hbd721342),
	.w3(32'h3ae8bf73),
	.w4(32'h3b39e979),
	.w5(32'hbd82a0e7),
	.w6(32'h3b4225b5),
	.w7(32'h3aacbc59),
	.w8(32'hbd3e5a24),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3e075),
	.w1(32'h3d060688),
	.w2(32'h3b28f231),
	.w3(32'h3d578457),
	.w4(32'h3dbfba58),
	.w5(32'hba9dfb40),
	.w6(32'h3d4e0fae),
	.w7(32'h3d976e4f),
	.w8(32'hb9225643),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53f9da),
	.w1(32'h3a1f8800),
	.w2(32'h3bd5f7b4),
	.w3(32'hbb5694b7),
	.w4(32'hbba1337e),
	.w5(32'hbb56f20b),
	.w6(32'hb96afae7),
	.w7(32'hbb2724c4),
	.w8(32'hbb80012d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c6dcc0),
	.w1(32'h3b5239f3),
	.w2(32'h3a9e660b),
	.w3(32'h39b780ba),
	.w4(32'h3b81c127),
	.w5(32'hbb19afac),
	.w6(32'h3b309621),
	.w7(32'h3b8265a5),
	.w8(32'hb77154a1),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b7781),
	.w1(32'h3bc215c7),
	.w2(32'h3b7be2f5),
	.w3(32'hbacd82bc),
	.w4(32'h3af20d00),
	.w5(32'hbb79ab41),
	.w6(32'hb82de57b),
	.w7(32'h3afd9385),
	.w8(32'hbb491477),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41b9b0),
	.w1(32'h3bcbada5),
	.w2(32'hba438168),
	.w3(32'h3c0d0493),
	.w4(32'h3bedc686),
	.w5(32'h3b248260),
	.w6(32'h3bb739d1),
	.w7(32'h3c13368e),
	.w8(32'h3b369ce2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a7f3b),
	.w1(32'h3ab19c3c),
	.w2(32'hbc6dc573),
	.w3(32'h3bfb4564),
	.w4(32'h3af7d129),
	.w5(32'hbc113c18),
	.w6(32'h3c227a23),
	.w7(32'h3b24f2f6),
	.w8(32'hbbf285f6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990d631),
	.w1(32'h3c137e24),
	.w2(32'h39214f71),
	.w3(32'h3c98f6e9),
	.w4(32'h3cef9235),
	.w5(32'hba53b666),
	.w6(32'h3c82cbd9),
	.w7(32'h3ca59ad3),
	.w8(32'h3a4d56c8),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8ae2b),
	.w1(32'hbbfa764c),
	.w2(32'hba1802fd),
	.w3(32'hbb0986b7),
	.w4(32'hbb30e134),
	.w5(32'hbb760395),
	.w6(32'h3b3fb35f),
	.w7(32'h3b2c631c),
	.w8(32'hba6776c8),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95063c),
	.w1(32'hbb940680),
	.w2(32'hbc1fa866),
	.w3(32'h3a99f532),
	.w4(32'h3b8ff50d),
	.w5(32'hbbe9ff02),
	.w6(32'hbbdd0ea0),
	.w7(32'hbb88253e),
	.w8(32'hbb9b5570),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19d7d3),
	.w1(32'hbb64585a),
	.w2(32'h3c7f1371),
	.w3(32'hbb9361ea),
	.w4(32'h3a938ec8),
	.w5(32'h3bd01853),
	.w6(32'hbaea7c5d),
	.w7(32'h3bcc71e5),
	.w8(32'h3bb001a2),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7dbf7),
	.w1(32'hbbe28c25),
	.w2(32'hba0bb6bf),
	.w3(32'hbbccc46c),
	.w4(32'hbc0a31a4),
	.w5(32'h3a92e3dd),
	.w6(32'hbb576c82),
	.w7(32'hbad08e67),
	.w8(32'h3b5096d9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9c989),
	.w1(32'hbb179453),
	.w2(32'hbd44ed66),
	.w3(32'h3b84f993),
	.w4(32'h3a59200a),
	.w5(32'hbd31cdac),
	.w6(32'h3b9474ad),
	.w7(32'h3a808820),
	.w8(32'hbd1572f9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe0053),
	.w1(32'h3d180b2f),
	.w2(32'h3b35133b),
	.w3(32'h3d72352a),
	.w4(32'h3dbc600f),
	.w5(32'h3afe4be4),
	.w6(32'h3d441595),
	.w7(32'h3d900592),
	.w8(32'hba96ed04),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38c355),
	.w1(32'hbb89733a),
	.w2(32'h3af39833),
	.w3(32'h3aa369c9),
	.w4(32'hbb87fe09),
	.w5(32'h3a7200d9),
	.w6(32'h3b47ffc6),
	.w7(32'h3b6fa2a4),
	.w8(32'hbab219de),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa96112),
	.w1(32'h3b9f7676),
	.w2(32'h39446197),
	.w3(32'h3b79b0f4),
	.w4(32'h399232d3),
	.w5(32'h3a3a5a1e),
	.w6(32'hbbad981c),
	.w7(32'hbbb0910c),
	.w8(32'hbb3ca5d4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91de31),
	.w1(32'h3b6e282a),
	.w2(32'hbac32192),
	.w3(32'hb9f8e26e),
	.w4(32'h3a5e8a6b),
	.w5(32'h3aac9403),
	.w6(32'hb9a1b22d),
	.w7(32'h3b5a1334),
	.w8(32'hbbb4c3af),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb300aae),
	.w1(32'h3b393627),
	.w2(32'h3b261714),
	.w3(32'hbb375461),
	.w4(32'h3b99d5cd),
	.w5(32'hbb570752),
	.w6(32'h3ada3690),
	.w7(32'hba4fb078),
	.w8(32'h3a4d1413),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af38c3c),
	.w1(32'hb9e2d414),
	.w2(32'hbba3b7bd),
	.w3(32'h3a520bfb),
	.w4(32'h3c227ca1),
	.w5(32'hbc15f1fc),
	.w6(32'hbb6292f7),
	.w7(32'h3ae02ffe),
	.w8(32'hbbe178c0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94aef7),
	.w1(32'hbbdf9856),
	.w2(32'h3ab3e155),
	.w3(32'hbade72d9),
	.w4(32'h3b8d3f37),
	.w5(32'hbb82ae85),
	.w6(32'hbb426d40),
	.w7(32'h3b8a762c),
	.w8(32'hbb48203a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06bc04),
	.w1(32'hbaa16942),
	.w2(32'h3a5228c1),
	.w3(32'hbbf14fbb),
	.w4(32'hb9ec1df2),
	.w5(32'h3b1f066e),
	.w6(32'hbb710995),
	.w7(32'hbb805db3),
	.w8(32'hbc253386),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902787a),
	.w1(32'h3b870069),
	.w2(32'h3a1f6ae8),
	.w3(32'hbb1ed6b3),
	.w4(32'hba8076f3),
	.w5(32'hbb8a21d2),
	.w6(32'hbc1048f3),
	.w7(32'hbad6d2f2),
	.w8(32'hbb46943b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c7b0c),
	.w1(32'h3a2f814c),
	.w2(32'hbb8e54f9),
	.w3(32'hbbb1e929),
	.w4(32'hbb28323e),
	.w5(32'hbad385b5),
	.w6(32'hbad8a742),
	.w7(32'hbb38af1c),
	.w8(32'hba9a2cbd),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c5311),
	.w1(32'h3aa02530),
	.w2(32'h3bf734e9),
	.w3(32'h3b639fbf),
	.w4(32'h3a9e2658),
	.w5(32'h3b4072fe),
	.w6(32'h3b973e1b),
	.w7(32'h3aac275b),
	.w8(32'h38f3322b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17884e),
	.w1(32'h3be1030f),
	.w2(32'h3b6b562e),
	.w3(32'h3c0195f9),
	.w4(32'h3bd1e5c9),
	.w5(32'hbb1557fb),
	.w6(32'h3bc210f8),
	.w7(32'h3af22aa3),
	.w8(32'h3b4100f1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7320a),
	.w1(32'h39ecdaae),
	.w2(32'h3915cb60),
	.w3(32'h3b240f26),
	.w4(32'hbad5d4b4),
	.w5(32'hb999e642),
	.w6(32'hbb1880a4),
	.w7(32'h3ae55a48),
	.w8(32'h3b235356),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4f871),
	.w1(32'h3c2ff195),
	.w2(32'hbbabb5cf),
	.w3(32'h3b9bebab),
	.w4(32'h3c2a6834),
	.w5(32'hbac4121b),
	.w6(32'h3b77de8b),
	.w7(32'h3c127e62),
	.w8(32'hbbb405bc),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4caac8),
	.w1(32'hbb775be3),
	.w2(32'h3aa9da45),
	.w3(32'hb9dd0143),
	.w4(32'h3ac39084),
	.w5(32'h3b89a773),
	.w6(32'hbb0fa561),
	.w7(32'hba2b6ca5),
	.w8(32'hbb0a218e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27ab83),
	.w1(32'h3b908d36),
	.w2(32'hbb180162),
	.w3(32'h3a147547),
	.w4(32'h3a1fe80d),
	.w5(32'hbbd8bd49),
	.w6(32'h39c23bff),
	.w7(32'h3b47164b),
	.w8(32'hbbae004e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fefbb),
	.w1(32'hba532ecd),
	.w2(32'h3aa47d82),
	.w3(32'hb8aae0ee),
	.w4(32'h3b94d8b7),
	.w5(32'hbb819ecc),
	.w6(32'hbaea72b6),
	.w7(32'h3aebbfa1),
	.w8(32'hbb7ab5ff),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d6f9e),
	.w1(32'h3b04b81f),
	.w2(32'hbb12ec4a),
	.w3(32'hbb9a17a5),
	.w4(32'hbacf09e4),
	.w5(32'h3ad309a7),
	.w6(32'hbb02b2f2),
	.w7(32'hb98021d1),
	.w8(32'hbb01d775),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91d718),
	.w1(32'h3b8bf1e0),
	.w2(32'h3a26ad30),
	.w3(32'hbaf90faa),
	.w4(32'h3bbf79bd),
	.w5(32'h39d85faa),
	.w6(32'hba7491d8),
	.w7(32'hb9aca044),
	.w8(32'hbb00f1ef),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cbabd),
	.w1(32'h3b9a6658),
	.w2(32'hbad01fe6),
	.w3(32'hbb637199),
	.w4(32'h3a2bd43f),
	.w5(32'hbb08fc6a),
	.w6(32'hbbb7d087),
	.w7(32'h3a993ab0),
	.w8(32'hbba621b3),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5a2a2),
	.w1(32'h3b29af25),
	.w2(32'hbaa36614),
	.w3(32'hb982990c),
	.w4(32'h3b921906),
	.w5(32'hbac51267),
	.w6(32'h3ac5020c),
	.w7(32'h3bbf91d1),
	.w8(32'hbb9dbcb7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ae5f2),
	.w1(32'h3bdc2bbe),
	.w2(32'h3b402a9f),
	.w3(32'h3ae8966e),
	.w4(32'h3b8bd7f9),
	.w5(32'h3a8877ab),
	.w6(32'hbb208615),
	.w7(32'h3b92760a),
	.w8(32'hbb300653),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d110e),
	.w1(32'hb964300b),
	.w2(32'h3b7e2918),
	.w3(32'hbb30e1b6),
	.w4(32'hbb31f638),
	.w5(32'h3949e17f),
	.w6(32'hb6995f6e),
	.w7(32'hbb336934),
	.w8(32'hbb955d27),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97ce14),
	.w1(32'hbb615a06),
	.w2(32'hb994b9c8),
	.w3(32'h397dc767),
	.w4(32'h3aa1655f),
	.w5(32'hbb3bd033),
	.w6(32'h3b92d3ff),
	.w7(32'h3bfca9a2),
	.w8(32'hbbb764d1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ccd43),
	.w1(32'h3af0ae62),
	.w2(32'hbad19932),
	.w3(32'h3a316ed1),
	.w4(32'h3ae030c4),
	.w5(32'hbbb312a5),
	.w6(32'hba793578),
	.w7(32'hba488585),
	.w8(32'h3a8f86c0),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1365fe),
	.w1(32'h3ab7df7f),
	.w2(32'h3a6b1449),
	.w3(32'h3b4fadc3),
	.w4(32'h3bc9ed2e),
	.w5(32'hb9a62d02),
	.w6(32'hbba1f865),
	.w7(32'hbb98a8b8),
	.w8(32'h3a35d128),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981aeba),
	.w1(32'h3b0168c5),
	.w2(32'hb9feeef9),
	.w3(32'h39374d8a),
	.w4(32'h3b6b4672),
	.w5(32'h3a80da1f),
	.w6(32'hbc163dcd),
	.w7(32'h3a8f9064),
	.w8(32'h3b89ebac),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b770ff5),
	.w1(32'hba8eacf5),
	.w2(32'h3c77883a),
	.w3(32'h3c0cf74e),
	.w4(32'h3b8d4477),
	.w5(32'h3c906f59),
	.w6(32'h3b84f1b1),
	.w7(32'h3b1abb0e),
	.w8(32'h3c8d4e03),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64ea5c),
	.w1(32'hbc19375c),
	.w2(32'h3c04ecfa),
	.w3(32'hbc3fea47),
	.w4(32'hbcd34642),
	.w5(32'h3bd4cb40),
	.w6(32'hbbe9e4ab),
	.w7(32'hbc88aebc),
	.w8(32'h3c2db863),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87d964),
	.w1(32'hbb8bc730),
	.w2(32'hbab7f5a8),
	.w3(32'hbbfc6778),
	.w4(32'hbbfc768d),
	.w5(32'hbb3e531a),
	.w6(32'hb99b12f5),
	.w7(32'hbaf595b8),
	.w8(32'h3a9e6d07),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d3a0c),
	.w1(32'hba9cd239),
	.w2(32'h3a17ce24),
	.w3(32'hbb2d6ed4),
	.w4(32'hbb27a3f7),
	.w5(32'hbab9d47e),
	.w6(32'hbb91235c),
	.w7(32'hbb750e80),
	.w8(32'hba7d8968),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45e4cf),
	.w1(32'h3bea0028),
	.w2(32'hbb876ebd),
	.w3(32'h3b7569c6),
	.w4(32'h3b12d068),
	.w5(32'hbad95ea5),
	.w6(32'h3b016ba2),
	.w7(32'h39c5853a),
	.w8(32'hbb2f6715),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08a562),
	.w1(32'h3c160881),
	.w2(32'h3a09efe4),
	.w3(32'h3b9a71a7),
	.w4(32'h3c26d059),
	.w5(32'hbabb2424),
	.w6(32'h3b857f62),
	.w7(32'h3a9a0070),
	.w8(32'hbb4d9d64),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab89771),
	.w1(32'h3b1defb5),
	.w2(32'hbad58478),
	.w3(32'hbb4c65be),
	.w4(32'h3b8b30b0),
	.w5(32'hbbaf1cc4),
	.w6(32'h3b2941dc),
	.w7(32'h3bba3d35),
	.w8(32'hbb2d1a85),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0341a0),
	.w1(32'h3bfc6e86),
	.w2(32'h3bb09637),
	.w3(32'hbb513a68),
	.w4(32'h3b793c8a),
	.w5(32'hbb491f8e),
	.w6(32'h39c788f4),
	.w7(32'h3b1cc733),
	.w8(32'hba1aea38),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule