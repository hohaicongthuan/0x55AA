module layer_10_featuremap_201(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961a487),
	.w1(32'h39c6e772),
	.w2(32'h3639847c),
	.w3(32'h39313060),
	.w4(32'h39b590e1),
	.w5(32'h39d1c70a),
	.w6(32'h398adddf),
	.w7(32'h3694213d),
	.w8(32'hb7db1538),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e0c11),
	.w1(32'hbad063fb),
	.w2(32'hb9b38a39),
	.w3(32'hbb15fc37),
	.w4(32'hbb6ea207),
	.w5(32'hbb074dd5),
	.w6(32'hbab6ca63),
	.w7(32'hbb3943e7),
	.w8(32'hbb17a7d9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381cddc3),
	.w1(32'hb952c144),
	.w2(32'hb95911f0),
	.w3(32'h381f6447),
	.w4(32'hb92853bc),
	.w5(32'hb93cdb4e),
	.w6(32'hb98340c2),
	.w7(32'hb9880a3d),
	.w8(32'hb928ea36),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e2251c),
	.w1(32'h3a87f620),
	.w2(32'h3a34bc4f),
	.w3(32'hb9db4b6e),
	.w4(32'h3a26996e),
	.w5(32'h39599284),
	.w6(32'h39e96b83),
	.w7(32'h3a1a0121),
	.w8(32'h39af55ac),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f89225),
	.w1(32'h39aca28e),
	.w2(32'h38890669),
	.w3(32'hb89ab9f1),
	.w4(32'h396b356c),
	.w5(32'h3987487d),
	.w6(32'h3963c38f),
	.w7(32'h38a3bee8),
	.w8(32'h394635c0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932a2a0),
	.w1(32'h397c4f06),
	.w2(32'h3982760a),
	.w3(32'h394acfd4),
	.w4(32'h395384b6),
	.w5(32'h398c0175),
	.w6(32'h39bf8ab2),
	.w7(32'h398bb25b),
	.w8(32'h39836a9a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43b3aa),
	.w1(32'h3b8da199),
	.w2(32'hbbdb7fdd),
	.w3(32'h3b789d2f),
	.w4(32'h3ba6bdeb),
	.w5(32'hbbd174dd),
	.w6(32'h3b13185d),
	.w7(32'h3b777db8),
	.w8(32'hbb9f709d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b140041),
	.w1(32'hbb3fc370),
	.w2(32'hbc383528),
	.w3(32'hbb953dbf),
	.w4(32'hbb8e63a0),
	.w5(32'hbb9f6ac2),
	.w6(32'hbacb019c),
	.w7(32'hbb5817c7),
	.w8(32'hbc332fca),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb830532d),
	.w1(32'h39cbdc04),
	.w2(32'h39ed698e),
	.w3(32'h390d2559),
	.w4(32'h395ead0c),
	.w5(32'h39cdb30d),
	.w6(32'h39034478),
	.w7(32'h38e05f60),
	.w8(32'h3867197a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacd6f0),
	.w1(32'h3a3f885a),
	.w2(32'hbc066f6b),
	.w3(32'hb912886b),
	.w4(32'h3aea02d7),
	.w5(32'hbbdd7d07),
	.w6(32'hb8db0cca),
	.w7(32'h3b3dbfd1),
	.w8(32'hbb8ff878),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9ee4f),
	.w1(32'hb9258565),
	.w2(32'hb8a69a3a),
	.w3(32'h387969b7),
	.w4(32'hb9650664),
	.w5(32'h3872844f),
	.w6(32'h38bc8941),
	.w7(32'hb8b0737e),
	.w8(32'h3962443a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e5bbb),
	.w1(32'h3c27877a),
	.w2(32'hbb8f49ee),
	.w3(32'h387b4d72),
	.w4(32'h3c27949e),
	.w5(32'hbb88ae06),
	.w6(32'h39b69df9),
	.w7(32'h3c080459),
	.w8(32'hbbc233b1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01a52f),
	.w1(32'h3b32c607),
	.w2(32'hbc07aabd),
	.w3(32'h3b0a96f8),
	.w4(32'h3b895981),
	.w5(32'hbbc4c814),
	.w6(32'h3aa394e7),
	.w7(32'h3b99c200),
	.w8(32'hbb9a81de),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af66b34),
	.w1(32'h3732a090),
	.w2(32'hbabfe064),
	.w3(32'h390db097),
	.w4(32'hbad6a450),
	.w5(32'hbb1afd6e),
	.w6(32'hb82f4069),
	.w7(32'hbab44b16),
	.w8(32'hbb195f7a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad63f04),
	.w1(32'hba0d6614),
	.w2(32'hba8c12e0),
	.w3(32'hbb0c6ff0),
	.w4(32'hbaebbc99),
	.w5(32'hbab4e5fd),
	.w6(32'hba8c7d9d),
	.w7(32'hba0f28cc),
	.w8(32'hba9a5be1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1035c6),
	.w1(32'hbba72f23),
	.w2(32'hbb845da3),
	.w3(32'hbaf48e85),
	.w4(32'hbbb0346b),
	.w5(32'hbbd2c91a),
	.w6(32'hbb864bfc),
	.w7(32'hbbb5c8e3),
	.w8(32'hbb83c136),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389b2727),
	.w1(32'hb95d40d0),
	.w2(32'h38eb029d),
	.w3(32'h386882b5),
	.w4(32'hb98d872c),
	.w5(32'h394f66d5),
	.w6(32'h38dca085),
	.w7(32'hb8366b67),
	.w8(32'h397033c0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b465c5f),
	.w1(32'h3a4659eb),
	.w2(32'hbc47c881),
	.w3(32'h3a995952),
	.w4(32'h3b192c79),
	.w5(32'hbc18dfaa),
	.w6(32'hbb0104ae),
	.w7(32'h3ab956b6),
	.w8(32'hbc0dc1db),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe3e12),
	.w1(32'h3ae1dfb5),
	.w2(32'hbbc2a964),
	.w3(32'h3a5a6afe),
	.w4(32'h3b1afd7e),
	.w5(32'hbb81bf20),
	.w6(32'hb9677873),
	.w7(32'h3b2133c3),
	.w8(32'hbb7419a5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb816776d),
	.w1(32'h38a660b6),
	.w2(32'hb881ed78),
	.w3(32'hb9044841),
	.w4(32'h38fa6cab),
	.w5(32'h388dbfaf),
	.w6(32'hb85418ea),
	.w7(32'hb8bacad8),
	.w8(32'hb8a35997),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb795cb82),
	.w1(32'h3a14d813),
	.w2(32'h39a475b8),
	.w3(32'h391d5f84),
	.w4(32'h396b0735),
	.w5(32'h3989318b),
	.w6(32'h39d85fe9),
	.w7(32'h3925c0a8),
	.w8(32'h37b68598),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a068055),
	.w1(32'h3a51a3f6),
	.w2(32'h391169fe),
	.w3(32'hb9afcec5),
	.w4(32'h39037dd7),
	.w5(32'hb7cca958),
	.w6(32'hb8e5e439),
	.w7(32'h39f1e876),
	.w8(32'h39441ace),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6242d),
	.w1(32'hbb00c48b),
	.w2(32'hbc2b933b),
	.w3(32'hbbdafe4b),
	.w4(32'hba8ecf53),
	.w5(32'hbc530371),
	.w6(32'hbc0940bf),
	.w7(32'h3b2258df),
	.w8(32'hbbeec18c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bbf97),
	.w1(32'h3a83354b),
	.w2(32'hbb5c2cfa),
	.w3(32'hbacdcd31),
	.w4(32'h3a8a0ecc),
	.w5(32'hbb31a01a),
	.w6(32'hbaaf10fc),
	.w7(32'h3b2164d7),
	.w8(32'hbab06222),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ce42a),
	.w1(32'h3ab6b1a8),
	.w2(32'h3b31cb38),
	.w3(32'hbbb1c027),
	.w4(32'hbb848d31),
	.w5(32'hba6ff35d),
	.w6(32'hbb2dc1af),
	.w7(32'hbb1f4c52),
	.w8(32'hbac9137c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96fac6e),
	.w1(32'hb9a511d7),
	.w2(32'hb9c037b8),
	.w3(32'h38174c5b),
	.w4(32'hb9dc2667),
	.w5(32'hba5ef8ba),
	.w6(32'hb958eb50),
	.w7(32'hb9c43546),
	.w8(32'hb9e869da),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75ec880),
	.w1(32'h38657913),
	.w2(32'h3802274a),
	.w3(32'hb5786d51),
	.w4(32'hb6be0ea5),
	.w5(32'h37fcc6fb),
	.w6(32'h391bd2f3),
	.w7(32'hb7c2b409),
	.w8(32'h36dff9e5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e9f77),
	.w1(32'h3b51e3aa),
	.w2(32'h3b707d8f),
	.w3(32'hbb2237ef),
	.w4(32'hbb237eaf),
	.w5(32'hbaf2b564),
	.w6(32'h3b29931d),
	.w7(32'h3bb4d875),
	.w8(32'h3b1a047c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c8bb0),
	.w1(32'h3932d715),
	.w2(32'h3a2ed5b8),
	.w3(32'hbb015324),
	.w4(32'hba366e1b),
	.w5(32'h376b5e71),
	.w6(32'hbad87089),
	.w7(32'hba10cfe4),
	.w8(32'hb93c730d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb078f11),
	.w1(32'h3b24afac),
	.w2(32'h3b8a011a),
	.w3(32'hbb005baf),
	.w4(32'hb9a4c56d),
	.w5(32'h399502ac),
	.w6(32'h3aaf5727),
	.w7(32'h3b168e1a),
	.w8(32'h3aab37ee),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d61b19),
	.w1(32'h390d6236),
	.w2(32'h388efe09),
	.w3(32'hb80c255b),
	.w4(32'h38dc2e0d),
	.w5(32'h38947861),
	.w6(32'h39188600),
	.w7(32'h37f69ac1),
	.w8(32'hb7b79072),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36acad1e),
	.w1(32'h388e1092),
	.w2(32'h381ec3ed),
	.w3(32'h38227564),
	.w4(32'h3841aa66),
	.w5(32'h37dfae78),
	.w6(32'h391eeb16),
	.w7(32'h38d640e2),
	.w8(32'h38ca13f2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e90189),
	.w1(32'h3a427ab4),
	.w2(32'hbb66e93e),
	.w3(32'h3915c946),
	.w4(32'h3a6e2152),
	.w5(32'hbb259396),
	.w6(32'hb992f93f),
	.w7(32'h3a830ea2),
	.w8(32'hbb1595e4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad59d99),
	.w1(32'h39a0b862),
	.w2(32'h3a565192),
	.w3(32'hbb1b1bad),
	.w4(32'hbaaad6b1),
	.w5(32'hb9e8583e),
	.w6(32'hba8076dc),
	.w7(32'hba8c4150),
	.w8(32'hba885ab6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d4e81),
	.w1(32'hb97e4aee),
	.w2(32'hba89ba28),
	.w3(32'h398640b2),
	.w4(32'h3919d4ce),
	.w5(32'hba943e14),
	.w6(32'h3a836c26),
	.w7(32'h392d1772),
	.w8(32'hba418791),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21b2ba),
	.w1(32'h3b297feb),
	.w2(32'hbb2621a8),
	.w3(32'h3ab15b42),
	.w4(32'h3ae7430d),
	.w5(32'hbb404ae5),
	.w6(32'hb97d38c3),
	.w7(32'h3ab36801),
	.w8(32'hbb3af252),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bd4e0),
	.w1(32'h3c71228b),
	.w2(32'hba36ff3b),
	.w3(32'hbc2cceb6),
	.w4(32'h3c3eeba0),
	.w5(32'hba9ef45e),
	.w6(32'hbc25ab0a),
	.w7(32'h3bd33e8c),
	.w8(32'hbb9b5913),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa6289),
	.w1(32'h3b8ad39c),
	.w2(32'h3c10ca1c),
	.w3(32'hbc066156),
	.w4(32'hbace31e9),
	.w5(32'h3bb56398),
	.w6(32'hbb0b2af8),
	.w7(32'h3b86a804),
	.w8(32'h3b61d393),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e4118),
	.w1(32'h3b88512f),
	.w2(32'h3c0b4586),
	.w3(32'hbb8f375f),
	.w4(32'hba8bea1e),
	.w5(32'h3b7c2b50),
	.w6(32'h3b56fd22),
	.w7(32'h3bd97839),
	.w8(32'h3ba5ac3f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5470c6),
	.w1(32'h3ac1cf3b),
	.w2(32'h3ab3aacb),
	.w3(32'hba92b39f),
	.w4(32'h3a1aea39),
	.w5(32'h3aad8a5a),
	.w6(32'hba47b46f),
	.w7(32'h3a8ff44d),
	.w8(32'h3a8206cc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913d8d8),
	.w1(32'hb970a58b),
	.w2(32'hb786c4a7),
	.w3(32'h38fe01ec),
	.w4(32'hb97577c2),
	.w5(32'h360718e1),
	.w6(32'hb8cf7f1a),
	.w7(32'hb824d4d4),
	.w8(32'hb82ca65e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896e14a),
	.w1(32'hb6f5f2f4),
	.w2(32'hb667bf05),
	.w3(32'hb83fc5a6),
	.w4(32'hb9824fbb),
	.w5(32'hb7d8e3e3),
	.w6(32'hb7a75908),
	.w7(32'hb93e71e6),
	.w8(32'hb9541f14),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1195bb),
	.w1(32'h3a192df4),
	.w2(32'h3b203d35),
	.w3(32'hbb05cc57),
	.w4(32'h39f0ae04),
	.w5(32'h3aa1869b),
	.w6(32'hbade3a52),
	.w7(32'hb9b7e178),
	.w8(32'h387c1a82),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1669c),
	.w1(32'hba6acc15),
	.w2(32'hbbc3f6bb),
	.w3(32'hbb727a72),
	.w4(32'hba3c209f),
	.w5(32'hbbc21ee2),
	.w6(32'hbba99923),
	.w7(32'hba334667),
	.w8(32'hbb4bd43b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70e627),
	.w1(32'h3a33f0ef),
	.w2(32'hba6f637a),
	.w3(32'hbb681600),
	.w4(32'hb9fa3a37),
	.w5(32'hba94406f),
	.w6(32'hbae5d6c6),
	.w7(32'h3ad2d968),
	.w8(32'h3931f492),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb641961),
	.w1(32'h3ae85715),
	.w2(32'hbb8509f9),
	.w3(32'hbb88f4c3),
	.w4(32'h3a17e098),
	.w5(32'hbb652e25),
	.w6(32'hbb8fd628),
	.w7(32'h3b1035cb),
	.w8(32'hbb411051),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e8a07),
	.w1(32'hba17b141),
	.w2(32'hb8dc2ff7),
	.w3(32'hbb85539b),
	.w4(32'hbaaca975),
	.w5(32'hba19401e),
	.w6(32'hba9b02d6),
	.w7(32'h39a568ac),
	.w8(32'h39f986eb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc025c),
	.w1(32'h3b8b8aff),
	.w2(32'hbc4701a4),
	.w3(32'h3b9d8933),
	.w4(32'h3b83efc1),
	.w5(32'hbc25b4ba),
	.w6(32'h3b1045f5),
	.w7(32'h3b93a8fb),
	.w8(32'hbc1ce6f3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c86d0),
	.w1(32'h38f6ad05),
	.w2(32'h382647e8),
	.w3(32'hb78e9413),
	.w4(32'h3890c624),
	.w5(32'hb84d2964),
	.w6(32'h387712b3),
	.w7(32'hb8affb63),
	.w8(32'h37c0510e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97bba13),
	.w1(32'h3962dfb9),
	.w2(32'h39aa772c),
	.w3(32'hb94bfdc7),
	.w4(32'h3819d2e3),
	.w5(32'h389eebc1),
	.w6(32'h3814513b),
	.w7(32'h38223aa2),
	.w8(32'hb77580e4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397ce0fe),
	.w1(32'hb8330d82),
	.w2(32'hb79e861a),
	.w3(32'h3907bc77),
	.w4(32'hb9356f5b),
	.w5(32'hb904da41),
	.w6(32'hb8c85865),
	.w7(32'hb94386fa),
	.w8(32'hb8afa6fc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e232f),
	.w1(32'hba848f4a),
	.w2(32'hbafee43e),
	.w3(32'hbaec4489),
	.w4(32'hb76e83ad),
	.w5(32'hbb1986db),
	.w6(32'hbb00d7fe),
	.w7(32'h3a87cfc7),
	.w8(32'hba596888),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba691231),
	.w1(32'hb89e15c4),
	.w2(32'hba384a08),
	.w3(32'hba7505f4),
	.w4(32'hba015d63),
	.w5(32'hba8a9d72),
	.w6(32'hbabd58ac),
	.w7(32'hba00d71f),
	.w8(32'hbabc81c7),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c9bc4),
	.w1(32'h3a9fc88b),
	.w2(32'hbc58c9b0),
	.w3(32'h3abfdefa),
	.w4(32'h3b50e6cf),
	.w5(32'hbc1c7964),
	.w6(32'h3b263547),
	.w7(32'h3b93c439),
	.w8(32'hbc050b15),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92be936),
	.w1(32'h39dc6bc6),
	.w2(32'hba102e48),
	.w3(32'hbad78cf4),
	.w4(32'hb9e19177),
	.w5(32'hb9843e58),
	.w6(32'hba47ad16),
	.w7(32'hba185404),
	.w8(32'hba9c6e49),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ebb50),
	.w1(32'hb76f1e13),
	.w2(32'h36a7f698),
	.w3(32'hb918582d),
	.w4(32'hb986ebb8),
	.w5(32'hb96e5108),
	.w6(32'h36c4f616),
	.w7(32'hb918e149),
	.w8(32'hb9d47f3f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8badfb6),
	.w1(32'hb8d30f12),
	.w2(32'h37d5c306),
	.w3(32'hb8dd32fc),
	.w4(32'hb968669b),
	.w5(32'hb91c76a4),
	.w6(32'hb8115418),
	.w7(32'hb725190e),
	.w8(32'hb80b4921),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d7e97),
	.w1(32'h394dfe09),
	.w2(32'h39b01f51),
	.w3(32'h395e6af5),
	.w4(32'h376182c1),
	.w5(32'h393de7d8),
	.w6(32'h3a1ae5fb),
	.w7(32'h398ee1bb),
	.w8(32'h399adef3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987bfb9),
	.w1(32'h39a4b5d0),
	.w2(32'h39ae5b1c),
	.w3(32'hba577a07),
	.w4(32'hb91d4a79),
	.w5(32'hb9248f17),
	.w6(32'hba29fb43),
	.w7(32'hb8925583),
	.w8(32'hb9325a3d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a51e2),
	.w1(32'h3996764d),
	.w2(32'h398ef36f),
	.w3(32'hb8d9201d),
	.w4(32'h3a23832b),
	.w5(32'hb8e273cb),
	.w6(32'h3a444fbe),
	.w7(32'h39e25c49),
	.w8(32'h391216a7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a852337),
	.w1(32'h39b7f55f),
	.w2(32'hbb8bdb2a),
	.w3(32'h39fcd104),
	.w4(32'h3a37c06a),
	.w5(32'hbb6e0bda),
	.w6(32'hba02c3d1),
	.w7(32'h3a86059f),
	.w8(32'hbb19f947),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48c269),
	.w1(32'hbba653e2),
	.w2(32'hbae18544),
	.w3(32'hbba1dc7a),
	.w4(32'hbb48db59),
	.w5(32'hbb0a9905),
	.w6(32'hbb684e4b),
	.w7(32'hbb463238),
	.w8(32'hbb10be49),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3828c5a9),
	.w1(32'hb804bd86),
	.w2(32'hba08e773),
	.w3(32'h3899e412),
	.w4(32'h382b9d8e),
	.w5(32'h38813f0c),
	.w6(32'hb94972e7),
	.w7(32'hb9e3ffc0),
	.w8(32'hb990669f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dd9fe),
	.w1(32'hb93729e2),
	.w2(32'hb968019a),
	.w3(32'hb98a3153),
	.w4(32'hb70f4a32),
	.w5(32'hb89e17a6),
	.w6(32'hb8f184e6),
	.w7(32'hb941d9fa),
	.w8(32'h38090abc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38440c26),
	.w1(32'hb92324de),
	.w2(32'hb984f644),
	.w3(32'h391a59d6),
	.w4(32'hb8d042db),
	.w5(32'hb9392b6c),
	.w6(32'hb91a9f61),
	.w7(32'hb923bef6),
	.w8(32'hb8823a37),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a38269),
	.w1(32'hb956f9a3),
	.w2(32'h38308e41),
	.w3(32'hb80cd1bd),
	.w4(32'hb98435d5),
	.w5(32'hb90e23f4),
	.w6(32'hb933155f),
	.w7(32'hb89c14e0),
	.w8(32'hb89d0bdc),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4df7e2),
	.w1(32'hbb6b15c1),
	.w2(32'hbc5cdb4c),
	.w3(32'h398490a9),
	.w4(32'hbb2cc64f),
	.w5(32'hbc45084e),
	.w6(32'h3bdb5716),
	.w7(32'h3af0e259),
	.w8(32'hbbc7f1e7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa72c3),
	.w1(32'h3b0a2065),
	.w2(32'hbbbfafed),
	.w3(32'hbb38be8d),
	.w4(32'hba27d8a2),
	.w5(32'hbbe7dcd5),
	.w6(32'hbc07ea6e),
	.w7(32'hbb3ae6df),
	.w8(32'hbc345daf),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb210b33),
	.w1(32'hbab114c1),
	.w2(32'hbb40cc04),
	.w3(32'hbb84c6b0),
	.w4(32'hbaabbe88),
	.w5(32'hbb824429),
	.w6(32'hbb8451cb),
	.w7(32'hba6c3559),
	.w8(32'hbb8e83f9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65be48),
	.w1(32'h3bd64480),
	.w2(32'h3b9c6bef),
	.w3(32'hbbac88d5),
	.w4(32'h39768bf1),
	.w5(32'h3b1c9b34),
	.w6(32'hba77e435),
	.w7(32'h3b505acf),
	.w8(32'h3adb0b7c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c42ca),
	.w1(32'hb931c69b),
	.w2(32'hb920a234),
	.w3(32'hb8b87776),
	.w4(32'hb8843727),
	.w5(32'hb88824a7),
	.w6(32'hb8cf5e69),
	.w7(32'hb91f064e),
	.w8(32'hb892ded6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382765c5),
	.w1(32'h38b5e7c8),
	.w2(32'h3921157e),
	.w3(32'h38a9c0d9),
	.w4(32'h38e35bdd),
	.w5(32'h39176a32),
	.w6(32'h3950e3e3),
	.w7(32'h381e1cf7),
	.w8(32'h38d52b37),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39432f80),
	.w1(32'h39273027),
	.w2(32'h39523209),
	.w3(32'h392b5b8a),
	.w4(32'h393b79b5),
	.w5(32'h3949fc3a),
	.w6(32'h397bc051),
	.w7(32'h3888dea8),
	.w8(32'h38dbe2a6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70b731),
	.w1(32'h39a8c189),
	.w2(32'hbb00941a),
	.w3(32'h39998f29),
	.w4(32'h3a3cc703),
	.w5(32'hbab4c487),
	.w6(32'h3a07eb32),
	.w7(32'h3a1b3d51),
	.w8(32'hbaf9bcb9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395931c4),
	.w1(32'hb835a178),
	.w2(32'hb8b917dc),
	.w3(32'h39057957),
	.w4(32'hb8d1c8dd),
	.w5(32'hb90cafdd),
	.w6(32'h34f6422d),
	.w7(32'hb905a88c),
	.w8(32'hb8c81cfa),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a5c4c),
	.w1(32'h3b33dc76),
	.w2(32'hbb9aa3f4),
	.w3(32'h3a717e60),
	.w4(32'h3aad4304),
	.w5(32'hbb36038c),
	.w6(32'h3b447408),
	.w7(32'h3b4bed85),
	.w8(32'hbb22c7ea),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa612d8),
	.w1(32'h3b7dc5bb),
	.w2(32'hbb802dc9),
	.w3(32'hb984f395),
	.w4(32'h3af1863d),
	.w5(32'hbb14a32f),
	.w6(32'hbb10f05b),
	.w7(32'h3b1c1ae4),
	.w8(32'hbb89b146),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb244d73),
	.w1(32'h39d4afa2),
	.w2(32'hbac9f8c1),
	.w3(32'hbacf2e8f),
	.w4(32'hba0b8dde),
	.w5(32'hbaaced47),
	.w6(32'h37cdbd9a),
	.w7(32'h3a9ccb80),
	.w8(32'hb9b70d79),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a03e6a),
	.w1(32'hba5a2afc),
	.w2(32'hbb8dbdab),
	.w3(32'hba8a5157),
	.w4(32'hba92aed6),
	.w5(32'hbb816e5b),
	.w6(32'hba6213ca),
	.w7(32'hba4ea7c7),
	.w8(32'hbb4d1eea),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e34d1),
	.w1(32'h3aa1cb1b),
	.w2(32'hbbcad0f1),
	.w3(32'h381b19c0),
	.w4(32'h3b07e5f3),
	.w5(32'hbb95456e),
	.w6(32'h3b8a27ff),
	.w7(32'h3b8c762d),
	.w8(32'hbadb3557),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab32ca1),
	.w1(32'hba6ea4bd),
	.w2(32'hb969e384),
	.w3(32'hbaab4436),
	.w4(32'hbaed40f1),
	.w5(32'hba99b056),
	.w6(32'h39e7f029),
	.w7(32'hb9e4d527),
	.w8(32'hba2a9522),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd8c67),
	.w1(32'h3b12451b),
	.w2(32'hbb8e35e5),
	.w3(32'h3ae035c8),
	.w4(32'h3b0e034a),
	.w5(32'hbb6d4bf5),
	.w6(32'h3aa7aa73),
	.w7(32'h3b287994),
	.w8(32'hbb35f69e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dc74c1),
	.w1(32'hb7f90d6d),
	.w2(32'hb830a6f2),
	.w3(32'h3847f82b),
	.w4(32'hb88e0260),
	.w5(32'hb8bf7104),
	.w6(32'h36eba818),
	.w7(32'hb8447eaf),
	.w8(32'hb803fee0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fd241c),
	.w1(32'h38511d09),
	.w2(32'h38758a3d),
	.w3(32'h371ea1bb),
	.w4(32'h3836aedf),
	.w5(32'h37cc8485),
	.w6(32'h385e0fe4),
	.w7(32'h37415a79),
	.w8(32'hb60daa23),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3875c7e0),
	.w1(32'hb90f530e),
	.w2(32'hb9500103),
	.w3(32'h3821e9aa),
	.w4(32'hb96260e1),
	.w5(32'hb7d048bd),
	.w6(32'hb7de5813),
	.w7(32'hb77423e6),
	.w8(32'hb906e073),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c3286),
	.w1(32'h3a3c7460),
	.w2(32'h3995e4b6),
	.w3(32'h3a1a2d03),
	.w4(32'h3a41e2be),
	.w5(32'h39f41219),
	.w6(32'h3a571aff),
	.w7(32'h3a6c7cd5),
	.w8(32'h39c30de5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac64c7),
	.w1(32'h391344f4),
	.w2(32'h3b428214),
	.w3(32'hbbae71ef),
	.w4(32'hbb0127a2),
	.w5(32'h3aa3e05c),
	.w6(32'hbb3f1b14),
	.w7(32'hb998118a),
	.w8(32'h3a838de7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74dd839),
	.w1(32'h3a109bf3),
	.w2(32'h3a018429),
	.w3(32'hb9a24ad2),
	.w4(32'h39b8ff33),
	.w5(32'h38d8b4d8),
	.w6(32'hb830f3ad),
	.w7(32'h39a0aa86),
	.w8(32'h387010c0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30c49a),
	.w1(32'hbaedec2c),
	.w2(32'hbb5fc999),
	.w3(32'hbb770387),
	.w4(32'hbb7da5bb),
	.w5(32'hbb51cd8b),
	.w6(32'hbb5c00a2),
	.w7(32'hbb0c3c41),
	.w8(32'hbb548c60),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e2bdb),
	.w1(32'h3a066289),
	.w2(32'hbbe388fe),
	.w3(32'hbadb77d0),
	.w4(32'hba8b1ec5),
	.w5(32'hbbe202b2),
	.w6(32'hbb1f248f),
	.w7(32'hba486d24),
	.w8(32'hbbf0b573),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5c110),
	.w1(32'h3b42f954),
	.w2(32'h3ba06524),
	.w3(32'hba89043e),
	.w4(32'h3aa9c158),
	.w5(32'h3b865cc7),
	.w6(32'h3b56204e),
	.w7(32'h3ba198be),
	.w8(32'h3baeeba7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb7994),
	.w1(32'h3b38fb64),
	.w2(32'hbbaba31a),
	.w3(32'h3afae57d),
	.w4(32'h3b95a690),
	.w5(32'hbbc18c11),
	.w6(32'h3a41b5d1),
	.w7(32'h3be76263),
	.w8(32'hbb32279b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52666d),
	.w1(32'h3b893a67),
	.w2(32'h3b2aea30),
	.w3(32'hb9cf2668),
	.w4(32'h3b7a63fa),
	.w5(32'h3b6ee5f4),
	.w6(32'h3b15e6b7),
	.w7(32'h3ba92a22),
	.w8(32'h3b9ebd89),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81430b),
	.w1(32'hbb305315),
	.w2(32'hbbdddaaf),
	.w3(32'hbb58cff2),
	.w4(32'hbb8da8e5),
	.w5(32'hbc1013b1),
	.w6(32'hbbad3a6f),
	.w7(32'hbb8abe41),
	.w8(32'hbc1656a6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb641717),
	.w1(32'hbb8a8482),
	.w2(32'hbb938251),
	.w3(32'hbb29eece),
	.w4(32'hbb6b368a),
	.w5(32'hbbbc8d14),
	.w6(32'hb989c654),
	.w7(32'hbaaba232),
	.w8(32'hbb2b9a09),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b75ce),
	.w1(32'h3a4e4af4),
	.w2(32'h3b3937d6),
	.w3(32'hba8ea3f5),
	.w4(32'hb96e4261),
	.w5(32'h3a908b1c),
	.w6(32'h3aa17ca4),
	.w7(32'h3b2a0dd7),
	.w8(32'h3b17e0f0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3f70f),
	.w1(32'h3985085a),
	.w2(32'h363d1f11),
	.w3(32'h397e2719),
	.w4(32'hb8bd1d66),
	.w5(32'hb9b19b2b),
	.w6(32'hb93629f5),
	.w7(32'hb93ecd76),
	.w8(32'hb936a1ec),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3836d669),
	.w1(32'h3afd8586),
	.w2(32'hbbec9fac),
	.w3(32'hba688217),
	.w4(32'h3aec1ffa),
	.w5(32'hbbc17851),
	.w6(32'hbb139755),
	.w7(32'h3ae259bb),
	.w8(32'hbbb5e1b8),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d9b32),
	.w1(32'h3a6fcf64),
	.w2(32'hbbcb02c8),
	.w3(32'h379959c4),
	.w4(32'h3b366bd5),
	.w5(32'hbb6cd7b3),
	.w6(32'h3bbfe2c5),
	.w7(32'h3bc8e54e),
	.w8(32'hba7f2d12),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32f135),
	.w1(32'h3c30e941),
	.w2(32'hbb3c6b7b),
	.w3(32'hbc0d1754),
	.w4(32'h3b99fc46),
	.w5(32'hbb9ed280),
	.w6(32'hbc3be226),
	.w7(32'h3b578b82),
	.w8(32'hbb6bdd50),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a4596),
	.w1(32'h3b8b90d8),
	.w2(32'h3c09e841),
	.w3(32'hbc3db471),
	.w4(32'hba4c2ddc),
	.w5(32'h3b40ade4),
	.w6(32'hbc058fbe),
	.w7(32'hb99c39a1),
	.w8(32'h3a837a0f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c48b1),
	.w1(32'h3b28d17b),
	.w2(32'hba8a9cf4),
	.w3(32'hbb2d1602),
	.w4(32'hba64f1ae),
	.w5(32'hbb0b0e89),
	.w6(32'hbb163551),
	.w7(32'h3a06b0e3),
	.w8(32'hbaf52df9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ff3701),
	.w1(32'h3bee23a5),
	.w2(32'hbb95dea6),
	.w3(32'hbb43a656),
	.w4(32'h3bea8f62),
	.w5(32'hbb7df891),
	.w6(32'hbac1faaf),
	.w7(32'h3bbaa683),
	.w8(32'hbb46f83f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7470f4d),
	.w1(32'h3936c03b),
	.w2(32'h39f2d4a2),
	.w3(32'h39ab4a21),
	.w4(32'hb8fe0fd7),
	.w5(32'hb8a2aff8),
	.w6(32'h388c1b18),
	.w7(32'hb92458a3),
	.w8(32'hb7b021f6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67a269),
	.w1(32'h3bb0ea42),
	.w2(32'hbbcf8da8),
	.w3(32'hbb704575),
	.w4(32'hba6c2208),
	.w5(32'hbb6b4e7e),
	.w6(32'hbb09eebe),
	.w7(32'h3b2e3c6f),
	.w8(32'hbb7cdd07),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db0272),
	.w1(32'h3ba20ff4),
	.w2(32'h3b641651),
	.w3(32'h3b59b443),
	.w4(32'h3bc07964),
	.w5(32'h3baa93f2),
	.w6(32'h3b22c1e9),
	.w7(32'h3baf2251),
	.w8(32'h3b83223f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb588540e),
	.w1(32'hb8855e05),
	.w2(32'hb979ae67),
	.w3(32'hb7d6817d),
	.w4(32'hb8949e3f),
	.w5(32'hb90fa5c9),
	.w6(32'hb9290ed0),
	.w7(32'hb79d0ec2),
	.w8(32'hb9050259),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba391603),
	.w1(32'hba0dcdd6),
	.w2(32'h38aa07f4),
	.w3(32'hba52fa2d),
	.w4(32'hb95db33a),
	.w5(32'hbad5883f),
	.w6(32'hba0c9591),
	.w7(32'hba41fb84),
	.w8(32'hbad88ef8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba009d88),
	.w1(32'h3aff4122),
	.w2(32'hbb4f10d0),
	.w3(32'hb917471f),
	.w4(32'h3b0d8384),
	.w5(32'hbb40428a),
	.w6(32'hbaad3ed8),
	.w7(32'h3ae0454c),
	.w8(32'hbb25a2a1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d50da4),
	.w1(32'h3b1b7d57),
	.w2(32'h3a638d26),
	.w3(32'hb996cefb),
	.w4(32'h3893fe10),
	.w5(32'hb94616d8),
	.w6(32'h39f70a8f),
	.w7(32'h3b0386c8),
	.w8(32'h3a7461d5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03e436),
	.w1(32'h38a040da),
	.w2(32'h3b4cb197),
	.w3(32'hb831f83b),
	.w4(32'hba142e08),
	.w5(32'h3ace9daf),
	.w6(32'h3b462ec6),
	.w7(32'h3b22acdb),
	.w8(32'h3b30d0e7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eb03d),
	.w1(32'hbac8cc94),
	.w2(32'hba9520fa),
	.w3(32'hbb1cb68f),
	.w4(32'hbae46590),
	.w5(32'hba96296c),
	.w6(32'hbad18a26),
	.w7(32'hbae91ad4),
	.w8(32'hbad8f3c9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26b004),
	.w1(32'h3b635239),
	.w2(32'h39f161d0),
	.w3(32'hbb3539f8),
	.w4(32'hba45ddab),
	.w5(32'hbb27bf56),
	.w6(32'hbba9e500),
	.w7(32'hbb37ec70),
	.w8(32'hbbbb5d02),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96eda0c),
	.w1(32'hbb381c37),
	.w2(32'hbbc7c487),
	.w3(32'hba34d75b),
	.w4(32'hbb28fa19),
	.w5(32'hbbe243fb),
	.w6(32'hbb1c3e59),
	.w7(32'hbb403c21),
	.w8(32'hbb89d459),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0d48b),
	.w1(32'h3a086811),
	.w2(32'hb9e6e60f),
	.w3(32'hbab99861),
	.w4(32'hb8a78947),
	.w5(32'hba294773),
	.w6(32'hba91e3af),
	.w7(32'h3a052947),
	.w8(32'hb9a7b945),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d4571),
	.w1(32'h396c6b7c),
	.w2(32'h39653a00),
	.w3(32'hb9a8962d),
	.w4(32'h393c98b5),
	.w5(32'h391b5923),
	.w6(32'h399b82ec),
	.w7(32'h3920ef09),
	.w8(32'h394c6f12),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b1010),
	.w1(32'hb9cb5f14),
	.w2(32'hb922f586),
	.w3(32'hb98fc934),
	.w4(32'hb6f8f848),
	.w5(32'hb9cb4190),
	.w6(32'h372faaa1),
	.w7(32'hb96e2229),
	.w8(32'hba484cbb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e7921e),
	.w1(32'h39432dd4),
	.w2(32'h392fc5f4),
	.w3(32'h3886e351),
	.w4(32'h392c98f0),
	.w5(32'h39206b5b),
	.w6(32'h398c5da4),
	.w7(32'h393a6549),
	.w8(32'h3920aa8d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f4b7c),
	.w1(32'hb70caf9b),
	.w2(32'h38cd8192),
	.w3(32'h39043a27),
	.w4(32'hb82e783a),
	.w5(32'hb8f25171),
	.w6(32'h37268807),
	.w7(32'hb8f115eb),
	.w8(32'h3892128d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26181b),
	.w1(32'h39e307be),
	.w2(32'hbab26626),
	.w3(32'hbb02f9b0),
	.w4(32'hb90c19d0),
	.w5(32'hbaa2ac32),
	.w6(32'hba95f170),
	.w7(32'h3a264c26),
	.w8(32'hba64183c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cfbf22),
	.w1(32'h38e2d230),
	.w2(32'hb4d5c51f),
	.w3(32'h381cf096),
	.w4(32'h392816ca),
	.w5(32'hb894b7b7),
	.w6(32'h37e2b107),
	.w7(32'h38cc4422),
	.w8(32'h38c1aadb),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d9b17),
	.w1(32'h3b13abd3),
	.w2(32'hbb51924e),
	.w3(32'h3ad20d9a),
	.w4(32'h3b0efcfd),
	.w5(32'hbb2e4508),
	.w6(32'h3b02e9a5),
	.w7(32'h3b125ce4),
	.w8(32'hbb141fb6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba58dc9),
	.w1(32'hbb380280),
	.w2(32'h3b03727c),
	.w3(32'hbb937781),
	.w4(32'hbbbebf14),
	.w5(32'hbaaf9408),
	.w6(32'hbb005718),
	.w7(32'hbb86dede),
	.w8(32'hbb56c2b5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3953132d),
	.w1(32'hb9825da9),
	.w2(32'h378ddac2),
	.w3(32'h392c4c8a),
	.w4(32'h376c787e),
	.w5(32'h3751dcf3),
	.w6(32'hb960e82e),
	.w7(32'hb8d500ce),
	.w8(32'hb97aad2e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fed036),
	.w1(32'h39a2c9d3),
	.w2(32'h3986a9a7),
	.w3(32'hb883a12d),
	.w4(32'h391cea1e),
	.w5(32'h395d5b28),
	.w6(32'h39a2619d),
	.w7(32'h38be97e1),
	.w8(32'hb6498436),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b5908),
	.w1(32'h394eace8),
	.w2(32'h3919310f),
	.w3(32'h3993ae58),
	.w4(32'h3934dfeb),
	.w5(32'h3916e948),
	.w6(32'h3944ec98),
	.w7(32'h37a745ee),
	.w8(32'hb7ba6336),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69064d),
	.w1(32'hb9dbc61f),
	.w2(32'hb8be80a4),
	.w3(32'hba510344),
	.w4(32'hb9eb04b5),
	.w5(32'h38a6718e),
	.w6(32'hba6f31f7),
	.w7(32'hb9cb266c),
	.w8(32'hb8d1c61f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbaa57d),
	.w1(32'h3bb5da0b),
	.w2(32'hbb9cef8d),
	.w3(32'h3a85825d),
	.w4(32'h3ad704cb),
	.w5(32'hbbf804e2),
	.w6(32'hbc1abe2f),
	.w7(32'h3857eb7c),
	.w8(32'hbbfc5d4a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56423c),
	.w1(32'hb99118e6),
	.w2(32'hbc07bed9),
	.w3(32'h3a1126bd),
	.w4(32'h3a878f15),
	.w5(32'hbbc52e2c),
	.w6(32'hb9a175d7),
	.w7(32'h3acd6acd),
	.w8(32'hbbaece34),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f088c0),
	.w1(32'h39791563),
	.w2(32'hba1b9100),
	.w3(32'h39900d40),
	.w4(32'h3962ae9d),
	.w5(32'hba022a9b),
	.w6(32'h3a4e3195),
	.w7(32'h3a3c5931),
	.w8(32'hb9c3d54c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba198b0f),
	.w1(32'hb9325159),
	.w2(32'hbafd7e8c),
	.w3(32'hbab0c0b2),
	.w4(32'hba29f6c9),
	.w5(32'hbacade67),
	.w6(32'hba8a3380),
	.w7(32'hbab03380),
	.w8(32'hbb3affcb),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfc595),
	.w1(32'hb964b7f1),
	.w2(32'hb8f29c19),
	.w3(32'hbacf9910),
	.w4(32'hb9a0b7a3),
	.w5(32'hba4b5e78),
	.w6(32'hba3b8197),
	.w7(32'h3982a088),
	.w8(32'hb909c769),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f0944),
	.w1(32'hba258a66),
	.w2(32'hbb15e6b9),
	.w3(32'hbaba5b0e),
	.w4(32'hba844280),
	.w5(32'hbb108560),
	.w6(32'hbaba5f37),
	.w7(32'hbaa9aaf3),
	.w8(32'hbb300228),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab42edd),
	.w1(32'hbb592aaf),
	.w2(32'hbab64f5f),
	.w3(32'hbae51b9f),
	.w4(32'hbb6bd97f),
	.w5(32'hbb6f138f),
	.w6(32'h397fb788),
	.w7(32'hbad36be5),
	.w8(32'hbae840a7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47c541),
	.w1(32'h3a9c759a),
	.w2(32'hbc35be59),
	.w3(32'h3b2675f7),
	.w4(32'h3b4ac835),
	.w5(32'hbc12a43e),
	.w6(32'h3ae23e29),
	.w7(32'h3b7dcff2),
	.w8(32'hbbbe4c44),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2be6b6),
	.w1(32'h39ab0912),
	.w2(32'h3aaddd62),
	.w3(32'hbb3f10f3),
	.w4(32'hbaee5248),
	.w5(32'hb92b4398),
	.w6(32'hbb0fcb7b),
	.w7(32'hba5fa158),
	.w8(32'hb9d84975),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb195d08),
	.w1(32'hbb06938b),
	.w2(32'hbba14271),
	.w3(32'hba220494),
	.w4(32'h391d1785),
	.w5(32'hbb41a8ac),
	.w6(32'hbac7b13b),
	.w7(32'hb99f8dce),
	.w8(32'hbb72e209),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68a91a),
	.w1(32'h3986899d),
	.w2(32'hbc16c5a4),
	.w3(32'h38b75322),
	.w4(32'h39a2d44a),
	.w5(32'hbc0a35a3),
	.w6(32'h39ebcc1d),
	.w7(32'h3b040697),
	.w8(32'hbbe82961),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb417517),
	.w1(32'h3ac448a4),
	.w2(32'h3b1211e8),
	.w3(32'hbb7155c3),
	.w4(32'hba53c6f5),
	.w5(32'h3a1f40b8),
	.w6(32'hbb92eb84),
	.w7(32'hba683be6),
	.w8(32'hb8d6361a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0b0f6),
	.w1(32'h3841c0e0),
	.w2(32'hbb854975),
	.w3(32'hbaaf82cb),
	.w4(32'h39293ba3),
	.w5(32'hbb67eb0f),
	.w6(32'hba85b1bb),
	.w7(32'h39a34270),
	.w8(32'hbb333e1e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993a636),
	.w1(32'h399b798d),
	.w2(32'hba3d6838),
	.w3(32'hb81d4f35),
	.w4(32'h39d57898),
	.w5(32'hb9d4373e),
	.w6(32'h38617864),
	.w7(32'h3a2f2b23),
	.w8(32'hb90370b8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba607189),
	.w1(32'h3b74f5de),
	.w2(32'h3b15b05a),
	.w3(32'hbb105933),
	.w4(32'hb9b3c940),
	.w5(32'hba8e6cab),
	.w6(32'h39f1a29d),
	.w7(32'h3b3ef2c8),
	.w8(32'h3a59b452),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac15272),
	.w1(32'hba913db8),
	.w2(32'h3970c979),
	.w3(32'hbaf1b616),
	.w4(32'hba7d01c2),
	.w5(32'hb8900470),
	.w6(32'hbaf078de),
	.w7(32'hb9dcaa67),
	.w8(32'hb9f20d51),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f59a54),
	.w1(32'h35f1c691),
	.w2(32'hb8df8d9b),
	.w3(32'h38e6ec19),
	.w4(32'h387ebdb6),
	.w5(32'hb88f06f2),
	.w6(32'h38e454ee),
	.w7(32'h3810a6ca),
	.w8(32'hb906d4fd),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c7b574),
	.w1(32'hb7da95fd),
	.w2(32'hb786f0b8),
	.w3(32'h37b42e12),
	.w4(32'hb842154d),
	.w5(32'hb851b305),
	.w6(32'h38cbdbd0),
	.w7(32'h38773c0a),
	.w8(32'h3613ee21),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17f381),
	.w1(32'h3a5c1b9d),
	.w2(32'h3a3708ce),
	.w3(32'h3a1c56f9),
	.w4(32'h3a09e49c),
	.w5(32'h3ac1004a),
	.w6(32'h3a9a1747),
	.w7(32'h39d510e2),
	.w8(32'h3ac5c117),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c559b),
	.w1(32'h3ad6f581),
	.w2(32'hb9cfb08e),
	.w3(32'hbb4cd324),
	.w4(32'hba5bc919),
	.w5(32'hba1c0f79),
	.w6(32'hbabec04d),
	.w7(32'h39f6f66a),
	.w8(32'hb9b164f5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b588a),
	.w1(32'h3b059639),
	.w2(32'hbba1ed71),
	.w3(32'h3a88d8c7),
	.w4(32'h3b33ec60),
	.w5(32'hbb5e9ef6),
	.w6(32'h3a9c2b89),
	.w7(32'h3b70486c),
	.w8(32'hbaff1842),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fe3400),
	.w1(32'hb7f428e4),
	.w2(32'hb6a9c667),
	.w3(32'h37d249a1),
	.w4(32'hb8056ad6),
	.w5(32'hb6dedb18),
	.w6(32'h36fea1f9),
	.w7(32'hb7ea47a7),
	.w8(32'hb792e229),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f1e5c),
	.w1(32'h3a09a5b9),
	.w2(32'hbbc55868),
	.w3(32'hba06a45d),
	.w4(32'h3a367c4a),
	.w5(32'hbba2a592),
	.w6(32'hb8f2b3b8),
	.w7(32'h3b165b28),
	.w8(32'hbb685ea5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffa9f9),
	.w1(32'h3910cbc8),
	.w2(32'hbad20a8f),
	.w3(32'hbaa05ee7),
	.w4(32'h3966d7ec),
	.w5(32'hbaaf3114),
	.w6(32'hbae2aca6),
	.w7(32'h391aaaf2),
	.w8(32'hba8b731f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3db6af),
	.w1(32'h3b38bcaa),
	.w2(32'hbbe7dcdc),
	.w3(32'h3b0b2bae),
	.w4(32'h3b8d0372),
	.w5(32'hbba94cd7),
	.w6(32'h3ab019b8),
	.w7(32'h3b969bac),
	.w8(32'hbb7005df),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd8b90),
	.w1(32'h3b12e3d5),
	.w2(32'h3af842bf),
	.w3(32'hbaa06fae),
	.w4(32'h3a2a661d),
	.w5(32'hba6ff651),
	.w6(32'h3bc353ca),
	.w7(32'h3bd8e574),
	.w8(32'h39583f83),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a155d),
	.w1(32'hbaa5597a),
	.w2(32'hb96fe036),
	.w3(32'hbb1b867a),
	.w4(32'hbb1e7fd6),
	.w5(32'hbadf2de9),
	.w6(32'hbb07355e),
	.w7(32'hbb1610fe),
	.w8(32'hbb0cddaa),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c35ead),
	.w1(32'h3898c4fc),
	.w2(32'h39902400),
	.w3(32'hb83fb9cf),
	.w4(32'hb7e63150),
	.w5(32'hb98e4159),
	.w6(32'hb98f26d5),
	.w7(32'hb97ad380),
	.w8(32'hb9836eae),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b1580),
	.w1(32'h3a7f4755),
	.w2(32'h3b143198),
	.w3(32'hbb36f908),
	.w4(32'hb9e74ee0),
	.w5(32'h3ab57af7),
	.w6(32'hbaff5dec),
	.w7(32'h3959756d),
	.w8(32'h3a1c6616),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc830),
	.w1(32'hbb0eece0),
	.w2(32'h3abc9e2a),
	.w3(32'hbbaa702f),
	.w4(32'hbb5ba8c2),
	.w5(32'h39a196f1),
	.w6(32'hbb149438),
	.w7(32'hbabbf2cc),
	.w8(32'hb9a1ed9a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba011e9b),
	.w1(32'h3aab7ac5),
	.w2(32'h3abf819f),
	.w3(32'hbab28d67),
	.w4(32'hb9eab3c0),
	.w5(32'h3a4fd4e8),
	.w6(32'hb9638f2f),
	.w7(32'h3a307ea9),
	.w8(32'h39dd137c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e55e8),
	.w1(32'h3a12ebc4),
	.w2(32'hbad7299f),
	.w3(32'h3a0ab0ef),
	.w4(32'h3a01edad),
	.w5(32'hbaa2500b),
	.w6(32'h3a6f25ed),
	.w7(32'h3a8bec19),
	.w8(32'hba59d8be),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97da519),
	.w1(32'hb98adbfd),
	.w2(32'hb92f7e25),
	.w3(32'hb9bf1c76),
	.w4(32'hb9aa2564),
	.w5(32'hb9d3b3b9),
	.w6(32'hb9d89714),
	.w7(32'hb9ca7dd3),
	.w8(32'hb9db0159),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ae096),
	.w1(32'h3a5df929),
	.w2(32'hbbb5ba50),
	.w3(32'hba1b6e5c),
	.w4(32'h3a6f131a),
	.w5(32'hbb8e1285),
	.w6(32'hbaa4438f),
	.w7(32'h3a436f75),
	.w8(32'hbb87e641),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa345c8),
	.w1(32'h3aed5c03),
	.w2(32'hba0e6493),
	.w3(32'h3ab594bd),
	.w4(32'h3b03ea87),
	.w5(32'hb9a5043f),
	.w6(32'h3af36a3f),
	.w7(32'h3af50b05),
	.w8(32'h3a0e96a4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb7b96),
	.w1(32'hb972fd0a),
	.w2(32'h395ecca1),
	.w3(32'hbb055d11),
	.w4(32'hbaa4fdff),
	.w5(32'hbaa0b1e7),
	.w6(32'hbaa05fb9),
	.w7(32'hba595fa8),
	.w8(32'hbad439fb),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3825ed73),
	.w1(32'h3947cf62),
	.w2(32'h3949b476),
	.w3(32'h379a24a3),
	.w4(32'h38d7f711),
	.w5(32'h39779838),
	.w6(32'h38ef37af),
	.w7(32'h38d8f848),
	.w8(32'h39323dc4),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77c0e3),
	.w1(32'h3b449481),
	.w2(32'hbaf74868),
	.w3(32'h3ae9f632),
	.w4(32'h3a94dff6),
	.w5(32'hbb562c8f),
	.w6(32'h393d681b),
	.w7(32'h39a7e400),
	.w8(32'hbb56f9e8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb858f85d),
	.w1(32'hb8795097),
	.w2(32'hb71a5b8c),
	.w3(32'hb81d81ad),
	.w4(32'hb882e89b),
	.w5(32'hb81f6dc4),
	.w6(32'hb6eaea8a),
	.w7(32'hb833bb6a),
	.w8(32'hb7badc74),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37958fe7),
	.w1(32'h38334b84),
	.w2(32'hb64d31bd),
	.w3(32'hb82f0a7d),
	.w4(32'hb7a1db13),
	.w5(32'hb8794311),
	.w6(32'h38283a41),
	.w7(32'hb898b6e8),
	.w8(32'hb97f0c94),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36b344),
	.w1(32'hb97f864d),
	.w2(32'h3a0e5ca8),
	.w3(32'hbb31175a),
	.w4(32'hbada1511),
	.w5(32'hb9f5ad9d),
	.w6(32'hbb28aba7),
	.w7(32'hba42ee15),
	.w8(32'hb9ee909e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4bee8),
	.w1(32'h3b590fc7),
	.w2(32'hbb7c7b73),
	.w3(32'hb997903a),
	.w4(32'h3a9081c9),
	.w5(32'hbb948368),
	.w6(32'hbb8a5549),
	.w7(32'h3a74f4b6),
	.w8(32'hbb9c10d0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f8425),
	.w1(32'h3a80826c),
	.w2(32'h3a42ee7e),
	.w3(32'hba8dd34c),
	.w4(32'h39f98169),
	.w5(32'h39b7f5f7),
	.w6(32'hba40874d),
	.w7(32'h39f1242d),
	.w8(32'h388e0c29),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab644a8),
	.w1(32'h3aaa44f8),
	.w2(32'h39c23c3e),
	.w3(32'hba833f33),
	.w4(32'hb9d306c5),
	.w5(32'hba54b81f),
	.w6(32'hba2524df),
	.w7(32'h3a29e71d),
	.w8(32'hb932d5c3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a48a3b),
	.w1(32'h3a3f5748),
	.w2(32'h3af63879),
	.w3(32'hb98fe485),
	.w4(32'h39e72544),
	.w5(32'h3a8f3bf0),
	.w6(32'h3a8bbe2c),
	.w7(32'h3abe5fd0),
	.w8(32'h3acf1690),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb277171),
	.w1(32'hbaa9a312),
	.w2(32'hbba9561e),
	.w3(32'hbb3f6060),
	.w4(32'hb91133ee),
	.w5(32'hbbaa5e64),
	.w6(32'hbb5b4304),
	.w7(32'h3aaab33e),
	.w8(32'hbb176376),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a605d5d),
	.w1(32'h3a003e75),
	.w2(32'hbb2a78b6),
	.w3(32'hba050062),
	.w4(32'hb99fd0c8),
	.w5(32'hbb08280c),
	.w6(32'h3a18300a),
	.w7(32'h3ad02557),
	.w8(32'hba729f4b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b9c5cc),
	.w1(32'hb9673194),
	.w2(32'hbc089812),
	.w3(32'hb812db9c),
	.w4(32'h39991c54),
	.w5(32'hbbe18778),
	.w6(32'hba108630),
	.w7(32'h3a6243d2),
	.w8(32'hbbb21c56),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8edbcaa),
	.w1(32'h381aa11b),
	.w2(32'h3913cf8f),
	.w3(32'hb949937b),
	.w4(32'hb82feddf),
	.w5(32'h38a7a32f),
	.w6(32'hb8e28081),
	.w7(32'hb8ecb061),
	.w8(32'h37c7ca56),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ac688),
	.w1(32'hbb2caf2b),
	.w2(32'hbb679c47),
	.w3(32'hbb156a01),
	.w4(32'hbb3e6608),
	.w5(32'hbb89c541),
	.w6(32'hbaaaeb58),
	.w7(32'hbabf8bf0),
	.w8(32'hbb4f4824),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385055c2),
	.w1(32'hb4b11870),
	.w2(32'hb7f3c949),
	.w3(32'h386bfc69),
	.w4(32'h3604a7a8),
	.w5(32'hb7d44b80),
	.w6(32'h384fc093),
	.w7(32'hb68895d8),
	.w8(32'hb7d51421),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78759eb),
	.w1(32'h3920dcbd),
	.w2(32'hb9f6f94c),
	.w3(32'h3a012127),
	.w4(32'h39675008),
	.w5(32'h38879821),
	.w6(32'h3a5066ea),
	.w7(32'h3a0abd98),
	.w8(32'h39450177),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982f980),
	.w1(32'h39c495f8),
	.w2(32'hb7cbb5e9),
	.w3(32'hb980df41),
	.w4(32'hb7598bcb),
	.w5(32'hb89a8fdf),
	.w6(32'hb69f0289),
	.w7(32'hb8c45fda),
	.w8(32'hb996cfd7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ab4cc),
	.w1(32'hbadf6c82),
	.w2(32'hbb32c0c4),
	.w3(32'hbae731b3),
	.w4(32'hbb1adadb),
	.w5(32'hbb707f0d),
	.w6(32'hba7ce575),
	.w7(32'hbaab27f9),
	.w8(32'hbb157966),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371d7a39),
	.w1(32'hb5a25b3e),
	.w2(32'h366b0008),
	.w3(32'h357b2fe0),
	.w4(32'hb6b594c1),
	.w5(32'h36f6bc25),
	.w6(32'h36624691),
	.w7(32'hb6b1c041),
	.w8(32'h36671858),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3694cfa9),
	.w1(32'h37060203),
	.w2(32'h37c6e193),
	.w3(32'h37fe470f),
	.w4(32'hb63eeb62),
	.w5(32'hb7250bc8),
	.w6(32'hb726e61c),
	.w7(32'hb84a3041),
	.w8(32'hb628234e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9990d),
	.w1(32'hba71033f),
	.w2(32'h3a3098a6),
	.w3(32'hbad655e1),
	.w4(32'hbaaf4bf0),
	.w5(32'hb9c562af),
	.w6(32'hba17744f),
	.w7(32'hba667ebb),
	.w8(32'hba962891),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae26c42),
	.w1(32'h3a56fb2c),
	.w2(32'hbad570f4),
	.w3(32'hb9fd0eb8),
	.w4(32'h3b3a4b27),
	.w5(32'hbb0db01f),
	.w6(32'h3aae1706),
	.w7(32'h3b2c335b),
	.w8(32'hba3e5f91),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41a6ae),
	.w1(32'h3b93a542),
	.w2(32'h39caa4b6),
	.w3(32'hbb5d35f7),
	.w4(32'h3b400226),
	.w5(32'h3ac67121),
	.w6(32'hbb1b61ce),
	.w7(32'h3ab4d0ed),
	.w8(32'h3a466f32),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37421712),
	.w1(32'h392fa257),
	.w2(32'hb98b9726),
	.w3(32'hb924178b),
	.w4(32'h371c3a26),
	.w5(32'hb98c32bc),
	.w6(32'hb983f46b),
	.w7(32'h392c57a4),
	.w8(32'hb94d968f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23dd98),
	.w1(32'h3b544571),
	.w2(32'hbc527748),
	.w3(32'h3b97f7b7),
	.w4(32'h3bd6c00f),
	.w5(32'hbc273885),
	.w6(32'h399a6d58),
	.w7(32'h3ba52259),
	.w8(32'hbc0fe46f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01dfbc),
	.w1(32'hbbc9e13c),
	.w2(32'h3b4df8a7),
	.w3(32'hbc07dc49),
	.w4(32'hbc1a6593),
	.w5(32'hbb1a2427),
	.w6(32'h39f7be2e),
	.w7(32'hb9aa239c),
	.w8(32'h3aafa86a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f13d1),
	.w1(32'h3ae36ab9),
	.w2(32'hba668a5e),
	.w3(32'h3a5fcfcc),
	.w4(32'h3aa5a03f),
	.w5(32'hba15adff),
	.w6(32'h3a6256da),
	.w7(32'h3a9a52be),
	.w8(32'hba82d98c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384d43e2),
	.w1(32'hb79d3588),
	.w2(32'hb831968d),
	.w3(32'h384018f1),
	.w4(32'hb7a56dd8),
	.w5(32'hb7a87d8b),
	.w6(32'h37e4bc41),
	.w7(32'hb7534725),
	.w8(32'hb7f113a4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385b76af),
	.w1(32'h3704612f),
	.w2(32'h383c51f3),
	.w3(32'h38f01b0f),
	.w4(32'h383d904b),
	.w5(32'h381782c8),
	.w6(32'h37f9c1a8),
	.w7(32'hb540d610),
	.w8(32'h37fe6a60),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380ea799),
	.w1(32'hb6374b5a),
	.w2(32'hb76a8727),
	.w3(32'h380aaefc),
	.w4(32'hb697e283),
	.w5(32'hb79ad956),
	.w6(32'h37c52d6b),
	.w7(32'hb736583b),
	.w8(32'hb77220d2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f91ed),
	.w1(32'h3b29bc57),
	.w2(32'hbb0b3756),
	.w3(32'h3ab06e8e),
	.w4(32'h3b2f6d03),
	.w5(32'hbb02d7e3),
	.w6(32'hb9e9f119),
	.w7(32'h3a9cdd53),
	.w8(32'hbb4ceabc),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb140531),
	.w1(32'hba625bcd),
	.w2(32'hbb458dca),
	.w3(32'hba723a58),
	.w4(32'h38a4a35c),
	.w5(32'hbb1dde55),
	.w6(32'hbb047984),
	.w7(32'hba9f839e),
	.w8(32'hbb2d31d5),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad543bb),
	.w1(32'h3aa2d97d),
	.w2(32'hb8dc6684),
	.w3(32'hbb04fefa),
	.w4(32'hba20d289),
	.w5(32'hba0ff597),
	.w6(32'hbac6b575),
	.w7(32'h3a7ad88f),
	.w8(32'hb9e27bbd),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea38a0),
	.w1(32'h39e7d3db),
	.w2(32'h39d87cfd),
	.w3(32'hba46af44),
	.w4(32'hb8d1e201),
	.w5(32'h39a17b95),
	.w6(32'hb9ed980f),
	.w7(32'h3783810f),
	.w8(32'hb8849528),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964342a),
	.w1(32'h3b24909c),
	.w2(32'hbba79ae7),
	.w3(32'h3a37a8e8),
	.w4(32'h3b576688),
	.w5(32'hbb6b0119),
	.w6(32'hb9151fdc),
	.w7(32'h3b647d12),
	.w8(32'hbb34431b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb908cb2f),
	.w1(32'h3b385d6e),
	.w2(32'h3af354ad),
	.w3(32'hba443020),
	.w4(32'h3b090c96),
	.w5(32'h3b049ea4),
	.w6(32'h39a570ec),
	.w7(32'h3ae0d9bb),
	.w8(32'h3af94d83),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a4ebe1),
	.w1(32'hb78eb4f1),
	.w2(32'hb68722db),
	.w3(32'h37c7f5ce),
	.w4(32'hb709a053),
	.w5(32'h36fd832d),
	.w6(32'h37dcce72),
	.w7(32'hb786f2c6),
	.w8(32'hb6b2d8d4),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e9db7),
	.w1(32'hbb2b0d78),
	.w2(32'hbaf0611d),
	.w3(32'hb9e57674),
	.w4(32'hbb2e4d40),
	.w5(32'hbb0b7999),
	.w6(32'hbae51f24),
	.w7(32'hbad0a8f0),
	.w8(32'hbb2e3543),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38929647),
	.w1(32'hb848192f),
	.w2(32'hb7a052c3),
	.w3(32'h38bf282c),
	.w4(32'hb829175d),
	.w5(32'hb709c90a),
	.w6(32'h38a7fbf4),
	.w7(32'hb8222bec),
	.w8(32'hb79846ab),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba649c32),
	.w1(32'h3b0bb616),
	.w2(32'hb9177a73),
	.w3(32'hba651279),
	.w4(32'h3b1ac637),
	.w5(32'hb9b7232b),
	.w6(32'hba750e85),
	.w7(32'h3b438ebf),
	.w8(32'h3a702fc2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d81c6),
	.w1(32'hba41085a),
	.w2(32'h3b20b7b0),
	.w3(32'hbbb84db3),
	.w4(32'hbb8035f8),
	.w5(32'h39862c44),
	.w6(32'hbb2f8174),
	.w7(32'hbaad5935),
	.w8(32'hb9e01d65),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d0875),
	.w1(32'h3a1dfb65),
	.w2(32'h3834bc8f),
	.w3(32'hbb68a2f9),
	.w4(32'hb903a456),
	.w5(32'hb94465c9),
	.w6(32'hbb2577c4),
	.w7(32'h3a412092),
	.w8(32'h39adb5c1),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba726087),
	.w1(32'h380e2945),
	.w2(32'h3a82afae),
	.w3(32'hbaa47438),
	.w4(32'hb9ae03fc),
	.w5(32'h39ffd5f3),
	.w6(32'hba922560),
	.w7(32'hb9e1f29f),
	.w8(32'h3905582b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ad227),
	.w1(32'hbaf81c26),
	.w2(32'h3a84f66a),
	.w3(32'hbbafccf9),
	.w4(32'hbb7dc34d),
	.w5(32'hba811858),
	.w6(32'hbb5ce287),
	.w7(32'hbb04b5c5),
	.w8(32'h396ae87c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3696eeda),
	.w1(32'h3786a222),
	.w2(32'hbb58b978),
	.w3(32'hb9e34e97),
	.w4(32'h37315eb8),
	.w5(32'hbb52ba2f),
	.w6(32'hba98242d),
	.w7(32'h394fbafc),
	.w8(32'hbb3eadc3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b14f3),
	.w1(32'h3aec1622),
	.w2(32'hbbb3e2ef),
	.w3(32'h3abb2ac7),
	.w4(32'h3b59f2dd),
	.w5(32'hbb4ac33c),
	.w6(32'h3b1b5a6c),
	.w7(32'h3b82bfbd),
	.w8(32'hbb3c6f88),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380b1e61),
	.w1(32'h36b22c74),
	.w2(32'hb7e8460c),
	.w3(32'h387304ef),
	.w4(32'h382fe176),
	.w5(32'h37c89929),
	.w6(32'h3902e5d2),
	.w7(32'h3842beef),
	.w8(32'h35fc5fbe),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390be19e),
	.w1(32'h384f0198),
	.w2(32'h37cd75b5),
	.w3(32'h390d0b26),
	.w4(32'h37a2895c),
	.w5(32'hb8b629dd),
	.w6(32'h38e64b49),
	.w7(32'hb5eb8947),
	.w8(32'h3832be96),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c5bbb),
	.w1(32'h3b87bfbf),
	.w2(32'hbab2ea34),
	.w3(32'hbaaedf4f),
	.w4(32'h3abcfedd),
	.w5(32'hba9a9083),
	.w6(32'hbb4ff773),
	.w7(32'h3a75930c),
	.w8(32'hbb77c693),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14ef65),
	.w1(32'h3a89f7a0),
	.w2(32'hbb9b1726),
	.w3(32'hb98a33e3),
	.w4(32'h39c99265),
	.w5(32'hbbb1c44f),
	.w6(32'hbb4ad05a),
	.w7(32'h39cb3856),
	.w8(32'hbb9878fd),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dd8c2),
	.w1(32'hba1b2571),
	.w2(32'hbacf4df8),
	.w3(32'hbb93a4c8),
	.w4(32'hbae208e7),
	.w5(32'hbadaf05a),
	.w6(32'hbb524bed),
	.w7(32'h390d2763),
	.w8(32'hbacd5020),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a099e9b),
	.w1(32'h3af84615),
	.w2(32'hbbec47ce),
	.w3(32'hbab0c121),
	.w4(32'h3b86f2e1),
	.w5(32'hbbcce6e2),
	.w6(32'h3ba55d77),
	.w7(32'h3bd88e0f),
	.w8(32'hbb12da3b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399801f3),
	.w1(32'hba7975da),
	.w2(32'hba950963),
	.w3(32'hb822067c),
	.w4(32'hba2a39ac),
	.w5(32'hba90453f),
	.w6(32'hba5999b3),
	.w7(32'hba6b121c),
	.w8(32'hba9768d7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4434f6),
	.w1(32'h390981d1),
	.w2(32'hba7a4e90),
	.w3(32'hb8a924e3),
	.w4(32'hba1530f1),
	.w5(32'hbac735f5),
	.w6(32'hba17ab85),
	.w7(32'hba042986),
	.w8(32'hbac567b6),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22a34e),
	.w1(32'h3c8dc731),
	.w2(32'hba69c1d3),
	.w3(32'hbaa6eb82),
	.w4(32'h3c611fe4),
	.w5(32'hbb1b92cc),
	.w6(32'hbbb39a56),
	.w7(32'h3c29e117),
	.w8(32'hbb9fecc0),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f2496),
	.w1(32'h3b51a78e),
	.w2(32'hbc27116c),
	.w3(32'h3b39506d),
	.w4(32'h3b9f4128),
	.w5(32'hbbee5b30),
	.w6(32'h39e2d4e7),
	.w7(32'h3b838109),
	.w8(32'hbbf44d52),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7f169),
	.w1(32'h3af841dc),
	.w2(32'hbb488b44),
	.w3(32'h38f9e7c1),
	.w4(32'h39a833d6),
	.w5(32'hbb2806a1),
	.w6(32'hb9d8fda5),
	.w7(32'h3b0d4bb7),
	.w8(32'hbaeee4bb),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa93338),
	.w1(32'h3ac0c0b5),
	.w2(32'h3b66aa77),
	.w3(32'hbb3cb790),
	.w4(32'hba336d10),
	.w5(32'h3b14e08f),
	.w6(32'hb9e56f62),
	.w7(32'h3a5d1caa),
	.w8(32'h3ad04a67),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15f356),
	.w1(32'hbad10ed0),
	.w2(32'h3aa222a1),
	.w3(32'hbb3ad417),
	.w4(32'hbb86b93f),
	.w5(32'hbaa45898),
	.w6(32'hb8ef044c),
	.w7(32'hbacd1fe0),
	.w8(32'hbae4f4f2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378315fb),
	.w1(32'h3637b14f),
	.w2(32'h3618734a),
	.w3(32'h3746d4c3),
	.w4(32'h36827e10),
	.w5(32'h36bd0ea0),
	.w6(32'h37580615),
	.w7(32'h35a9d32e),
	.w8(32'h357e1a5a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3818c26b),
	.w1(32'h36d4201d),
	.w2(32'h3701d568),
	.w3(32'h3822c9fc),
	.w4(32'h372f8b0a),
	.w5(32'h373b7310),
	.w6(32'h3800c329),
	.w7(32'h363f921f),
	.w8(32'h359c1602),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78d4f9),
	.w1(32'h3a030282),
	.w2(32'hba97db8b),
	.w3(32'h39dbe6ad),
	.w4(32'h39b8623b),
	.w5(32'hbae4cf11),
	.w6(32'hba5ed580),
	.w7(32'hba3d2b6f),
	.w8(32'hbab6a9be),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38125b33),
	.w1(32'hb7019b9b),
	.w2(32'hb7a4e24a),
	.w3(32'h3838d330),
	.w4(32'hb6488c41),
	.w5(32'hb7670868),
	.w6(32'h380563b0),
	.w7(32'hb7993007),
	.w8(32'hb7c7fd7d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2eb310),
	.w1(32'h3b23226a),
	.w2(32'hba173ef2),
	.w3(32'h3b1292d0),
	.w4(32'h3ac46fdb),
	.w5(32'hb98310c0),
	.w6(32'h3a7cc660),
	.w7(32'h3a9d4dcc),
	.w8(32'hba65d15c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e447eb),
	.w1(32'h3a8822f7),
	.w2(32'hbba59084),
	.w3(32'hbb02b2f3),
	.w4(32'hb93d4e86),
	.w5(32'hbbfab64e),
	.w6(32'hbbde041c),
	.w7(32'hbb01cf72),
	.w8(32'hbbd5dae9),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb318a27),
	.w1(32'hb942a991),
	.w2(32'hba5190a3),
	.w3(32'hbb233d27),
	.w4(32'hba1fd242),
	.w5(32'hba7656bb),
	.w6(32'hbb07c4bd),
	.w7(32'hb9ea0b66),
	.w8(32'hba6ff004),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb505c221),
	.w1(32'hb751728e),
	.w2(32'hb6f789dd),
	.w3(32'hb4c0d73e),
	.w4(32'hb753fcb7),
	.w5(32'hb70a99e8),
	.w6(32'h37859736),
	.w7(32'hb688124e),
	.w8(32'hb6ecd5e2),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c90da),
	.w1(32'h3baf488b),
	.w2(32'hbb977fe0),
	.w3(32'h3914070e),
	.w4(32'h3b4b1f63),
	.w5(32'hbbaf11a4),
	.w6(32'hbb2778a3),
	.w7(32'h3b22531b),
	.w8(32'hbb791efc),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a944b8b),
	.w1(32'h3a6a7360),
	.w2(32'hbb8c0018),
	.w3(32'h3ab44355),
	.w4(32'h3a65246e),
	.w5(32'hbb796a51),
	.w6(32'hb8e0bf40),
	.w7(32'h3a954bf7),
	.w8(32'hbb450b95),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3888765e),
	.w1(32'hb8a862de),
	.w2(32'hb83990f2),
	.w3(32'hb5c50f7a),
	.w4(32'hb90e4c4d),
	.w5(32'hb886e728),
	.w6(32'hb8855b70),
	.w7(32'hb9069f26),
	.w8(32'hb85fad5c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f7beb),
	.w1(32'h3b3e209a),
	.w2(32'hbb6e117e),
	.w3(32'h3af5361a),
	.w4(32'h3b1bb085),
	.w5(32'hbb4f6136),
	.w6(32'h3a9d03ad),
	.w7(32'h3b25fdc8),
	.w8(32'hbb47e9c5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77f7995),
	.w1(32'hb6c0a1a9),
	.w2(32'hb7acb44c),
	.w3(32'hb69bff01),
	.w4(32'hb794ccc3),
	.w5(32'hb8001b57),
	.w6(32'hb7791861),
	.w7(32'hb80a29f6),
	.w8(32'hb7ddb38d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9294394),
	.w1(32'h3941c1da),
	.w2(32'h363a777e),
	.w3(32'hb95e85ac),
	.w4(32'hb6740aa2),
	.w5(32'hb8d56591),
	.w6(32'hb9288f91),
	.w7(32'h37991499),
	.w8(32'hb982f1a5),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3514155d),
	.w1(32'hb5ba9cea),
	.w2(32'h3714f97c),
	.w3(32'h36487745),
	.w4(32'h378de9f6),
	.w5(32'h37c4db7d),
	.w6(32'h37d9f08d),
	.w7(32'h37a85313),
	.w8(32'h38218acc),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385dc045),
	.w1(32'h389e6b4f),
	.w2(32'hb75715c1),
	.w3(32'h37558905),
	.w4(32'h383d73ee),
	.w5(32'hb8019b56),
	.w6(32'h38cfd071),
	.w7(32'h3845096f),
	.w8(32'hb7b11a19),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e63d91),
	.w1(32'h3a8f3db9),
	.w2(32'h3aa8c311),
	.w3(32'hbac5e435),
	.w4(32'hb945fab0),
	.w5(32'h39d1b3ef),
	.w6(32'hb989b305),
	.w7(32'h3743aa00),
	.w8(32'h3a3351c3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e10a78),
	.w1(32'hbaa29e1b),
	.w2(32'hbc1088a2),
	.w3(32'h3ac6befb),
	.w4(32'h399d146f),
	.w5(32'hbc0a8051),
	.w6(32'h3b43bd2f),
	.w7(32'h3b31be70),
	.w8(32'hbb87cc61),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c5ef2),
	.w1(32'h3b004c4d),
	.w2(32'hbba2f1d6),
	.w3(32'h3a1aaa98),
	.w4(32'h3ad6b00b),
	.w5(32'hbb90a5cf),
	.w6(32'hb90d68f6),
	.w7(32'h3ae2caf0),
	.w8(32'hbb81e578),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a887a49),
	.w1(32'h39dfea6d),
	.w2(32'hbbeb4a56),
	.w3(32'h3ab668fe),
	.w4(32'h3af8e187),
	.w5(32'hbbc452cb),
	.w6(32'h3ae30976),
	.w7(32'h3b692541),
	.w8(32'hbb521bc2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86770a9),
	.w1(32'h378f6ba4),
	.w2(32'h38c89e0a),
	.w3(32'hb910ae4b),
	.w4(32'hb8496906),
	.w5(32'h38abc3bb),
	.w6(32'hb8d195f1),
	.w7(32'hb22edd71),
	.w8(32'h3889f5b5),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394966e7),
	.w1(32'hb933cfef),
	.w2(32'hb9056665),
	.w3(32'hb853d4f8),
	.w4(32'hb77b3509),
	.w5(32'hb965e7e2),
	.w6(32'hb9b2a1e4),
	.w7(32'hb99e5348),
	.w8(32'hba213c99),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379834e2),
	.w1(32'hb7831500),
	.w2(32'hb6b9ced5),
	.w3(32'h381fdea6),
	.w4(32'h34beb219),
	.w5(32'h37580f0d),
	.w6(32'h3725a7e7),
	.w7(32'hb624109a),
	.w8(32'hb6959c0f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37469d3c),
	.w1(32'h372860c7),
	.w2(32'h37ab4725),
	.w3(32'h3747f55a),
	.w4(32'h379601ca),
	.w5(32'h37e99dcb),
	.w6(32'h37adcdf4),
	.w7(32'h377c8ed3),
	.w8(32'h3713a16a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86045b),
	.w1(32'hbb3f78bf),
	.w2(32'hbbbeb219),
	.w3(32'hbb3ed3dc),
	.w4(32'hbb439c3f),
	.w5(32'hbba62483),
	.w6(32'hbb44004f),
	.w7(32'hbb26e530),
	.w8(32'hbba230b5),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3878f108),
	.w1(32'h383de1f4),
	.w2(32'h38737075),
	.w3(32'h38bdcee5),
	.w4(32'h38ae7a67),
	.w5(32'h3861ff79),
	.w6(32'h38817634),
	.w7(32'h38471523),
	.w8(32'h386a706e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9ab0b),
	.w1(32'h3982bf98),
	.w2(32'h3a762a4d),
	.w3(32'hba48af9c),
	.w4(32'h38a7d3d7),
	.w5(32'h39fe0b2b),
	.w6(32'hba1e319b),
	.w7(32'hb869b766),
	.w8(32'h371a56a4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9f8bc),
	.w1(32'hba668f7a),
	.w2(32'h3a5fb68c),
	.w3(32'hba81da16),
	.w4(32'hba508ba6),
	.w5(32'h38c42889),
	.w6(32'hba08039c),
	.w7(32'hb998a094),
	.w8(32'hb9249f89),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38822a2a),
	.w1(32'h35e94571),
	.w2(32'h37b501fa),
	.w3(32'h389e0479),
	.w4(32'h380b8221),
	.w5(32'h37a99a02),
	.w6(32'h37c6ca0a),
	.w7(32'h37e78673),
	.w8(32'h378e1a77),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393bd113),
	.w1(32'h3a1424a9),
	.w2(32'hbadeb074),
	.w3(32'h39b0e851),
	.w4(32'h3a814340),
	.w5(32'hbaa031eb),
	.w6(32'h390747ef),
	.w7(32'h3a99ca5c),
	.w8(32'hba98188e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390715bd),
	.w1(32'hb8b3729c),
	.w2(32'hb9f4ff84),
	.w3(32'h37be716c),
	.w4(32'hb8abff4a),
	.w5(32'hba0f55d3),
	.w6(32'hb9814c23),
	.w7(32'hb9956eeb),
	.w8(32'hb9f0abae),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9566d2),
	.w1(32'hbba2e332),
	.w2(32'hbbc52271),
	.w3(32'hbad2e41b),
	.w4(32'hbbac0c19),
	.w5(32'hbc0d893b),
	.w6(32'hbb482551),
	.w7(32'hbb919b41),
	.w8(32'hbba482b1),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389195ba),
	.w1(32'hbabbae3b),
	.w2(32'hb938d20e),
	.w3(32'h37ba490f),
	.w4(32'hbab0847c),
	.w5(32'hbac8b96d),
	.w6(32'hb9aa3418),
	.w7(32'hb9ae190f),
	.w8(32'hbac10899),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb955624),
	.w1(32'h3acd4d82),
	.w2(32'h3ab8afd8),
	.w3(32'hbbd2aedc),
	.w4(32'hbadd11f5),
	.w5(32'h3995e132),
	.w6(32'hbb832eaa),
	.w7(32'hbb447544),
	.w8(32'hbae13e35),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule