module layer_10_featuremap_347(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a779174),
	.w1(32'h3a2f18e6),
	.w2(32'h3a8fedb2),
	.w3(32'hb99f79f8),
	.w4(32'hba25ea91),
	.w5(32'hba39450a),
	.w6(32'h3a0f8f88),
	.w7(32'hb8a4eef0),
	.w8(32'hba3c4055),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80027f),
	.w1(32'hbadd3510),
	.w2(32'h39a5bccb),
	.w3(32'h3a13ae6d),
	.w4(32'hba213ce9),
	.w5(32'h3bcc99c8),
	.w6(32'h3ab9a3ca),
	.w7(32'hbac7aef1),
	.w8(32'hba024b90),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0e191),
	.w1(32'h3ba81190),
	.w2(32'h3b933f2f),
	.w3(32'h3b242b33),
	.w4(32'h3ad898e3),
	.w5(32'hbae41855),
	.w6(32'h3a0b5cdd),
	.w7(32'h3a020975),
	.w8(32'hbae14c13),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0db0e7),
	.w1(32'h398b2eb2),
	.w2(32'hbaa01f39),
	.w3(32'hbaca4e05),
	.w4(32'hbababf2a),
	.w5(32'hbb1ed18e),
	.w6(32'hba531f07),
	.w7(32'hbacda994),
	.w8(32'hbb7f6388),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b53b3),
	.w1(32'hbb939e0e),
	.w2(32'hba1b6cf3),
	.w3(32'hbb6aeac3),
	.w4(32'hbb046ce7),
	.w5(32'hba30ab0f),
	.w6(32'hbb8be683),
	.w7(32'hbafa0b24),
	.w8(32'hba90d643),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4dfbe0),
	.w1(32'hba89ffe7),
	.w2(32'hba6104ea),
	.w3(32'hbabd5c2c),
	.w4(32'hbac25f32),
	.w5(32'hbb048d93),
	.w6(32'hba9bb94a),
	.w7(32'hba986c25),
	.w8(32'hbb11db10),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25d999),
	.w1(32'hbbc1c5fe),
	.w2(32'hbbc2e85b),
	.w3(32'hbb74ccac),
	.w4(32'hbbe63fe6),
	.w5(32'hbbd7bb5c),
	.w6(32'h39e08f6b),
	.w7(32'hbb9d975c),
	.w8(32'hbbe473e2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8b6a8),
	.w1(32'hbba6878b),
	.w2(32'hbb371694),
	.w3(32'hbbeebf0e),
	.w4(32'hbb27e515),
	.w5(32'h39f05800),
	.w6(32'h3a81a246),
	.w7(32'hba25246a),
	.w8(32'h3b633124),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeae58b),
	.w1(32'hbb338922),
	.w2(32'hbb2eda7e),
	.w3(32'hbb20a007),
	.w4(32'hbab9b805),
	.w5(32'hb94d9fab),
	.w6(32'hbb1de9c9),
	.w7(32'hba91d0f0),
	.w8(32'hb9811d64),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab90b81),
	.w1(32'h3a6ed27b),
	.w2(32'hbb04eaec),
	.w3(32'hbc0fcf1f),
	.w4(32'hbbc34f76),
	.w5(32'hbbc6777d),
	.w6(32'hbbb40475),
	.w7(32'hbaf835df),
	.w8(32'hbab6cc6b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad67376),
	.w1(32'hbaadf2d9),
	.w2(32'hbac9fafe),
	.w3(32'hba832b38),
	.w4(32'hbaee07c5),
	.w5(32'h3a0e6089),
	.w6(32'hb8e189b7),
	.w7(32'hbab24ba7),
	.w8(32'h3b851f4d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f8be3),
	.w1(32'h3bcd310f),
	.w2(32'h3b605b73),
	.w3(32'h3b151d5d),
	.w4(32'h3b4337d4),
	.w5(32'hbb03331e),
	.w6(32'h3c3a6893),
	.w7(32'h3c134797),
	.w8(32'hbab2d9a6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb463a),
	.w1(32'h3b5a9593),
	.w2(32'hba15f455),
	.w3(32'hbbb188a3),
	.w4(32'h385e5a7c),
	.w5(32'hbbd1ef7a),
	.w6(32'h3a4af27a),
	.w7(32'h3b781741),
	.w8(32'hbb791da9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97917d),
	.w1(32'hbb9146e1),
	.w2(32'h3a293972),
	.w3(32'hbaec8373),
	.w4(32'hbb15b4c5),
	.w5(32'hbb7e29f6),
	.w6(32'hbb46fb38),
	.w7(32'hbad6e387),
	.w8(32'hba708c36),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d4d2d),
	.w1(32'h3a4195a9),
	.w2(32'hba8daa1d),
	.w3(32'hbb641099),
	.w4(32'h3a9c4b27),
	.w5(32'h39fcab4d),
	.w6(32'hbb3704db),
	.w7(32'h3ac317b6),
	.w8(32'h39cb7e28),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b2c06),
	.w1(32'hb9ea2d15),
	.w2(32'h3ab8a08c),
	.w3(32'hbb78737f),
	.w4(32'h3a1280c6),
	.w5(32'h3a543d54),
	.w6(32'hbb828322),
	.w7(32'hb9af6888),
	.w8(32'h3b1ad097),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88f2b6),
	.w1(32'h3a3692df),
	.w2(32'h3a91a5fe),
	.w3(32'h3a5dff73),
	.w4(32'hb9522c2f),
	.w5(32'hbb29dd0e),
	.w6(32'hb88353b2),
	.w7(32'hba32253a),
	.w8(32'hbafb1d2e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18affc),
	.w1(32'hbb3de3c9),
	.w2(32'hbaf157ca),
	.w3(32'hbbd0998d),
	.w4(32'hbb302f7f),
	.w5(32'hbb05d9f2),
	.w6(32'hb911704c),
	.w7(32'h3aa96591),
	.w8(32'h3b0e7da7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ca82a),
	.w1(32'hbaec33c7),
	.w2(32'hbabd7cd7),
	.w3(32'h39a98662),
	.w4(32'hb7f78d66),
	.w5(32'hbb18a068),
	.w6(32'h3a49cf8d),
	.w7(32'h39e2c3bb),
	.w8(32'hb9eb23c4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60f5a7),
	.w1(32'hbb334dc2),
	.w2(32'hb9eb7cf6),
	.w3(32'hbb1c78d3),
	.w4(32'hbacb0d69),
	.w5(32'h3ac46254),
	.w6(32'hbb92cb72),
	.w7(32'hbaeb40d1),
	.w8(32'h3a3858bf),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374cea8e),
	.w1(32'hba4b6af2),
	.w2(32'h3a2281c0),
	.w3(32'h3aca2113),
	.w4(32'h3b88cc6f),
	.w5(32'hbb635d12),
	.w6(32'hb986878e),
	.w7(32'h398a30fa),
	.w8(32'hbb26572f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefb731),
	.w1(32'hba8fd8e2),
	.w2(32'hbb030bfd),
	.w3(32'hba913529),
	.w4(32'hbacdfd1a),
	.w5(32'hba50500b),
	.w6(32'hbab540d3),
	.w7(32'hbaf52c33),
	.w8(32'h38754e44),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e6c92),
	.w1(32'hbb677291),
	.w2(32'hba8823c4),
	.w3(32'hbc0e5253),
	.w4(32'h3a034e52),
	.w5(32'h3a6c1320),
	.w6(32'hbb0bed7e),
	.w7(32'h3a98a224),
	.w8(32'h3bac0a90),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992ae32),
	.w1(32'hba7d4b12),
	.w2(32'hb8b80734),
	.w3(32'hbbbcc08c),
	.w4(32'h3a36ac34),
	.w5(32'h3b4ccd4d),
	.w6(32'hbae464a5),
	.w7(32'h3b37e4ec),
	.w8(32'hbacc2476),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ccbfa),
	.w1(32'hba2cf6db),
	.w2(32'h3a1409ae),
	.w3(32'hbb4f480e),
	.w4(32'h3a896e74),
	.w5(32'h3ad2aaff),
	.w6(32'hbb20ec09),
	.w7(32'h3a4551c2),
	.w8(32'hba5da80e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb0458),
	.w1(32'h3acb1258),
	.w2(32'h3b33f365),
	.w3(32'hbb40d149),
	.w4(32'hba5056ac),
	.w5(32'h3a052f79),
	.w6(32'hbb277720),
	.w7(32'hb89aa798),
	.w8(32'hba786792),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9bd24),
	.w1(32'hb9555e9b),
	.w2(32'h3ad64337),
	.w3(32'hba15f582),
	.w4(32'hba99fceb),
	.w5(32'hbaa939be),
	.w6(32'hbb150732),
	.w7(32'hb9da1040),
	.w8(32'hbb22f335),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95eb67),
	.w1(32'hbbc2b0fa),
	.w2(32'hbb106da4),
	.w3(32'hbbb2ded2),
	.w4(32'hbc011251),
	.w5(32'h3b43ee55),
	.w6(32'hbbc0f74e),
	.w7(32'hbb2134a6),
	.w8(32'h3ac7e496),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a091358),
	.w1(32'hbae22ea2),
	.w2(32'hbb190a82),
	.w3(32'h3ae9b290),
	.w4(32'hba581847),
	.w5(32'h3b3dba6f),
	.w6(32'hbb02575b),
	.w7(32'hbaa29f85),
	.w8(32'h3b0fbfe4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eac9d6),
	.w1(32'h3ad99127),
	.w2(32'h39ed7989),
	.w3(32'hbbe61cf3),
	.w4(32'hbbb9d8d7),
	.w5(32'hbbc9d925),
	.w6(32'hbc01da87),
	.w7(32'hbb12332e),
	.w8(32'h3b88275b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6318dd),
	.w1(32'hbb46dd6a),
	.w2(32'hb9ef2e90),
	.w3(32'h3a9897b2),
	.w4(32'hba44c349),
	.w5(32'h3a86cdec),
	.w6(32'h3be6d9ae),
	.w7(32'hb9e25a5c),
	.w8(32'hb9e9b98a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c6e39e),
	.w1(32'hbaa6cecc),
	.w2(32'h395fe1f8),
	.w3(32'h3a44cad6),
	.w4(32'h387c2819),
	.w5(32'hba023965),
	.w6(32'hbaeb5689),
	.w7(32'h3ab6cae1),
	.w8(32'hbb29ff91),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba076e81),
	.w1(32'h39146e34),
	.w2(32'h3a3a1ba3),
	.w3(32'h39cf47a8),
	.w4(32'hbb218058),
	.w5(32'hbba9a727),
	.w6(32'hbafbb81c),
	.w7(32'h3a6075a5),
	.w8(32'hba9b51c9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba866098),
	.w1(32'hbabc02c1),
	.w2(32'hbb83efb1),
	.w3(32'hbb6143f5),
	.w4(32'hba66817a),
	.w5(32'hbaf58827),
	.w6(32'hbad60ba3),
	.w7(32'hba87072b),
	.w8(32'hbb0a8372),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c47cb2),
	.w1(32'hbb2e2289),
	.w2(32'hba1707a8),
	.w3(32'hbbb070ca),
	.w4(32'hbb555d90),
	.w5(32'hb7da3352),
	.w6(32'hbb65d080),
	.w7(32'hbab67fdb),
	.w8(32'hba1da2e4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace2552),
	.w1(32'hbbd83dbe),
	.w2(32'hbb43bc09),
	.w3(32'hbb09b736),
	.w4(32'h3b031764),
	.w5(32'hbaeff87b),
	.w6(32'h3b6d61cf),
	.w7(32'hbb4e4766),
	.w8(32'hb9fd3f42),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ae16c),
	.w1(32'h398e0552),
	.w2(32'h3a662698),
	.w3(32'hbb880b99),
	.w4(32'hbb8a1a15),
	.w5(32'hbb356acf),
	.w6(32'hbbde916c),
	.w7(32'h3b03e53f),
	.w8(32'hbba47ab4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc783ea9),
	.w1(32'hbba8d641),
	.w2(32'hbab0e1af),
	.w3(32'hbb979877),
	.w4(32'hb98b2bd8),
	.w5(32'h3b80fe79),
	.w6(32'hbb0b384e),
	.w7(32'h3a4f39fe),
	.w8(32'h3b1335aa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb772d98),
	.w1(32'hbb85eff9),
	.w2(32'h3afb9c00),
	.w3(32'h3a95e026),
	.w4(32'hb9ca8ad7),
	.w5(32'h3b97f692),
	.w6(32'h3ad28d4a),
	.w7(32'hbaa19d66),
	.w8(32'h3babd54f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2b199),
	.w1(32'hbbca6f86),
	.w2(32'hbbca4e53),
	.w3(32'hbb66f4d6),
	.w4(32'hbb75c6d5),
	.w5(32'h3b08cd10),
	.w6(32'hbb7f400b),
	.w7(32'hbb4b257e),
	.w8(32'h3b91c793),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b897b44),
	.w1(32'h3b19e187),
	.w2(32'hb93db080),
	.w3(32'h3b43bd14),
	.w4(32'h3b0cd115),
	.w5(32'h386cb5ad),
	.w6(32'h3bb475d8),
	.w7(32'h3b0121a9),
	.w8(32'hba711ac2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10b30f),
	.w1(32'h38c23524),
	.w2(32'h3a90f045),
	.w3(32'hba9e0312),
	.w4(32'hba9fcc65),
	.w5(32'h3b081611),
	.w6(32'hb714dd6e),
	.w7(32'hba69373b),
	.w8(32'h3bc12657),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91a18b),
	.w1(32'h3bbde12a),
	.w2(32'h3bb4fb08),
	.w3(32'h3bd97c9b),
	.w4(32'h3bc084dd),
	.w5(32'h3b656620),
	.w6(32'h3b9cb44a),
	.w7(32'h3bea597c),
	.w8(32'h3aea371d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a687ed),
	.w1(32'hbbb9f0a2),
	.w2(32'hbb12ff16),
	.w3(32'hbbcc2bd3),
	.w4(32'hbb89a991),
	.w5(32'hbab45c58),
	.w6(32'hba0c3686),
	.w7(32'h3ab1f5d9),
	.w8(32'h3b8c2ec0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb737919),
	.w1(32'hbaf42a2d),
	.w2(32'hbabf54c2),
	.w3(32'hbae93977),
	.w4(32'hbaf5c61c),
	.w5(32'h3a571c71),
	.w6(32'hbbc44dfb),
	.w7(32'hbb4f11d6),
	.w8(32'h3b0a33ca),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac832c),
	.w1(32'h3aef752c),
	.w2(32'h398fcac4),
	.w3(32'hbac89bcb),
	.w4(32'hbb063bf9),
	.w5(32'hba993227),
	.w6(32'h3b098660),
	.w7(32'h3b0cc4af),
	.w8(32'h39ac7031),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf978b),
	.w1(32'hbaf20fe4),
	.w2(32'hba41922e),
	.w3(32'hbb2c2cc0),
	.w4(32'hbac12cf8),
	.w5(32'hb9b98ed6),
	.w6(32'hbb6e4bc4),
	.w7(32'hbac9c733),
	.w8(32'h3a043da9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dd37c),
	.w1(32'hbac3d7f8),
	.w2(32'hbaebd899),
	.w3(32'hbb31f721),
	.w4(32'hbbaf6ee0),
	.w5(32'hbbe94a57),
	.w6(32'h3ac42dc5),
	.w7(32'h3a8fc223),
	.w8(32'h3ab230cc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba994da),
	.w1(32'h3b32001f),
	.w2(32'h3a0abfc9),
	.w3(32'h3ae1e511),
	.w4(32'h3b8d4342),
	.w5(32'hbb3dca3b),
	.w6(32'h3b9319e8),
	.w7(32'h3b6bb1c6),
	.w8(32'hbae8f2cb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb195e53),
	.w1(32'hb9ed300f),
	.w2(32'hbaafbf7b),
	.w3(32'hbb4175ae),
	.w4(32'hbad7a411),
	.w5(32'hbb01d442),
	.w6(32'hbb3359a2),
	.w7(32'hbab705d2),
	.w8(32'hbbb361ff),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb968435),
	.w1(32'hbb015d4c),
	.w2(32'h3b55944b),
	.w3(32'hbace262f),
	.w4(32'h382f8fbe),
	.w5(32'hb93bd7a0),
	.w6(32'hbb5a2f9e),
	.w7(32'h3a4995a8),
	.w8(32'h39f3e4c7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad25310),
	.w1(32'hbaa07204),
	.w2(32'hba0c9961),
	.w3(32'hb8f4c133),
	.w4(32'hba718cd5),
	.w5(32'hba6725f4),
	.w6(32'h3a843726),
	.w7(32'hba3f1588),
	.w8(32'h3b8bddcc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89bf717),
	.w1(32'hba44620b),
	.w2(32'h3b11bc96),
	.w3(32'h3a939c82),
	.w4(32'hbb0d6348),
	.w5(32'h37ba7142),
	.w6(32'h3b7b2184),
	.w7(32'h3adef0dc),
	.w8(32'hb996d42b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb018a5),
	.w1(32'hba874c23),
	.w2(32'hba5ed6e3),
	.w3(32'hbc2064ac),
	.w4(32'hbbdb7238),
	.w5(32'h382509c0),
	.w6(32'hbab8089a),
	.w7(32'h3b3f32db),
	.w8(32'h3b7d0f83),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb338b24),
	.w1(32'hbb8f98ed),
	.w2(32'hbb07c74e),
	.w3(32'hba8002dc),
	.w4(32'h38aeb668),
	.w5(32'h3a5054df),
	.w6(32'hbb1f30dd),
	.w7(32'hbae4dfde),
	.w8(32'hb992b010),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b0e6b),
	.w1(32'h3a92f93c),
	.w2(32'h3b0c7a70),
	.w3(32'hbafbc666),
	.w4(32'hbaed8c60),
	.w5(32'hb9a1de5c),
	.w6(32'hbb66569b),
	.w7(32'hbb22108e),
	.w8(32'h398b33eb),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ecb5c),
	.w1(32'h3a1c5c4f),
	.w2(32'hba6a4f67),
	.w3(32'h3ad92c20),
	.w4(32'h3a26bea5),
	.w5(32'hba64d34b),
	.w6(32'h39c5bb98),
	.w7(32'hbad2423e),
	.w8(32'hbac48cc1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb106628),
	.w1(32'hba4bbeac),
	.w2(32'hbab2db6e),
	.w3(32'hba8ed26a),
	.w4(32'hbb22088e),
	.w5(32'hbaf89488),
	.w6(32'h38a68186),
	.w7(32'hba7e5b86),
	.w8(32'hbb0f766e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd8c25),
	.w1(32'hba5226a8),
	.w2(32'hbacbd513),
	.w3(32'hbae11fcd),
	.w4(32'hba81c527),
	.w5(32'hba2fd115),
	.w6(32'hbac3c3ec),
	.w7(32'hba8d3b39),
	.w8(32'hbaba21b5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62b64c),
	.w1(32'hb8ded1ce),
	.w2(32'hbb20e146),
	.w3(32'hba3b1075),
	.w4(32'hbba372ca),
	.w5(32'hba614c2c),
	.w6(32'h3991a24b),
	.w7(32'hbb35ea82),
	.w8(32'hbad4c18e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab32f29),
	.w1(32'hbb1e782b),
	.w2(32'hb907983a),
	.w3(32'hbb4a9ead),
	.w4(32'hbb46c71a),
	.w5(32'hbb471e44),
	.w6(32'hbab92f28),
	.w7(32'hbaaa3946),
	.w8(32'hbac2b92b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57ceed),
	.w1(32'hba051b84),
	.w2(32'hba59dd7c),
	.w3(32'hbbd33fe2),
	.w4(32'hbafccf8b),
	.w5(32'hbb812371),
	.w6(32'hbaee4890),
	.w7(32'hb93016b8),
	.w8(32'hb9923046),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1d08d),
	.w1(32'hba071d2d),
	.w2(32'h3a608979),
	.w3(32'hbb27f636),
	.w4(32'hbb3c9fe5),
	.w5(32'hba48ab43),
	.w6(32'hbaaaf0a9),
	.w7(32'hbae080d8),
	.w8(32'hb95e499f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17672b),
	.w1(32'hbaf6c9f7),
	.w2(32'hba04220e),
	.w3(32'hb90c58bd),
	.w4(32'hb9efcb3c),
	.w5(32'hbb2995a6),
	.w6(32'hbaf2b179),
	.w7(32'hbaeed362),
	.w8(32'hbae53213),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae58038),
	.w1(32'hbb5a7386),
	.w2(32'hbb051e12),
	.w3(32'hbb307814),
	.w4(32'hb9cd7747),
	.w5(32'h3aad3416),
	.w6(32'hbb6b9386),
	.w7(32'hba9ac084),
	.w8(32'h3b5c80d2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cbda6),
	.w1(32'hba9471e4),
	.w2(32'h39b1551b),
	.w3(32'h3adac70d),
	.w4(32'h3b1cdae1),
	.w5(32'h395347dc),
	.w6(32'h3b77b4e2),
	.w7(32'h3afdcd10),
	.w8(32'hbad72c95),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ca660),
	.w1(32'hb714afd0),
	.w2(32'h3a17aae2),
	.w3(32'hbb5e97b0),
	.w4(32'hbbb8d4ce),
	.w5(32'h398c95fa),
	.w6(32'h39119639),
	.w7(32'hbb12ccd7),
	.w8(32'h3b8b9178),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937496f),
	.w1(32'hbb34f396),
	.w2(32'h3a58f783),
	.w3(32'h3a40ad1d),
	.w4(32'h3a5d4c79),
	.w5(32'hbb30051a),
	.w6(32'h3b2edec8),
	.w7(32'h3b6e9621),
	.w8(32'hb9d4c871),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb4eac),
	.w1(32'hbbddbfaa),
	.w2(32'hb890da22),
	.w3(32'hbb4526bf),
	.w4(32'hba475cd6),
	.w5(32'h3bb7124c),
	.w6(32'h36beab94),
	.w7(32'h3a2b3ec8),
	.w8(32'h3c00f772),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb627b77),
	.w1(32'hba94b4cf),
	.w2(32'hbbb65982),
	.w3(32'hbaa0f774),
	.w4(32'h3c04c172),
	.w5(32'h3b29da2c),
	.w6(32'h3b953327),
	.w7(32'hba4cd01d),
	.w8(32'h3b7c487f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ac6872),
	.w1(32'hb93103c3),
	.w2(32'h3ab69613),
	.w3(32'h3a9e1a80),
	.w4(32'hba2a7fa8),
	.w5(32'h3ade3c99),
	.w6(32'h3a19ac61),
	.w7(32'h3a4412e8),
	.w8(32'h39cfde05),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32715e),
	.w1(32'h3984949f),
	.w2(32'h3af83337),
	.w3(32'h3a42cad7),
	.w4(32'h3b354533),
	.w5(32'hbb1396de),
	.w6(32'h3b2c7b5b),
	.w7(32'hb9b6270d),
	.w8(32'h3ad99bae),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb215b24),
	.w1(32'hbae56447),
	.w2(32'hb8b56180),
	.w3(32'hbacff892),
	.w4(32'hbac45798),
	.w5(32'hba6af1fa),
	.w6(32'h3b1b535b),
	.w7(32'hbb8057da),
	.w8(32'h3b37211a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b954e6d),
	.w1(32'h3b4c011a),
	.w2(32'h3a8baf9f),
	.w3(32'h3aa1b506),
	.w4(32'h3b3eede4),
	.w5(32'h3ac2739f),
	.w6(32'h3bf8e913),
	.w7(32'h3b9e6c0c),
	.w8(32'hbab341ff),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba666190),
	.w1(32'hba884ad4),
	.w2(32'hba64f1ae),
	.w3(32'hb84e3fa2),
	.w4(32'hba2f53f1),
	.w5(32'h3a85d47d),
	.w6(32'h3a672406),
	.w7(32'hba4baef1),
	.w8(32'h3b4b2963),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be54119),
	.w1(32'h3b23682a),
	.w2(32'h3ac80680),
	.w3(32'h3b46ba3d),
	.w4(32'h3b8f8930),
	.w5(32'hbb4f0bce),
	.w6(32'h3b9a6959),
	.w7(32'h3b8d7e55),
	.w8(32'h3af20a18),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3088e7),
	.w1(32'hbb1a2dd2),
	.w2(32'hbb0e0517),
	.w3(32'hb9bf9aa4),
	.w4(32'hbab1982f),
	.w5(32'hbb47a8e5),
	.w6(32'h3be6c875),
	.w7(32'h3b164d93),
	.w8(32'h3ad3a49d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba915cb3),
	.w1(32'hbaf9c6e0),
	.w2(32'hbad7017b),
	.w3(32'h3afc3a17),
	.w4(32'h3b4fbfb2),
	.w5(32'hbb2952e0),
	.w6(32'h3b10079c),
	.w7(32'hb935889d),
	.w8(32'hbad8af5a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae70c49),
	.w1(32'h38071ccf),
	.w2(32'hbb2b0f50),
	.w3(32'hba62c146),
	.w4(32'h3934f869),
	.w5(32'hba5e1e12),
	.w6(32'h3b89ba48),
	.w7(32'h3ad02a1a),
	.w8(32'hbad81e24),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3957cdc6),
	.w1(32'hbb0c2448),
	.w2(32'hbab2f2a8),
	.w3(32'hbb44f08a),
	.w4(32'hbb9a25e2),
	.w5(32'hb98c5ad6),
	.w6(32'hba18a665),
	.w7(32'hbb048dee),
	.w8(32'h3b538a79),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c130af4),
	.w1(32'h3bc256ad),
	.w2(32'h3b59912d),
	.w3(32'h3ae3a856),
	.w4(32'h3bb7c47e),
	.w5(32'hbb1be2e3),
	.w6(32'h3af063f5),
	.w7(32'h3bb13bcb),
	.w8(32'h3a9cf599),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a199e),
	.w1(32'h3b079ba0),
	.w2(32'hba390623),
	.w3(32'h3a917767),
	.w4(32'h3b827354),
	.w5(32'hbb40d1cf),
	.w6(32'h3baeeda3),
	.w7(32'h3b224005),
	.w8(32'hbabab9ff),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a973660),
	.w1(32'hba167ff8),
	.w2(32'h3a0448c6),
	.w3(32'h39957c80),
	.w4(32'hbaef83fe),
	.w5(32'h3b4088f8),
	.w6(32'h38df72b1),
	.w7(32'hbab3c297),
	.w8(32'h3b51ef8c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a985642),
	.w1(32'h3b346817),
	.w2(32'h3b521ee8),
	.w3(32'h3b183597),
	.w4(32'h39d37db1),
	.w5(32'h3aa4f80c),
	.w6(32'h3aceea1b),
	.w7(32'h3b072c5d),
	.w8(32'h39e8cae1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af70c81),
	.w1(32'h3af078f4),
	.w2(32'h3b5e6ce7),
	.w3(32'h3978c355),
	.w4(32'hb9236b5b),
	.w5(32'h3968b65b),
	.w6(32'h3b13d9d2),
	.w7(32'h3ab1f30a),
	.w8(32'hbb01a2da),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69f7a5),
	.w1(32'hbb7cb1bc),
	.w2(32'hb9ad86c3),
	.w3(32'hb9ea057c),
	.w4(32'h3936d522),
	.w5(32'h3ac79267),
	.w6(32'h3a26bd7c),
	.w7(32'h395f34e0),
	.w8(32'h3a2035a8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb965d07),
	.w1(32'hbae4c6d4),
	.w2(32'hbb1b5738),
	.w3(32'hbb13760f),
	.w4(32'h39b35f17),
	.w5(32'h3ad03ee3),
	.w6(32'hbb626b0c),
	.w7(32'hbabc1c42),
	.w8(32'hba921121),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ff4648),
	.w1(32'hb9847899),
	.w2(32'h3b080d05),
	.w3(32'hb9fd875e),
	.w4(32'hbaf99b9d),
	.w5(32'hbaa72a72),
	.w6(32'hbb048606),
	.w7(32'hbade4866),
	.w8(32'hbad5fc7d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ce4c2),
	.w1(32'hbb6dd735),
	.w2(32'hbb454973),
	.w3(32'hbb90bf7a),
	.w4(32'hbb37f0d0),
	.w5(32'h3a451c71),
	.w6(32'hbb95cc7e),
	.w7(32'hbaa70685),
	.w8(32'h3acfaab8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cee50),
	.w1(32'h3b402ed1),
	.w2(32'hb9aba507),
	.w3(32'h3a667669),
	.w4(32'h39f636a9),
	.w5(32'hba0ff083),
	.w6(32'h3b8c6940),
	.w7(32'h3b0193e9),
	.w8(32'h39d462e3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5c618),
	.w1(32'h38f0936f),
	.w2(32'h3af525b0),
	.w3(32'h3a648963),
	.w4(32'h3aa297c4),
	.w5(32'h3b78a92b),
	.w6(32'h3998a14d),
	.w7(32'h3b2955f0),
	.w8(32'h3add2072),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02f10b),
	.w1(32'hbae30086),
	.w2(32'hb8317614),
	.w3(32'hbbf3e9ee),
	.w4(32'hbb7ea31b),
	.w5(32'hba9a4d54),
	.w6(32'hbb895be8),
	.w7(32'h3b5116ab),
	.w8(32'hbb13a3d7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd48646),
	.w1(32'hbb98eeaa),
	.w2(32'h3ac8145c),
	.w3(32'hbae011d4),
	.w4(32'hbabff6d3),
	.w5(32'h3b085548),
	.w6(32'hbbb7dbef),
	.w7(32'h39ca1fb8),
	.w8(32'h3a75f183),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a6db8),
	.w1(32'hbba0218a),
	.w2(32'hba8ba9b9),
	.w3(32'hbb6fccbe),
	.w4(32'hbaf85c09),
	.w5(32'h3b8dbc8c),
	.w6(32'hba7895ba),
	.w7(32'hba4811f6),
	.w8(32'h3b85293d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f8267),
	.w1(32'h3b05d57a),
	.w2(32'h3b29a382),
	.w3(32'h3ab1a969),
	.w4(32'h3b42cea8),
	.w5(32'h3b8dcf9a),
	.w6(32'h3b420a6f),
	.w7(32'h3b08c991),
	.w8(32'h3b1b17eb),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99dd92),
	.w1(32'hb9d32740),
	.w2(32'h3b8a0082),
	.w3(32'h38c826ce),
	.w4(32'h3aeb191b),
	.w5(32'h3b2459c2),
	.w6(32'hba419f27),
	.w7(32'h3bc5d757),
	.w8(32'h3bc9921d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40681d),
	.w1(32'h3accb443),
	.w2(32'h3a357e68),
	.w3(32'h3b909b0b),
	.w4(32'hba3e81be),
	.w5(32'hbb0b30d0),
	.w6(32'h3b61ace4),
	.w7(32'h3acb2c5b),
	.w8(32'h3b5ecde9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b691cb),
	.w1(32'hbb4c18aa),
	.w2(32'hbac8e47a),
	.w3(32'hbb913a06),
	.w4(32'h3ace487f),
	.w5(32'hba32f0d8),
	.w6(32'h3b120bc6),
	.w7(32'h3ad2ea00),
	.w8(32'hba386613),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9630de),
	.w1(32'hbb527c9b),
	.w2(32'h39ac0836),
	.w3(32'hbbc680aa),
	.w4(32'h3b352372),
	.w5(32'hbb6d7d43),
	.w6(32'hbb895841),
	.w7(32'h3bacf9af),
	.w8(32'hb9a9d0c8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8544d),
	.w1(32'hbc07d3e5),
	.w2(32'h3a1f2e09),
	.w3(32'h3a8c1fc8),
	.w4(32'hbb3adf62),
	.w5(32'hbbf9d9f6),
	.w6(32'h3c0a937d),
	.w7(32'h3a3cdcf9),
	.w8(32'h3b02230f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78e021),
	.w1(32'hbc5eb8cc),
	.w2(32'hbbe6dfbc),
	.w3(32'hbc272196),
	.w4(32'h3bba96ad),
	.w5(32'h3ba4f5f7),
	.w6(32'hbc831ca5),
	.w7(32'h3c228dd8),
	.w8(32'h3b674a4d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44ef99),
	.w1(32'hbc744c98),
	.w2(32'hbc647157),
	.w3(32'hbc491714),
	.w4(32'hb9dcef47),
	.w5(32'hbb384ccc),
	.w6(32'hbc5386f3),
	.w7(32'hbb6410f2),
	.w8(32'h3b2e1629),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e2a87),
	.w1(32'hbb4043a4),
	.w2(32'hba85ce9a),
	.w3(32'hbc2384aa),
	.w4(32'h3a4256a6),
	.w5(32'hbab5cf15),
	.w6(32'hbbe558fb),
	.w7(32'h3b62d5cf),
	.w8(32'h3c2a407b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20bb92),
	.w1(32'h3b171145),
	.w2(32'hbb6aae9e),
	.w3(32'hbc43da3d),
	.w4(32'hbb893688),
	.w5(32'hbbd163ea),
	.w6(32'hbaac9137),
	.w7(32'hbc2534c7),
	.w8(32'hbb3c89c3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36f824),
	.w1(32'hbb76dbda),
	.w2(32'hbbb268f4),
	.w3(32'h3afcbc26),
	.w4(32'h3b97b87c),
	.w5(32'hbba9bad3),
	.w6(32'hbc229a68),
	.w7(32'h3c3ba883),
	.w8(32'h3b241aa1),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dc649),
	.w1(32'h3b2f799e),
	.w2(32'hbb716b68),
	.w3(32'hbabb3dde),
	.w4(32'hbc064233),
	.w5(32'hbb515056),
	.w6(32'h3ac1ad55),
	.w7(32'hbbec813d),
	.w8(32'hbba49be4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadeca99),
	.w1(32'h3aee8fb7),
	.w2(32'h3ac2099c),
	.w3(32'h3b007a2c),
	.w4(32'h3c0c866a),
	.w5(32'hb9ff82f9),
	.w6(32'hb93ec980),
	.w7(32'h3bca70d2),
	.w8(32'h3915b2b2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4760dd),
	.w1(32'hbb3839bf),
	.w2(32'hbb93fc36),
	.w3(32'hba562f81),
	.w4(32'hbadc5805),
	.w5(32'hb8bf98bb),
	.w6(32'hbb43c774),
	.w7(32'hbb48136b),
	.w8(32'hbb2006a3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e91be),
	.w1(32'h3a0366b0),
	.w2(32'h39af5f73),
	.w3(32'hbc062e19),
	.w4(32'h3b56e865),
	.w5(32'h3b924cfa),
	.w6(32'hbb955e3c),
	.w7(32'h3b5f8ce6),
	.w8(32'h3b4a88ce),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4723f1),
	.w1(32'h3bb2899f),
	.w2(32'h3aaa6548),
	.w3(32'hbb80377e),
	.w4(32'hbb0eff79),
	.w5(32'hbbd53f9f),
	.w6(32'h380b1cec),
	.w7(32'h3abb0a59),
	.w8(32'hbb6e385f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc346a86),
	.w1(32'hbbcf0d48),
	.w2(32'hb8c4a00c),
	.w3(32'hbb9b64f9),
	.w4(32'h3a23e50e),
	.w5(32'h3c19c37c),
	.w6(32'hbab49f1e),
	.w7(32'h3b772c2a),
	.w8(32'h3b22499b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9c05d),
	.w1(32'h3c892876),
	.w2(32'hbbfb235b),
	.w3(32'h3b83144f),
	.w4(32'hbc6d7573),
	.w5(32'h3ba57474),
	.w6(32'h3c5d7587),
	.w7(32'hbc9ec7c4),
	.w8(32'h3b644fb7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39deaf20),
	.w1(32'hbad49bf0),
	.w2(32'h3af25cf2),
	.w3(32'h3c082caa),
	.w4(32'h3bca3621),
	.w5(32'h3c169bf1),
	.w6(32'h3b880512),
	.w7(32'h3c1a42cb),
	.w8(32'h3cdb15d9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba963bfb),
	.w1(32'h3c202ad3),
	.w2(32'h3bd9612a),
	.w3(32'hbc8bd56e),
	.w4(32'hbc71c8bb),
	.w5(32'hb7e34455),
	.w6(32'h3bf09327),
	.w7(32'hbc306f7c),
	.w8(32'hbbad76a7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99bfd0),
	.w1(32'h3b5f9b89),
	.w2(32'hba56824b),
	.w3(32'hbaa71739),
	.w4(32'hba790fb8),
	.w5(32'hbbde5908),
	.w6(32'h3b1e5d9b),
	.w7(32'h3ad74965),
	.w8(32'hbbee26eb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb936309f),
	.w1(32'h3ba72f8a),
	.w2(32'hbbbcba82),
	.w3(32'h3b8a7472),
	.w4(32'h3b304e9c),
	.w5(32'hb95da7a4),
	.w6(32'hbaa8d0aa),
	.w7(32'hbc1867c6),
	.w8(32'h3ac3e4ec),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b0236),
	.w1(32'h3aa78687),
	.w2(32'hba1150de),
	.w3(32'h3b1b06cf),
	.w4(32'h3b5a13ea),
	.w5(32'h3b0bfb69),
	.w6(32'hb6cc348a),
	.w7(32'hb790b902),
	.w8(32'hbbc508b1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2a0d3),
	.w1(32'hbb5a64dc),
	.w2(32'h3a245db4),
	.w3(32'h3b9be74c),
	.w4(32'hb9301b1f),
	.w5(32'hbb34982c),
	.w6(32'h3c14426a),
	.w7(32'h3ba5cfe3),
	.w8(32'hbba5866c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47d44b),
	.w1(32'hbbb0849d),
	.w2(32'hba8a64be),
	.w3(32'hbb4b9448),
	.w4(32'h3b190928),
	.w5(32'h3beadbc5),
	.w6(32'hbc06165e),
	.w7(32'h3ab02f3a),
	.w8(32'h3c40a00b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fa644),
	.w1(32'h3b1679ee),
	.w2(32'hbb198efd),
	.w3(32'hbb2fa8d9),
	.w4(32'hbbc294e7),
	.w5(32'hbb18e1d1),
	.w6(32'h39766476),
	.w7(32'hbc0bf887),
	.w8(32'hbc004bb0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7644dd),
	.w1(32'h3c08f395),
	.w2(32'h3b0609bf),
	.w3(32'h3c9c6822),
	.w4(32'hb9b75907),
	.w5(32'hbb2778b5),
	.w6(32'hbaf8d2ca),
	.w7(32'hbbda146e),
	.w8(32'hbbad335c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ba7c6),
	.w1(32'hbb28e71b),
	.w2(32'hb96f2516),
	.w3(32'h39cf0e9c),
	.w4(32'h3bb11e47),
	.w5(32'hb79dd8c1),
	.w6(32'h3ae5f274),
	.w7(32'h3bfb40ff),
	.w8(32'h3b01cfd2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eaae2),
	.w1(32'hbbf5a498),
	.w2(32'h3b9d2862),
	.w3(32'h3b13a835),
	.w4(32'h3ba94be8),
	.w5(32'h3b85480c),
	.w6(32'hbb6ff75e),
	.w7(32'h3b0beda9),
	.w8(32'hbba4b123),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b0c22),
	.w1(32'hbac383e0),
	.w2(32'h3be4899a),
	.w3(32'h3bdcac22),
	.w4(32'h39f03eae),
	.w5(32'h3b5b54e3),
	.w6(32'h3bbcb8c7),
	.w7(32'h3c16f33a),
	.w8(32'hbb058189),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3de694),
	.w1(32'hbac36677),
	.w2(32'h3c0bf9ca),
	.w3(32'hbb3acdbc),
	.w4(32'hba26ba95),
	.w5(32'h3c9a586f),
	.w6(32'hba373c08),
	.w7(32'h3b2a62cf),
	.w8(32'h3c895faa),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92d400),
	.w1(32'h3c5d7ece),
	.w2(32'h3c5a99d6),
	.w3(32'hbbba7f0f),
	.w4(32'hbcda711c),
	.w5(32'h3b5e0fdd),
	.w6(32'h3d6bf01f),
	.w7(32'hbbdb3a98),
	.w8(32'hbafb9155),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3ed11),
	.w1(32'hba5afbdc),
	.w2(32'h3bcbd512),
	.w3(32'h3bade595),
	.w4(32'h3aabe34f),
	.w5(32'h3c049cf7),
	.w6(32'h39ecd270),
	.w7(32'h3be08680),
	.w8(32'h3c031234),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba90f48),
	.w1(32'hbb2c8f26),
	.w2(32'hbbff086d),
	.w3(32'hbbc76c7b),
	.w4(32'hbc454757),
	.w5(32'hbb9be90d),
	.w6(32'h3c5952a2),
	.w7(32'hb9c85d5a),
	.w8(32'h3b570c68),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b7da6),
	.w1(32'hbb212a91),
	.w2(32'hbb6ddeef),
	.w3(32'hbc4e05b8),
	.w4(32'hbc49505e),
	.w5(32'h3bbbb9ec),
	.w6(32'hbb87ddc7),
	.w7(32'hbb5a5242),
	.w8(32'h3920efca),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaac34d),
	.w1(32'hbac45df8),
	.w2(32'h3b8715e7),
	.w3(32'hb7214821),
	.w4(32'h3a8088a9),
	.w5(32'hbc27e310),
	.w6(32'hbad1edf3),
	.w7(32'h3b4a14e0),
	.w8(32'h3a5f2bad),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05d787),
	.w1(32'hbb84316b),
	.w2(32'hbbb29019),
	.w3(32'h3a8e5021),
	.w4(32'h3b1389f5),
	.w5(32'hbbabfd4e),
	.w6(32'h3a1c4dc3),
	.w7(32'h3b8e50b2),
	.w8(32'hbbbb7f26),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5089de),
	.w1(32'hbbd55acc),
	.w2(32'hb82a2e01),
	.w3(32'hbab50c4c),
	.w4(32'h3b9482b0),
	.w5(32'hbaa94366),
	.w6(32'hb9ae7e1a),
	.w7(32'h3ba1bbdd),
	.w8(32'hbc8229d4),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd02c1d),
	.w1(32'hbca17b7c),
	.w2(32'hbb68ec5d),
	.w3(32'hbc1e7b3a),
	.w4(32'h3bd8c927),
	.w5(32'h3ad70ca2),
	.w6(32'hbca40670),
	.w7(32'hbb516ce1),
	.w8(32'hba2d0a62),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb988e),
	.w1(32'hbb80f202),
	.w2(32'hbbc048ca),
	.w3(32'h39b23509),
	.w4(32'hb8b3cdfe),
	.w5(32'hbb09a3a5),
	.w6(32'h3932fc60),
	.w7(32'hbb2806e6),
	.w8(32'hba6eb01a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17862b),
	.w1(32'h39ff38ff),
	.w2(32'hba9292d2),
	.w3(32'hbb8eb050),
	.w4(32'hbb60c739),
	.w5(32'hbbd82c90),
	.w6(32'hba643087),
	.w7(32'h3a82fecb),
	.w8(32'hbb696b18),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc101695),
	.w1(32'hbc08ead6),
	.w2(32'hbc5f67e1),
	.w3(32'hb9f57654),
	.w4(32'h3b492dd5),
	.w5(32'h3b25725c),
	.w6(32'hbbe70db8),
	.w7(32'hbb2390ef),
	.w8(32'h3ab1c2eb),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad442cd),
	.w1(32'h3ac5a02b),
	.w2(32'h3a5df065),
	.w3(32'hbb15d0e8),
	.w4(32'hbabc6b07),
	.w5(32'h3b2d23e3),
	.w6(32'hba7ee57f),
	.w7(32'hb893d6c7),
	.w8(32'h3a589b97),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d97a2),
	.w1(32'hbb2e7d0e),
	.w2(32'hbb30e64f),
	.w3(32'hbb311c5e),
	.w4(32'hba36478b),
	.w5(32'hbbbb1f61),
	.w6(32'h3856a671),
	.w7(32'hba662e29),
	.w8(32'hbb49ba39),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8263e6),
	.w1(32'hbbe5e00e),
	.w2(32'hbc031bf6),
	.w3(32'hbb072a10),
	.w4(32'h3b787a1f),
	.w5(32'hbb89fce4),
	.w6(32'hbb9a7e05),
	.w7(32'hbb42b5b8),
	.w8(32'h3be0ff0c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba39cc0),
	.w1(32'hbabe7c3d),
	.w2(32'hbbb44e53),
	.w3(32'hbbfd0fde),
	.w4(32'hbb15864b),
	.w5(32'h3c113c8f),
	.w6(32'hbc5a4e27),
	.w7(32'hb97c034f),
	.w8(32'h3c121f8f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0e3d0),
	.w1(32'h3b9bf9ee),
	.w2(32'hbb865384),
	.w3(32'hbb914987),
	.w4(32'hbc108976),
	.w5(32'h3b15a5b2),
	.w6(32'h3a9910fd),
	.w7(32'hbba55b4c),
	.w8(32'h3b3e1e93),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc727c27),
	.w1(32'h3bdc27fe),
	.w2(32'hb965d0e2),
	.w3(32'hbc7af9af),
	.w4(32'hbcaa4e84),
	.w5(32'hbb2ea762),
	.w6(32'h3cbdff27),
	.w7(32'hbc757930),
	.w8(32'hbb733f6b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad0a59),
	.w1(32'hbb9fa917),
	.w2(32'hbb493cde),
	.w3(32'hbb18c6b9),
	.w4(32'hba049238),
	.w5(32'h3bc21d69),
	.w6(32'hba869522),
	.w7(32'hba4111cb),
	.w8(32'hbae2a927),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b66a9),
	.w1(32'hbb654070),
	.w2(32'h3b648d02),
	.w3(32'h3bcd5b67),
	.w4(32'h3c110ec3),
	.w5(32'h3b1ba5b9),
	.w6(32'h3b0d538b),
	.w7(32'h3c03340c),
	.w8(32'hba8148e0),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0448bd),
	.w1(32'hbbe5d434),
	.w2(32'hbbbd6acc),
	.w3(32'hb99da052),
	.w4(32'hb9f682aa),
	.w5(32'h3af0a380),
	.w6(32'hbb87f3ba),
	.w7(32'hbb76bd91),
	.w8(32'h3aba9f95),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cccee),
	.w1(32'hbad2ca5a),
	.w2(32'hba862376),
	.w3(32'hbb5006da),
	.w4(32'h399d5a1f),
	.w5(32'hba79e854),
	.w6(32'hbaac1879),
	.w7(32'h3b33bca7),
	.w8(32'h3ab4964e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f8f19),
	.w1(32'hbb415393),
	.w2(32'h3b9ab154),
	.w3(32'hbb883f02),
	.w4(32'h3b2b325b),
	.w5(32'h3c7cdfb4),
	.w6(32'hbb962aba),
	.w7(32'hbad35789),
	.w8(32'h3b2cc7c6),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62c4e2),
	.w1(32'h3c561223),
	.w2(32'h3c1affe1),
	.w3(32'hba213a23),
	.w4(32'hbc97f83a),
	.w5(32'hbb55b64c),
	.w6(32'h3d33f2fe),
	.w7(32'hbb1f69c3),
	.w8(32'hbb5bd4eb),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea6fce),
	.w1(32'hba80c6b1),
	.w2(32'h3b96cec4),
	.w3(32'h3bba0e8b),
	.w4(32'h3bc5a24c),
	.w5(32'h3aff2ffb),
	.w6(32'h3bbafc38),
	.w7(32'h3b14e6a5),
	.w8(32'h3b3580b5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89a2b8),
	.w1(32'h3a2c9651),
	.w2(32'h3a8eaa73),
	.w3(32'hbb363170),
	.w4(32'hbac29341),
	.w5(32'hbb971db8),
	.w6(32'hbb17b041),
	.w7(32'h3a9f3d1f),
	.w8(32'h3c052eb5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99fa91),
	.w1(32'hbbc92a0c),
	.w2(32'h3a01e21d),
	.w3(32'hbc5ac81a),
	.w4(32'hbbc5deaa),
	.w5(32'hbbc61599),
	.w6(32'hbc5c4da6),
	.w7(32'hbb81165c),
	.w8(32'h3aa7f7a6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dad69),
	.w1(32'hbb1b546a),
	.w2(32'hbb093789),
	.w3(32'hbb666b5c),
	.w4(32'hba31a420),
	.w5(32'hbc444a96),
	.w6(32'hbb39f3fc),
	.w7(32'h3a16913f),
	.w8(32'hbb1bd7dd),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b364e99),
	.w1(32'hbb1d8158),
	.w2(32'hbc0f8e62),
	.w3(32'hbbe4c793),
	.w4(32'hbaa1eb1a),
	.w5(32'hbb0817ce),
	.w6(32'hbc1863e3),
	.w7(32'hbc08294b),
	.w8(32'h39b6beb6),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaeeb4),
	.w1(32'hbc208883),
	.w2(32'hbb5b6cca),
	.w3(32'hb9a0ac72),
	.w4(32'hba0e8325),
	.w5(32'hbb0f94e2),
	.w6(32'hba1cc66a),
	.w7(32'hb9dbaa46),
	.w8(32'h38f3f7b8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cff42),
	.w1(32'hba525a23),
	.w2(32'h39aa71e2),
	.w3(32'h39beb11a),
	.w4(32'h3ba35807),
	.w5(32'h3c49f6c5),
	.w6(32'hbb662fdd),
	.w7(32'h3b9cd9cb),
	.w8(32'h3be95f00),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbfda8),
	.w1(32'h3c06d32c),
	.w2(32'h3baf4ff7),
	.w3(32'hba6027ae),
	.w4(32'hbb7a5ab4),
	.w5(32'hbad22f9a),
	.w6(32'h3a52ce12),
	.w7(32'hbab5475d),
	.w8(32'hbc46b116),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc8b2c6),
	.w1(32'hbc8ade2a),
	.w2(32'hbb232bbf),
	.w3(32'hbc12ed09),
	.w4(32'hbc190132),
	.w5(32'h3bb9ff29),
	.w6(32'h3ca2ab18),
	.w7(32'h3aa5f349),
	.w8(32'hbb6f5e24),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9101e7),
	.w1(32'h3b1c6907),
	.w2(32'h3bc421c6),
	.w3(32'h3b154aef),
	.w4(32'h3bab8836),
	.w5(32'h3b4f5c91),
	.w6(32'h3c0defdc),
	.w7(32'h3bbaa0ee),
	.w8(32'hbaccba95),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7949ba2),
	.w1(32'h3b80dc70),
	.w2(32'h3ba1ad58),
	.w3(32'hbc20679e),
	.w4(32'h3b0137b1),
	.w5(32'hbbba5f00),
	.w6(32'h3bc55670),
	.w7(32'h3b66f3db),
	.w8(32'h3b1e58ed),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57afcc),
	.w1(32'hbab55d43),
	.w2(32'hb9616bc8),
	.w3(32'hbbae7ab8),
	.w4(32'hbc033744),
	.w5(32'hba215dac),
	.w6(32'h3b5149c5),
	.w7(32'hbb22f3bc),
	.w8(32'h3b897f4a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42a9cf),
	.w1(32'hbb5bd215),
	.w2(32'hba96ffae),
	.w3(32'hbb8de0e5),
	.w4(32'hbb95877a),
	.w5(32'h3b85efc7),
	.w6(32'hbb438949),
	.w7(32'h3a602219),
	.w8(32'h3b6455bf),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a0e5b),
	.w1(32'h3b26e139),
	.w2(32'h3a6decb5),
	.w3(32'h3b5e5675),
	.w4(32'hbbbb8c6e),
	.w5(32'hbc0a6941),
	.w6(32'h3bf76f2a),
	.w7(32'hb968129b),
	.w8(32'h3b4fe2e2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d42cb),
	.w1(32'h3af1c679),
	.w2(32'hbbb6495b),
	.w3(32'hbbe69bf3),
	.w4(32'h3c054e6d),
	.w5(32'hbb938226),
	.w6(32'h3a482e4c),
	.w7(32'hbb9276ed),
	.w8(32'hbb09dcc0),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01487b),
	.w1(32'hbb137b5e),
	.w2(32'hba872d4d),
	.w3(32'h3a213c39),
	.w4(32'hba7838ba),
	.w5(32'hbb054f80),
	.w6(32'hbb32969e),
	.w7(32'hbb1a3bff),
	.w8(32'h39321fe5),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c278bd1),
	.w1(32'hbba1eeff),
	.w2(32'hba96b91e),
	.w3(32'hb95a2a78),
	.w4(32'h3b707733),
	.w5(32'h380ae1cc),
	.w6(32'h3b8dc0e2),
	.w7(32'h3b89e71b),
	.w8(32'h3b1d70c7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e1a3b),
	.w1(32'h3a05df7c),
	.w2(32'hbc13a3f8),
	.w3(32'h3b0b1e7c),
	.w4(32'hba7f395d),
	.w5(32'hb919fc86),
	.w6(32'h3b3a63d6),
	.w7(32'hbb278310),
	.w8(32'hbc0309aa),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac39c67),
	.w1(32'hbb8e15f7),
	.w2(32'hba5db61c),
	.w3(32'h3a1d530f),
	.w4(32'h3ad183c7),
	.w5(32'h39b150ff),
	.w6(32'hbbabbcd1),
	.w7(32'hbba82fe1),
	.w8(32'h3b76a8f1),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aa83f),
	.w1(32'h3aa2fd98),
	.w2(32'hbb023b00),
	.w3(32'hbb683ebc),
	.w4(32'hbbf53099),
	.w5(32'hbacbce5e),
	.w6(32'hbb4dce76),
	.w7(32'hbb52e0c9),
	.w8(32'hb862fe0c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d8039),
	.w1(32'h3b3a2a92),
	.w2(32'hbaa734ba),
	.w3(32'hbc3b91f3),
	.w4(32'hb9c8213f),
	.w5(32'hbb8b3726),
	.w6(32'hbc1aa70c),
	.w7(32'hbae37494),
	.w8(32'hbb44078d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa18141),
	.w1(32'hbbb44c52),
	.w2(32'hbb507fcc),
	.w3(32'h3bbbc36f),
	.w4(32'h3ac5797a),
	.w5(32'hba345357),
	.w6(32'hba85a7d0),
	.w7(32'h3b4eab2a),
	.w8(32'h3b207adc),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7f4f5),
	.w1(32'h39b5e115),
	.w2(32'hb9026d73),
	.w3(32'hbaf13b7c),
	.w4(32'hb87000c3),
	.w5(32'hbbf6b8ec),
	.w6(32'h39f764a6),
	.w7(32'hba5f1466),
	.w8(32'hbc7b09f4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5521d5),
	.w1(32'hbc06fb7e),
	.w2(32'h3b9a6686),
	.w3(32'hbac75778),
	.w4(32'h3b9f2fe9),
	.w5(32'hbb8f4af8),
	.w6(32'hbbbb4960),
	.w7(32'h3c26a287),
	.w8(32'hbb39cdcb),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcaf34),
	.w1(32'hbbb92481),
	.w2(32'hb831308e),
	.w3(32'h3af3a7be),
	.w4(32'h3ad58937),
	.w5(32'h3b4b0834),
	.w6(32'hbc1d6c85),
	.w7(32'h3b868b06),
	.w8(32'h3b9a4eab),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb901553),
	.w1(32'h3affcb51),
	.w2(32'h3b58c2e1),
	.w3(32'h3bbf0f91),
	.w4(32'h3b3d5b00),
	.w5(32'h3ad16e08),
	.w6(32'hb9a4caff),
	.w7(32'hb950e7f2),
	.w8(32'h3a8412ff),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7451ad),
	.w1(32'hbb00c6a5),
	.w2(32'h3b6216de),
	.w3(32'h3b92ba4d),
	.w4(32'h3b942dad),
	.w5(32'hbab10789),
	.w6(32'hbaaec4b8),
	.w7(32'h3bc57521),
	.w8(32'h3af7247c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbdabc),
	.w1(32'hbabded8a),
	.w2(32'hbaa4072a),
	.w3(32'h3ad4b948),
	.w4(32'h3b1f4d7c),
	.w5(32'h384db35b),
	.w6(32'hbb2f6215),
	.w7(32'h3b2a9256),
	.w8(32'h3bdaedf0),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6337f),
	.w1(32'h3a9a89df),
	.w2(32'hbac71538),
	.w3(32'hbbcc2837),
	.w4(32'hbb9e1669),
	.w5(32'h3b3b8f5d),
	.w6(32'hbb16672b),
	.w7(32'hbb449e4e),
	.w8(32'h3b54adcd),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96dfcce),
	.w1(32'hbb55c12e),
	.w2(32'h3ab7b509),
	.w3(32'h3b5a7c1d),
	.w4(32'h3b82aa5f),
	.w5(32'hbabd5766),
	.w6(32'hb9c7d803),
	.w7(32'h3ba0859e),
	.w8(32'hbc4fd535),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafb517),
	.w1(32'hbb36b930),
	.w2(32'h3b10de9b),
	.w3(32'h3c13386b),
	.w4(32'hbab222a6),
	.w5(32'hbaa0f804),
	.w6(32'h3b37b12f),
	.w7(32'hbb2290d3),
	.w8(32'hbb939550),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02badd),
	.w1(32'hbb400ce6),
	.w2(32'hb8f058a6),
	.w3(32'hbb411996),
	.w4(32'h3b255877),
	.w5(32'hbbfc5fca),
	.w6(32'h3b00502d),
	.w7(32'h3ba0cabf),
	.w8(32'hbc2bc101),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb22901),
	.w1(32'hbb482bf0),
	.w2(32'hbc86dbec),
	.w3(32'hbb8104c0),
	.w4(32'hbbd8acd4),
	.w5(32'hbb75dafb),
	.w6(32'hbbd1aa72),
	.w7(32'hbc83204c),
	.w8(32'h3b2c51b9),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dbb0b),
	.w1(32'h3b3e2613),
	.w2(32'hba99863e),
	.w3(32'h3c51c7e0),
	.w4(32'h3ab461a4),
	.w5(32'h3b9462e4),
	.w6(32'h3b9d70b5),
	.w7(32'h397ef3ac),
	.w8(32'h3bb67c49),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ecd17),
	.w1(32'h3b2ffaf9),
	.w2(32'h3a93ac67),
	.w3(32'hbb15e53d),
	.w4(32'hbb2ed0c2),
	.w5(32'hbb80df85),
	.w6(32'h3be5e960),
	.w7(32'h3b0beae4),
	.w8(32'hbba6e6f8),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1179f2),
	.w1(32'hbb9e8fc9),
	.w2(32'hbb8d8862),
	.w3(32'hbb289b6d),
	.w4(32'hba93162c),
	.w5(32'hbb9975e6),
	.w6(32'h3b87b3e4),
	.w7(32'hb8553a95),
	.w8(32'h3b3472de),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ff9c2),
	.w1(32'hb9b23a25),
	.w2(32'hbabc06af),
	.w3(32'hbbe27906),
	.w4(32'hb9e4ba1a),
	.w5(32'h3bc0c742),
	.w6(32'h3a960722),
	.w7(32'hbb69cf48),
	.w8(32'hba62de72),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6f485),
	.w1(32'hbabfd383),
	.w2(32'hbc2580a2),
	.w3(32'hbc349237),
	.w4(32'hbb96470b),
	.w5(32'hbb814ee0),
	.w6(32'h3a167cc5),
	.w7(32'hbbc94f2a),
	.w8(32'h38f4ed2f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed1d29),
	.w1(32'hbbb1f21d),
	.w2(32'hbb31b7ac),
	.w3(32'h3a7cc634),
	.w4(32'h3a40bd80),
	.w5(32'h3b54f294),
	.w6(32'h3a1ad3ea),
	.w7(32'h3ad894b2),
	.w8(32'h3c0a71b4),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4f152),
	.w1(32'hbc5b861e),
	.w2(32'hbb14006a),
	.w3(32'hbb887709),
	.w4(32'hbb166677),
	.w5(32'hbc78e91c),
	.w6(32'hbbb4ec00),
	.w7(32'h3a696fdc),
	.w8(32'hbc4c15e6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8926d),
	.w1(32'hbbbd5ae6),
	.w2(32'hbaeea095),
	.w3(32'hbb6d25da),
	.w4(32'h3b8c7fb4),
	.w5(32'h3aac2b12),
	.w6(32'hbb937053),
	.w7(32'h3ac0445e),
	.w8(32'h3a27a0f5),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6186e),
	.w1(32'hbbf9b591),
	.w2(32'hba2f51f1),
	.w3(32'h3bd28a34),
	.w4(32'h3b4e8f9f),
	.w5(32'hbc06291b),
	.w6(32'h39e6db84),
	.w7(32'h3bd3c959),
	.w8(32'h3af9adcf),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8faf6f),
	.w1(32'hbb329b74),
	.w2(32'hbb9e8bce),
	.w3(32'hbab6b729),
	.w4(32'h3c605eea),
	.w5(32'hbb4b3b89),
	.w6(32'hbc1149b5),
	.w7(32'hbc296bad),
	.w8(32'hba35da04),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c337430),
	.w1(32'h39ee4450),
	.w2(32'hbb81dad1),
	.w3(32'hbba9838e),
	.w4(32'hba6b9ff2),
	.w5(32'hb95ba5d0),
	.w6(32'h3abeed8c),
	.w7(32'hbbaa8880),
	.w8(32'h3b1f0934),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7419c3),
	.w1(32'hba89f0d7),
	.w2(32'h3a93816a),
	.w3(32'hbba1874f),
	.w4(32'h3a822775),
	.w5(32'hbb94ef29),
	.w6(32'h3bbd0dd7),
	.w7(32'hbac8f796),
	.w8(32'h39b61afc),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e6fd6),
	.w1(32'hbc34e06b),
	.w2(32'hbbe151cb),
	.w3(32'hbabdb8e5),
	.w4(32'h3a916b5b),
	.w5(32'hbc24246c),
	.w6(32'hbbf80a3c),
	.w7(32'h3b20b752),
	.w8(32'hbbbf2d3a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31c92b),
	.w1(32'hbb74faa3),
	.w2(32'hbb483506),
	.w3(32'h3a2c72b1),
	.w4(32'h3b4151eb),
	.w5(32'hbb9e7a33),
	.w6(32'hbb1c27d7),
	.w7(32'hbad45c4d),
	.w8(32'hbbab7f11),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc406894),
	.w1(32'hbbc1c658),
	.w2(32'hbb3accc4),
	.w3(32'hbb9cf4be),
	.w4(32'hba2ff1f0),
	.w5(32'hbbbe2984),
	.w6(32'hbbc110b7),
	.w7(32'h3aa81dbc),
	.w8(32'hbb1db5e6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02a3ff),
	.w1(32'hbc3f1dbc),
	.w2(32'hbc32ec07),
	.w3(32'hbc12c07e),
	.w4(32'h3af10863),
	.w5(32'hbb1ccec9),
	.w6(32'hbc2c72c5),
	.w7(32'hba93cf9e),
	.w8(32'hbb1b112c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82db45),
	.w1(32'h3b263d7b),
	.w2(32'hbafc3c9e),
	.w3(32'hba8f36bd),
	.w4(32'hbb0938a9),
	.w5(32'hbbaaa4b5),
	.w6(32'h3a0118b0),
	.w7(32'h3b837789),
	.w8(32'h3a838ead),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e76b9),
	.w1(32'h3b884ffd),
	.w2(32'hb9a811a1),
	.w3(32'h3ba5e4ba),
	.w4(32'h3ba7ee0b),
	.w5(32'h3ac191cc),
	.w6(32'hba56fd54),
	.w7(32'h3bedfa6e),
	.w8(32'hba167588),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b900e94),
	.w1(32'h3be0ebc8),
	.w2(32'hbbc5ffdb),
	.w3(32'hba355aa9),
	.w4(32'hbb7bd37b),
	.w5(32'hba4f35a0),
	.w6(32'h3ade9e30),
	.w7(32'hbba7296c),
	.w8(32'hbba55545),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfd3da),
	.w1(32'hbbe11003),
	.w2(32'hbbb0b55a),
	.w3(32'hbb212f4a),
	.w4(32'hbb61d029),
	.w5(32'h3ba399ea),
	.w6(32'h38ef9e13),
	.w7(32'h3c1b2610),
	.w8(32'h3bc6dd94),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0ec0e),
	.w1(32'h3b9b6fa9),
	.w2(32'h3ac29db8),
	.w3(32'hbbb85670),
	.w4(32'hbc02084e),
	.w5(32'hbac5fb47),
	.w6(32'h3bc1a42c),
	.w7(32'hbc331545),
	.w8(32'h3b9450bf),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf58e31),
	.w1(32'hbbf3e8ae),
	.w2(32'hbb5c0523),
	.w3(32'hbb71601b),
	.w4(32'hbb665f56),
	.w5(32'h3bc7b521),
	.w6(32'hbb1388c7),
	.w7(32'h3a84e736),
	.w8(32'h3c7d1cf9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfee7da),
	.w1(32'h3b8f4afc),
	.w2(32'hbbbf5d4e),
	.w3(32'hbbecefe3),
	.w4(32'hbc0a45e9),
	.w5(32'h3b084532),
	.w6(32'h3b8b5e39),
	.w7(32'hbc568ccd),
	.w8(32'h3ba8c2d3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba019277),
	.w1(32'hbc194dc3),
	.w2(32'hbbbdcb90),
	.w3(32'hbc1f2992),
	.w4(32'hbb06b84f),
	.w5(32'h3b22e950),
	.w6(32'hbc69868e),
	.w7(32'hbb906739),
	.w8(32'hba9b549f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b4161),
	.w1(32'hbb4c00e2),
	.w2(32'h3b1b5cd0),
	.w3(32'h3c3ae690),
	.w4(32'h3be94879),
	.w5(32'hbb3b51ee),
	.w6(32'h3c268b32),
	.w7(32'h3c32e6b7),
	.w8(32'h3c384086),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97d3c5),
	.w1(32'hba82d904),
	.w2(32'hbbca907f),
	.w3(32'hbc21aba0),
	.w4(32'hbb2eeba4),
	.w5(32'h3a219cf8),
	.w6(32'hbbc1b440),
	.w7(32'hbb757f7f),
	.w8(32'hb9ff3d77),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e4ba1e),
	.w1(32'h3aadb97c),
	.w2(32'hba6b7f2d),
	.w3(32'hbab40463),
	.w4(32'hbb133d5c),
	.w5(32'hbb8f5ca9),
	.w6(32'hbbc50e10),
	.w7(32'h3a198d0a),
	.w8(32'h3c89cf32),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2d2b3),
	.w1(32'h3c458776),
	.w2(32'hbb8e762a),
	.w3(32'hbc309f91),
	.w4(32'hbc16a358),
	.w5(32'h3b8e5d48),
	.w6(32'h3ba2c4e0),
	.w7(32'hbc182628),
	.w8(32'h3bd2dbb1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9563308),
	.w1(32'h3af97349),
	.w2(32'hbb2bdf10),
	.w3(32'hbb42de94),
	.w4(32'hbc1dcccc),
	.w5(32'h3b0b26cc),
	.w6(32'h3b867a2f),
	.w7(32'hbbc55b90),
	.w8(32'h3c86b664),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c620ba4),
	.w1(32'hba3a2236),
	.w2(32'hbb15487d),
	.w3(32'hbc1e816e),
	.w4(32'hbb17b658),
	.w5(32'hbb310aa1),
	.w6(32'hbb851765),
	.w7(32'hbb242f14),
	.w8(32'hbad7aad0),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba98792),
	.w1(32'hbb6da3c0),
	.w2(32'hbb832b92),
	.w3(32'hbbd5e21a),
	.w4(32'h3c34dafa),
	.w5(32'hbb4372b3),
	.w6(32'hbc015d7e),
	.w7(32'h3c129f1a),
	.w8(32'h3c9809d3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b0d56),
	.w1(32'hbbbeb444),
	.w2(32'hbb0eb87d),
	.w3(32'hbca4f695),
	.w4(32'hbc09eb14),
	.w5(32'hbb77694c),
	.w6(32'hbc3de71b),
	.w7(32'hbbde236a),
	.w8(32'h3a546602),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5a660),
	.w1(32'hbb26591e),
	.w2(32'hb96b6b0d),
	.w3(32'hbb22dc29),
	.w4(32'h3b77b0c1),
	.w5(32'hbbc58162),
	.w6(32'hbb859906),
	.w7(32'hba8fe8ad),
	.w8(32'hba36a129),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba253a90),
	.w1(32'hbb5d93d9),
	.w2(32'h3b625042),
	.w3(32'h3ba7a6fe),
	.w4(32'h3b96f005),
	.w5(32'h3bf9271f),
	.w6(32'hba7a1087),
	.w7(32'h3b3f7e79),
	.w8(32'hbba581c3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78cd5c),
	.w1(32'hbbe65ac9),
	.w2(32'h3c19de18),
	.w3(32'hbad4b2c2),
	.w4(32'hbc39d653),
	.w5(32'h3b64da19),
	.w6(32'h3c974378),
	.w7(32'h3b6f199e),
	.w8(32'h3ac0b9fd),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0ce38),
	.w1(32'hbb1d1cc5),
	.w2(32'hbad9c769),
	.w3(32'h3b04dda0),
	.w4(32'h3ac611e1),
	.w5(32'h3a756a8d),
	.w6(32'h3a46cb44),
	.w7(32'h3a209c82),
	.w8(32'hbbc01c22),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebb481),
	.w1(32'hbbb4c875),
	.w2(32'h3abc5bbc),
	.w3(32'h3bcc5193),
	.w4(32'h3b5b62a8),
	.w5(32'hbc3e4c07),
	.w6(32'h3bb2e934),
	.w7(32'h3c3aba57),
	.w8(32'hba91a4d2),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f5cb8),
	.w1(32'hbba61487),
	.w2(32'hbb987f1e),
	.w3(32'hbbe5b3b5),
	.w4(32'hbc318bd4),
	.w5(32'hbc75be31),
	.w6(32'h3ae5b987),
	.w7(32'hbb2afa88),
	.w8(32'hbc52d049),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc292b4a),
	.w1(32'hbc9c05d8),
	.w2(32'hbbbcc32c),
	.w3(32'hbbe05e28),
	.w4(32'h3b82e682),
	.w5(32'h3ad02e8f),
	.w6(32'hbc1496f8),
	.w7(32'h3bbcca14),
	.w8(32'hbb290012),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3081ae),
	.w1(32'hbc3d37e9),
	.w2(32'hbad269e7),
	.w3(32'hbbac07a4),
	.w4(32'h3bb211b4),
	.w5(32'h3b214669),
	.w6(32'hbb3cbef7),
	.w7(32'h3b140556),
	.w8(32'h3b77855b),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7783d),
	.w1(32'hbb6e8d89),
	.w2(32'hbafa264f),
	.w3(32'hbbbf7e52),
	.w4(32'hba392769),
	.w5(32'hba8797e0),
	.w6(32'hbbec12c8),
	.w7(32'h3aeb8b34),
	.w8(32'hbb3735d2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ee473),
	.w1(32'h39edcc31),
	.w2(32'hbb143e1e),
	.w3(32'h3a22fb42),
	.w4(32'h3aa6f04b),
	.w5(32'hbbd83475),
	.w6(32'h3aa24dae),
	.w7(32'h3aa37cad),
	.w8(32'hbaba0c25),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b2def),
	.w1(32'hbac73945),
	.w2(32'hbb5cf676),
	.w3(32'hba704585),
	.w4(32'h3b8b579f),
	.w5(32'h3a345842),
	.w6(32'hbb1d0f8d),
	.w7(32'h39cf7c62),
	.w8(32'h3c2c118c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ed812),
	.w1(32'hbb18f272),
	.w2(32'h3a12d0ed),
	.w3(32'hbbe4dbc6),
	.w4(32'hbbaeceb7),
	.w5(32'h3b5cbdb9),
	.w6(32'hba115814),
	.w7(32'hbc18f6d1),
	.w8(32'hba7f66db),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b81e8),
	.w1(32'hbb5368ba),
	.w2(32'hbb897d98),
	.w3(32'hbbf020e6),
	.w4(32'hbb5979a8),
	.w5(32'h3b660778),
	.w6(32'hba9c00a3),
	.w7(32'hbbc76e9f),
	.w8(32'h3bc769c9),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba6bdc),
	.w1(32'h3a5c740a),
	.w2(32'h3b22fa27),
	.w3(32'h3b68fe1d),
	.w4(32'h3a9115aa),
	.w5(32'h3a3800d1),
	.w6(32'h3b99d94f),
	.w7(32'h3b99e37c),
	.w8(32'hbb067ed5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d834f),
	.w1(32'hbaf25f76),
	.w2(32'hbb1c0340),
	.w3(32'hbb2c76ef),
	.w4(32'hbb5de13a),
	.w5(32'h3b82021c),
	.w6(32'hb86e3076),
	.w7(32'hbb8fae74),
	.w8(32'h3befce54),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f80e4),
	.w1(32'h3afbc38e),
	.w2(32'h3b4ca718),
	.w3(32'h3b0aa052),
	.w4(32'h3b664b27),
	.w5(32'hbb959ce1),
	.w6(32'h3af2d773),
	.w7(32'h3bebf326),
	.w8(32'hbaee3a3a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4148ae),
	.w1(32'hbb98c49c),
	.w2(32'hbb051512),
	.w3(32'hbba4fede),
	.w4(32'hbb30b91b),
	.w5(32'h39de5ba9),
	.w6(32'hbb0d5859),
	.w7(32'hbb05c07e),
	.w8(32'hba946f6e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e3478),
	.w1(32'hbb916f67),
	.w2(32'hbb75691d),
	.w3(32'hbb9a5845),
	.w4(32'hbb86a915),
	.w5(32'hb996c8db),
	.w6(32'hb97fa515),
	.w7(32'h3aa0f46d),
	.w8(32'h3b58a192),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06c0d2),
	.w1(32'h3aa8356d),
	.w2(32'h3b91a959),
	.w3(32'hba8964e0),
	.w4(32'h3a48d4cd),
	.w5(32'hbb238343),
	.w6(32'h3adec3b9),
	.w7(32'h3b83237f),
	.w8(32'h3bb6062f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba453a4),
	.w1(32'h3b15cf35),
	.w2(32'hb7cb0078),
	.w3(32'h3aedd280),
	.w4(32'hbb0786f7),
	.w5(32'hbb73d742),
	.w6(32'h3c20fc91),
	.w7(32'h3b0ff210),
	.w8(32'hbb6eef02),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70ba02),
	.w1(32'hbb7ecac3),
	.w2(32'hbb8bfee1),
	.w3(32'hbaf3633d),
	.w4(32'hbb323602),
	.w5(32'h3a97655d),
	.w6(32'hba10eb12),
	.w7(32'hba7cfa18),
	.w8(32'h3b1a1e6d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5249df),
	.w1(32'hbace882a),
	.w2(32'hbb87494b),
	.w3(32'hbab2af7b),
	.w4(32'hbb4cf31b),
	.w5(32'h3981ed5d),
	.w6(32'hbac832e7),
	.w7(32'h37d39234),
	.w8(32'hba622d6f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d442b0),
	.w1(32'h3960584c),
	.w2(32'hb91394aa),
	.w3(32'hba634ca1),
	.w4(32'h39d1d19a),
	.w5(32'hbb2bc751),
	.w6(32'hba05b8dc),
	.w7(32'hba318e6f),
	.w8(32'h3aeb3271),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76965b),
	.w1(32'hbb63c889),
	.w2(32'hba405aa9),
	.w3(32'hbb5710e4),
	.w4(32'hbb850838),
	.w5(32'hba2ba207),
	.w6(32'hbb1b3f12),
	.w7(32'h385390a4),
	.w8(32'hbab6bf91),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac78c29),
	.w1(32'hbb2cb3e9),
	.w2(32'hbb321dee),
	.w3(32'hbaf48b3a),
	.w4(32'hbab7a82d),
	.w5(32'h3bc4b262),
	.w6(32'hbae5d4a4),
	.w7(32'hbae4aff2),
	.w8(32'h3ad9fc84),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb821c86),
	.w1(32'hbaab1d20),
	.w2(32'hbb3a1c7d),
	.w3(32'hbab43638),
	.w4(32'hba8bce57),
	.w5(32'h3a93d5d3),
	.w6(32'h3925fef3),
	.w7(32'hb8ccd864),
	.w8(32'hba157952),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41f476),
	.w1(32'h3a8d2fcb),
	.w2(32'hbb0e0524),
	.w3(32'hbb93d2a0),
	.w4(32'hbb84a08c),
	.w5(32'hbb23321e),
	.w6(32'hbb890ca3),
	.w7(32'hbb3bd6e3),
	.w8(32'hbaf4cde4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e71b2),
	.w1(32'hbba471e4),
	.w2(32'hbb657b42),
	.w3(32'hbb7ce74a),
	.w4(32'hb9c903d5),
	.w5(32'h3a9ea5f4),
	.w6(32'hbb1a25be),
	.w7(32'h392d49e7),
	.w8(32'h3a86bce5),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac06b8),
	.w1(32'h3abf34a9),
	.w2(32'h3b06c079),
	.w3(32'hbb0f9e5a),
	.w4(32'hbb14e9c2),
	.w5(32'hb958042d),
	.w6(32'hbb55a726),
	.w7(32'h3a38a215),
	.w8(32'h3b3d2e60),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb637c1d),
	.w1(32'h3bb05ad4),
	.w2(32'h3b105211),
	.w3(32'h3b06b170),
	.w4(32'h3b41f5ed),
	.w5(32'hb9e5b155),
	.w6(32'h3b7ce8d8),
	.w7(32'h392f2ffd),
	.w8(32'hbae5669b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9e4be),
	.w1(32'hbb08fb9f),
	.w2(32'hbb6ce970),
	.w3(32'hb9fece1d),
	.w4(32'hbae55639),
	.w5(32'h3b7217b2),
	.w6(32'h3947f97d),
	.w7(32'hbaea2026),
	.w8(32'h3b662295),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d990e),
	.w1(32'h3b9ae634),
	.w2(32'h3bac5838),
	.w3(32'h3b7c12de),
	.w4(32'h3b9a822e),
	.w5(32'hbb64f999),
	.w6(32'h3b8780c8),
	.w7(32'h3ba3aaa0),
	.w8(32'h3afbb082),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2556a),
	.w1(32'h3913ee9d),
	.w2(32'h3ba0b5fe),
	.w3(32'h3afaea10),
	.w4(32'hbaa3509f),
	.w5(32'h3ac97b25),
	.w6(32'h3c0e22d8),
	.w7(32'h3aadfc79),
	.w8(32'h3ba828e2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17d03d),
	.w1(32'hbb7f5e19),
	.w2(32'hba8fc0b4),
	.w3(32'hbb3fb6b4),
	.w4(32'hbb5e5956),
	.w5(32'h3bff3db7),
	.w6(32'h3a25b2fb),
	.w7(32'h3a2f600e),
	.w8(32'h3c508c84),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4f715),
	.w1(32'h3b3ed9b8),
	.w2(32'h3bac6758),
	.w3(32'h3bb4188a),
	.w4(32'h3b2c9a65),
	.w5(32'hbb19794b),
	.w6(32'h3b6c2269),
	.w7(32'h3c0a8160),
	.w8(32'hbb5975e1),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebbaa7),
	.w1(32'h39ad8938),
	.w2(32'hbb01d550),
	.w3(32'h3b91cd9e),
	.w4(32'hb8e28bc8),
	.w5(32'h3a121978),
	.w6(32'h3ba2538e),
	.w7(32'h3a55b2f0),
	.w8(32'hba110b1f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb249f19),
	.w1(32'hba9d558c),
	.w2(32'hbae62b51),
	.w3(32'h3a1b5b19),
	.w4(32'hba8cddce),
	.w5(32'hbb17e69d),
	.w6(32'hba85ba9c),
	.w7(32'hbb004875),
	.w8(32'h3a7f12d3),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a506524),
	.w1(32'hbab93594),
	.w2(32'hb9eb53e9),
	.w3(32'hba67dc1d),
	.w4(32'hb7ae6605),
	.w5(32'hba725daf),
	.w6(32'h39325875),
	.w7(32'h3aaf3b60),
	.w8(32'hbaeec433),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddb308),
	.w1(32'hbb08a246),
	.w2(32'hbada68cf),
	.w3(32'hb9f90ccb),
	.w4(32'hba9a9c5b),
	.w5(32'hbb2801ed),
	.w6(32'hba77be05),
	.w7(32'hba9a5a7d),
	.w8(32'hb7b12c74),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ee11a),
	.w1(32'hbac80518),
	.w2(32'hbaad5578),
	.w3(32'hba3b80c3),
	.w4(32'h395ea1d0),
	.w5(32'hba9b3c9a),
	.w6(32'hbac9aa6e),
	.w7(32'hba982db2),
	.w8(32'hba8101f7),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb727ec2),
	.w1(32'hba81da75),
	.w2(32'hbb163834),
	.w3(32'hbb963e18),
	.w4(32'hbb78bc49),
	.w5(32'hbb24fee7),
	.w6(32'hba9e2b69),
	.w7(32'hbaccc348),
	.w8(32'h3b5a6c6b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b006e2c),
	.w1(32'hb9672f95),
	.w2(32'hbacd3ad2),
	.w3(32'hbb059629),
	.w4(32'hb96cac47),
	.w5(32'h39f88022),
	.w6(32'h37d82398),
	.w7(32'hb91ebc54),
	.w8(32'hba1fbf93),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc77286),
	.w1(32'hbaae5af0),
	.w2(32'hbb091afd),
	.w3(32'hbaf16c80),
	.w4(32'h3b3e63a4),
	.w5(32'hbaafdcdc),
	.w6(32'hba970e77),
	.w7(32'h3b8ee08f),
	.w8(32'hbb0e5741),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule