module layer_8_featuremap_137(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4137ff),
	.w1(32'hbc286356),
	.w2(32'h3b450963),
	.w3(32'hbbba9a2a),
	.w4(32'hbbe76111),
	.w5(32'hbb854595),
	.w6(32'h3afdfe15),
	.w7(32'h3c39f5dd),
	.w8(32'h3c580ee5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb357ffa),
	.w1(32'hbc2f22d9),
	.w2(32'h3c124ff2),
	.w3(32'hbcee0a15),
	.w4(32'hbc13b4a3),
	.w5(32'hbc57b7ae),
	.w6(32'hbc9c6f09),
	.w7(32'hbc094bfa),
	.w8(32'h3b9cfa14),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7e0e6),
	.w1(32'h3bdcdcf0),
	.w2(32'h3c884110),
	.w3(32'h3bd4af3e),
	.w4(32'h3c12a0db),
	.w5(32'hbb2d3cd4),
	.w6(32'h3bc443e9),
	.w7(32'hbc2e21b5),
	.w8(32'hba3aba3b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f8545),
	.w1(32'hbc8df8d3),
	.w2(32'hbc2dfd3a),
	.w3(32'hbbe7bd57),
	.w4(32'h3c882f9e),
	.w5(32'h3c3855d9),
	.w6(32'hbbe4d33b),
	.w7(32'h3cee5503),
	.w8(32'h3ba74da5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc473836),
	.w1(32'h3bd7a695),
	.w2(32'hbc42a7c5),
	.w3(32'hbca42586),
	.w4(32'h3b7926df),
	.w5(32'h3b2149d5),
	.w6(32'hbc820e11),
	.w7(32'h3c96c296),
	.w8(32'h3b6f40a8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2aaca3),
	.w1(32'hbc332d4e),
	.w2(32'h3c0a4e77),
	.w3(32'h38f2dcf7),
	.w4(32'h3b9d7ddf),
	.w5(32'hbcf8b6d2),
	.w6(32'hbc0eb2f5),
	.w7(32'hbabd1d6d),
	.w8(32'hbcfff370),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb367174),
	.w1(32'hbbd7d8eb),
	.w2(32'hbc635ea2),
	.w3(32'hbc979a05),
	.w4(32'hbc4d04d1),
	.w5(32'hbc192d0a),
	.w6(32'hbc51e6f7),
	.w7(32'hbc8c6a88),
	.w8(32'hbc3a8062),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa4039),
	.w1(32'hbb10dad1),
	.w2(32'hbc60467b),
	.w3(32'hbcacc741),
	.w4(32'h3bcb1624),
	.w5(32'hbc88c5bc),
	.w6(32'hbb3280bc),
	.w7(32'hbc53015e),
	.w8(32'hb97a9063),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a66f9),
	.w1(32'h3c2f4628),
	.w2(32'hbb2e9971),
	.w3(32'hbc67b5fc),
	.w4(32'hb9481f0e),
	.w5(32'hbbf9f65c),
	.w6(32'h39b7476f),
	.w7(32'hbb946b66),
	.w8(32'hbca89d45),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ee5ac),
	.w1(32'hbbf034f3),
	.w2(32'h3bfd411e),
	.w3(32'hbd12b30f),
	.w4(32'h3b21c40a),
	.w5(32'hbb4727cd),
	.w6(32'hbcf9d8fb),
	.w7(32'h3b1a95f1),
	.w8(32'hbc1fa7cf),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c645406),
	.w1(32'hbbf0e30c),
	.w2(32'h3b994ef4),
	.w3(32'hbb96de19),
	.w4(32'h3c5162b1),
	.w5(32'h3d1cd874),
	.w6(32'hbc939bf3),
	.w7(32'hbc852729),
	.w8(32'hbb713eec),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced20f8),
	.w1(32'hbcc25c6b),
	.w2(32'hbc85c116),
	.w3(32'hba75733c),
	.w4(32'h3b2f8560),
	.w5(32'hbc6a3fd7),
	.w6(32'hbc358fbb),
	.w7(32'hbc143a46),
	.w8(32'hbc19545a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc40d53),
	.w1(32'hbbcd1a43),
	.w2(32'h3b60d3d0),
	.w3(32'hbc0a0c0b),
	.w4(32'h3b168ae9),
	.w5(32'hba983f87),
	.w6(32'hbb9ba411),
	.w7(32'h3ad7e8ed),
	.w8(32'h3b249f3d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c282029),
	.w1(32'h3b6ba19b),
	.w2(32'h3b802116),
	.w3(32'hb98a3889),
	.w4(32'h3aafa2a7),
	.w5(32'hba5712e1),
	.w6(32'h3a4537a1),
	.w7(32'h3b59a8a7),
	.w8(32'h398255e0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b044ca1),
	.w1(32'h3b79d766),
	.w2(32'h3acac0e4),
	.w3(32'h3a1bba4c),
	.w4(32'h3a8b7a1b),
	.w5(32'hbb1f2017),
	.w6(32'h3ad74813),
	.w7(32'h3af2d0d4),
	.w8(32'hba888642),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c7eae),
	.w1(32'h3b15df23),
	.w2(32'hbaf9880f),
	.w3(32'hba7f017e),
	.w4(32'hbb9caf4b),
	.w5(32'hbbe15834),
	.w6(32'hb69eb7cf),
	.w7(32'hbb897123),
	.w8(32'hbc18f3f2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe685f),
	.w1(32'h3a633661),
	.w2(32'h3acea5eb),
	.w3(32'hbc160533),
	.w4(32'hbb4b34cd),
	.w5(32'hbc4e0f35),
	.w6(32'hbc192a34),
	.w7(32'h37be3851),
	.w8(32'hbb5d57b3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e6bde),
	.w1(32'hb8e90353),
	.w2(32'hbbacf63a),
	.w3(32'hbc319040),
	.w4(32'hbc26ee3a),
	.w5(32'hbbb8d57a),
	.w6(32'hba4bc424),
	.w7(32'hbb894d43),
	.w8(32'hbbb3af37),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce47ead),
	.w1(32'hbd18f2d7),
	.w2(32'h3bcf5f0f),
	.w3(32'hbd1f4cbb),
	.w4(32'hbc6fab70),
	.w5(32'h3d05b782),
	.w6(32'hbc930f2a),
	.w7(32'h3c42bab6),
	.w8(32'h3d2cbb73),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ebcbc),
	.w1(32'hbc903a34),
	.w2(32'hbbbd331b),
	.w3(32'h3b53058c),
	.w4(32'h3b739324),
	.w5(32'h3c03e366),
	.w6(32'h394f4c50),
	.w7(32'h3b66cb2b),
	.w8(32'h3b5d8a79),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4376f),
	.w1(32'h3b413b6a),
	.w2(32'hbc34b7dc),
	.w3(32'h3bc127fb),
	.w4(32'hbc753446),
	.w5(32'hbb40c598),
	.w6(32'h3c54571a),
	.w7(32'hbc8ec12e),
	.w8(32'hbc18b176),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63e8aa),
	.w1(32'hbbd614b4),
	.w2(32'hbba1bcc8),
	.w3(32'h3b4011b2),
	.w4(32'hbb9c4096),
	.w5(32'hbc942add),
	.w6(32'hbb94fbef),
	.w7(32'hbc33ac90),
	.w8(32'hbc945631),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43ee5e),
	.w1(32'hbbbf2c00),
	.w2(32'h3b59fa29),
	.w3(32'hbc8e7f7c),
	.w4(32'h3b5d1061),
	.w5(32'h3d096695),
	.w6(32'hbacc9cb1),
	.w7(32'h3ca9a11e),
	.w8(32'h3d295793),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b296cb1),
	.w1(32'h39de066b),
	.w2(32'hb9998c4c),
	.w3(32'h3bcf6fad),
	.w4(32'h3c778ca7),
	.w5(32'hbb20807c),
	.w6(32'h3bc9f9d9),
	.w7(32'h3b523597),
	.w8(32'hbbdb004c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0571de),
	.w1(32'h3beb508e),
	.w2(32'h3a7bfe09),
	.w3(32'hbb5638b2),
	.w4(32'h3b2feab1),
	.w5(32'hbb13479d),
	.w6(32'h3a71a7a4),
	.w7(32'hba1c609a),
	.w8(32'hbc1b6dcd),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ae317),
	.w1(32'hbc1bca58),
	.w2(32'hbbcb4a04),
	.w3(32'hbbc56e42),
	.w4(32'hbaafed3f),
	.w5(32'h3bd270c9),
	.w6(32'hb92c854f),
	.w7(32'h3b35e96b),
	.w8(32'h3be83d3c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b873cfa),
	.w1(32'hbb6bc9f6),
	.w2(32'hbabf53ba),
	.w3(32'h3c301c87),
	.w4(32'h3b83cc53),
	.w5(32'h3b39e266),
	.w6(32'h39c7b9fc),
	.w7(32'h3b81c6aa),
	.w8(32'h3b6ee20a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c88f8),
	.w1(32'h3d52af6c),
	.w2(32'hbdc6ecf2),
	.w3(32'hbd5bd94e),
	.w4(32'hbd714e24),
	.w5(32'hbd8a50b9),
	.w6(32'h3d4b47eb),
	.w7(32'hbd6fc143),
	.w8(32'hbcd3f848),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2273e0),
	.w1(32'hbcc524d6),
	.w2(32'h3959aa3e),
	.w3(32'hbcf0469e),
	.w4(32'hbc292a50),
	.w5(32'h3b6cc67f),
	.w6(32'hbc4b619d),
	.w7(32'hbaa74024),
	.w8(32'h3bcc1d38),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0275f4),
	.w1(32'h3b0eaa1d),
	.w2(32'hb8a69282),
	.w3(32'h3a69ebd9),
	.w4(32'hbb38aeb7),
	.w5(32'hbb9017cd),
	.w6(32'hba8d0e05),
	.w7(32'hbb83fa18),
	.w8(32'hbbc6f4ad),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19823e),
	.w1(32'h3c0f4f82),
	.w2(32'h3a03fe29),
	.w3(32'hbc385b83),
	.w4(32'hbb0a52d5),
	.w5(32'hba4613d2),
	.w6(32'hbc152e38),
	.w7(32'hb81e7cae),
	.w8(32'h3b17fd86),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0383d1),
	.w1(32'h3bd6853a),
	.w2(32'h3b62e22d),
	.w3(32'h3b8dccb1),
	.w4(32'h3a542f26),
	.w5(32'hbb0f4042),
	.w6(32'h3ba2f042),
	.w7(32'hba13c93c),
	.w8(32'h3bba46af),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be96454),
	.w1(32'h3aaec52b),
	.w2(32'h3d0081d3),
	.w3(32'hbb66fc7a),
	.w4(32'hbb8873a1),
	.w5(32'h3cc07a2f),
	.w6(32'hbaa36cb0),
	.w7(32'hbbfe30e2),
	.w8(32'h3cabf785),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4ecb0d),
	.w1(32'h3c8df4f6),
	.w2(32'hbb97de23),
	.w3(32'h3c024043),
	.w4(32'hba517257),
	.w5(32'hba9d4e57),
	.w6(32'hba0f8046),
	.w7(32'h3a5d4d57),
	.w8(32'h3ac48ccf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4ca91),
	.w1(32'h3b550d7e),
	.w2(32'hba9ff4a2),
	.w3(32'h3c7b305d),
	.w4(32'h3c09b3a5),
	.w5(32'h3aa0b339),
	.w6(32'h3bfd817d),
	.w7(32'h3b0b1343),
	.w8(32'hbb7a3e28),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8aba3),
	.w1(32'hbc44b8ad),
	.w2(32'hbc0de2ed),
	.w3(32'hbc3dbe56),
	.w4(32'hbc0d534f),
	.w5(32'hb94fbe58),
	.w6(32'hbb9b56c5),
	.w7(32'hbb998dd9),
	.w8(32'hb9bd0ea6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf48e0),
	.w1(32'hbc23ce78),
	.w2(32'hbb82bf4c),
	.w3(32'hbc0902d8),
	.w4(32'hbb62c5bb),
	.w5(32'h3bb4f653),
	.w6(32'hbc196d1d),
	.w7(32'hbc8d0b3e),
	.w8(32'hbba670e6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2174fe),
	.w1(32'hbb8cfc06),
	.w2(32'h3ab85a76),
	.w3(32'hba5d7076),
	.w4(32'hbb8625b7),
	.w5(32'hbc2d4f64),
	.w6(32'hbc31848f),
	.w7(32'hb9d8d76f),
	.w8(32'hbc5713c3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bbe2b),
	.w1(32'hbc056603),
	.w2(32'hbc394132),
	.w3(32'hbb3e988e),
	.w4(32'hbbd5232b),
	.w5(32'hbace2e58),
	.w6(32'hbb93e517),
	.w7(32'hbc13a288),
	.w8(32'hbb10c0c4),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada2ca4),
	.w1(32'hbbe36ff2),
	.w2(32'hbb3c6ab3),
	.w3(32'hbc1d3f9f),
	.w4(32'h3975dd59),
	.w5(32'h39cdb6f5),
	.w6(32'hbbe75694),
	.w7(32'hbafaead2),
	.w8(32'hba9a784b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8cc0c),
	.w1(32'hbc8c9339),
	.w2(32'hbccfcc0f),
	.w3(32'hbcd1464a),
	.w4(32'hbc589b31),
	.w5(32'hbca2267c),
	.w6(32'hbbbf054d),
	.w7(32'h3c25029f),
	.w8(32'hbc0d9e60),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61b008),
	.w1(32'hba1f048b),
	.w2(32'hbc5d711a),
	.w3(32'hbbea9cb3),
	.w4(32'hbb41b687),
	.w5(32'hb92f874d),
	.w6(32'hbb3984a1),
	.w7(32'hbc6b574a),
	.w8(32'hbc2038d7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb299a11),
	.w1(32'h3a790274),
	.w2(32'hbc2837ab),
	.w3(32'hbbbff068),
	.w4(32'hbc4fcbeb),
	.w5(32'hbbe73d49),
	.w6(32'hbbc33283),
	.w7(32'hbc8b40a7),
	.w8(32'hbc75a7f6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59252f),
	.w1(32'hbc4bc87c),
	.w2(32'h3b2328e7),
	.w3(32'hbc87b0cf),
	.w4(32'hbb8360a0),
	.w5(32'hbb2408a4),
	.w6(32'hbc3f0175),
	.w7(32'h39bd7aa3),
	.w8(32'h3bdca867),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a866a),
	.w1(32'hbc066d3d),
	.w2(32'h3abee1db),
	.w3(32'hbc77ee74),
	.w4(32'hbc2d7208),
	.w5(32'h3bf8c313),
	.w6(32'hbb5fc07b),
	.w7(32'h3a95e156),
	.w8(32'h3c8dca75),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37f229),
	.w1(32'hbbd01c6c),
	.w2(32'hbbf27425),
	.w3(32'hbc0cbe46),
	.w4(32'hbbd41443),
	.w5(32'h3b5f31b5),
	.w6(32'hbb52bca5),
	.w7(32'hbbc5a3a8),
	.w8(32'h3b0145b2),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae954ec),
	.w1(32'h3a8f6467),
	.w2(32'hbb70a8da),
	.w3(32'hbbcce47e),
	.w4(32'hbc03b70b),
	.w5(32'hbbcf036f),
	.w6(32'hbc101675),
	.w7(32'hbae7e532),
	.w8(32'h3a027ced),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f92a6),
	.w1(32'hbc03e9c4),
	.w2(32'hbb33bed7),
	.w3(32'hbc39e583),
	.w4(32'hbbc8c3dd),
	.w5(32'h3b04a79e),
	.w6(32'h395e46aa),
	.w7(32'h399473f1),
	.w8(32'h3c5c2365),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc130702),
	.w1(32'hbb25abae),
	.w2(32'hbbfa57e2),
	.w3(32'hb99e8010),
	.w4(32'hbb52f925),
	.w5(32'hbc2d6d42),
	.w6(32'hba26afd1),
	.w7(32'hbba04408),
	.w8(32'hbc65a614),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b0306),
	.w1(32'hbb33817b),
	.w2(32'hbbd77d2a),
	.w3(32'hbcaa7f71),
	.w4(32'hbb667a05),
	.w5(32'hbc2c60ac),
	.w6(32'hbbf82c9c),
	.w7(32'hbad541c6),
	.w8(32'hbc0fb9ce),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5a404),
	.w1(32'h3b9901f7),
	.w2(32'h3be675c4),
	.w3(32'hbc6a84bc),
	.w4(32'h3cae5890),
	.w5(32'h3b12f743),
	.w6(32'hbb8bad49),
	.w7(32'h3ce39c0d),
	.w8(32'h3b073a36),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd36f62),
	.w1(32'h3c62141a),
	.w2(32'h3c13855c),
	.w3(32'hbca51cd0),
	.w4(32'hbbc2fdb6),
	.w5(32'h3c25bbe8),
	.w6(32'h3c1a7e28),
	.w7(32'h3cbb72db),
	.w8(32'h3d3a539e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fd75d),
	.w1(32'h3c50b4ab),
	.w2(32'h3b94cfa0),
	.w3(32'h3c8b4a6f),
	.w4(32'h3c02964f),
	.w5(32'h3ba6cd0b),
	.w6(32'h3cd67448),
	.w7(32'h3c48f560),
	.w8(32'h3c0ef487),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9902b3),
	.w1(32'hbcc5595f),
	.w2(32'hbaf1edd0),
	.w3(32'hbc565dff),
	.w4(32'hbbaf0f54),
	.w5(32'h3ba8cdf9),
	.w6(32'hbc2394f1),
	.w7(32'h3b685bf1),
	.w8(32'h3c1002b5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7c519),
	.w1(32'h3b4af71d),
	.w2(32'hbb083844),
	.w3(32'hbab2bc5b),
	.w4(32'h3ba51a5b),
	.w5(32'h3bc3e20a),
	.w6(32'hb91127ea),
	.w7(32'hbb35f25a),
	.w8(32'hbb77c8e6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0a481),
	.w1(32'hbcc5ced7),
	.w2(32'hbbf2d0a1),
	.w3(32'hbbcadf70),
	.w4(32'hbc6660f6),
	.w5(32'h3c09570f),
	.w6(32'hbc44f437),
	.w7(32'hbafa2aa2),
	.w8(32'h3c3de511),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7edee5),
	.w1(32'h3b118c5b),
	.w2(32'h3ae75497),
	.w3(32'hbc03e58f),
	.w4(32'h3b469a0e),
	.w5(32'hbbbe2ba4),
	.w6(32'hbb6548ef),
	.w7(32'h3bfddc0c),
	.w8(32'h3b4b1535),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fdd59),
	.w1(32'h3bec30ad),
	.w2(32'hbcc9c50f),
	.w3(32'hbca8c0b3),
	.w4(32'hbcaa3bf5),
	.w5(32'hbcd103fe),
	.w6(32'hbb02ea81),
	.w7(32'hbc6e410b),
	.w8(32'hbc8b223a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd14da8a),
	.w1(32'hbce9e318),
	.w2(32'h3a823cfb),
	.w3(32'hbcbeed81),
	.w4(32'hbc39b4a6),
	.w5(32'hbb437820),
	.w6(32'hbca61809),
	.w7(32'hbbb88dff),
	.w8(32'h3bc0f53c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc12b9),
	.w1(32'hb9e1b964),
	.w2(32'hbc8cacf0),
	.w3(32'hbbabd9af),
	.w4(32'hbc4bc792),
	.w5(32'hbb9252d6),
	.w6(32'hbb8d7f0f),
	.w7(32'hbc347298),
	.w8(32'hb9f4da5d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb395a90),
	.w1(32'hbc5fab00),
	.w2(32'hbc1bcc9d),
	.w3(32'h3b0f591d),
	.w4(32'hbac8df25),
	.w5(32'hbbc08622),
	.w6(32'hbb0d52ac),
	.w7(32'hbbf24a33),
	.w8(32'hbbb9873f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c321a),
	.w1(32'h3c10e41c),
	.w2(32'hbc4d9a94),
	.w3(32'h3bed2848),
	.w4(32'hbbefd138),
	.w5(32'hbc5ac251),
	.w6(32'h3babcf65),
	.w7(32'hbc6a1d93),
	.w8(32'hbc877616),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce17bc9),
	.w1(32'hbc91bb12),
	.w2(32'hbc96247e),
	.w3(32'hbccff013),
	.w4(32'hbc55e09e),
	.w5(32'hbc2dcef6),
	.w6(32'hbc24dae9),
	.w7(32'h3b8aa7a6),
	.w8(32'h3b5aac48),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe1f1e),
	.w1(32'hbc1ca059),
	.w2(32'h3afc9f0d),
	.w3(32'hbbe309a1),
	.w4(32'hbb2d18cd),
	.w5(32'h3b9a9900),
	.w6(32'hbbe45a53),
	.w7(32'hbbb7c508),
	.w8(32'h3b7bba81),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0168d4),
	.w1(32'h3baa350b),
	.w2(32'hbc098082),
	.w3(32'h3b074340),
	.w4(32'hbb8a00e7),
	.w5(32'hbbc0496f),
	.w6(32'h3b1a1e64),
	.w7(32'hbbaaab6b),
	.w8(32'hbbc0e19c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10c156),
	.w1(32'hbbc4deec),
	.w2(32'hbb2758bd),
	.w3(32'hbc0d50a1),
	.w4(32'h3b32bcce),
	.w5(32'hbbd97d76),
	.w6(32'hbbc566cc),
	.w7(32'h3b8cc6a6),
	.w8(32'hbab6a318),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37b741),
	.w1(32'h3b79b814),
	.w2(32'hbc1b4275),
	.w3(32'hbbfc90c2),
	.w4(32'hbaa4ab4d),
	.w5(32'h3b84cb86),
	.w6(32'h39b80a88),
	.w7(32'hbb7b5c8e),
	.w8(32'h3af355d6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eee28),
	.w1(32'hbc423bef),
	.w2(32'h3c313fc8),
	.w3(32'hbb80ffe1),
	.w4(32'hbbbf3ee2),
	.w5(32'h3c263fc9),
	.w6(32'h3a9c16f0),
	.w7(32'hbba33bbc),
	.w8(32'h3c44d670),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf86657),
	.w1(32'h3b3afcb5),
	.w2(32'h3acece85),
	.w3(32'hbb1e058c),
	.w4(32'hbb7bd70e),
	.w5(32'hbc106928),
	.w6(32'hbc058940),
	.w7(32'hbbda4595),
	.w8(32'hbbb06570),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a21de),
	.w1(32'hbc59dc38),
	.w2(32'h3b53cdf7),
	.w3(32'hbcb3a105),
	.w4(32'hbccf2113),
	.w5(32'h3bb3bfcf),
	.w6(32'hbc5b3d07),
	.w7(32'hbb516c09),
	.w8(32'h3ca84562),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a4047),
	.w1(32'h3c2e9e64),
	.w2(32'hbbf10aaa),
	.w3(32'h3be2bb40),
	.w4(32'hbb9b6924),
	.w5(32'hbbf5f900),
	.w6(32'h3bafe827),
	.w7(32'hbc15c22e),
	.w8(32'hbbf3ed02),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98f5ef),
	.w1(32'h3b311cae),
	.w2(32'hbbcf5cd0),
	.w3(32'hbc0315d5),
	.w4(32'hbc0d4b6d),
	.w5(32'hbb0e1cfd),
	.w6(32'hba3780a2),
	.w7(32'hbb80ba1e),
	.w8(32'h3c12e16c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aba68),
	.w1(32'hbb4a1220),
	.w2(32'hbb2cea10),
	.w3(32'h3bd8cedc),
	.w4(32'h3b75072e),
	.w5(32'hbb2a7ec0),
	.w6(32'h3a9110c4),
	.w7(32'hbc1128a9),
	.w8(32'hbc2c327a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbec1fc),
	.w1(32'hbc545548),
	.w2(32'hbba8f199),
	.w3(32'hbca8b9eb),
	.w4(32'h3af5c5d5),
	.w5(32'h3bb44e82),
	.w6(32'hbc946042),
	.w7(32'hbbfeb3d0),
	.w8(32'hbba644c1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf53c89),
	.w1(32'hbc664972),
	.w2(32'hb8ac872a),
	.w3(32'hbba41b22),
	.w4(32'h3a313ac1),
	.w5(32'hbb02ba8a),
	.w6(32'hbbb40c61),
	.w7(32'h388d0639),
	.w8(32'hbad72119),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1c3a7),
	.w1(32'h3c42af0e),
	.w2(32'hbab9c284),
	.w3(32'hb981d829),
	.w4(32'hba06f4ae),
	.w5(32'hb99f0951),
	.w6(32'h3c3c9fe7),
	.w7(32'hba8f6007),
	.w8(32'h3b56aa56),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae6ff1),
	.w1(32'h3ab826ed),
	.w2(32'h379f0393),
	.w3(32'hbbde86ca),
	.w4(32'hb80585fd),
	.w5(32'h370dba4c),
	.w6(32'hbbabcb93),
	.w7(32'h3598437a),
	.w8(32'h3777eb36),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbdb85),
	.w1(32'hbbebfc42),
	.w2(32'hbb9654eb),
	.w3(32'hbc1b5cde),
	.w4(32'hbbe0741d),
	.w5(32'h3b82d6cc),
	.w6(32'hbb32ca44),
	.w7(32'h3ad280de),
	.w8(32'h3c192cef),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30eed5),
	.w1(32'hbbf61e07),
	.w2(32'h3a5fbade),
	.w3(32'hbbd3a191),
	.w4(32'hbb865a5e),
	.w5(32'h3baca11f),
	.w6(32'hbb5d5746),
	.w7(32'h3ab37bce),
	.w8(32'h3be65f93),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea0d3c),
	.w1(32'h3a28b42f),
	.w2(32'h39f1cebe),
	.w3(32'h39887fd7),
	.w4(32'h39c1c9c3),
	.w5(32'h39e49d65),
	.w6(32'h3a28dfdc),
	.w7(32'h3a05b96f),
	.w8(32'h39a3ecbf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f429ae),
	.w1(32'h371ecf91),
	.w2(32'h393eee0d),
	.w3(32'hb7e5f6c9),
	.w4(32'h37b8643f),
	.w5(32'h3954121d),
	.w6(32'hb79eac8d),
	.w7(32'h38824e80),
	.w8(32'h393a1325),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5d517),
	.w1(32'h3a80ca3f),
	.w2(32'hbafed48f),
	.w3(32'h3ada323f),
	.w4(32'hbaf75bd8),
	.w5(32'hbba68527),
	.w6(32'hbb825931),
	.w7(32'hbc24678a),
	.w8(32'hbbdedbbd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8da26d),
	.w1(32'hbbb428e5),
	.w2(32'hbba00d8f),
	.w3(32'hbc1c4b7e),
	.w4(32'hbbfbd788),
	.w5(32'h3ac55062),
	.w6(32'h3a6eb175),
	.w7(32'h3b8394d9),
	.w8(32'h3c16a24e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc937f04),
	.w1(32'hbca4311e),
	.w2(32'hbcf9f87e),
	.w3(32'hbc8c4f8c),
	.w4(32'hbba86a61),
	.w5(32'hbc72367d),
	.w6(32'h3b5bf17c),
	.w7(32'h3cc275ec),
	.w8(32'hbbd6ec5d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77e9c2),
	.w1(32'hbc9bfda5),
	.w2(32'hbbfe5b5c),
	.w3(32'hbcc49a77),
	.w4(32'hbc7820a1),
	.w5(32'h3be6eeab),
	.w6(32'h3a0bb6d0),
	.w7(32'h3bf9a3da),
	.w8(32'h3ca5d7ad),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7ea2b),
	.w1(32'h38f8bd72),
	.w2(32'hbabd51e7),
	.w3(32'hbb578849),
	.w4(32'hbb2ab605),
	.w5(32'hbb419255),
	.w6(32'h3a84413f),
	.w7(32'hbb36822f),
	.w8(32'h3b9c5b77),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b2c2c),
	.w1(32'hb735cc5a),
	.w2(32'h39337a6b),
	.w3(32'h383f273c),
	.w4(32'h392809f1),
	.w5(32'h3945af40),
	.w6(32'hb81e8dac),
	.w7(32'h389c527c),
	.w8(32'hb830bbb8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89b778c),
	.w1(32'hb8ff7262),
	.w2(32'hb811a08f),
	.w3(32'hb8c0ba3e),
	.w4(32'hb8c7baa3),
	.w5(32'h35796282),
	.w6(32'hb8d74899),
	.w7(32'hb8a6514e),
	.w8(32'hb79700c8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f889c4),
	.w1(32'h381ca8b9),
	.w2(32'h36cf57ac),
	.w3(32'h39050169),
	.w4(32'hb88e8b4d),
	.w5(32'h364b0d6c),
	.w6(32'h38da44ec),
	.w7(32'hb8631c88),
	.w8(32'h37d4072a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c7a84),
	.w1(32'hb8ee7420),
	.w2(32'h3a19b9b0),
	.w3(32'hbac01733),
	.w4(32'hbb0d4ef1),
	.w5(32'h39925953),
	.w6(32'hb9dc1f11),
	.w7(32'hba339ddf),
	.w8(32'h3a72b634),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83a5d4),
	.w1(32'hbb35680c),
	.w2(32'hbb439c40),
	.w3(32'hbb92386a),
	.w4(32'hbb22235e),
	.w5(32'hbb3f1e9f),
	.w6(32'h3a5563ba),
	.w7(32'hb93f4775),
	.w8(32'hba7c5318),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39574de0),
	.w1(32'h3989415d),
	.w2(32'h38ae1a13),
	.w3(32'h39905f7b),
	.w4(32'h399421ab),
	.w5(32'h39b8dca1),
	.w6(32'h39a9bb97),
	.w7(32'h399dcd18),
	.w8(32'h39b27a1a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddbf00),
	.w1(32'h3bc90135),
	.w2(32'h3b087303),
	.w3(32'h3b501b25),
	.w4(32'h3b224f80),
	.w5(32'hba438565),
	.w6(32'hb9b222f9),
	.w7(32'h3ab7ac26),
	.w8(32'hba556c8f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11f95f),
	.w1(32'hbb0ec254),
	.w2(32'hba67386c),
	.w3(32'hbb3acbad),
	.w4(32'hbac89881),
	.w5(32'h3b2a9723),
	.w6(32'h3abaf1a1),
	.w7(32'h3b6dffea),
	.w8(32'h3bbba450),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ff0e6),
	.w1(32'hb9c73c1f),
	.w2(32'h3a8cf95b),
	.w3(32'h3af268d6),
	.w4(32'h3b4cdeb6),
	.w5(32'h3b0732af),
	.w6(32'h3b17cd93),
	.w7(32'h3b1db690),
	.w8(32'hb794bff4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b785725),
	.w1(32'hbb2fe97a),
	.w2(32'hbb1c9cdc),
	.w3(32'h3b826c1a),
	.w4(32'hba65e700),
	.w5(32'h3b1c8f4a),
	.w6(32'h3bbfebd7),
	.w7(32'h3b4d442e),
	.w8(32'h3c0b1cb8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18d0ae),
	.w1(32'h3a94458b),
	.w2(32'h3b1eb300),
	.w3(32'hbb7174b0),
	.w4(32'h3a1db5cb),
	.w5(32'h3b46fe2e),
	.w6(32'h3b6926e5),
	.w7(32'h3bb7beba),
	.w8(32'h3be2d1eb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a2aaa),
	.w1(32'hb905046e),
	.w2(32'h38842cc1),
	.w3(32'hb8a645c1),
	.w4(32'hb8e8e9d3),
	.w5(32'h388242e8),
	.w6(32'hb8fdfb55),
	.w7(32'hb90840f5),
	.w8(32'h388b6158),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394258fc),
	.w1(32'h37d64b59),
	.w2(32'h38f41cc9),
	.w3(32'h391bd5d0),
	.w4(32'hb8958de5),
	.w5(32'hb7b80db6),
	.w6(32'h370d45a5),
	.w7(32'hb9685f6e),
	.w8(32'hb8655e6b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39136065),
	.w1(32'h383f8044),
	.w2(32'h381b9898),
	.w3(32'h38fce4bd),
	.w4(32'hb856d87b),
	.w5(32'hb8574329),
	.w6(32'h3781c015),
	.w7(32'hb903a0f5),
	.w8(32'hb8c535ed),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a7d13),
	.w1(32'hb98cfb3d),
	.w2(32'hb99fe168),
	.w3(32'hb91d082c),
	.w4(32'hb9a055c6),
	.w5(32'hb9a42f8d),
	.w6(32'hb8b814b4),
	.w7(32'hb919a28e),
	.w8(32'hb9390153),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62b243),
	.w1(32'hba8157e5),
	.w2(32'h3a2f6a37),
	.w3(32'hba0728d6),
	.w4(32'h3b239f0a),
	.w5(32'h3b783373),
	.w6(32'hbb07caef),
	.w7(32'hb84b64cc),
	.w8(32'h3af25662),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e93623),
	.w1(32'h39c37eed),
	.w2(32'h395ca6aa),
	.w3(32'h3a38fb28),
	.w4(32'h3a59f19d),
	.w5(32'h3a831e5e),
	.w6(32'h3a7c2b5e),
	.w7(32'h3a618a13),
	.w8(32'h3a8bf5e9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e9a05),
	.w1(32'h3b8fa968),
	.w2(32'h3acd4724),
	.w3(32'h3bb4bf7c),
	.w4(32'h3bb33ca9),
	.w5(32'h3ab6a82f),
	.w6(32'hbb1dfd96),
	.w7(32'hbb6d2919),
	.w8(32'hbbba2ae3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ac939),
	.w1(32'h3ad5640d),
	.w2(32'h3aadfbad),
	.w3(32'h3b54e473),
	.w4(32'h3b3f43e3),
	.w5(32'h3a80a18e),
	.w6(32'h3a467386),
	.w7(32'h3915621a),
	.w8(32'hba7b77f8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1878dc),
	.w1(32'hbba3178b),
	.w2(32'h3a03d493),
	.w3(32'hbc3b3bde),
	.w4(32'hbc4f1f12),
	.w5(32'h3b934f30),
	.w6(32'hbb187055),
	.w7(32'hbb905ea1),
	.w8(32'h3c09aac4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe1db2),
	.w1(32'h3a6dc05c),
	.w2(32'hb9d37c98),
	.w3(32'h3aba4e11),
	.w4(32'h396466a9),
	.w5(32'h3a6b5695),
	.w6(32'h3b0c2ce7),
	.w7(32'h38eeaa9d),
	.w8(32'h3a589512),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8df8ff),
	.w1(32'h3b57a45c),
	.w2(32'h3b0b2e04),
	.w3(32'h3b7996b7),
	.w4(32'h3b203bcc),
	.w5(32'h38bfdb96),
	.w6(32'h3b39f820),
	.w7(32'h3b02354b),
	.w8(32'h39b21992),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dca7b3),
	.w1(32'hb96c1e9f),
	.w2(32'hb9b2c321),
	.w3(32'h39d10b22),
	.w4(32'h39c8da80),
	.w5(32'hba5c96ae),
	.w6(32'hbac7205a),
	.w7(32'hbac44c02),
	.w8(32'hbb07f08d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf05b68),
	.w1(32'h3b15d624),
	.w2(32'h3b9aec98),
	.w3(32'hbb31ecbc),
	.w4(32'h3a890a18),
	.w5(32'h3b4d07bd),
	.w6(32'hbb29e67a),
	.w7(32'h3a5f8be8),
	.w8(32'h3b87f847),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45018f),
	.w1(32'hba14ee68),
	.w2(32'hb9bd4b54),
	.w3(32'hba1e6ab1),
	.w4(32'hba7dd24c),
	.w5(32'hbac9598d),
	.w6(32'h3b65a431),
	.w7(32'h3b8daef1),
	.w8(32'h3a3bcf4d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b1bfc),
	.w1(32'hbb540486),
	.w2(32'hbb96c3ae),
	.w3(32'hbb24adda),
	.w4(32'hba8eace3),
	.w5(32'hbb350b0d),
	.w6(32'h3aaae389),
	.w7(32'hb9268a8b),
	.w8(32'hbb28c54a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae46e13),
	.w1(32'h3b6ca535),
	.w2(32'h3b944317),
	.w3(32'h3ae3c12a),
	.w4(32'h3b870d7e),
	.w5(32'h3b1ca322),
	.w6(32'hbad70df1),
	.w7(32'hb9faf75f),
	.w8(32'hbac7e699),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9651b55),
	.w1(32'hb9a4db8c),
	.w2(32'h37d64999),
	.w3(32'hba1aec20),
	.w4(32'hb708db0e),
	.w5(32'hb99a80ba),
	.w6(32'hb95a0ad6),
	.w7(32'hb8d44b04),
	.w8(32'hb919e293),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cca5f),
	.w1(32'hbae61cab),
	.w2(32'hba962bd4),
	.w3(32'hbb23c55f),
	.w4(32'hbae68bb2),
	.w5(32'hbaa62624),
	.w6(32'hbb283a06),
	.w7(32'hbaaa4e07),
	.w8(32'hba0b6473),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa52185),
	.w1(32'hbaaddd94),
	.w2(32'hb93638ec),
	.w3(32'hba878f46),
	.w4(32'hbab33941),
	.w5(32'h399e6679),
	.w6(32'hb918e893),
	.w7(32'hb970df60),
	.w8(32'h3a983e75),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a859d26),
	.w1(32'h3ac97ffe),
	.w2(32'h3a4f7608),
	.w3(32'h3a90a608),
	.w4(32'hbadf6255),
	.w5(32'hbb2271fc),
	.w6(32'h3b0844c7),
	.w7(32'h3a0881b5),
	.w8(32'h3a84241d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fb9d2),
	.w1(32'hbb6327f2),
	.w2(32'hbb509d0c),
	.w3(32'hbc23d519),
	.w4(32'hbc06c7e8),
	.w5(32'hba20b971),
	.w6(32'hbb83d09e),
	.w7(32'h38a0f83f),
	.w8(32'h3b7e96d0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387d57d5),
	.w1(32'h38287003),
	.w2(32'h38413da4),
	.w3(32'h38848fdd),
	.w4(32'h38041ace),
	.w5(32'h37d314b3),
	.w6(32'h37f5e462),
	.w7(32'hb625006a),
	.w8(32'h3764d7b3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ab99f),
	.w1(32'hba3c1be2),
	.w2(32'h389f7005),
	.w3(32'hb936dee6),
	.w4(32'h39cc7e4f),
	.w5(32'h3a7e66eb),
	.w6(32'h39c780af),
	.w7(32'h3a736549),
	.w8(32'h3a94f347),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ed268),
	.w1(32'hbaadd526),
	.w2(32'h3a7cd41e),
	.w3(32'hbb699660),
	.w4(32'hbbe077fc),
	.w5(32'hbb2a37d7),
	.w6(32'hba464b5b),
	.w7(32'h3a314b6e),
	.w8(32'h3bf32c27),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03fcdb),
	.w1(32'h3a9ecf85),
	.w2(32'hbaf6816c),
	.w3(32'h3b33341b),
	.w4(32'h3c04e77e),
	.w5(32'h3afd8cae),
	.w6(32'h3b0d3baa),
	.w7(32'h3b813237),
	.w8(32'hbaa931f4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e30cea),
	.w1(32'hb9abccde),
	.w2(32'hb81157d1),
	.w3(32'h39f97e3b),
	.w4(32'hb9276fef),
	.w5(32'hb9d9f7f6),
	.w6(32'h393bd05a),
	.w7(32'hb925286b),
	.w8(32'hb9eb4ffd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ca16b),
	.w1(32'h3a13c984),
	.w2(32'h38bc48fc),
	.w3(32'h3b111844),
	.w4(32'h3ac2430d),
	.w5(32'h39076c94),
	.w6(32'h3b186d4f),
	.w7(32'h3b0dd42a),
	.w8(32'h3a7e3b15),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9db823),
	.w1(32'h39728b55),
	.w2(32'h391f69a9),
	.w3(32'hbaaf0e89),
	.w4(32'h399a4f1d),
	.w5(32'h3a106405),
	.w6(32'hb9874cc6),
	.w7(32'h3a53e60c),
	.w8(32'h3ac8f839),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8bb55),
	.w1(32'hbb3c8ecf),
	.w2(32'hbb871312),
	.w3(32'hbb0005de),
	.w4(32'hbb98f423),
	.w5(32'hbacc5bf0),
	.w6(32'hbb3cf851),
	.w7(32'hbaf3b5f8),
	.w8(32'h3b129691),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb104453),
	.w1(32'h3aa80452),
	.w2(32'h3b3a79cb),
	.w3(32'h3a678fb4),
	.w4(32'h3b57e3f5),
	.w5(32'h3b7bd51f),
	.w6(32'h3b4481c2),
	.w7(32'h3b8c7e60),
	.w8(32'h3b1c9a91),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d46ff),
	.w1(32'hbbb3e762),
	.w2(32'hbb3b17b6),
	.w3(32'hba9321f2),
	.w4(32'hbbe4bfb3),
	.w5(32'hbad686d3),
	.w6(32'hbb206919),
	.w7(32'hbb544744),
	.w8(32'h3b8cb955),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule