module layer_8_featuremap_76(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebea32),
	.w1(32'hb9255c2c),
	.w2(32'h3c43869a),
	.w3(32'hbc347abe),
	.w4(32'hbae473d1),
	.w5(32'h3bdad881),
	.w6(32'hbbd89709),
	.w7(32'hbb702391),
	.w8(32'h3b9f44ee),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb143a2e),
	.w1(32'hbb70e897),
	.w2(32'hbba5b4de),
	.w3(32'hbb8a1649),
	.w4(32'hbae1eea6),
	.w5(32'hbbe46794),
	.w6(32'hbbfd24e8),
	.w7(32'hba37e5a2),
	.w8(32'hbb31e36a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2835a),
	.w1(32'h3ba27c2b),
	.w2(32'h3b45e11b),
	.w3(32'h3b5625d7),
	.w4(32'h3b16290b),
	.w5(32'hbb095c4f),
	.w6(32'h3b0e4ed5),
	.w7(32'h3bcc886b),
	.w8(32'h39d40388),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb35778),
	.w1(32'h3b00d4eb),
	.w2(32'hbc2714b5),
	.w3(32'hbbf27f3c),
	.w4(32'h3bfe8d56),
	.w5(32'hbc8353ff),
	.w6(32'hbba9e812),
	.w7(32'hbab6d850),
	.w8(32'hbbe41c6a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c9bac),
	.w1(32'hbbead3a6),
	.w2(32'hbb450862),
	.w3(32'hbbebb367),
	.w4(32'hba9d1b02),
	.w5(32'hbb1052e0),
	.w6(32'hbc14e9f5),
	.w7(32'hbbca8a50),
	.w8(32'hbba85c8b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2435ac),
	.w1(32'h3b0eac87),
	.w2(32'hbd44442e),
	.w3(32'h3d6ef818),
	.w4(32'h3d84b944),
	.w5(32'h3c243e4e),
	.w6(32'hbd4916d1),
	.w7(32'hbd39b1cd),
	.w8(32'hbc4b995c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94c406),
	.w1(32'hbb81759f),
	.w2(32'hbba400db),
	.w3(32'hbc0dc786),
	.w4(32'hbb63cc33),
	.w5(32'hbb8abbfc),
	.w6(32'hbbd691f5),
	.w7(32'hbb842d0a),
	.w8(32'hba2a731c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba219d9e),
	.w1(32'hba29362a),
	.w2(32'h3c1d9265),
	.w3(32'hbc3062dd),
	.w4(32'hbae382ae),
	.w5(32'h3baf393b),
	.w6(32'hbc30013a),
	.w7(32'hbb5b7667),
	.w8(32'h3b08e135),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14de1b),
	.w1(32'hbbc67b31),
	.w2(32'hbb04d790),
	.w3(32'hbc3a0ea5),
	.w4(32'hbbbb0a6b),
	.w5(32'hbadd8cee),
	.w6(32'hbbc5b7b4),
	.w7(32'hba81ed2d),
	.w8(32'hbb86457c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc56c4d),
	.w1(32'hbbae95d6),
	.w2(32'hbb8ecd0c),
	.w3(32'hbbc4e439),
	.w4(32'hbc00a3da),
	.w5(32'hbc02571b),
	.w6(32'hbc882d8b),
	.w7(32'h3b67d161),
	.w8(32'h3ae5bf28),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e8bee),
	.w1(32'h3ad88925),
	.w2(32'h3c48823c),
	.w3(32'hbc9afc70),
	.w4(32'hbbc3fa5b),
	.w5(32'h3c67c3a4),
	.w6(32'hbbc7b9a1),
	.w7(32'hbbbb67f9),
	.w8(32'h3b9d1740),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9db65),
	.w1(32'hbb6ffaa8),
	.w2(32'hb98e9102),
	.w3(32'hbc1a24f5),
	.w4(32'hbbf5d7fb),
	.w5(32'hbbb7b688),
	.w6(32'hbbbddf54),
	.w7(32'hbb2b3991),
	.w8(32'hbb755801),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdc6d5),
	.w1(32'hbc274fdb),
	.w2(32'hbc233e75),
	.w3(32'hbbfc5905),
	.w4(32'hbba04354),
	.w5(32'hbbf34f66),
	.w6(32'hbbed2784),
	.w7(32'hbb3c882d),
	.w8(32'hbc39ed09),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d072b13),
	.w1(32'hbb643f64),
	.w2(32'hbd2768c7),
	.w3(32'h3d802596),
	.w4(32'h3d8df883),
	.w5(32'h3ca06bb4),
	.w6(32'hbd507250),
	.w7(32'hbd309642),
	.w8(32'hbb8a405e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9db20a),
	.w1(32'hbba80ddf),
	.w2(32'hbcfde40f),
	.w3(32'h3cf78fc8),
	.w4(32'h3d1a747d),
	.w5(32'h3b7b5d93),
	.w6(32'hbd0de126),
	.w7(32'hbcf56770),
	.w8(32'hbb2f6bd5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f3302),
	.w1(32'hbb0c1ec9),
	.w2(32'hb99e8dff),
	.w3(32'h3a96301d),
	.w4(32'h3b3f6d91),
	.w5(32'hba69b2e7),
	.w6(32'hbc03bb85),
	.w7(32'h3afe0e0e),
	.w8(32'hbcacf093),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc711893),
	.w1(32'h3bfa8cb6),
	.w2(32'h3c12b891),
	.w3(32'hba7fc4b1),
	.w4(32'h3991efa6),
	.w5(32'hbc2d60cf),
	.w6(32'hbbfe68b6),
	.w7(32'hb8b557a8),
	.w8(32'h3b68a36b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67e5d6),
	.w1(32'hbb5f1426),
	.w2(32'h3bdf6cc8),
	.w3(32'hbc026053),
	.w4(32'hbb91735f),
	.w5(32'h3aa3ca2e),
	.w6(32'h3b992db6),
	.w7(32'h3bad7c3d),
	.w8(32'h3b485625),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88079c),
	.w1(32'h3bda88bf),
	.w2(32'h3d427ea8),
	.w3(32'hbcccde1a),
	.w4(32'h3ac11c98),
	.w5(32'h3d128d70),
	.w6(32'hbc364c69),
	.w7(32'hbc32c92c),
	.w8(32'hb9ca7cf6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70f7e9),
	.w1(32'hbcabc3da),
	.w2(32'h3d093b73),
	.w3(32'hbc2bc51e),
	.w4(32'hbd0c4d99),
	.w5(32'hbc059b69),
	.w6(32'hbca184e2),
	.w7(32'h3c926cfb),
	.w8(32'h3a976b45),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2608e2),
	.w1(32'h3c76b287),
	.w2(32'h3cb16b00),
	.w3(32'hbc88da1d),
	.w4(32'hbc1a6c49),
	.w5(32'hbb3e87d1),
	.w6(32'h3d2cc531),
	.w7(32'h3cf3e9e6),
	.w8(32'hbc204f46),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91842e),
	.w1(32'hbb297a65),
	.w2(32'hbbff8e8a),
	.w3(32'h3ab95547),
	.w4(32'h3bde7470),
	.w5(32'hbb4e5c50),
	.w6(32'hbbb86713),
	.w7(32'hbb8fb9e9),
	.w8(32'h3be0e7eb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd73def0),
	.w1(32'hbb882699),
	.w2(32'h3d4be12a),
	.w3(32'hbd71c8df),
	.w4(32'hbd695303),
	.w5(32'h3c77ed99),
	.w6(32'h3d2bac77),
	.w7(32'h3caa06b9),
	.w8(32'h38c87167),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88e444c),
	.w1(32'hbb803a3b),
	.w2(32'h3b7ae782),
	.w3(32'h3bc21239),
	.w4(32'h3bee8754),
	.w5(32'h39f1cd43),
	.w6(32'hbb5027de),
	.w7(32'h3c3521fb),
	.w8(32'hba0d4a5e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc39106),
	.w1(32'h3b9ae9f8),
	.w2(32'h3c9da9e1),
	.w3(32'hbc1b67c0),
	.w4(32'hbcc0850b),
	.w5(32'hba7371ae),
	.w6(32'h3c25f9d8),
	.w7(32'h3b3a5522),
	.w8(32'h3badf801),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd300c90),
	.w1(32'hbb7f8f51),
	.w2(32'h3ce40d15),
	.w3(32'hbd2de1c4),
	.w4(32'hbd4a2d40),
	.w5(32'hbb6f38bd),
	.w6(32'h3d1858f5),
	.w7(32'h3c97c1a2),
	.w8(32'hbbba113d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce0fa66),
	.w1(32'h3af24c8b),
	.w2(32'h3cae006c),
	.w3(32'hbccc0012),
	.w4(32'hbce7a597),
	.w5(32'h39a6f951),
	.w6(32'h3d19a2f9),
	.w7(32'h3cd98712),
	.w8(32'h3ad8132c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8e94ef),
	.w1(32'hbc11c46c),
	.w2(32'h3db805dd),
	.w3(32'hbdb91c25),
	.w4(32'hbd68389a),
	.w5(32'h3db6fba1),
	.w6(32'h3d774d77),
	.w7(32'h3c6d3793),
	.w8(32'hbdce9764),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c9daa),
	.w1(32'hb9f04f21),
	.w2(32'h3cb272e5),
	.w3(32'h3a66b755),
	.w4(32'hbc33a138),
	.w5(32'hbcbf2f12),
	.w6(32'hbcb87149),
	.w7(32'h3cca3021),
	.w8(32'hbb1e3a29),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20f4fd),
	.w1(32'hbb6b965c),
	.w2(32'hbb919bb3),
	.w3(32'hb991c74b),
	.w4(32'h3a0d17f1),
	.w5(32'hba718c2d),
	.w6(32'hbbe6831f),
	.w7(32'hbb5ecd6a),
	.w8(32'h3bc54f95),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ed279),
	.w1(32'hbc505976),
	.w2(32'hbca255b2),
	.w3(32'hbd269dc0),
	.w4(32'hbc549a32),
	.w5(32'hbb7ec9c2),
	.w6(32'hbc6b34bf),
	.w7(32'hbc963c95),
	.w8(32'h3be7ee08),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb13c8d),
	.w1(32'h3c564d79),
	.w2(32'h3cd89a6a),
	.w3(32'hbd12080c),
	.w4(32'hbcd2b743),
	.w5(32'hbb8b99af),
	.w6(32'h3d1b25d3),
	.w7(32'h3c61d1c7),
	.w8(32'hbbaec692),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1583fb),
	.w1(32'hbcb12880),
	.w2(32'hbd4df26a),
	.w3(32'hbc646ae6),
	.w4(32'hbbbe8a9e),
	.w5(32'hbd049c71),
	.w6(32'hbbf8e243),
	.w7(32'hbaf5cfc8),
	.w8(32'hbabf1979),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8d778),
	.w1(32'hbc00636c),
	.w2(32'h3beb9c04),
	.w3(32'hbc10af97),
	.w4(32'hbc0ead0d),
	.w5(32'hbc57b07c),
	.w6(32'h3bc621c7),
	.w7(32'h3b992a28),
	.w8(32'hbbb81cb9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdfe9bc),
	.w1(32'hbbc43f86),
	.w2(32'hbd21ebe6),
	.w3(32'h3d7b4cc7),
	.w4(32'h3d7ff973),
	.w5(32'h3c5fafc7),
	.w6(32'hbd31ea25),
	.w7(32'hbd0bedac),
	.w8(32'hba07f8a5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdfefd),
	.w1(32'hba7f9d80),
	.w2(32'h3ca59c51),
	.w3(32'hbbc4b97e),
	.w4(32'h3bb452dd),
	.w5(32'h3b952c4f),
	.w6(32'hbbe6c9a6),
	.w7(32'h3b571b77),
	.w8(32'h3ba96219),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc214117),
	.w1(32'h3bc12963),
	.w2(32'h3c65aa6b),
	.w3(32'hbcc7041f),
	.w4(32'hbc79a55a),
	.w5(32'h382cd6ac),
	.w6(32'h3cc84314),
	.w7(32'hb88c65bd),
	.w8(32'h3af10c9d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefd235),
	.w1(32'hbb9de287),
	.w2(32'hbb2b4598),
	.w3(32'hbad53b6f),
	.w4(32'hbb1cabc8),
	.w5(32'hba8776d1),
	.w6(32'hbbd1cd79),
	.w7(32'hbacff038),
	.w8(32'hbc153d69),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d10c6ce),
	.w1(32'hbc17d5d7),
	.w2(32'hbd79c569),
	.w3(32'h3d42b3d4),
	.w4(32'h3d8ad9b3),
	.w5(32'h3af4122c),
	.w6(32'hbd7c1b13),
	.w7(32'hbd6948ab),
	.w8(32'h3a1c5127),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7be452),
	.w1(32'h3a88ffa7),
	.w2(32'h3c3c4222),
	.w3(32'hbcd77c6c),
	.w4(32'hbca2e76d),
	.w5(32'hbb93273c),
	.w6(32'h3c90a242),
	.w7(32'h3bc197ba),
	.w8(32'h3b00781a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb67412),
	.w1(32'hbba3eeec),
	.w2(32'h3c2a5b02),
	.w3(32'hbd148700),
	.w4(32'hbd09dc43),
	.w5(32'hbc8aac26),
	.w6(32'h3b8d2b30),
	.w7(32'h3aebda21),
	.w8(32'hbc0fac08),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05bd5b),
	.w1(32'h3ba07a48),
	.w2(32'h3c1d522a),
	.w3(32'h3b536310),
	.w4(32'h3bbf60fe),
	.w5(32'h3bf1e6eb),
	.w6(32'h3c22ad9e),
	.w7(32'h3bbef7cb),
	.w8(32'hb96bf3d5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebe094),
	.w1(32'hbc51595c),
	.w2(32'h3c3ccb1a),
	.w3(32'h3b9d562f),
	.w4(32'hbc40bc9b),
	.w5(32'h3c156f28),
	.w6(32'hbc8d226d),
	.w7(32'h3c6eca29),
	.w8(32'h3ab56606),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac74aa),
	.w1(32'h3b19b8fd),
	.w2(32'h3c2b57b5),
	.w3(32'hbba17817),
	.w4(32'h3a801c70),
	.w5(32'h3c1bfe96),
	.w6(32'hb95e5b3d),
	.w7(32'hb98af2b7),
	.w8(32'hbb184fd9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ab9ec),
	.w1(32'h3bec363d),
	.w2(32'h3c502b90),
	.w3(32'hbc843b9b),
	.w4(32'hbbb05194),
	.w5(32'h3c3d1ff9),
	.w6(32'hb9a313cb),
	.w7(32'hbc45e3e2),
	.w8(32'hbbfae69f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d9097),
	.w1(32'hbc545cd2),
	.w2(32'hbbe03810),
	.w3(32'hbc29c7d5),
	.w4(32'hbc7095dd),
	.w5(32'hb8cfe712),
	.w6(32'hbb3b5030),
	.w7(32'hbbbab087),
	.w8(32'h3c46f18d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c1410),
	.w1(32'hbc5ac215),
	.w2(32'hbbc81057),
	.w3(32'h3b76f7cd),
	.w4(32'h3b9413a1),
	.w5(32'h3ca34d2d),
	.w6(32'hbc17cab3),
	.w7(32'hbb08c81d),
	.w8(32'hbbb0cb70),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99a330),
	.w1(32'hbc8d0c59),
	.w2(32'h3bd97fc1),
	.w3(32'hbbffdca6),
	.w4(32'hbc2dfdc4),
	.w5(32'h3b26302d),
	.w6(32'hbb6f2825),
	.w7(32'hbbd832c9),
	.w8(32'hb68786a4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93e675),
	.w1(32'h375bfee0),
	.w2(32'h3b6bd112),
	.w3(32'hba2de2ce),
	.w4(32'hbb96e800),
	.w5(32'hba98428a),
	.w6(32'hba0092da),
	.w7(32'h3b8c5522),
	.w8(32'hba392131),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80a9e1),
	.w1(32'h3ad71a83),
	.w2(32'h3918e8d6),
	.w3(32'hbc47731e),
	.w4(32'hbbdcc898),
	.w5(32'h3b07fe1f),
	.w6(32'hbb3132f1),
	.w7(32'hbc42eb5f),
	.w8(32'hbbd03bc5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61bafe),
	.w1(32'hbbae0ee4),
	.w2(32'hbc9df796),
	.w3(32'h3bc1ed38),
	.w4(32'hbbcd7743),
	.w5(32'hbcac011d),
	.w6(32'h3c49a268),
	.w7(32'h3b6b9868),
	.w8(32'hbc661dbe),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1177c1),
	.w1(32'h3c9be73c),
	.w2(32'h3cb9dc93),
	.w3(32'hbccf8a7e),
	.w4(32'hba30ea6a),
	.w5(32'h3cab0b71),
	.w6(32'hbc5d9390),
	.w7(32'hbceb1220),
	.w8(32'h3c65563d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bca15),
	.w1(32'hbc8b7f1c),
	.w2(32'h3b8952af),
	.w3(32'hbc8fa926),
	.w4(32'hbcc0546c),
	.w5(32'hbb9fcc9b),
	.w6(32'hbcd34374),
	.w7(32'hbba881fd),
	.w8(32'hbbf32590),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf52792),
	.w1(32'hbb83abdc),
	.w2(32'h3ba7f671),
	.w3(32'hbc0a2f2e),
	.w4(32'hbc05b84e),
	.w5(32'hbb8fb122),
	.w6(32'hbbb9147a),
	.w7(32'h3b4d384a),
	.w8(32'h3c437f03),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01bd8a),
	.w1(32'hbc4e33e7),
	.w2(32'h3c54e498),
	.w3(32'hbbd934d1),
	.w4(32'hbc3fbda3),
	.w5(32'h3c694210),
	.w6(32'hbc321353),
	.w7(32'h3c389e48),
	.w8(32'h3bb959a6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd74b35),
	.w1(32'hbd060306),
	.w2(32'h3b5d89dc),
	.w3(32'hbc91d28a),
	.w4(32'hbd01f9c8),
	.w5(32'hbbb5ffa5),
	.w6(32'hbc2e5641),
	.w7(32'hbca8ccf0),
	.w8(32'h3ac227ce),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d4aee),
	.w1(32'hbc4d1dbb),
	.w2(32'hbad3f634),
	.w3(32'hba8ea0d2),
	.w4(32'hbc60a84d),
	.w5(32'h3bbf95c1),
	.w6(32'hb975607b),
	.w7(32'h3be9a309),
	.w8(32'h3b649ee7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9756f4),
	.w1(32'h3ba4fef6),
	.w2(32'h3d17911e),
	.w3(32'hbc28259c),
	.w4(32'hbbe0512c),
	.w5(32'h3c70a4a2),
	.w6(32'hbb379bee),
	.w7(32'h3ca13ebb),
	.w8(32'h3c408ff6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0747fa),
	.w1(32'h3b130c6b),
	.w2(32'h3c0544a6),
	.w3(32'hbb5ea42b),
	.w4(32'hbb105197),
	.w5(32'h3bac86fe),
	.w6(32'h3b1ca1d7),
	.w7(32'h39853667),
	.w8(32'h3a8f3a05),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1a648),
	.w1(32'hbbba2e5f),
	.w2(32'hbb9a229c),
	.w3(32'hbc06d52b),
	.w4(32'hbbdc2fde),
	.w5(32'hbb96e98b),
	.w6(32'hbc07c6d0),
	.w7(32'hba242985),
	.w8(32'h3baabf19),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd88eee),
	.w1(32'hbcd4cef9),
	.w2(32'hbc8ce72a),
	.w3(32'hbbedabf0),
	.w4(32'hbc8d0e0d),
	.w5(32'h3c82071f),
	.w6(32'hbc40ed9e),
	.w7(32'hbbe9c8b4),
	.w8(32'hbc183b6c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc894f0a),
	.w1(32'hbc92ec53),
	.w2(32'hbc319407),
	.w3(32'hbc272046),
	.w4(32'hbbf92aed),
	.w5(32'hbb6b9301),
	.w6(32'hbc50a4fa),
	.w7(32'hbc16bf36),
	.w8(32'h3a76fb2a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11f123),
	.w1(32'h3c07f4da),
	.w2(32'h3c236a72),
	.w3(32'hbc742f7b),
	.w4(32'hbc39de00),
	.w5(32'hbbc47ab2),
	.w6(32'hba9a85f9),
	.w7(32'hbba58d15),
	.w8(32'hbbfdcf98),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbec3e6),
	.w1(32'hbc521041),
	.w2(32'hbbf9d76d),
	.w3(32'h3ba265ed),
	.w4(32'h3a9bb252),
	.w5(32'hbbb95404),
	.w6(32'hbb0cf000),
	.w7(32'h3cb7d61c),
	.w8(32'h3bde0f31),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a84589),
	.w1(32'hba5d69c2),
	.w2(32'hba53f81f),
	.w3(32'h3b0c8241),
	.w4(32'h3a654164),
	.w5(32'h3af13e04),
	.w6(32'h3a4cbc71),
	.w7(32'h399df021),
	.w8(32'h3aa253db),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29fc08),
	.w1(32'h3bcd7fa0),
	.w2(32'h3c5ace65),
	.w3(32'hb93e3696),
	.w4(32'h3b2c9aa2),
	.w5(32'h3bf6f0ac),
	.w6(32'h3b79260e),
	.w7(32'h3b3ee042),
	.w8(32'h3915e4b9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3498cd),
	.w1(32'h3ab78438),
	.w2(32'hbb3debdf),
	.w3(32'hba9c1f60),
	.w4(32'hba530537),
	.w5(32'hbb3f8a62),
	.w6(32'h3b7ad3ca),
	.w7(32'h3b002eb6),
	.w8(32'hbbc1df44),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77645c),
	.w1(32'hbc89f100),
	.w2(32'hbc01614a),
	.w3(32'h3b18f407),
	.w4(32'hbb1b696c),
	.w5(32'h3a661cf9),
	.w6(32'hbb419e94),
	.w7(32'hbb50dfd2),
	.w8(32'hbc1253f3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc3c13),
	.w1(32'h3b1edc23),
	.w2(32'hb62975c0),
	.w3(32'hbab22261),
	.w4(32'h3b038898),
	.w5(32'h3ab20d42),
	.w6(32'hba32a630),
	.w7(32'hbb0ceec6),
	.w8(32'hb923bbed),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc933d76),
	.w1(32'h3b53a827),
	.w2(32'h3c8f230b),
	.w3(32'hbc965854),
	.w4(32'h3b0cd519),
	.w5(32'h3ca482d5),
	.w6(32'h3c38a74b),
	.w7(32'hbbb230fd),
	.w8(32'hbb29def3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c703b),
	.w1(32'h3b85b98f),
	.w2(32'h3bbf2020),
	.w3(32'h3b987b1b),
	.w4(32'h3bad61f2),
	.w5(32'h3baa0fb6),
	.w6(32'h3bc70a67),
	.w7(32'h3ba242cd),
	.w8(32'hbada4b20),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb414fa9),
	.w1(32'h3b5dbe44),
	.w2(32'h3b75f569),
	.w3(32'hbbbe4e28),
	.w4(32'hba1fd083),
	.w5(32'h3aec68a4),
	.w6(32'h3ab28409),
	.w7(32'h3b7d9e66),
	.w8(32'h3c374924),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6e088),
	.w1(32'h3bf42185),
	.w2(32'h3c1d7c8b),
	.w3(32'h3bac57f8),
	.w4(32'h3be23483),
	.w5(32'h3c0c7b05),
	.w6(32'h3bde8112),
	.w7(32'h3bd681a8),
	.w8(32'hbc3fba97),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb38af7),
	.w1(32'hbcc2cb77),
	.w2(32'hbb96ee52),
	.w3(32'h3b445e4c),
	.w4(32'h3be20146),
	.w5(32'h3b0185ae),
	.w6(32'hbb748234),
	.w7(32'h3c883c44),
	.w8(32'hbbdfa88d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcde420),
	.w1(32'hbb98336a),
	.w2(32'hbb3351df),
	.w3(32'hbb418643),
	.w4(32'hbad41259),
	.w5(32'hba8448a4),
	.w6(32'hbb594f3d),
	.w7(32'hb90e7dca),
	.w8(32'h3b230486),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba832d85),
	.w1(32'h3abe96be),
	.w2(32'h3b82276d),
	.w3(32'hbb983caf),
	.w4(32'hbb43e514),
	.w5(32'h3baed1ff),
	.w6(32'hbb7ce604),
	.w7(32'hbbca0ac9),
	.w8(32'hbb81df75),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45de45),
	.w1(32'hbb2d3c09),
	.w2(32'h3a22919d),
	.w3(32'hb813275b),
	.w4(32'h3ac219a7),
	.w5(32'h3b028c66),
	.w6(32'hbaeeaf8b),
	.w7(32'h3a087160),
	.w8(32'h3a07e214),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e2aa6),
	.w1(32'h3c080968),
	.w2(32'h3c9965b8),
	.w3(32'hbc818dba),
	.w4(32'hbb46b228),
	.w5(32'h3c0cb16c),
	.w6(32'h394bb176),
	.w7(32'hbc26dd99),
	.w8(32'hbbf9fdb4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5b92d),
	.w1(32'h3b25a98a),
	.w2(32'h3c3f1504),
	.w3(32'hbc021073),
	.w4(32'hbb4e8fbc),
	.w5(32'h3abf9d40),
	.w6(32'hb9a4ee9b),
	.w7(32'hbbb6bab0),
	.w8(32'h3886ba6c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba374e34),
	.w1(32'hba560a53),
	.w2(32'h3b48dbed),
	.w3(32'h3b585344),
	.w4(32'h3b3cfb15),
	.w5(32'h3b6bfb77),
	.w6(32'hbacb9091),
	.w7(32'h3b81c05b),
	.w8(32'h3be04298),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3458c3),
	.w1(32'hbc2fb8e8),
	.w2(32'hbc5fe819),
	.w3(32'h3bf42025),
	.w4(32'h3bbacca9),
	.w5(32'h3c0c0fe8),
	.w6(32'h3bee3e29),
	.w7(32'hba454953),
	.w8(32'hbad94eea),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c8bf1),
	.w1(32'h39ec8ed4),
	.w2(32'hbb3d34d6),
	.w3(32'hbc1d3e81),
	.w4(32'hbac3c1e8),
	.w5(32'h3b750a19),
	.w6(32'hbbc62ae5),
	.w7(32'hbbdcbebd),
	.w8(32'hbc5d4e49),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdcce2e),
	.w1(32'hbc426c32),
	.w2(32'hb8987fd9),
	.w3(32'hbcd08bdb),
	.w4(32'hbc91fa66),
	.w5(32'hbab1e9ef),
	.w6(32'hbc8fa1dd),
	.w7(32'hbc85ee2d),
	.w8(32'h3cf26a38),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac5b1d),
	.w1(32'hbca8d9d4),
	.w2(32'hbce8981b),
	.w3(32'hbce3d4a0),
	.w4(32'hbcf4867b),
	.w5(32'hbc8c2f39),
	.w6(32'hbd186146),
	.w7(32'hbcd7d4e7),
	.w8(32'hbcb1afa8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb65765),
	.w1(32'hbba41e38),
	.w2(32'h3c7878d8),
	.w3(32'hbd0d682e),
	.w4(32'hbcc49034),
	.w5(32'h3b9694a7),
	.w6(32'hbb972e7d),
	.w7(32'hbc73a340),
	.w8(32'hbc305061),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ce281),
	.w1(32'h39b82388),
	.w2(32'hbb3dd7b1),
	.w3(32'hbcd8b425),
	.w4(32'hbc2655ab),
	.w5(32'h3a55cbeb),
	.w6(32'hbc6b86b4),
	.w7(32'hbca7b960),
	.w8(32'h3bfffbbe),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b253b98),
	.w1(32'hbc07041f),
	.w2(32'hbb31eb27),
	.w3(32'hbb084856),
	.w4(32'hbc2a43a5),
	.w5(32'hbba749e7),
	.w6(32'hbadf86c3),
	.w7(32'h3b0b97d3),
	.w8(32'h3c0503f0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8353da),
	.w1(32'hbb680d75),
	.w2(32'h39b9d6bf),
	.w3(32'h3b3c6271),
	.w4(32'hbb14898e),
	.w5(32'h3b90665c),
	.w6(32'h3aaeae56),
	.w7(32'hbabb24e7),
	.w8(32'hba64ee29),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaed488),
	.w1(32'hbbb79e12),
	.w2(32'hbabe5d0f),
	.w3(32'hbbcda37d),
	.w4(32'hbb91dcae),
	.w5(32'h39ba4d9b),
	.w6(32'hbb6bbdac),
	.w7(32'hba462123),
	.w8(32'h3b57eee8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a9cea),
	.w1(32'hbc17747b),
	.w2(32'hbb4558e7),
	.w3(32'hbbc73666),
	.w4(32'hbc43203f),
	.w5(32'hbbaead48),
	.w6(32'hbb19c0eb),
	.w7(32'h399289fa),
	.w8(32'h3b7f5626),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6265f2),
	.w1(32'hbbf71b5f),
	.w2(32'hbbc42f5c),
	.w3(32'hbbf7755c),
	.w4(32'hbc61d74e),
	.w5(32'hbbe3303d),
	.w6(32'hbb4ec6fc),
	.w7(32'h3a54c355),
	.w8(32'hbb89f36c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f1c48),
	.w1(32'hbab4d63c),
	.w2(32'hba66d747),
	.w3(32'hbb4eb044),
	.w4(32'hbac96b2a),
	.w5(32'hba87e7f2),
	.w6(32'hbabb16c6),
	.w7(32'hb9b8c734),
	.w8(32'h3c98c525),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a2214),
	.w1(32'hbc438fa7),
	.w2(32'hbb9b4f11),
	.w3(32'h3c33b8a0),
	.w4(32'h3969836c),
	.w5(32'hbbc4e029),
	.w6(32'hbc55c26e),
	.w7(32'h3b5a37c3),
	.w8(32'h3ab363a6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71c7b03),
	.w1(32'h3bb361d6),
	.w2(32'h3be59c9c),
	.w3(32'hbb2c3db5),
	.w4(32'h3922d412),
	.w5(32'h3b2d0831),
	.w6(32'h3ac549c5),
	.w7(32'h3a0cd6cd),
	.w8(32'h3ca1ead0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2069a6),
	.w1(32'hbc8528b7),
	.w2(32'hbc2c0712),
	.w3(32'hbb35c461),
	.w4(32'hbc1d1877),
	.w5(32'hbbace414),
	.w6(32'h3ca83ccb),
	.w7(32'h3c67f2ce),
	.w8(32'hbbb85ced),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb867a7e),
	.w1(32'hba86e343),
	.w2(32'h3b894eb1),
	.w3(32'hbb89a320),
	.w4(32'hbb9627a0),
	.w5(32'hbacd84a2),
	.w6(32'hba4b0a17),
	.w7(32'hba007b78),
	.w8(32'h3ca09b33),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc018ca7),
	.w1(32'hbca20cb0),
	.w2(32'h3982c037),
	.w3(32'hbc47c717),
	.w4(32'hbc64d47a),
	.w5(32'hbba2b8fe),
	.w6(32'hbb8a8ed9),
	.w7(32'hbbf285f0),
	.w8(32'h3c05881a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc709eda),
	.w1(32'hbc937d66),
	.w2(32'hbc502f87),
	.w3(32'hbb469e3b),
	.w4(32'h39077629),
	.w5(32'h3ae465d9),
	.w6(32'hbabd1ecb),
	.w7(32'h3b17008d),
	.w8(32'h39ec3c2f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c3189),
	.w1(32'h3c14309a),
	.w2(32'h3bc8a244),
	.w3(32'hbb1d7954),
	.w4(32'h3b20366b),
	.w5(32'hba953e58),
	.w6(32'h3b5145f5),
	.w7(32'hbad6ea67),
	.w8(32'h3a8ddfd4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae78c2b),
	.w1(32'hbb212128),
	.w2(32'h3b5776a4),
	.w3(32'hba870398),
	.w4(32'hb9bee701),
	.w5(32'h3ba30f6e),
	.w6(32'hba1c0ddd),
	.w7(32'h399aa34b),
	.w8(32'hbb51e9eb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00d0c3),
	.w1(32'hbc0385d3),
	.w2(32'hba5770f0),
	.w3(32'hbbf3a232),
	.w4(32'hbbfa56d3),
	.w5(32'h3adb0e6a),
	.w6(32'hbbf71e9c),
	.w7(32'h3a243105),
	.w8(32'h3823fdd1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d01e4),
	.w1(32'h383191bd),
	.w2(32'hb8f63b2e),
	.w3(32'h38ac42ed),
	.w4(32'h3ac39978),
	.w5(32'h3b22b64e),
	.w6(32'h3b227d15),
	.w7(32'h39a91df1),
	.w8(32'h3978d037),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f8eb1),
	.w1(32'h3c6d1fa0),
	.w2(32'h3c111f98),
	.w3(32'hbab50aeb),
	.w4(32'h3c1260f9),
	.w5(32'h3a17aeee),
	.w6(32'h3c09b374),
	.w7(32'hbb16ad5e),
	.w8(32'hbb827bba),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d6d98),
	.w1(32'hb88dae2f),
	.w2(32'hbac7b4a6),
	.w3(32'hbbcac8ad),
	.w4(32'h3bbf99ea),
	.w5(32'h3b2c5743),
	.w6(32'hba612c36),
	.w7(32'h3c04b4b0),
	.w8(32'h3bffda24),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82661e),
	.w1(32'h380dbd79),
	.w2(32'h39d4119e),
	.w3(32'h3ba73e51),
	.w4(32'h3b09e400),
	.w5(32'h3a4c2250),
	.w6(32'h3b00af1a),
	.w7(32'h3ba401c7),
	.w8(32'h3bc27a07),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb89888),
	.w1(32'h3bce3b7c),
	.w2(32'h3c870b70),
	.w3(32'hbc40e56c),
	.w4(32'hbb8b215c),
	.w5(32'h3c5dba6e),
	.w6(32'h3bdacc6a),
	.w7(32'hbb7e7024),
	.w8(32'h3add2e03),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa16f2e),
	.w1(32'hbb395de2),
	.w2(32'h3bef8bdf),
	.w3(32'h3aa2b341),
	.w4(32'hbb38e149),
	.w5(32'h3b9d5125),
	.w6(32'h382dbdad),
	.w7(32'h3b871b70),
	.w8(32'h399b8c05),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf0d1c),
	.w1(32'h3ba16473),
	.w2(32'h3b1af59d),
	.w3(32'h3a59bd55),
	.w4(32'h3b9793f5),
	.w5(32'h3a54de3a),
	.w6(32'h3bc37836),
	.w7(32'h3bed5330),
	.w8(32'h3bf3bfe3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c042b75),
	.w1(32'h3c15fc51),
	.w2(32'h3bd67fdb),
	.w3(32'h3bc27592),
	.w4(32'h3c037dac),
	.w5(32'h3baceae8),
	.w6(32'h3bab50fc),
	.w7(32'h3c09f429),
	.w8(32'h3a7940c8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41f264),
	.w1(32'hbab45605),
	.w2(32'hba08eeef),
	.w3(32'hbb96db54),
	.w4(32'hbbc1354c),
	.w5(32'hbb850b6b),
	.w6(32'h39c117fe),
	.w7(32'h3afa31c0),
	.w8(32'hbb048f0d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a059d47),
	.w1(32'hb8bc7702),
	.w2(32'h3a51439d),
	.w3(32'h3b6d86f4),
	.w4(32'hba8087f1),
	.w5(32'hbc0101f1),
	.w6(32'h3a328a96),
	.w7(32'h3b4a2664),
	.w8(32'hbb37d178),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad40f62),
	.w1(32'h3bc66cdf),
	.w2(32'hbb02c78d),
	.w3(32'hbbb0c3b4),
	.w4(32'hb72b656a),
	.w5(32'hba8e441f),
	.w6(32'h390f05cb),
	.w7(32'hbbdf35cb),
	.w8(32'hbbe60787),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bf137),
	.w1(32'h3b68d80f),
	.w2(32'hb88fe505),
	.w3(32'h3bee54ec),
	.w4(32'h3bc1a90e),
	.w5(32'h3b97d6ce),
	.w6(32'h3ab96009),
	.w7(32'h3b188ab6),
	.w8(32'h3be4a12b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24373b),
	.w1(32'h3b93cfc7),
	.w2(32'h3b260699),
	.w3(32'hbaa4ea76),
	.w4(32'h3aa86f90),
	.w5(32'hb9b01e44),
	.w6(32'h3b1bbf7a),
	.w7(32'h3b623273),
	.w8(32'hbac7a2ab),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a6709),
	.w1(32'hbb70f91a),
	.w2(32'hbb8e06e6),
	.w3(32'hbbab22df),
	.w4(32'hbba313e4),
	.w5(32'hbb94b62c),
	.w6(32'hbbb03340),
	.w7(32'hbba28427),
	.w8(32'hbb51e609),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69be10),
	.w1(32'hbaefc126),
	.w2(32'hbb37bd09),
	.w3(32'hbbba0d2f),
	.w4(32'hbb94cb90),
	.w5(32'hbb577891),
	.w6(32'h39dac664),
	.w7(32'hbafab874),
	.w8(32'h3b01ca84),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc05db1),
	.w1(32'h3aff4774),
	.w2(32'h3bd31f79),
	.w3(32'h3aebf52b),
	.w4(32'hba4dedda),
	.w5(32'h3b074bda),
	.w6(32'h3bb9a016),
	.w7(32'h3c074d96),
	.w8(32'hb9da2d3c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b8414),
	.w1(32'h3a582a4a),
	.w2(32'h3aecff4d),
	.w3(32'hbc19dc47),
	.w4(32'hbbf495dd),
	.w5(32'hbb0dd8b2),
	.w6(32'hbbdc30c7),
	.w7(32'hbc0d3ddd),
	.w8(32'hbc0d763b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33c428),
	.w1(32'h37e5c8a0),
	.w2(32'h3ad25086),
	.w3(32'hbae54423),
	.w4(32'h39e62299),
	.w5(32'hbb3a8082),
	.w6(32'hba8671e1),
	.w7(32'h3a3ec553),
	.w8(32'hbbcc2ebf),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf16b20),
	.w1(32'hbba19153),
	.w2(32'h3aa692fa),
	.w3(32'hbb86343f),
	.w4(32'hba95b079),
	.w5(32'h3ad76e85),
	.w6(32'hbbaee56c),
	.w7(32'h3a27f0bb),
	.w8(32'hbb5bb911),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a8d2f),
	.w1(32'hbb733546),
	.w2(32'hbb52901d),
	.w3(32'hbbe8751b),
	.w4(32'hbbd500f8),
	.w5(32'hbbfb6ffc),
	.w6(32'h3ad59a14),
	.w7(32'h3c56d983),
	.w8(32'h3c57cd3b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaea3ce),
	.w1(32'hba9f75a5),
	.w2(32'h3bd57309),
	.w3(32'hbbab8788),
	.w4(32'hbb4ed081),
	.w5(32'h3b10b6c6),
	.w6(32'hbc1f9de2),
	.w7(32'hbc4194bd),
	.w8(32'hb9a48ea5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b794d),
	.w1(32'h3b2b3efd),
	.w2(32'h3b0fe3e7),
	.w3(32'h3b46ba75),
	.w4(32'h3a8a3aaf),
	.w5(32'h39ed8eee),
	.w6(32'h3b693e09),
	.w7(32'h3b6676af),
	.w8(32'hbaee6c17),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b9aba),
	.w1(32'hba3f99f3),
	.w2(32'h3aa249a6),
	.w3(32'h3b293e99),
	.w4(32'h3b0835d6),
	.w5(32'h3b576c77),
	.w6(32'hbb05b82a),
	.w7(32'h3b0a890b),
	.w8(32'h3bce526c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24943b),
	.w1(32'hbbaec165),
	.w2(32'hbb6bd49a),
	.w3(32'h3b7b52a1),
	.w4(32'hba4561a9),
	.w5(32'hba98e22b),
	.w6(32'h3ab09ace),
	.w7(32'h3b1d31cf),
	.w8(32'hbb9b02a3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7bcf3),
	.w1(32'h392a19fd),
	.w2(32'hbb9df2e0),
	.w3(32'hbb9e3581),
	.w4(32'hbbaa92ae),
	.w5(32'hbc17625d),
	.w6(32'hba85d03b),
	.w7(32'hbab43028),
	.w8(32'h3c4962f5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cb372),
	.w1(32'h3c4fe8b0),
	.w2(32'h3c9c3703),
	.w3(32'h3c2b2848),
	.w4(32'h3c154899),
	.w5(32'h3c521183),
	.w6(32'h3c843680),
	.w7(32'h3c90e4b5),
	.w8(32'h3a5a4234),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b433bcb),
	.w1(32'hbbb133c5),
	.w2(32'h3b79988d),
	.w3(32'h3b7f47bc),
	.w4(32'h399ef51b),
	.w5(32'h3b728e82),
	.w6(32'h3b9a50bf),
	.w7(32'hba6bf813),
	.w8(32'h3a6607ce),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule