module layer_10_featuremap_236(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4e7db),
	.w1(32'hbad911a3),
	.w2(32'hb8808635),
	.w3(32'hbab60d98),
	.w4(32'hba56ab2d),
	.w5(32'h3b21886e),
	.w6(32'hbaf49027),
	.w7(32'hbac132dd),
	.w8(32'hb9e30ce3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba020c51),
	.w1(32'h39e6b43b),
	.w2(32'hba080c2d),
	.w3(32'hba0225eb),
	.w4(32'hba042b5e),
	.w5(32'hbb3767dd),
	.w6(32'h3a0ad454),
	.w7(32'hba6bcfbf),
	.w8(32'hbb88cd58),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378ef641),
	.w1(32'h3a813803),
	.w2(32'h39d991b6),
	.w3(32'hbaea4611),
	.w4(32'hbab33bc6),
	.w5(32'hb914c102),
	.w6(32'h3acca4e1),
	.w7(32'h3a8acec5),
	.w8(32'h38f7ed02),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4e139),
	.w1(32'h3a55602d),
	.w2(32'h3a08ffdc),
	.w3(32'hba083d07),
	.w4(32'hb8c5df72),
	.w5(32'hba2b8995),
	.w6(32'h398d1043),
	.w7(32'h3a407d3f),
	.w8(32'hb9f54b6c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa63d9),
	.w1(32'hbb2830c7),
	.w2(32'hbac3c98e),
	.w3(32'hbaf8c0f0),
	.w4(32'hba9c3f2d),
	.w5(32'hbb2152d1),
	.w6(32'hba689401),
	.w7(32'hbaa4d8b7),
	.w8(32'hbae99614),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7dca8),
	.w1(32'hba13dcde),
	.w2(32'hb9d50865),
	.w3(32'hbab300aa),
	.w4(32'hbab2ae89),
	.w5(32'hba8ca6d4),
	.w6(32'h36ddce4e),
	.w7(32'hb9f5c58e),
	.w8(32'hbac14153),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd94f2),
	.w1(32'hbb91ed4b),
	.w2(32'hbbbd8c05),
	.w3(32'h3993f4a9),
	.w4(32'hbba642ef),
	.w5(32'hbbe17c15),
	.w6(32'h3b0e9b70),
	.w7(32'hbb334aff),
	.w8(32'hbb8bf960),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc446fae),
	.w1(32'hbc26bf40),
	.w2(32'hbbf8deec),
	.w3(32'hbc1427b8),
	.w4(32'hbbaedddd),
	.w5(32'hba9deec3),
	.w6(32'hbc0555a9),
	.w7(32'hbb41045d),
	.w8(32'hbb69b43c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca8060),
	.w1(32'hba50425c),
	.w2(32'hba9ef5af),
	.w3(32'hba9b6344),
	.w4(32'hba5580dc),
	.w5(32'hbb12cecd),
	.w6(32'hbac1e604),
	.w7(32'hba922abb),
	.w8(32'hbade6408),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb660ed0),
	.w1(32'hbb94388c),
	.w2(32'hbc191421),
	.w3(32'hbb27c8df),
	.w4(32'hbb77aa4b),
	.w5(32'hbbdc0ce6),
	.w6(32'hb9fc9a57),
	.w7(32'hbb0f4128),
	.w8(32'hbbc55293),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b1fac),
	.w1(32'hb9ce3266),
	.w2(32'hba583e24),
	.w3(32'h391a2512),
	.w4(32'hb91dcf7d),
	.w5(32'h3a6e565a),
	.w6(32'h3b034dfc),
	.w7(32'h3acfbb6d),
	.w8(32'hbac5c0f3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfc4f4),
	.w1(32'h39b677a3),
	.w2(32'hbb23ae51),
	.w3(32'h3b3ad465),
	.w4(32'hb9c09d88),
	.w5(32'hbb848cc8),
	.w6(32'h3ac67478),
	.w7(32'h3a9a946b),
	.w8(32'hbb0a18d8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb144d45),
	.w1(32'hbb9a97e0),
	.w2(32'hbbe3b969),
	.w3(32'h3a6c61bb),
	.w4(32'hba25eca1),
	.w5(32'hbbbf35fb),
	.w6(32'hbb0c635d),
	.w7(32'hbb38dd17),
	.w8(32'hbbb05d35),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb069a5b),
	.w1(32'hbbcdc06e),
	.w2(32'hbbf36a8b),
	.w3(32'hba580453),
	.w4(32'hbabb955f),
	.w5(32'hbb6d7e1f),
	.w6(32'hb870f58e),
	.w7(32'hbad7505a),
	.w8(32'hbb475068),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a7e8e),
	.w1(32'hb904ab29),
	.w2(32'hbb049d0c),
	.w3(32'hb8d89de0),
	.w4(32'h3b09447a),
	.w5(32'hbb06e13f),
	.w6(32'hb9617f6a),
	.w7(32'hba6aac09),
	.w8(32'hbb685df5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd59ef8),
	.w1(32'hbc13298f),
	.w2(32'hbc23a462),
	.w3(32'hbbe43eba),
	.w4(32'hbb97f06a),
	.w5(32'hbbf4d6e7),
	.w6(32'hbbc64848),
	.w7(32'hbb7a1723),
	.w8(32'hbbdf3580),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d0e61),
	.w1(32'hbb0b32bc),
	.w2(32'hbb0f0ded),
	.w3(32'hbb12fa4d),
	.w4(32'hbacc724c),
	.w5(32'hba90aad5),
	.w6(32'hb938154b),
	.w7(32'hbabc5dcd),
	.w8(32'h388a5d6c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cb5b4),
	.w1(32'hbbe1c0d7),
	.w2(32'hbbdf1da2),
	.w3(32'hbb912c4f),
	.w4(32'hbb7f0e20),
	.w5(32'hbba5f43b),
	.w6(32'hbb49c05e),
	.w7(32'h397f1297),
	.w8(32'h3ad3723d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb683dac),
	.w1(32'hbb7278dc),
	.w2(32'hbb70fc5f),
	.w3(32'hbb3cac43),
	.w4(32'hbb28230a),
	.w5(32'hbb494657),
	.w6(32'h39ee803c),
	.w7(32'hb9f60f1b),
	.w8(32'hbb1c5fa1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7c1b0),
	.w1(32'hb93c1f16),
	.w2(32'hba5b1457),
	.w3(32'h39c52177),
	.w4(32'h394634ec),
	.w5(32'hbad88bf2),
	.w6(32'hb9669032),
	.w7(32'h3865a4a6),
	.w8(32'hbabd9808),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac128e),
	.w1(32'hbb0505e1),
	.w2(32'hba4d39d3),
	.w3(32'hbb1eaadd),
	.w4(32'hba240662),
	.w5(32'hb9102710),
	.w6(32'hbadc3b18),
	.w7(32'h3953a168),
	.w8(32'h3a16a709),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a310005),
	.w1(32'h3a11245e),
	.w2(32'hb9aa9be0),
	.w3(32'hb967bc3d),
	.w4(32'h3aad9526),
	.w5(32'h3ab4ec79),
	.w6(32'hba982c37),
	.w7(32'h3ac45de6),
	.w8(32'h39752218),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02ca3a),
	.w1(32'hbba4dfd7),
	.w2(32'hbbd61046),
	.w3(32'hbb2fc3e2),
	.w4(32'h3a99c183),
	.w5(32'hbbc8534c),
	.w6(32'hbacfced0),
	.w7(32'hbab131c9),
	.w8(32'hbbaeb5fe),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24b290),
	.w1(32'hbb4e79ac),
	.w2(32'hbc189ffc),
	.w3(32'h39f92b7f),
	.w4(32'h37eed3b9),
	.w5(32'hbb87d6ae),
	.w6(32'hba08883a),
	.w7(32'hbae2ddb5),
	.w8(32'hbbb82616),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50f272),
	.w1(32'h39adb32a),
	.w2(32'hbb253dae),
	.w3(32'hbb31a3b4),
	.w4(32'h3a9f5a79),
	.w5(32'hbb2756a4),
	.w6(32'hbb008498),
	.w7(32'hbabaaa0c),
	.w8(32'hbc052ad6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6aedd),
	.w1(32'hbad7a45a),
	.w2(32'hbab67c91),
	.w3(32'hba64ba42),
	.w4(32'hbaa3de4b),
	.w5(32'hbb00cfa0),
	.w6(32'h3aaa2c0c),
	.w7(32'hba087851),
	.w8(32'hbae3aacf),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63652a),
	.w1(32'hbb1d2dfb),
	.w2(32'hbab1b332),
	.w3(32'hbb7b74d0),
	.w4(32'hbaa24b6a),
	.w5(32'hbb381ea0),
	.w6(32'hbb1cb003),
	.w7(32'hbaf1731b),
	.w8(32'hbb3c638d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f70c8),
	.w1(32'hbb53dc83),
	.w2(32'hbb036819),
	.w3(32'hbb93a256),
	.w4(32'hbbb7ce7f),
	.w5(32'hbb93bdfe),
	.w6(32'hbb065261),
	.w7(32'hba8a90af),
	.w8(32'h3a880907),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381f4f6a),
	.w1(32'h3acad0c3),
	.w2(32'h3b13633f),
	.w3(32'h39419b1a),
	.w4(32'h3ad89441),
	.w5(32'hba57866b),
	.w6(32'h3a2df27c),
	.w7(32'h3ade9ea5),
	.w8(32'hbaf2fe8d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b285a6c),
	.w1(32'hb95ec8cb),
	.w2(32'hbb0f65c0),
	.w3(32'hb99ec053),
	.w4(32'hbba1ca38),
	.w5(32'hbb90f555),
	.w6(32'h3a000a06),
	.w7(32'hbba5bae4),
	.w8(32'hbba9a3e5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea12cb),
	.w1(32'h3aab5c64),
	.w2(32'h3a8e2142),
	.w3(32'h3b372013),
	.w4(32'h3aa2b4ab),
	.w5(32'h3af10bde),
	.w6(32'h3b8f79d0),
	.w7(32'h3b21d567),
	.w8(32'h3b35c8f9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f9b72),
	.w1(32'h3ae7a378),
	.w2(32'h3a887256),
	.w3(32'h3b0712cb),
	.w4(32'h3a13c6bb),
	.w5(32'hbaf26f50),
	.w6(32'h3b4a9c72),
	.w7(32'h3a2e49c5),
	.w8(32'hb9ef1bec),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd4778),
	.w1(32'hbb75ec77),
	.w2(32'hbb9c42fc),
	.w3(32'h3a2af366),
	.w4(32'hba56b992),
	.w5(32'hbb9f946d),
	.w6(32'h3a09435e),
	.w7(32'hbb1555c9),
	.w8(32'hbb8dc479),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f2146),
	.w1(32'hbaea3fd6),
	.w2(32'hbb7ec3bf),
	.w3(32'hbb402f78),
	.w4(32'hbb422121),
	.w5(32'hb8b64579),
	.w6(32'hbabb601b),
	.w7(32'hbb748eed),
	.w8(32'hbb19ed81),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38468a33),
	.w1(32'hb9e802b2),
	.w2(32'h399c2748),
	.w3(32'h3a9bac91),
	.w4(32'h3a8b7ad0),
	.w5(32'hb9d38db8),
	.w6(32'h3987001c),
	.w7(32'h3a83f2cc),
	.w8(32'h3b1bee46),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2f91c),
	.w1(32'hba32f99a),
	.w2(32'hbb324241),
	.w3(32'h39666656),
	.w4(32'hba793d3b),
	.w5(32'hbaa275bf),
	.w6(32'h3b4b309a),
	.w7(32'h384bf4fc),
	.w8(32'hba1151a3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2085ea),
	.w1(32'hbaf5e928),
	.w2(32'hbbd2a030),
	.w3(32'hbaad6ed6),
	.w4(32'h3aa755f7),
	.w5(32'hbb82013c),
	.w6(32'h3afaafb5),
	.w7(32'h3b9f6a63),
	.w8(32'hbb1cd31d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a665e7a),
	.w1(32'h3b92dfca),
	.w2(32'h3a86e616),
	.w3(32'hbb627789),
	.w4(32'h3ba63671),
	.w5(32'hba6d4d0d),
	.w6(32'hbb8f335a),
	.w7(32'h3b23ac36),
	.w8(32'hbbd37783),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff17e1),
	.w1(32'h3bc651a1),
	.w2(32'h3acbe0b2),
	.w3(32'h3a05e3c4),
	.w4(32'h3a989459),
	.w5(32'hbbc441d7),
	.w6(32'hbab31180),
	.w7(32'hb8a1e0a2),
	.w8(32'hbbb13cd1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcb45c),
	.w1(32'h3aea8e8d),
	.w2(32'h39afeb09),
	.w3(32'h399ab017),
	.w4(32'h3accf7fa),
	.w5(32'h3ae1a20f),
	.w6(32'hba7ac81c),
	.w7(32'h3a800f4c),
	.w8(32'hba754b54),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397438c9),
	.w1(32'h39c28b7e),
	.w2(32'h3af1ad05),
	.w3(32'hb89be52b),
	.w4(32'h3a392120),
	.w5(32'hba945207),
	.w6(32'hba57ab83),
	.w7(32'h3aa41d7c),
	.w8(32'hba94fa7b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc5a74),
	.w1(32'hbab0ab4c),
	.w2(32'hbaae84eb),
	.w3(32'hb97e9ce1),
	.w4(32'hba532d93),
	.w5(32'h3b0c37cd),
	.w6(32'h3a60976d),
	.w7(32'hb95aeea2),
	.w8(32'h3b3c18bc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa83e3),
	.w1(32'h3a97e555),
	.w2(32'h3b77cd3f),
	.w3(32'h3a8e3bb3),
	.w4(32'h3b44fec3),
	.w5(32'hb8a80639),
	.w6(32'h3ad59562),
	.w7(32'h3b67132f),
	.w8(32'hbb2e8016),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3562c),
	.w1(32'hbbc610be),
	.w2(32'hbc24eacf),
	.w3(32'hbbb841d5),
	.w4(32'hbb7c24d1),
	.w5(32'hbc2832b5),
	.w6(32'hbb2a9642),
	.w7(32'hbb83c51f),
	.w8(32'hbbd9b182),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac57f5),
	.w1(32'hbb8c387a),
	.w2(32'hbbe83c0d),
	.w3(32'hbb8fd728),
	.w4(32'hbb1ef5c1),
	.w5(32'hbbe8dda4),
	.w6(32'hbbc43b4e),
	.w7(32'hbb8c2a5a),
	.w8(32'hbc103c5e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe27b9d),
	.w1(32'hbb9aa208),
	.w2(32'hbc113dff),
	.w3(32'hbb295fd0),
	.w4(32'hbb1fe635),
	.w5(32'hbbc88782),
	.w6(32'hbb67f0d2),
	.w7(32'hbbb1e687),
	.w8(32'hbc189ff3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd119f5),
	.w1(32'hbbaa3793),
	.w2(32'hbbf1cacf),
	.w3(32'hbbdf351d),
	.w4(32'hbb80aa46),
	.w5(32'hba825079),
	.w6(32'hbb943619),
	.w7(32'hbb60cf70),
	.w8(32'hbb13b560),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cf8c4),
	.w1(32'hbb99e052),
	.w2(32'hbbb05928),
	.w3(32'hba9a395c),
	.w4(32'hbaacd91c),
	.w5(32'hbb2806c3),
	.w6(32'hbb08bd93),
	.w7(32'h39fd5070),
	.w8(32'hbab40df5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82f318),
	.w1(32'h3ab753b7),
	.w2(32'h3a140e29),
	.w3(32'h3af59710),
	.w4(32'h3a9612b5),
	.w5(32'h397f8e8e),
	.w6(32'hb7aa2a36),
	.w7(32'hb9751d02),
	.w8(32'h3a7841a3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e30ee),
	.w1(32'hba47b5e4),
	.w2(32'h3925f3e3),
	.w3(32'hba183b7a),
	.w4(32'hb9f1c9c3),
	.w5(32'hbb07988d),
	.w6(32'hba1bf9a8),
	.w7(32'hba0639f1),
	.w8(32'hbb1074da),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8554071),
	.w1(32'hb9ec4884),
	.w2(32'h398385e8),
	.w3(32'hbb3891a8),
	.w4(32'hba148642),
	.w5(32'hb88f44cb),
	.w6(32'hbaf4ca15),
	.w7(32'hb65272dd),
	.w8(32'h39ebe4ae),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0f737),
	.w1(32'hbb7e229a),
	.w2(32'hbb5c2131),
	.w3(32'hbb454bcf),
	.w4(32'hba9b0325),
	.w5(32'hba8fcbe3),
	.w6(32'h3a2eff02),
	.w7(32'hb924b47e),
	.w8(32'hbaebf5a5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada1dac),
	.w1(32'hba4c1502),
	.w2(32'hbb0f6361),
	.w3(32'hba773f1f),
	.w4(32'hba938634),
	.w5(32'hbb13ebbe),
	.w6(32'h392436db),
	.w7(32'hbaa92b8c),
	.w8(32'hbb07541b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc050309),
	.w1(32'hbc01f577),
	.w2(32'hbc2364a0),
	.w3(32'hbba42f58),
	.w4(32'hbb95d39f),
	.w5(32'hbbe05537),
	.w6(32'hbab1075d),
	.w7(32'hbacc4164),
	.w8(32'hbb3da051),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902d4c2),
	.w1(32'h39660e47),
	.w2(32'hbafca6a4),
	.w3(32'hb96dad12),
	.w4(32'hba552ff9),
	.w5(32'hbabd61fb),
	.w6(32'hba23c6d7),
	.w7(32'h3919d1bd),
	.w8(32'hbafcb09a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad97bc5),
	.w1(32'hbae75fae),
	.w2(32'hba24d9b3),
	.w3(32'hbab3e8a8),
	.w4(32'hba18dafe),
	.w5(32'h3a6f5e12),
	.w6(32'hba14911b),
	.w7(32'hb9d63de5),
	.w8(32'hb9fcc625),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28282d),
	.w1(32'hba1bbabe),
	.w2(32'h3a4a5ae5),
	.w3(32'hb995d2ac),
	.w4(32'h3aae9d1f),
	.w5(32'hba1a3bf2),
	.w6(32'hba4d156f),
	.w7(32'h3ac4273f),
	.w8(32'hba2cec25),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8003217),
	.w1(32'h39dca089),
	.w2(32'h39bbf8f3),
	.w3(32'h3a3ea754),
	.w4(32'h3a834997),
	.w5(32'h39ceaced),
	.w6(32'h3a695404),
	.w7(32'h3a9de525),
	.w8(32'h39969e6a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e80ba6),
	.w1(32'hb9037bbf),
	.w2(32'hb9a01e3c),
	.w3(32'h3985c7a5),
	.w4(32'h3ac622a8),
	.w5(32'hb9004c85),
	.w6(32'h38b8867b),
	.w7(32'h3adb1517),
	.w8(32'h39f0524a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fe45d7),
	.w1(32'hbb128a4a),
	.w2(32'hb8a87fe6),
	.w3(32'hbacd29b7),
	.w4(32'hba6b5be4),
	.w5(32'hb8e955e0),
	.w6(32'hb77e9863),
	.w7(32'hb96d91ed),
	.w8(32'hb9dbf956),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10a0fe),
	.w1(32'hbad15de8),
	.w2(32'hbb3adcf3),
	.w3(32'hbaa5fcbc),
	.w4(32'hba422542),
	.w5(32'hbb44d9b1),
	.w6(32'hba8f0af4),
	.w7(32'hb9cbabee),
	.w8(32'hbb14bf82),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf560eb),
	.w1(32'hbb89cf51),
	.w2(32'hbba75044),
	.w3(32'hbb5ebd11),
	.w4(32'hbb34d6e0),
	.w5(32'hba579b4d),
	.w6(32'h3ad09226),
	.w7(32'hb8fa2daf),
	.w8(32'h3ae1981b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a584549),
	.w1(32'h3a41d63c),
	.w2(32'h3ac5b8f7),
	.w3(32'h39262b54),
	.w4(32'hb969cd0f),
	.w5(32'h3a5ef8c1),
	.w6(32'h3b0c4a46),
	.w7(32'h3aa4ef62),
	.w8(32'hb9cb3384),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa17346),
	.w1(32'hba9a09ab),
	.w2(32'h394cf9aa),
	.w3(32'hba6213a5),
	.w4(32'h39cf2367),
	.w5(32'h3a5eb4e5),
	.w6(32'hb9d86f92),
	.w7(32'h3a45830a),
	.w8(32'h39f7bf26),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89cce11),
	.w1(32'h3aa589c6),
	.w2(32'h38992486),
	.w3(32'h39ec82b4),
	.w4(32'hbad1be3e),
	.w5(32'hb9b749e6),
	.w6(32'h381b34e8),
	.w7(32'hb960e6f7),
	.w8(32'h3a3e4789),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b031226),
	.w1(32'h3b03c93f),
	.w2(32'h3afa850f),
	.w3(32'h3808df70),
	.w4(32'hb96f05ef),
	.w5(32'hb9f6ede5),
	.w6(32'h3ae3123d),
	.w7(32'h3a88d74c),
	.w8(32'h3aa5b14a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85e3d6),
	.w1(32'hbbcd5920),
	.w2(32'hbc1d75b8),
	.w3(32'hbb533af6),
	.w4(32'hbbb73fc6),
	.w5(32'hbbb008ec),
	.w6(32'h3a854ef4),
	.w7(32'h37fdfc12),
	.w8(32'hb96f1f89),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e98a4),
	.w1(32'hbbd08df8),
	.w2(32'hbc15288c),
	.w3(32'h3adcd8ea),
	.w4(32'h3ad385be),
	.w5(32'hbbd8db05),
	.w6(32'hbbe39473),
	.w7(32'hbb9b77fe),
	.w8(32'hbc3af08d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbfc7b),
	.w1(32'hbbb7c642),
	.w2(32'hbbf7bb0c),
	.w3(32'hbb9c97df),
	.w4(32'hba39b8f9),
	.w5(32'hbb0a1582),
	.w6(32'hbb4d0366),
	.w7(32'h3a06020e),
	.w8(32'hbafe1055),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379ac09c),
	.w1(32'h3b11c1ea),
	.w2(32'hbb7a1746),
	.w3(32'hbb3dc423),
	.w4(32'h3b38c15d),
	.w5(32'hbb22cb5a),
	.w6(32'hbb644979),
	.w7(32'hbb0812cf),
	.w8(32'hbc03aa59),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5f5cc),
	.w1(32'h3a127d80),
	.w2(32'h3aee993a),
	.w3(32'h3a13e19d),
	.w4(32'h3ae77901),
	.w5(32'hb9636f17),
	.w6(32'hb8cf7646),
	.w7(32'h3aff6518),
	.w8(32'hbae3d58f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb016bc8),
	.w1(32'h3a1b6fe7),
	.w2(32'h39a9e825),
	.w3(32'h390982d4),
	.w4(32'h3a0844eb),
	.w5(32'h3a8b71e1),
	.w6(32'h3a499480),
	.w7(32'hb9c50c4d),
	.w8(32'h3b1798cc),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5bd5d),
	.w1(32'h3b0d2e9d),
	.w2(32'h3afeeb1e),
	.w3(32'hb8a5b638),
	.w4(32'h3a9e7da2),
	.w5(32'h3ace381f),
	.w6(32'h3b8d1c60),
	.w7(32'h3b860003),
	.w8(32'hb881428c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba827168),
	.w1(32'hb9931cd5),
	.w2(32'h3a8a63e8),
	.w3(32'h3a25df5b),
	.w4(32'hb9b1d369),
	.w5(32'hba0a7def),
	.w6(32'h3b1b90d8),
	.w7(32'h3ae46e46),
	.w8(32'h3a56039b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78c1ef),
	.w1(32'h39512a17),
	.w2(32'h3909ec01),
	.w3(32'h3acfb23f),
	.w4(32'h3a6562c7),
	.w5(32'h3a3964e0),
	.w6(32'h39c21a1f),
	.w7(32'hba7b86df),
	.w8(32'h3a273d90),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f7eb4),
	.w1(32'hbb11d538),
	.w2(32'h37ee9ed8),
	.w3(32'hba93e112),
	.w4(32'hba013eba),
	.w5(32'h3920b510),
	.w6(32'h39cc228e),
	.w7(32'h3ae017ac),
	.w8(32'h3aced8b3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee2cd4),
	.w1(32'hbb79f67e),
	.w2(32'hbb98bc39),
	.w3(32'hbb831895),
	.w4(32'hba03611a),
	.w5(32'hbb94f8d9),
	.w6(32'hbb658caf),
	.w7(32'h39714458),
	.w8(32'hbae4834a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9601d9),
	.w1(32'hbb5e4b3f),
	.w2(32'hbba28fbb),
	.w3(32'hbb60686b),
	.w4(32'hbab18456),
	.w5(32'hbadc1543),
	.w6(32'hbb4c2a0d),
	.w7(32'hbb318ce6),
	.w8(32'hba87e0d5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb612b9b),
	.w1(32'hb8d18fce),
	.w2(32'hbb3f028b),
	.w3(32'h3a747424),
	.w4(32'hb91cb1c7),
	.w5(32'hbb6e1f24),
	.w6(32'h3ab8eb2c),
	.w7(32'h3a6806c4),
	.w8(32'hbb4b9fc9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9182c9),
	.w1(32'hbb2377df),
	.w2(32'hbb8a6623),
	.w3(32'hbaea1904),
	.w4(32'hbb8fa734),
	.w5(32'h3b03d0fe),
	.w6(32'h3a911705),
	.w7(32'hbaa16d92),
	.w8(32'h3b527edf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add9981),
	.w1(32'h3a5311e6),
	.w2(32'h39ebf8d4),
	.w3(32'h3b3c5171),
	.w4(32'h3af18dbf),
	.w5(32'hbb39fb52),
	.w6(32'h3a385b6e),
	.w7(32'h3ad61f0d),
	.w8(32'hba590ea2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbae83),
	.w1(32'hba898660),
	.w2(32'hba510bed),
	.w3(32'h39a92c76),
	.w4(32'hb92a999d),
	.w5(32'hba99b868),
	.w6(32'h3affc1dd),
	.w7(32'h3b05b543),
	.w8(32'hba7b6be8),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7d2d8),
	.w1(32'h39b63d00),
	.w2(32'hba3b71c9),
	.w3(32'hba531262),
	.w4(32'hbaac11d1),
	.w5(32'h3ae7f21e),
	.w6(32'h38a14ed9),
	.w7(32'hba1f5740),
	.w8(32'h3a72ba45),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7f9fd),
	.w1(32'h39a3a066),
	.w2(32'hba59a130),
	.w3(32'hb999fe47),
	.w4(32'hba8be7f5),
	.w5(32'h3a150dc3),
	.w6(32'h3a2ed085),
	.w7(32'hbb2c0f26),
	.w8(32'h3a14d989),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fccefc),
	.w1(32'h3a950122),
	.w2(32'h3960b4a1),
	.w3(32'h39c3bbc6),
	.w4(32'h39987b6f),
	.w5(32'hbb08735a),
	.w6(32'h3a868c1c),
	.w7(32'h37b9a9f2),
	.w8(32'hbac9d5a8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cc671),
	.w1(32'h3a29756d),
	.w2(32'h3a3a91f9),
	.w3(32'hb8543e3a),
	.w4(32'hba5e085c),
	.w5(32'hbaaedcd1),
	.w6(32'h3af10407),
	.w7(32'h3a89f715),
	.w8(32'hbb4db892),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb955ae1),
	.w1(32'hbada6418),
	.w2(32'hbba49d79),
	.w3(32'hbb7c0440),
	.w4(32'h38618c74),
	.w5(32'hbaadfb34),
	.w6(32'hbb375da2),
	.w7(32'hbae05c70),
	.w8(32'hbb089092),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a186f),
	.w1(32'h3aa8abe1),
	.w2(32'h3aecff65),
	.w3(32'h3a70cafe),
	.w4(32'h3b0d42b5),
	.w5(32'hbad02e53),
	.w6(32'h3b1190f6),
	.w7(32'h3b13a49d),
	.w8(32'hbad15822),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cfb4a),
	.w1(32'hbb427f33),
	.w2(32'hbb5ee360),
	.w3(32'hbb393844),
	.w4(32'hbac2d0ee),
	.w5(32'h396d5320),
	.w6(32'hbb5cc162),
	.w7(32'hbb3eec3a),
	.w8(32'hbb4da549),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf184d),
	.w1(32'h3906b98a),
	.w2(32'hbb449888),
	.w3(32'hba3ea977),
	.w4(32'h3aad1f53),
	.w5(32'h3a128c84),
	.w6(32'h3a817e43),
	.w7(32'h3b14e2c2),
	.w8(32'h3996a31d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f4eab),
	.w1(32'h3b4a2e57),
	.w2(32'h3a2e742f),
	.w3(32'hba079bd0),
	.w4(32'hba2444a0),
	.w5(32'hbb060858),
	.w6(32'h3a189171),
	.w7(32'hb805c4ca),
	.w8(32'hbb037ef3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e22ec),
	.w1(32'hbb6233d2),
	.w2(32'hbbe266f9),
	.w3(32'hb982b7b6),
	.w4(32'hbb1279da),
	.w5(32'hbc29b7fc),
	.w6(32'h3ba7c556),
	.w7(32'hba225e21),
	.w8(32'hbbad214d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f372b),
	.w1(32'h3b0a6f5e),
	.w2(32'h3988f040),
	.w3(32'hbac4cd5d),
	.w4(32'h3a9508d3),
	.w5(32'hba48f8e9),
	.w6(32'hbadd0134),
	.w7(32'h390318bd),
	.w8(32'hbaa00ef0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb09310),
	.w1(32'hbbbb5602),
	.w2(32'hbc0f5ae6),
	.w3(32'hba92b84d),
	.w4(32'hbb0854a6),
	.w5(32'hbb658ae6),
	.w6(32'hbb00c2f9),
	.w7(32'hbae21f0f),
	.w8(32'hbba0cda9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e7b5d),
	.w1(32'hba62ba32),
	.w2(32'hba938321),
	.w3(32'h3a8896a0),
	.w4(32'hb9748328),
	.w5(32'hbaeb1616),
	.w6(32'h3acf1968),
	.w7(32'h3b03ce9f),
	.w8(32'h3a05480d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba664492),
	.w1(32'h3acc9230),
	.w2(32'h3a610282),
	.w3(32'hba5262dd),
	.w4(32'h3ae7bb67),
	.w5(32'hba566973),
	.w6(32'hba0afa7c),
	.w7(32'h3a77b239),
	.w8(32'h3a6a4da7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9afa0),
	.w1(32'h3b155f72),
	.w2(32'h3add0bf3),
	.w3(32'h3b2a43fb),
	.w4(32'h39918c19),
	.w5(32'h3acfea34),
	.w6(32'h3b865245),
	.w7(32'h3b3cc85d),
	.w8(32'h3ab834ad),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad95153),
	.w1(32'hbb6b1564),
	.w2(32'hbbbaed36),
	.w3(32'h3925fb8b),
	.w4(32'hbae9d944),
	.w5(32'hbba28f21),
	.w6(32'hba4c5618),
	.w7(32'hbaeaceb3),
	.w8(32'hbbc10779),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fee647),
	.w1(32'hbb0c6674),
	.w2(32'hbb17b6d7),
	.w3(32'hb9f4f3a9),
	.w4(32'hba01fa43),
	.w5(32'hbb81d70f),
	.w6(32'h3b81459e),
	.w7(32'h3b0b9f21),
	.w8(32'h3a54725f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa7419),
	.w1(32'hbbb8faeb),
	.w2(32'hbb897a19),
	.w3(32'hbbd5f57f),
	.w4(32'h3ab62e2b),
	.w5(32'hbb0c4fbb),
	.w6(32'hbbd76019),
	.w7(32'h3b1ab1e0),
	.w8(32'h39fbed86),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba577e72),
	.w1(32'h3ace956d),
	.w2(32'hbbae899e),
	.w3(32'hbbb112a1),
	.w4(32'h3aab193f),
	.w5(32'hb9cc09e3),
	.w6(32'hbb2abf51),
	.w7(32'hbabb4149),
	.w8(32'hbadf13b4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a509eab),
	.w1(32'hbb9395ac),
	.w2(32'hbbd076e4),
	.w3(32'hba9f8ac9),
	.w4(32'h3a5bbecd),
	.w5(32'hbb484c75),
	.w6(32'hbb7e22d9),
	.w7(32'hbbd1bb4d),
	.w8(32'hbbdd8677),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb014724),
	.w1(32'hbb111f27),
	.w2(32'h3a03a544),
	.w3(32'hbb09df7e),
	.w4(32'hbabe7ee6),
	.w5(32'hbbd6342b),
	.w6(32'h3b234b9a),
	.w7(32'h3be7ceed),
	.w8(32'hbb0875fa),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870c6f),
	.w1(32'hbb15edab),
	.w2(32'hba8d88ba),
	.w3(32'hbac41d37),
	.w4(32'hbab0d357),
	.w5(32'h3bacf5d6),
	.w6(32'hbaa893b3),
	.w7(32'hba9817c9),
	.w8(32'h3a88e9ac),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a3e6f),
	.w1(32'hbbe86f6c),
	.w2(32'hbbf6477b),
	.w3(32'hbbbb0963),
	.w4(32'h3b871f9d),
	.w5(32'h3a28338b),
	.w6(32'hbb1a77ab),
	.w7(32'h3b9dfe45),
	.w8(32'h3a1ead70),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac42735),
	.w1(32'hbaefadc4),
	.w2(32'hbb98c88a),
	.w3(32'hbab7c566),
	.w4(32'hba524b86),
	.w5(32'hbbc84320),
	.w6(32'hb9886e76),
	.w7(32'hbba44483),
	.w8(32'hbb950987),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14388d),
	.w1(32'hbaa8f643),
	.w2(32'h3a8766b7),
	.w3(32'hb95bc44d),
	.w4(32'h3a260ba5),
	.w5(32'hba98d60e),
	.w6(32'hbb3be6bc),
	.w7(32'hb9a7c5ff),
	.w8(32'hb9904013),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f42e0),
	.w1(32'h39968a3a),
	.w2(32'h3a074048),
	.w3(32'hbb7deb94),
	.w4(32'hbb1a6196),
	.w5(32'hbab5508d),
	.w6(32'hbb609f05),
	.w7(32'hba9835e8),
	.w8(32'hb9c8ea1f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cacf3a),
	.w1(32'hbb2dcfb1),
	.w2(32'hbbae56c6),
	.w3(32'h3b239ec1),
	.w4(32'h3a14e405),
	.w5(32'hbb8f9ae8),
	.w6(32'h3a3fe081),
	.w7(32'hbae1a7a2),
	.w8(32'hbbba94cf),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98e371),
	.w1(32'hbab3d66e),
	.w2(32'hbb605b6f),
	.w3(32'hbb96b882),
	.w4(32'hbb78dbb0),
	.w5(32'hba71b569),
	.w6(32'hbbb81abf),
	.w7(32'hbbc6eba5),
	.w8(32'hba7bb810),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b635ed2),
	.w1(32'h3afffb68),
	.w2(32'h3aa8e09b),
	.w3(32'hba9b4c43),
	.w4(32'h3b0eaaa4),
	.w5(32'h3b1908a9),
	.w6(32'h39d9de96),
	.w7(32'h3b116a9c),
	.w8(32'h3b9924eb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01054a),
	.w1(32'h3b533c4b),
	.w2(32'hb924e2a0),
	.w3(32'h3a05d93d),
	.w4(32'hbaa7a055),
	.w5(32'h3b5375eb),
	.w6(32'hba7c3eda),
	.w7(32'hbafe1dfd),
	.w8(32'hba735e40),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3adead),
	.w1(32'h38d5990d),
	.w2(32'hbb05793f),
	.w3(32'h3a741d7f),
	.w4(32'h398e5c4d),
	.w5(32'hb9874cc9),
	.w6(32'hbba29219),
	.w7(32'hbb92a786),
	.w8(32'hbb2c151f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7b354),
	.w1(32'hbc021d80),
	.w2(32'hbc0e10dc),
	.w3(32'hbc144fce),
	.w4(32'hbbb1ac7f),
	.w5(32'hbb8612d8),
	.w6(32'hbc057fc4),
	.w7(32'hbb109f54),
	.w8(32'hbb50c66b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39c651),
	.w1(32'hb9bcb356),
	.w2(32'hbae3e85d),
	.w3(32'hb9f24000),
	.w4(32'h39a4b36e),
	.w5(32'h3a7b261d),
	.w6(32'hbb0a5ae5),
	.w7(32'hbb0f4ab3),
	.w8(32'h3b6e4fd5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b6afe),
	.w1(32'h393c0c88),
	.w2(32'h3a053e59),
	.w3(32'h3a8144e8),
	.w4(32'hbac2d3d9),
	.w5(32'hb9c9270f),
	.w6(32'h3943f393),
	.w7(32'hbac5c561),
	.w8(32'h3a895462),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adec215),
	.w1(32'h3a8a235f),
	.w2(32'h398b6790),
	.w3(32'h3a3fb891),
	.w4(32'h3a0a9570),
	.w5(32'h3af441ee),
	.w6(32'h3af8c3c8),
	.w7(32'h3ad349f5),
	.w8(32'hb8baba4c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb451f),
	.w1(32'hba70203e),
	.w2(32'hba031be4),
	.w3(32'h3a0ffcab),
	.w4(32'h3a8489f4),
	.w5(32'hbae8a800),
	.w6(32'h3a0be32d),
	.w7(32'hba0f0ba5),
	.w8(32'hbb14ff5f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2daa3d),
	.w1(32'hba17263f),
	.w2(32'h3a387d39),
	.w3(32'hbae08198),
	.w4(32'hba324850),
	.w5(32'hbb67db0c),
	.w6(32'hba9eefc1),
	.w7(32'h39da47b1),
	.w8(32'hbb754db1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9c37f),
	.w1(32'hbb9df9d5),
	.w2(32'hbb9b2ada),
	.w3(32'hbb3baca7),
	.w4(32'hbb10cfeb),
	.w5(32'hbbce2cc5),
	.w6(32'hbb9b6412),
	.w7(32'hbb5195d1),
	.w8(32'hbbe47b68),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5650a3),
	.w1(32'h3b239cbe),
	.w2(32'h3ae3ddc4),
	.w3(32'hbab29427),
	.w4(32'hbb6c6132),
	.w5(32'h3bad0bea),
	.w6(32'hba2f28fe),
	.w7(32'hbaa7269b),
	.w8(32'h3bb5a7ef),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26b213),
	.w1(32'h3b3b2e0d),
	.w2(32'hbaefd9f1),
	.w3(32'h3b96c1b1),
	.w4(32'hbb91fbb2),
	.w5(32'h3b7c9606),
	.w6(32'h3b8163cf),
	.w7(32'hbb46bd5d),
	.w8(32'h39701868),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb289415),
	.w1(32'hbbc9a3d8),
	.w2(32'hbba886d4),
	.w3(32'h39e03ce3),
	.w4(32'h3b0884cc),
	.w5(32'hbb00b9db),
	.w6(32'hbbe8ae36),
	.w7(32'hbbc37214),
	.w8(32'hbb6fdaf8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f23e4),
	.w1(32'hbaa02977),
	.w2(32'hbac57b21),
	.w3(32'hbb3d763a),
	.w4(32'hbb80f666),
	.w5(32'h3b0cd76b),
	.w6(32'hbb4e5a35),
	.w7(32'hbb7fc568),
	.w8(32'h3ae341c9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba626f99),
	.w1(32'hbba9fd60),
	.w2(32'hbb305ba8),
	.w3(32'h3a019d46),
	.w4(32'h3aa1f3fe),
	.w5(32'hba5dadc8),
	.w6(32'hbb474898),
	.w7(32'hba08f5a0),
	.w8(32'hbaca612b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab39d35),
	.w1(32'hbadbc5f8),
	.w2(32'hba22aa06),
	.w3(32'hbb0f8ef9),
	.w4(32'hb85f8ac7),
	.w5(32'hba1aad67),
	.w6(32'hbbbeaccd),
	.w7(32'hbaacdbfb),
	.w8(32'hbb212086),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc3a0d),
	.w1(32'hbacf3be7),
	.w2(32'h38d3b74d),
	.w3(32'hbb548877),
	.w4(32'hba2bd91b),
	.w5(32'hb9f7ee37),
	.w6(32'hbbb66ea7),
	.w7(32'hbb87c0a9),
	.w8(32'hba42c729),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8d079),
	.w1(32'hbba35e68),
	.w2(32'hbbe9003b),
	.w3(32'h3a9f88ae),
	.w4(32'hbb2b88cc),
	.w5(32'hb91f2974),
	.w6(32'hbb2f8b91),
	.w7(32'hbb7ff040),
	.w8(32'hbaafa32b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af57417),
	.w1(32'h39367124),
	.w2(32'h3aa9d2ff),
	.w3(32'hb762c3ba),
	.w4(32'hba6f87b9),
	.w5(32'hbb06030e),
	.w6(32'hbada44c1),
	.w7(32'h3aafccc2),
	.w8(32'hbad36a37),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1bffd),
	.w1(32'h3ae574da),
	.w2(32'h3acc4fcc),
	.w3(32'h3a39d28b),
	.w4(32'h3ad939f3),
	.w5(32'h3b8d86e5),
	.w6(32'hb96d50a7),
	.w7(32'h3a1f5124),
	.w8(32'h3c24a771),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05ec1b),
	.w1(32'hbb3ba50a),
	.w2(32'hbbd6d565),
	.w3(32'h3b6c0dc1),
	.w4(32'hbaf1430c),
	.w5(32'hbb1a4338),
	.w6(32'h3b5d61a3),
	.w7(32'hbb49a55d),
	.w8(32'hbb85fb13),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16453a),
	.w1(32'hb9d0359a),
	.w2(32'hbb084f39),
	.w3(32'hbb08a46b),
	.w4(32'hbb088a8d),
	.w5(32'hbb319ac4),
	.w6(32'hba441f41),
	.w7(32'hbb1fb86c),
	.w8(32'hbabf30c3),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e447e6),
	.w1(32'h3a66538a),
	.w2(32'h3adfdc44),
	.w3(32'hbb493219),
	.w4(32'h3a408203),
	.w5(32'h39ee54f8),
	.w6(32'hbbcc35ec),
	.w7(32'hb8abb37d),
	.w8(32'hba56d248),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb300bc4),
	.w1(32'hbb7f520c),
	.w2(32'hbb8b652f),
	.w3(32'hbbc14fa0),
	.w4(32'hbb889437),
	.w5(32'h3ada739f),
	.w6(32'hbb6bb152),
	.w7(32'hbb308daf),
	.w8(32'h3a98ba05),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c615b),
	.w1(32'hbb2a88a2),
	.w2(32'hbb7317c0),
	.w3(32'hba4ede87),
	.w4(32'hbb41d9e7),
	.w5(32'hbba32b85),
	.w6(32'h39f33d71),
	.w7(32'hba11177d),
	.w8(32'h39132ef6),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03c268),
	.w1(32'hba017b54),
	.w2(32'h3a870559),
	.w3(32'hbb698f7c),
	.w4(32'hbac4dde2),
	.w5(32'h3abf51e1),
	.w6(32'hbb7b0e51),
	.w7(32'hbaa2d4e7),
	.w8(32'h360f9128),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988b11c),
	.w1(32'hbb23a9a9),
	.w2(32'hbb8ad922),
	.w3(32'hba4f997f),
	.w4(32'hba89cfeb),
	.w5(32'hbae9e854),
	.w6(32'hbab46362),
	.w7(32'hba9a18fb),
	.w8(32'hbb420bff),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48f236),
	.w1(32'hbb8f07fa),
	.w2(32'hbb3b06c5),
	.w3(32'hbbc1d2c2),
	.w4(32'hbbab4010),
	.w5(32'hb86377b5),
	.w6(32'hbb8984a1),
	.w7(32'hbb228e7c),
	.w8(32'h3b00e59a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88613f0),
	.w1(32'h3aef69ba),
	.w2(32'h3ad0a22a),
	.w3(32'hb72dcd11),
	.w4(32'h3ac8aacf),
	.w5(32'hbac75992),
	.w6(32'hbb159549),
	.w7(32'hb9dc22b7),
	.w8(32'hbabc53f2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fa6fc),
	.w1(32'hbacd1d01),
	.w2(32'hbbb1726d),
	.w3(32'hbac9d31f),
	.w4(32'hbb0f3720),
	.w5(32'hbbdf92af),
	.w6(32'hbac4785a),
	.w7(32'hba8e211f),
	.w8(32'hbbeb41a6),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7405d),
	.w1(32'hbaa1732a),
	.w2(32'h3ab96162),
	.w3(32'hba9c61de),
	.w4(32'h3b94b495),
	.w5(32'hbb92b407),
	.w6(32'hbb7aef70),
	.w7(32'h3a0f6ccf),
	.w8(32'hbb973fd0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61db96),
	.w1(32'hb9ea2ee8),
	.w2(32'h3afaf117),
	.w3(32'hbb86fddd),
	.w4(32'hbb90bb58),
	.w5(32'hbb221a3b),
	.w6(32'hbb876158),
	.w7(32'hbb508709),
	.w8(32'hbb7fc61d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0dce23),
	.w1(32'h3adf0d38),
	.w2(32'h3b0497d9),
	.w3(32'hb7d804e1),
	.w4(32'h3a7e9e44),
	.w5(32'hbb56befa),
	.w6(32'h3aa5dfcf),
	.w7(32'h3a32932a),
	.w8(32'hbb99fcd5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac93e21),
	.w1(32'h3a768bfc),
	.w2(32'h3be6fd3e),
	.w3(32'hbabb5e14),
	.w4(32'h3b719a13),
	.w5(32'h3bc26083),
	.w6(32'hbb2063ec),
	.w7(32'h3ba3cd9f),
	.w8(32'h3b998dfb),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89eff6),
	.w1(32'hba817ca0),
	.w2(32'h3ada22a3),
	.w3(32'h3ad171b1),
	.w4(32'h3b1f7724),
	.w5(32'hba803515),
	.w6(32'hbacd092b),
	.w7(32'hba042435),
	.w8(32'hbacb59b4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22564b),
	.w1(32'hba301f60),
	.w2(32'hbb10c746),
	.w3(32'hbade3189),
	.w4(32'hba955fab),
	.w5(32'h39f7e400),
	.w6(32'hba2e1d84),
	.w7(32'hba55bb77),
	.w8(32'hb90529de),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39d1a8),
	.w1(32'hbad13d31),
	.w2(32'h3aadfe7c),
	.w3(32'hbb1c9aff),
	.w4(32'h3aacc9f0),
	.w5(32'h3bc4c974),
	.w6(32'hbb51a158),
	.w7(32'h3a57945b),
	.w8(32'h3b5cbf94),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9acf7d),
	.w1(32'h3b12d4d6),
	.w2(32'hbb7cc4ab),
	.w3(32'h3a43ecba),
	.w4(32'hb9e8f957),
	.w5(32'hbb8b2360),
	.w6(32'hbba8b774),
	.w7(32'hbb06704c),
	.w8(32'hbba82863),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25e5c7),
	.w1(32'hbb553051),
	.w2(32'h3b878caa),
	.w3(32'hbb30f894),
	.w4(32'h3b4ddf72),
	.w5(32'hba940a2a),
	.w6(32'hbb60cc9a),
	.w7(32'h3b42f35b),
	.w8(32'hba03eb8d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83b8de),
	.w1(32'hbb4a413a),
	.w2(32'hbbdfce26),
	.w3(32'hbaac05f6),
	.w4(32'hbae0a1d1),
	.w5(32'hbbedf1b7),
	.w6(32'hba19b6c4),
	.w7(32'hbb2bb92f),
	.w8(32'hbbf406ed),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cbff4),
	.w1(32'hbb486715),
	.w2(32'hbaaddb03),
	.w3(32'hbb3a474b),
	.w4(32'h394b2fdb),
	.w5(32'hbbfc0db6),
	.w6(32'hbbbc6c96),
	.w7(32'hba939470),
	.w8(32'hbc01faca),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d37ea),
	.w1(32'h3b52666e),
	.w2(32'h3c1c995f),
	.w3(32'hbb7515ca),
	.w4(32'h3ac74d88),
	.w5(32'hba9b6167),
	.w6(32'hb749a5dd),
	.w7(32'h3c2c035d),
	.w8(32'h3b8f3002),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12b50b),
	.w1(32'hbb60e7ba),
	.w2(32'h3a0fd22a),
	.w3(32'hb92551ba),
	.w4(32'hba4faef3),
	.w5(32'hbadb5585),
	.w6(32'h3a9ca5e7),
	.w7(32'hba803782),
	.w8(32'hbaf7f488),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1861ab),
	.w1(32'hbb8b4d45),
	.w2(32'hbb81d405),
	.w3(32'hbbab4cab),
	.w4(32'hbb4684c2),
	.w5(32'hba42d7b7),
	.w6(32'hbbc8e3fb),
	.w7(32'hbbc4ca6d),
	.w8(32'hba6d8ae6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35bb02),
	.w1(32'h3a26ca77),
	.w2(32'h3a3f2a8f),
	.w3(32'h3b331584),
	.w4(32'h3b103135),
	.w5(32'h3b8276f8),
	.w6(32'h3b6c9dab),
	.w7(32'h3b0333c7),
	.w8(32'h3b3fad67),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74bb95),
	.w1(32'h3974b7ff),
	.w2(32'hb9cf82f6),
	.w3(32'h384d5324),
	.w4(32'h3a83e963),
	.w5(32'hbb2b66e0),
	.w6(32'hbb4752f2),
	.w7(32'hbb27b8ac),
	.w8(32'hbbbd288b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f42f6),
	.w1(32'h3a0fc5cb),
	.w2(32'hba8d6cb8),
	.w3(32'h39253620),
	.w4(32'h3b7df4e1),
	.w5(32'h3c2c0586),
	.w6(32'hbb1c09ce),
	.w7(32'h3b09a507),
	.w8(32'h3c22a20c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05c014),
	.w1(32'h3c1c8e72),
	.w2(32'h3b06d47f),
	.w3(32'h3c007515),
	.w4(32'h3a8840f7),
	.w5(32'hbb80ca69),
	.w6(32'h3bbb7239),
	.w7(32'h3a2f24bd),
	.w8(32'hbb652308),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef67b7),
	.w1(32'h3bd68c79),
	.w2(32'h3ba82ef4),
	.w3(32'hbb980a35),
	.w4(32'hba947a85),
	.w5(32'h3b24797f),
	.w6(32'hbb359317),
	.w7(32'h3b79cba9),
	.w8(32'h3b7d9ba9),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17ecf0),
	.w1(32'hbb426c20),
	.w2(32'hb80ed1be),
	.w3(32'h3b62e28f),
	.w4(32'h3a35b2db),
	.w5(32'h37c32b57),
	.w6(32'h3a59ec4c),
	.w7(32'hb9b22e75),
	.w8(32'h3ab89ebe),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a316774),
	.w1(32'hbba838e7),
	.w2(32'hbba9dc17),
	.w3(32'hbae23386),
	.w4(32'hbb5d76e5),
	.w5(32'hbbd254a6),
	.w6(32'hbb355ddf),
	.w7(32'hbb6de473),
	.w8(32'hbba353cb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb078493),
	.w1(32'hb96e526a),
	.w2(32'h3a135bd5),
	.w3(32'hbac4a31c),
	.w4(32'hbb1eadb1),
	.w5(32'hbaf1d6a0),
	.w6(32'hba230c2a),
	.w7(32'hb948b86b),
	.w8(32'hbb8176ae),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bd86d),
	.w1(32'hba9a8d12),
	.w2(32'h3b2c2ae5),
	.w3(32'h3aece31d),
	.w4(32'h3ab4f771),
	.w5(32'hb9c80852),
	.w6(32'hbb35ac9f),
	.w7(32'h3a49625b),
	.w8(32'hbb17da1d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04e060),
	.w1(32'hbb2c6ccc),
	.w2(32'h3bb4fb87),
	.w3(32'hbb923331),
	.w4(32'h395a54bd),
	.w5(32'h3aaca867),
	.w6(32'hbb95bf5e),
	.w7(32'h39031c07),
	.w8(32'h39ccc224),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aaf1ca),
	.w1(32'hbb2ed351),
	.w2(32'hbb0d075c),
	.w3(32'h3b3ceff9),
	.w4(32'h3a5bbc4e),
	.w5(32'h3a8335e8),
	.w6(32'hbab997e4),
	.w7(32'hbb0900ca),
	.w8(32'hbae6a850),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc236b),
	.w1(32'hbb36a26a),
	.w2(32'hba7b6377),
	.w3(32'hbaa63df5),
	.w4(32'hba9d260f),
	.w5(32'hb97e4a1e),
	.w6(32'hba3ace27),
	.w7(32'h3905f2fa),
	.w8(32'hba490e50),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67d81a),
	.w1(32'h3b49ef94),
	.w2(32'h3b5c17ef),
	.w3(32'hbba7146c),
	.w4(32'hbb85860c),
	.w5(32'hbb0b80cf),
	.w6(32'hbb6f8813),
	.w7(32'hb9f3b7cb),
	.w8(32'hbba9001c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3af0ad),
	.w1(32'h3b15f162),
	.w2(32'hbad4c8dc),
	.w3(32'hb9c4cdc6),
	.w4(32'h3b164454),
	.w5(32'hbbf2c102),
	.w6(32'h3a40927c),
	.w7(32'h3a13d5bf),
	.w8(32'hbbf49641),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0f8a8),
	.w1(32'h3b41616c),
	.w2(32'hbaecea66),
	.w3(32'hba3f08cc),
	.w4(32'h3b1a892e),
	.w5(32'hbbcd2120),
	.w6(32'hbb4d657f),
	.w7(32'h3b92b3cd),
	.w8(32'hbbab82da),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a1c345),
	.w1(32'hb96fd0dc),
	.w2(32'h3a542e95),
	.w3(32'hbb882cd4),
	.w4(32'hbaa1d5dc),
	.w5(32'h3b1abad6),
	.w6(32'hbb853cb0),
	.w7(32'hbb2655a8),
	.w8(32'h3a605b86),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ded1ac),
	.w1(32'hba68def8),
	.w2(32'hbb8c00c2),
	.w3(32'hba2a77c5),
	.w4(32'hba0acb8b),
	.w5(32'h38c84434),
	.w6(32'h3a2ec61a),
	.w7(32'hbb1b9975),
	.w8(32'hbb303e8c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9da92),
	.w1(32'hb9eac903),
	.w2(32'h3aa7f437),
	.w3(32'hba3fc1b7),
	.w4(32'hba2bf98a),
	.w5(32'hbbad077f),
	.w6(32'hbaad0076),
	.w7(32'hba6df79b),
	.w8(32'hbb676c33),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32141a),
	.w1(32'hbc0c83a4),
	.w2(32'hbc37c2a4),
	.w3(32'hbbeea357),
	.w4(32'hbb9b19c9),
	.w5(32'hbbace768),
	.w6(32'hbbb459f9),
	.w7(32'hbb90e56e),
	.w8(32'hbbb8d97c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85deb1),
	.w1(32'h3aa56095),
	.w2(32'hbb17b8b0),
	.w3(32'hb9366ab5),
	.w4(32'h3ae59b0a),
	.w5(32'hbb469fcb),
	.w6(32'hba4b153a),
	.w7(32'hb892fb7f),
	.w8(32'hbb065a5e),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9da51e),
	.w1(32'hbb6f57e1),
	.w2(32'hbbd796ba),
	.w3(32'hbab66b37),
	.w4(32'hbb32e5b2),
	.w5(32'hbb53f18c),
	.w6(32'hbb06f0e6),
	.w7(32'hbb142817),
	.w8(32'hbb166105),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2702fe),
	.w1(32'h398dd106),
	.w2(32'hba751aec),
	.w3(32'h397579d7),
	.w4(32'hb9d6a3cf),
	.w5(32'hbb8ed2e3),
	.w6(32'h3a178e92),
	.w7(32'hb9d411ed),
	.w8(32'hbbac0bc3),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba7983),
	.w1(32'hbb915d17),
	.w2(32'hbb8d46f1),
	.w3(32'hbbc92fdc),
	.w4(32'hbb5471e7),
	.w5(32'hba164abf),
	.w6(32'hbba68f6f),
	.w7(32'hbb3fbe9c),
	.w8(32'h3a7f82d1),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae1b31),
	.w1(32'hba386a33),
	.w2(32'hbaa623de),
	.w3(32'h3aecf9b4),
	.w4(32'h3a210b5e),
	.w5(32'hbbb83eb7),
	.w6(32'h3aa8f8a8),
	.w7(32'hba4afaa4),
	.w8(32'hbb07bc40),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45a9fd),
	.w1(32'h38967bf8),
	.w2(32'h3b18c130),
	.w3(32'hba0fad39),
	.w4(32'h3a802ee7),
	.w5(32'h3ac76f85),
	.w6(32'hbadc30fe),
	.w7(32'h3a206093),
	.w8(32'hb9f07f35),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d15ce),
	.w1(32'h3906680c),
	.w2(32'hb78e635b),
	.w3(32'hba9537e0),
	.w4(32'h3a8c1552),
	.w5(32'hbbe0e64b),
	.w6(32'hb98d6848),
	.w7(32'hba0ea4c7),
	.w8(32'hbba72274),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28eee0),
	.w1(32'h3b2efb82),
	.w2(32'h3a772109),
	.w3(32'hbbc4ddd3),
	.w4(32'hbb79fc85),
	.w5(32'hbb5d2300),
	.w6(32'hbb8e1085),
	.w7(32'h3b239a6a),
	.w8(32'hbbba29ea),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7e49d),
	.w1(32'h3c0eea4a),
	.w2(32'h3b15829d),
	.w3(32'h3ba82ac1),
	.w4(32'hbafc5ab3),
	.w5(32'h3acd52a6),
	.w6(32'h3b841051),
	.w7(32'hb9a279d9),
	.w8(32'hbb05455a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa92db2),
	.w1(32'hba40661c),
	.w2(32'hbacab3bc),
	.w3(32'hbabe4ef2),
	.w4(32'hba33d332),
	.w5(32'hba2767e2),
	.w6(32'hbbafaca0),
	.w7(32'hbb0c4a5e),
	.w8(32'hbac5d215),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab9942),
	.w1(32'hbabc1386),
	.w2(32'h3b2550af),
	.w3(32'h3b3b7005),
	.w4(32'h3bc3e7ec),
	.w5(32'hbb5359fc),
	.w6(32'h39784f24),
	.w7(32'h3b8ce27d),
	.w8(32'hbb517ba8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c4fdf),
	.w1(32'hb9e066f3),
	.w2(32'h3acd0ce3),
	.w3(32'h3b06c2e2),
	.w4(32'h3b937086),
	.w5(32'h3adb89f7),
	.w6(32'h3baaada2),
	.w7(32'h3c1b402f),
	.w8(32'h3a96308b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969902a),
	.w1(32'h3ac2c8d1),
	.w2(32'hba746717),
	.w3(32'hbaf865d0),
	.w4(32'hbabbd8ee),
	.w5(32'h3b02d123),
	.w6(32'hbb008949),
	.w7(32'hbaa17b2c),
	.w8(32'h3b046a5f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24af45),
	.w1(32'h3a1ff993),
	.w2(32'hb9cf0571),
	.w3(32'h3a91d370),
	.w4(32'h38051795),
	.w5(32'h3a2adf28),
	.w6(32'h3ae3be01),
	.w7(32'hb9bb733c),
	.w8(32'h3ac68705),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb83661),
	.w1(32'hbc17b84c),
	.w2(32'hbc88c155),
	.w3(32'h3a089c07),
	.w4(32'hbb69272a),
	.w5(32'hbb037d6f),
	.w6(32'h395fe280),
	.w7(32'hbb8575a4),
	.w8(32'hba37ce84),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c4ba0),
	.w1(32'h3bacf4b1),
	.w2(32'hba444f02),
	.w3(32'hbbb08e92),
	.w4(32'hbb080dc4),
	.w5(32'hbba13f2a),
	.w6(32'h3a404d9b),
	.w7(32'h3b8a06ca),
	.w8(32'hbb5ec3f3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d486fd),
	.w1(32'hbb33fe06),
	.w2(32'hba70537d),
	.w3(32'hbb2771c3),
	.w4(32'hbada164c),
	.w5(32'hbbb59a30),
	.w6(32'hbbaef374),
	.w7(32'hbb530aa8),
	.w8(32'hbba790ea),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba696e0d),
	.w1(32'h3b40a0af),
	.w2(32'h3b939b06),
	.w3(32'hbb0c5120),
	.w4(32'hb9e0f386),
	.w5(32'hbb5d1c2a),
	.w6(32'hbba1d446),
	.w7(32'h39e86992),
	.w8(32'hbb3f1879),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29815e),
	.w1(32'hbad982c5),
	.w2(32'h3b154823),
	.w3(32'hba963991),
	.w4(32'hba4deef8),
	.w5(32'hbb4b6b4c),
	.w6(32'hbb25b148),
	.w7(32'h3b463175),
	.w8(32'hbbaf5dae),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab949b),
	.w1(32'hba72ffcc),
	.w2(32'hba27f9b3),
	.w3(32'hba331a25),
	.w4(32'hbab018c3),
	.w5(32'hba45903f),
	.w6(32'hbb5a15eb),
	.w7(32'h386fbd93),
	.w8(32'hbb8a600f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a5e5e),
	.w1(32'h3ac70f32),
	.w2(32'hbb1eab19),
	.w3(32'hb9b968cd),
	.w4(32'hbaabfffb),
	.w5(32'h3aa2644d),
	.w6(32'hbb9b7623),
	.w7(32'hb820fd14),
	.w8(32'h3acd1a19),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bed1dc),
	.w1(32'hbabc7cc6),
	.w2(32'hbb08fbde),
	.w3(32'h39595de3),
	.w4(32'hbb26d417),
	.w5(32'hbbb4f6b0),
	.w6(32'hbb76153c),
	.w7(32'hbb92fa85),
	.w8(32'hbbe30933),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65bcbf),
	.w1(32'hbb5edc0d),
	.w2(32'hbbc21f6d),
	.w3(32'hbc0f12f3),
	.w4(32'hbbbc23ed),
	.w5(32'hbbbab0ca),
	.w6(32'hbbff2145),
	.w7(32'hbc0642fd),
	.w8(32'hbc1df209),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbeaa35),
	.w1(32'hbb155198),
	.w2(32'hbaeb73bb),
	.w3(32'hbb784056),
	.w4(32'hbb22476a),
	.w5(32'h3b56af62),
	.w6(32'hbbbea043),
	.w7(32'hbb28cb63),
	.w8(32'h3ad9dab0),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cc7b8),
	.w1(32'hbbc1bf01),
	.w2(32'hbbca0b82),
	.w3(32'h3a8e802c),
	.w4(32'h3a8b7e76),
	.w5(32'hbb8e6ada),
	.w6(32'h36972986),
	.w7(32'hbb37d985),
	.w8(32'hbba72e33),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15ccbf),
	.w1(32'hbb9f2852),
	.w2(32'hbb970221),
	.w3(32'hbaeeb7fa),
	.w4(32'hbaf2664b),
	.w5(32'hbba6d5c8),
	.w6(32'hbb149da0),
	.w7(32'hbb4d31c7),
	.w8(32'hbbddd7c6),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c5bbb),
	.w1(32'h3a8d0080),
	.w2(32'h3bf0e555),
	.w3(32'hbba1e125),
	.w4(32'h3ab632bb),
	.w5(32'hbadcedc8),
	.w6(32'hbb5a25ef),
	.w7(32'h3b4994f3),
	.w8(32'hbb48fd54),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ad2d4),
	.w1(32'hbbb20a00),
	.w2(32'hbb9ae09d),
	.w3(32'hbbdd4892),
	.w4(32'hbbe535f3),
	.w5(32'h38a86059),
	.w6(32'hbb9ff457),
	.w7(32'hbb8afba2),
	.w8(32'hba075e98),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0aa9e),
	.w1(32'h3aef203e),
	.w2(32'h39d23a9b),
	.w3(32'hb983cca7),
	.w4(32'hbb4b8b27),
	.w5(32'h3a8ca4b2),
	.w6(32'hb8c58d27),
	.w7(32'hbb1bb3d0),
	.w8(32'hb907142d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba15e8),
	.w1(32'hb816b3c5),
	.w2(32'hbb0d396a),
	.w3(32'h39fd4b1e),
	.w4(32'hba89578d),
	.w5(32'hbb81de2f),
	.w6(32'hba4b56e5),
	.w7(32'hbae1a7c9),
	.w8(32'hbb9fbab5),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaa2c3),
	.w1(32'h3a253195),
	.w2(32'hba162ee6),
	.w3(32'hbb825617),
	.w4(32'h3b3f3e59),
	.w5(32'hbad31407),
	.w6(32'hbb5462ac),
	.w7(32'h3b02ce81),
	.w8(32'hbb65b937),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d71ec),
	.w1(32'h3bbad8f4),
	.w2(32'h3b2ff9fb),
	.w3(32'hba4e4bf1),
	.w4(32'h3b3526f4),
	.w5(32'hbb1ffa44),
	.w6(32'hbb51579e),
	.w7(32'h3bafda46),
	.w8(32'hbb873880),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d0d05),
	.w1(32'hba6e4a9b),
	.w2(32'h3ad69c07),
	.w3(32'hba8328a4),
	.w4(32'h3af5a8e5),
	.w5(32'hbaf7431c),
	.w6(32'hba2089d4),
	.w7(32'h3aa68c54),
	.w8(32'hbb39d10e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34bdbd),
	.w1(32'hbade13ac),
	.w2(32'hbb9d8861),
	.w3(32'hbb29306b),
	.w4(32'hba168903),
	.w5(32'hbac285c3),
	.w6(32'hbb695d0a),
	.w7(32'hbb1bcc2f),
	.w8(32'hbbae3bb2),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9ca3b),
	.w1(32'h3a8d9c3d),
	.w2(32'h39987bcc),
	.w3(32'hbb1b4e88),
	.w4(32'hba87832d),
	.w5(32'hbb88d4c6),
	.w6(32'hbb96b55b),
	.w7(32'hbb2de0d9),
	.w8(32'hb898db48),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb878a39e),
	.w1(32'h3aa269e4),
	.w2(32'hbb08cce0),
	.w3(32'hba9afc8a),
	.w4(32'hba637a3e),
	.w5(32'hbb9ffbca),
	.w6(32'h3ae01508),
	.w7(32'h3b1e748f),
	.w8(32'hbbcd8224),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9374b47),
	.w1(32'hba3ab0e3),
	.w2(32'hba16ca20),
	.w3(32'hbad81242),
	.w4(32'hbab12416),
	.w5(32'hb98efb5a),
	.w6(32'hbad72d12),
	.w7(32'hbafac2f8),
	.w8(32'hb9e18eac),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdfdf0),
	.w1(32'h3b3eb417),
	.w2(32'h3ba9839f),
	.w3(32'h399abd44),
	.w4(32'h3b33404d),
	.w5(32'h3b367db2),
	.w6(32'h3a025e93),
	.w7(32'h3b922d28),
	.w8(32'h3b749014),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b526265),
	.w1(32'h3a6f451e),
	.w2(32'hbb910cc9),
	.w3(32'h3b8bd0ff),
	.w4(32'h3b4797ab),
	.w5(32'hbae3e6a6),
	.w6(32'h3a93f466),
	.w7(32'h38ef36ab),
	.w8(32'hbbb4d518),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85fb5d),
	.w1(32'hbbb1be78),
	.w2(32'hbbc69669),
	.w3(32'hba9e4bcf),
	.w4(32'h3ad9fce8),
	.w5(32'hbbb6d090),
	.w6(32'hbb668eef),
	.w7(32'hbaba9856),
	.w8(32'hbbc8ea74),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea176f),
	.w1(32'hba988e7f),
	.w2(32'hba7745e5),
	.w3(32'hbb79a77d),
	.w4(32'hba17246e),
	.w5(32'h3b111067),
	.w6(32'hbc1dbffb),
	.w7(32'hbb18f465),
	.w8(32'h3b0c0bbf),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b779563),
	.w1(32'h3b0a8a91),
	.w2(32'h3aa2a27d),
	.w3(32'h3b4163c2),
	.w4(32'hbb309cae),
	.w5(32'hbbcb1d56),
	.w6(32'h3c2526b9),
	.w7(32'h3b8dc2d2),
	.w8(32'h3ad48fb6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53ce24),
	.w1(32'h3b836ec9),
	.w2(32'h3b1d6c9b),
	.w3(32'hbb08a1b9),
	.w4(32'h398e94a6),
	.w5(32'h3b893f64),
	.w6(32'hbb401734),
	.w7(32'h3ae8b016),
	.w8(32'h3b3a7636),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31e46d),
	.w1(32'hbab4fb5e),
	.w2(32'hba05925e),
	.w3(32'h3ad10f74),
	.w4(32'h3aa65910),
	.w5(32'hba5bf800),
	.w6(32'hb9762e97),
	.w7(32'hba1247e7),
	.w8(32'h3abc47d3),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af01e69),
	.w1(32'hbb9ece4c),
	.w2(32'hbbcd5d72),
	.w3(32'hbb81d285),
	.w4(32'hbb44c315),
	.w5(32'hbbc3177a),
	.w6(32'hbbd0b428),
	.w7(32'hbb0f3969),
	.w8(32'hbbc1f487),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd76ef),
	.w1(32'hbabf8056),
	.w2(32'hbb8972f7),
	.w3(32'h3a4c87bc),
	.w4(32'hbac868b4),
	.w5(32'hba09c8bb),
	.w6(32'hbaacbcc2),
	.w7(32'h3983d0da),
	.w8(32'h3a705c98),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22aaf0),
	.w1(32'hbba6f8c5),
	.w2(32'hbbdea75c),
	.w3(32'hbb40a068),
	.w4(32'hbbc1d769),
	.w5(32'hbb30ae56),
	.w6(32'hbb45d079),
	.w7(32'hbba2c593),
	.w8(32'hba25ce8a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aafbc),
	.w1(32'h39dc7ec6),
	.w2(32'h3b1323c2),
	.w3(32'h3b1535ee),
	.w4(32'h3b6ad5fa),
	.w5(32'h38036960),
	.w6(32'hbb044a59),
	.w7(32'h3b3ac4f2),
	.w8(32'hbaec2350),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a54e8),
	.w1(32'hbb009812),
	.w2(32'hbbc8faf3),
	.w3(32'hbaa5400d),
	.w4(32'hbb049fe5),
	.w5(32'hbac6d425),
	.w6(32'hbacbb605),
	.w7(32'hbb3d4df8),
	.w8(32'hbb162198),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a398d17),
	.w1(32'hbaf06d6a),
	.w2(32'h3b035da8),
	.w3(32'hbb8285cc),
	.w4(32'hbb1224a9),
	.w5(32'h3b9818c5),
	.w6(32'hbb3fc479),
	.w7(32'h38e32955),
	.w8(32'h3b8f4ca7),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afd3c7),
	.w1(32'hbac91e98),
	.w2(32'h3b066730),
	.w3(32'h3ac47fee),
	.w4(32'hb921076a),
	.w5(32'hbb04db60),
	.w6(32'h3aef0d87),
	.w7(32'hb9e33ebe),
	.w8(32'hbb37467d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ecf456),
	.w1(32'hb92710ab),
	.w2(32'hba56b01d),
	.w3(32'h3a02ac12),
	.w4(32'hbb09c658),
	.w5(32'hbb864d8f),
	.w6(32'h38d36fec),
	.w7(32'hbaa5e49b),
	.w8(32'hbaadfa5a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21651b),
	.w1(32'h3c4651d8),
	.w2(32'h3c5494e8),
	.w3(32'h3ae13f53),
	.w4(32'h3bd076fc),
	.w5(32'hb9c3b1c2),
	.w6(32'h3a9070d4),
	.w7(32'h3c651852),
	.w8(32'hba0e0a19),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e97af6),
	.w1(32'hbb0ab1f9),
	.w2(32'hbb62caf4),
	.w3(32'hb96c5bac),
	.w4(32'hbace357d),
	.w5(32'hbb7d08f0),
	.w6(32'hbaf7f6fd),
	.w7(32'hbb34ff5f),
	.w8(32'hbb3626b3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55765f),
	.w1(32'hbb823e77),
	.w2(32'hbbe8db53),
	.w3(32'h3a293d04),
	.w4(32'hbb0427b1),
	.w5(32'hbb7d2f68),
	.w6(32'hba5ec16e),
	.w7(32'hbadd1aeb),
	.w8(32'hbb903071),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba313c54),
	.w1(32'hbadc4a44),
	.w2(32'hbb65cc4e),
	.w3(32'hb963f983),
	.w4(32'hba35ebff),
	.w5(32'hbb02fe67),
	.w6(32'hbb2131ec),
	.w7(32'hbb3279fc),
	.w8(32'hbb87792f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9106d4f),
	.w1(32'hbab157ea),
	.w2(32'hba89396a),
	.w3(32'hba533d3c),
	.w4(32'h39c52ffd),
	.w5(32'h3a23e437),
	.w6(32'h39efeaba),
	.w7(32'hba389ad1),
	.w8(32'h3a5379cf),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba09972),
	.w1(32'hbbb4ed6b),
	.w2(32'hbbd47855),
	.w3(32'hbaec5602),
	.w4(32'hbb0bf3a2),
	.w5(32'hbb334913),
	.w6(32'hb9aa5b78),
	.w7(32'hba428b70),
	.w8(32'h39df31c7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad932c0),
	.w1(32'hbaa0190a),
	.w2(32'hb9a0ca53),
	.w3(32'hb99ea2a6),
	.w4(32'hbac006b9),
	.w5(32'hbaa41623),
	.w6(32'hbabecdee),
	.w7(32'hb86b77ca),
	.w8(32'hbb1d4613),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea5bf5),
	.w1(32'hbb661518),
	.w2(32'hbb8217cf),
	.w3(32'hbab9695d),
	.w4(32'hbb38be7c),
	.w5(32'hb9dd96f1),
	.w6(32'h39545d05),
	.w7(32'hba3addee),
	.w8(32'hba60da07),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f8e0c),
	.w1(32'hbb2f1ae0),
	.w2(32'hbb006b77),
	.w3(32'hba274f5d),
	.w4(32'hba6bdae6),
	.w5(32'hbb36ebb4),
	.w6(32'hba64e847),
	.w7(32'hb826f3b7),
	.w8(32'hba998532),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa759c),
	.w1(32'hb983292b),
	.w2(32'hba164e60),
	.w3(32'hb90a3479),
	.w4(32'hb9597819),
	.w5(32'h3a2195d5),
	.w6(32'hba86907a),
	.w7(32'hb99972be),
	.w8(32'h3a2f6930),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ed4a61),
	.w1(32'h391dafe1),
	.w2(32'hb96ac3e9),
	.w3(32'h39ca1ed9),
	.w4(32'h3982c5bb),
	.w5(32'hbb3f35d0),
	.w6(32'h3a85d0fc),
	.w7(32'h3a291934),
	.w8(32'hbb52c6f2),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19044f),
	.w1(32'hbb374fdb),
	.w2(32'hbb36ebc9),
	.w3(32'hbb038161),
	.w4(32'hbb01cc93),
	.w5(32'h384213b9),
	.w6(32'hbb61f8aa),
	.w7(32'hbb5428f2),
	.w8(32'hb99bf2bd),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374dbf8a),
	.w1(32'hba67290e),
	.w2(32'hba3fec93),
	.w3(32'h38d4db66),
	.w4(32'h3a6a2f91),
	.w5(32'hbb187d2f),
	.w6(32'hb9e6910a),
	.w7(32'hb9b4eeba),
	.w8(32'hbb033272),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a911b4a),
	.w1(32'h3b14b1dd),
	.w2(32'hba81f316),
	.w3(32'hba444c09),
	.w4(32'h3aad0ff8),
	.w5(32'hba155a34),
	.w6(32'hbb0cd7af),
	.w7(32'hba969a36),
	.w8(32'h3963f54f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f94d2),
	.w1(32'hbba248be),
	.w2(32'hbbf508c1),
	.w3(32'hbb60aaf9),
	.w4(32'hbb91fb61),
	.w5(32'hbc07eb7f),
	.w6(32'hb9d7d426),
	.w7(32'hbae84f85),
	.w8(32'hbb8d07c4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850bfa),
	.w1(32'hbba8e37c),
	.w2(32'hbbd91ec5),
	.w3(32'hba8b129a),
	.w4(32'hba73a956),
	.w5(32'hbb3d99aa),
	.w6(32'hbad139eb),
	.w7(32'hbb1b2bfe),
	.w8(32'hba794857),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37ce98),
	.w1(32'hbba54919),
	.w2(32'hbbb90fce),
	.w3(32'hbb320fdc),
	.w4(32'hbb5dcbe0),
	.w5(32'hbba4f62f),
	.w6(32'hb96f1dfa),
	.w7(32'hbafa0cff),
	.w8(32'hbacc8842),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a614016),
	.w1(32'hb889446a),
	.w2(32'h3a98497d),
	.w3(32'hba890038),
	.w4(32'h3aa6a51c),
	.w5(32'hbab0e030),
	.w6(32'hba7dfd76),
	.w7(32'hb956117c),
	.w8(32'hb8e609df),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cdcca),
	.w1(32'hba940083),
	.w2(32'hb91fd4ce),
	.w3(32'hba693ccc),
	.w4(32'hba1b67c2),
	.w5(32'h3b10562b),
	.w6(32'h39b60141),
	.w7(32'hba3cccc5),
	.w8(32'h3aed14f3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc41e5),
	.w1(32'h3a32398c),
	.w2(32'h3a24216d),
	.w3(32'h3ab9ad48),
	.w4(32'h3ad81950),
	.w5(32'h3b10e014),
	.w6(32'h3aa3a6e3),
	.w7(32'h3ad7a955),
	.w8(32'h3a8d63ab),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a082f),
	.w1(32'hba906f09),
	.w2(32'h3998fda7),
	.w3(32'h3aa58ead),
	.w4(32'hba0178c4),
	.w5(32'hb9cd2baf),
	.w6(32'h3ac4afe5),
	.w7(32'h3a9c7184),
	.w8(32'hb9e64124),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc52297),
	.w1(32'hbbe3c772),
	.w2(32'hbbf9ba50),
	.w3(32'hbb5ffb22),
	.w4(32'hbb26a80a),
	.w5(32'hbb871beb),
	.w6(32'hbb8ce6ed),
	.w7(32'hbb108762),
	.w8(32'hbb2a2587),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba063d3d),
	.w1(32'hbb19253e),
	.w2(32'hbb26d61d),
	.w3(32'hba3ff741),
	.w4(32'hb98e01b5),
	.w5(32'hba97a50e),
	.w6(32'hbb08916d),
	.w7(32'hbae4bb12),
	.w8(32'h39cdde00),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385a846a),
	.w1(32'h39d0e260),
	.w2(32'hba0e7a03),
	.w3(32'hba149d01),
	.w4(32'h39f31384),
	.w5(32'hbaa8b4a6),
	.w6(32'h3aca6f15),
	.w7(32'h3a1b4e5d),
	.w8(32'hba673c13),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb992cb9),
	.w1(32'hbb5051b7),
	.w2(32'hbabbb74e),
	.w3(32'hbb368537),
	.w4(32'hbac6f14c),
	.w5(32'hbb90614a),
	.w6(32'hbad4ddca),
	.w7(32'hba4fafac),
	.w8(32'hbb733b74),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4e09e),
	.w1(32'hbae4176e),
	.w2(32'hba42ddd4),
	.w3(32'hbb2c9a95),
	.w4(32'hbacf78b4),
	.w5(32'hba4da4bb),
	.w6(32'hbaad3194),
	.w7(32'hbacb5bbd),
	.w8(32'hb9f2117e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebf537),
	.w1(32'hba8fb42e),
	.w2(32'hbae6824f),
	.w3(32'hba7d288e),
	.w4(32'h39d59a29),
	.w5(32'hbb0c3a46),
	.w6(32'hba605fa3),
	.w7(32'hbabeea85),
	.w8(32'hbb69fdf0),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1a89f),
	.w1(32'hba64ba27),
	.w2(32'hb9d163ae),
	.w3(32'hba378973),
	.w4(32'hb98f1a0c),
	.w5(32'hb848f31d),
	.w6(32'hba8b542a),
	.w7(32'hba9f537a),
	.w8(32'hb90df7fb),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3b2ae),
	.w1(32'hbbd04b44),
	.w2(32'hbc090d10),
	.w3(32'hbbd7af69),
	.w4(32'hbb8b160e),
	.w5(32'hbb751c11),
	.w6(32'hba857dd5),
	.w7(32'h3b3bde7a),
	.w8(32'h3a9ca3fc),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7efff),
	.w1(32'hb9869f62),
	.w2(32'hb8e80203),
	.w3(32'h3a17b638),
	.w4(32'h3accf145),
	.w5(32'h39b313b4),
	.w6(32'h3a37ce0b),
	.w7(32'h3abbc7c8),
	.w8(32'h3a5c8f95),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00b7dd),
	.w1(32'h3b99eb64),
	.w2(32'h3ae2f238),
	.w3(32'h3b2a66bb),
	.w4(32'h3b689936),
	.w5(32'h3b435c9d),
	.w6(32'hbad5b1af),
	.w7(32'h395b1bb7),
	.w8(32'hba33b470),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule