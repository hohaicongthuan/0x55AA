module layer_10_featuremap_44(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affe2e9),
	.w1(32'h3bfc0b80),
	.w2(32'hbb49b095),
	.w3(32'hba79eec2),
	.w4(32'h3ad12a1f),
	.w5(32'hbbc22cf6),
	.w6(32'hbb01bb7e),
	.w7(32'hbb5fa15c),
	.w8(32'hbc102a58),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96228e),
	.w1(32'h395b723c),
	.w2(32'hbc104f4d),
	.w3(32'h3b1042da),
	.w4(32'hbae78eba),
	.w5(32'hbbe02b32),
	.w6(32'hbba25791),
	.w7(32'hbb7a8cf3),
	.w8(32'hbc209366),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dbf16),
	.w1(32'h396938c7),
	.w2(32'h3b81475e),
	.w3(32'hbacb4acf),
	.w4(32'hb8ca8ba5),
	.w5(32'hbafd25fd),
	.w6(32'hbb092d27),
	.w7(32'hb954b640),
	.w8(32'h3b17102f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f143a),
	.w1(32'h3b5dd16e),
	.w2(32'hbb1319e4),
	.w3(32'h3ad54d83),
	.w4(32'hb9bb88f2),
	.w5(32'hbbccc984),
	.w6(32'hbbe84989),
	.w7(32'hbb858ba7),
	.w8(32'hba986c2d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6203a),
	.w1(32'hbae33b93),
	.w2(32'hbb9e0876),
	.w3(32'hbba85aba),
	.w4(32'hbbca9376),
	.w5(32'hbc15a746),
	.w6(32'hbbada793),
	.w7(32'hbb3c535a),
	.w8(32'hbc1f14a0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9cd55),
	.w1(32'h3bc21642),
	.w2(32'hbc62b486),
	.w3(32'hbba9ee32),
	.w4(32'hba8c4124),
	.w5(32'h3a20d2bb),
	.w6(32'hbbb1be62),
	.w7(32'h3b709132),
	.w8(32'hb9bd21b9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc874a1d),
	.w1(32'hbccea3c4),
	.w2(32'h3c094fa8),
	.w3(32'h3c158ca7),
	.w4(32'hbbbecf62),
	.w5(32'h3c1db5a7),
	.w6(32'hbb77362f),
	.w7(32'hbb0f9bfa),
	.w8(32'h3c25befa),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7be4b),
	.w1(32'h3be46a48),
	.w2(32'h3c2cb648),
	.w3(32'h3b2176ab),
	.w4(32'hbcaa0859),
	.w5(32'hbbac9ff6),
	.w6(32'hbc3087de),
	.w7(32'h3c4c3657),
	.w8(32'hbced3801),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d70f0),
	.w1(32'h3c348595),
	.w2(32'h3b10cace),
	.w3(32'h3c3c1722),
	.w4(32'h3b5e0c51),
	.w5(32'h3adcf62b),
	.w6(32'h3babe2f7),
	.w7(32'h3a294c45),
	.w8(32'h3b7442a6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb209d8b),
	.w1(32'h3bdb2fbf),
	.w2(32'h3c03b286),
	.w3(32'hbb77d4b4),
	.w4(32'hbad19057),
	.w5(32'hbaf964a0),
	.w6(32'hba76c910),
	.w7(32'hbb82ccac),
	.w8(32'h3c8bf4ff),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce93ebe),
	.w1(32'hbc9fab98),
	.w2(32'h3b268155),
	.w3(32'hbd26e87e),
	.w4(32'hbd0065fc),
	.w5(32'hbaad72f3),
	.w6(32'hbc00352d),
	.w7(32'hbad52784),
	.w8(32'hbbab9461),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a2c44),
	.w1(32'h3b95acc3),
	.w2(32'h3cd5f428),
	.w3(32'hbc22aadb),
	.w4(32'hbbaa7d78),
	.w5(32'h3c602ce7),
	.w6(32'hbc9548be),
	.w7(32'hbb9611de),
	.w8(32'h3bad748e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca875d5),
	.w1(32'h3cd76de8),
	.w2(32'h3c4fd065),
	.w3(32'h3cd128cf),
	.w4(32'h3cddd569),
	.w5(32'h3c06d48a),
	.w6(32'h3c060415),
	.w7(32'h3c16f7e4),
	.w8(32'h3bbd5d9b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb409e86),
	.w1(32'h39f8f157),
	.w2(32'h3bb2b757),
	.w3(32'h3bb73483),
	.w4(32'h3bf4ce02),
	.w5(32'hbb3a1f94),
	.w6(32'h3b92d9fa),
	.w7(32'h3c0323a1),
	.w8(32'h3a3eeb12),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23ec9a),
	.w1(32'hba85dd22),
	.w2(32'hbc0fb1ec),
	.w3(32'hbc0e4d64),
	.w4(32'hbc048f12),
	.w5(32'hbc07ce49),
	.w6(32'hbbc223c9),
	.w7(32'hbbd31d32),
	.w8(32'hbb71d301),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37270f),
	.w1(32'h3b1f0deb),
	.w2(32'hbb36bb1e),
	.w3(32'hbc0418c6),
	.w4(32'hbb4664f4),
	.w5(32'hbc22e6e2),
	.w6(32'hba5c70b4),
	.w7(32'hbc37776b),
	.w8(32'h3c4417b2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0fd4bb),
	.w1(32'hbce252fb),
	.w2(32'h3958c85b),
	.w3(32'hbd403c94),
	.w4(32'hbd20af62),
	.w5(32'h3b1c4659),
	.w6(32'hbc4f4ef8),
	.w7(32'hbc09bc23),
	.w8(32'h3a1bb682),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f36d30),
	.w1(32'h3c85de09),
	.w2(32'h3d02b64a),
	.w3(32'hbb87bded),
	.w4(32'h3c0134e6),
	.w5(32'h3caed67d),
	.w6(32'hbb0be8c7),
	.w7(32'h3adc511d),
	.w8(32'h3b455fab),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb644572),
	.w1(32'h3b81c168),
	.w2(32'h3c5cbf19),
	.w3(32'hbb43b3ad),
	.w4(32'hbaa46071),
	.w5(32'h3c896d2d),
	.w6(32'h39f5c24e),
	.w7(32'h3b7e0451),
	.w8(32'h3b92f1cc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5d268),
	.w1(32'h3bb8a7e0),
	.w2(32'hbb2afd1c),
	.w3(32'hbb97e39a),
	.w4(32'h3ab7f59b),
	.w5(32'hbb9066ab),
	.w6(32'hbb0ca4c2),
	.w7(32'h3b0032ee),
	.w8(32'hbbc4c94d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0b2ec),
	.w1(32'hba80a24b),
	.w2(32'h3acaf008),
	.w3(32'hbb86ff4e),
	.w4(32'hbab6a8dd),
	.w5(32'hbb7b4301),
	.w6(32'hbbae8992),
	.w7(32'hbba4f857),
	.w8(32'hbba91ae3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb639ab2),
	.w1(32'hbb5cb749),
	.w2(32'hbbbbd84d),
	.w3(32'hbbaeee13),
	.w4(32'hbaaaa608),
	.w5(32'hbb634554),
	.w6(32'hbbdfe5d4),
	.w7(32'hbb3b4d63),
	.w8(32'h3b0bd02c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7de6fd),
	.w1(32'h3c218aea),
	.w2(32'h3cf70de8),
	.w3(32'hbc428e16),
	.w4(32'hba6d8a30),
	.w5(32'h3bd2e9c4),
	.w6(32'hbc91b260),
	.w7(32'hbc5a4a7a),
	.w8(32'h3c38b4ad),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7c264),
	.w1(32'h3c89ba60),
	.w2(32'h3a37685b),
	.w3(32'hbab4a52d),
	.w4(32'h3bc83ec7),
	.w5(32'h3b199fc3),
	.w6(32'h3a9131e2),
	.w7(32'h3c087034),
	.w8(32'hbaae6c0e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab53e59),
	.w1(32'hbc4f5318),
	.w2(32'hbd01f5b4),
	.w3(32'hbac808f8),
	.w4(32'hba8e0e20),
	.w5(32'hbc70f38f),
	.w6(32'hbb29aa77),
	.w7(32'hbb7d3b36),
	.w8(32'hbb35e304),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02d785),
	.w1(32'hbb8d9fa1),
	.w2(32'h3a15e83f),
	.w3(32'hbba323d2),
	.w4(32'hbbb4efa4),
	.w5(32'h3b9c0918),
	.w6(32'h39fc6820),
	.w7(32'hbbae8bd4),
	.w8(32'hba199d93),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d48945),
	.w1(32'h3b1bd60a),
	.w2(32'h38e6770e),
	.w3(32'hbacc77fd),
	.w4(32'h3acf7c2e),
	.w5(32'hb8894b01),
	.w6(32'hbb8f9049),
	.w7(32'hba999400),
	.w8(32'h3a6045a3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d2b76),
	.w1(32'h3cd85214),
	.w2(32'h3c8b02d7),
	.w3(32'hbbae7321),
	.w4(32'h3c390143),
	.w5(32'h3ce22f97),
	.w6(32'h3cdcdce8),
	.w7(32'h3c52c67b),
	.w8(32'h3ce0d492),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ce0d7),
	.w1(32'h3b0e6206),
	.w2(32'hbb0611de),
	.w3(32'hbb57f476),
	.w4(32'hbc2a9f8e),
	.w5(32'hba8e5f49),
	.w6(32'hbb9f2c84),
	.w7(32'hbbd9c419),
	.w8(32'hbb1285b0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e4845),
	.w1(32'h3b21450b),
	.w2(32'hbc05992c),
	.w3(32'hbbfadfd1),
	.w4(32'h3ba4b532),
	.w5(32'h3bc38e3a),
	.w6(32'h3c377b3f),
	.w7(32'h3bcce2fd),
	.w8(32'h3be163f5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f89d9),
	.w1(32'hbbc01f1a),
	.w2(32'h3bafe676),
	.w3(32'h3aa89f26),
	.w4(32'hbb96ff49),
	.w5(32'h3c4502b1),
	.w6(32'h3b182ee8),
	.w7(32'hbb5faf17),
	.w8(32'hbb26d883),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8281b),
	.w1(32'h3c3d763a),
	.w2(32'hbbbebaea),
	.w3(32'h3c154c18),
	.w4(32'h3b4979e4),
	.w5(32'h3b962204),
	.w6(32'h3bd18da8),
	.w7(32'hba9a3d72),
	.w8(32'h3b798128),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc287161),
	.w1(32'hbb3fc0ab),
	.w2(32'h3c393c0c),
	.w3(32'hbbab6250),
	.w4(32'h3be5fbf3),
	.w5(32'h3c6a3eae),
	.w6(32'h3c2a84a2),
	.w7(32'h3be9d34f),
	.w8(32'h3c2b7b18),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c004684),
	.w1(32'h3b669657),
	.w2(32'hbbf0da85),
	.w3(32'h3bbbcd47),
	.w4(32'h3b2d8607),
	.w5(32'hbc2775ad),
	.w6(32'h3b9abf03),
	.w7(32'h3ad96252),
	.w8(32'h3b9fb45e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72817c),
	.w1(32'hbc868a13),
	.w2(32'h3b55d9e6),
	.w3(32'hbc548884),
	.w4(32'hbc2242ae),
	.w5(32'h3ad318b8),
	.w6(32'h3b8cf6de),
	.w7(32'hbbc1b2ab),
	.w8(32'h3ad58cd5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba041e60),
	.w1(32'h3b02c0ac),
	.w2(32'h3c8f663f),
	.w3(32'hba7deecb),
	.w4(32'h3b69f70d),
	.w5(32'h3badd44a),
	.w6(32'hbc2e6cb9),
	.w7(32'h3a01d5ca),
	.w8(32'hbb763b2c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a0b92),
	.w1(32'hbcd18e71),
	.w2(32'h3c4ee1d0),
	.w3(32'hbbde8282),
	.w4(32'hbcc07814),
	.w5(32'hbca591eb),
	.w6(32'hbcb26f7c),
	.w7(32'hbc1b3d0c),
	.w8(32'hbbc7b4d8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1c57a),
	.w1(32'h3bb61cef),
	.w2(32'hbd10a63b),
	.w3(32'hbc9ad6ac),
	.w4(32'h3b3a5145),
	.w5(32'hbca7a7ed),
	.w6(32'hbc1a7d78),
	.w7(32'h3aa254de),
	.w8(32'hbc3bc61c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca25393),
	.w1(32'h3c2b4b30),
	.w2(32'h3c089e91),
	.w3(32'hba70685c),
	.w4(32'h3c98ddaa),
	.w5(32'h3c96f87c),
	.w6(32'h3bbd15e0),
	.w7(32'h3c2812ac),
	.w8(32'h3c36fa44),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2122d9),
	.w1(32'hbc4879f4),
	.w2(32'hbc22e11d),
	.w3(32'h3cc867fb),
	.w4(32'hba2f0146),
	.w5(32'hbba40caa),
	.w6(32'h3ca143bb),
	.w7(32'h3c03b63d),
	.w8(32'hbaf5dda6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea59b1),
	.w1(32'hbc3a76aa),
	.w2(32'h3b33b5d0),
	.w3(32'h3b817c43),
	.w4(32'hbc49abc7),
	.w5(32'h3af08420),
	.w6(32'h3b8d7553),
	.w7(32'hbbc406b6),
	.w8(32'h3bac412e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba23223),
	.w1(32'h3b241f90),
	.w2(32'hba54e018),
	.w3(32'h3be00a4e),
	.w4(32'h3c237b45),
	.w5(32'hbbb87b9a),
	.w6(32'h3b8297fe),
	.w7(32'h3c5dd6c6),
	.w8(32'hbb4945d2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae9931),
	.w1(32'hbbef59f9),
	.w2(32'h3b9b17d2),
	.w3(32'h3bb6ad4b),
	.w4(32'h3b986f23),
	.w5(32'h3a44203f),
	.w6(32'hbb4a9082),
	.w7(32'h3b929003),
	.w8(32'h3b3f07d2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41e9cf),
	.w1(32'h3cd5a740),
	.w2(32'h3c852573),
	.w3(32'hbbc65d93),
	.w4(32'h3c80add2),
	.w5(32'h3c8e8161),
	.w6(32'h3baeefab),
	.w7(32'h38e31980),
	.w8(32'h3c16afbb),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec1693),
	.w1(32'hbc0fc74a),
	.w2(32'hbbca163c),
	.w3(32'hbc1e5b0a),
	.w4(32'hbc9a640d),
	.w5(32'h3ba89ee3),
	.w6(32'hbbf8054b),
	.w7(32'hbcb588eb),
	.w8(32'h3c34ff1b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd565fb),
	.w1(32'hbb13c02b),
	.w2(32'hb9068250),
	.w3(32'h3c6737f6),
	.w4(32'h3bde9d48),
	.w5(32'h3b13bce3),
	.w6(32'hbb6f72bd),
	.w7(32'hbb1d507d),
	.w8(32'hbc85b02e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56db78),
	.w1(32'hbaefd9b2),
	.w2(32'hbc90fc9d),
	.w3(32'h3c26c71c),
	.w4(32'h3bbceaa1),
	.w5(32'hbc922d1c),
	.w6(32'h3c178279),
	.w7(32'hbbb61658),
	.w8(32'hbcc44f4c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc8d9fe),
	.w1(32'h3b21cb16),
	.w2(32'h3d113d40),
	.w3(32'hbbe03e03),
	.w4(32'h3c295f2a),
	.w5(32'h3cabd532),
	.w6(32'hbc0219f8),
	.w7(32'h3b5654c3),
	.w8(32'h3bb9a04b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1cc00),
	.w1(32'h3bffcb26),
	.w2(32'hba41e9d8),
	.w3(32'hba1c7fc9),
	.w4(32'h3be3b1ef),
	.w5(32'hbc81234d),
	.w6(32'h3b5367c4),
	.w7(32'h3bee0e12),
	.w8(32'hbc10b5a6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02d889),
	.w1(32'h3bfe6dd1),
	.w2(32'h3ae77515),
	.w3(32'hb8e117d1),
	.w4(32'h3c029a6f),
	.w5(32'h3b502fb2),
	.w6(32'hbab22ef9),
	.w7(32'h3b92f6b9),
	.w8(32'h38182cf7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d96d3),
	.w1(32'hbb1ec871),
	.w2(32'hbc3cd6bb),
	.w3(32'hbbdce51e),
	.w4(32'h39836f14),
	.w5(32'hbc8fd5e3),
	.w6(32'h3ad2d912),
	.w7(32'h3a47efb9),
	.w8(32'hbb890a57),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c125d8f),
	.w1(32'h39761539),
	.w2(32'h3b40574d),
	.w3(32'h3c1b0e3a),
	.w4(32'h3b3f29f1),
	.w5(32'h3b910ea0),
	.w6(32'h3ba6e931),
	.w7(32'hbc0d5f39),
	.w8(32'h3bbbbcef),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba28ba5),
	.w1(32'h3b09f620),
	.w2(32'h3b05157d),
	.w3(32'h3b764f77),
	.w4(32'h3c54cd80),
	.w5(32'h3bc46161),
	.w6(32'h3a9a1383),
	.w7(32'h3c19e35e),
	.w8(32'h3a86ce04),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c732d),
	.w1(32'h3c94cc68),
	.w2(32'h3d27ed34),
	.w3(32'h39ac6285),
	.w4(32'h3b83fa88),
	.w5(32'h3c7c657a),
	.w6(32'hbb5c6ea1),
	.w7(32'hbbbe8292),
	.w8(32'h3bd26ce0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef8bfd),
	.w1(32'h3bdb3638),
	.w2(32'h3bd62bab),
	.w3(32'hbc2ba20a),
	.w4(32'hbc71ee66),
	.w5(32'h3be8f369),
	.w6(32'h38de7359),
	.w7(32'h39e3134f),
	.w8(32'hb7b84672),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1422ad),
	.w1(32'hbc231a34),
	.w2(32'hbbab8d20),
	.w3(32'h3ba80a71),
	.w4(32'hba44f109),
	.w5(32'h3c163a65),
	.w6(32'h3a01e4f9),
	.w7(32'hb9f5e2b7),
	.w8(32'h3b4226a7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb399d0),
	.w1(32'hbbf56918),
	.w2(32'h3bc930fc),
	.w3(32'h3ab3c8d6),
	.w4(32'hbbc57935),
	.w5(32'h3b35b475),
	.w6(32'h3b191b5f),
	.w7(32'hbb9dc5a9),
	.w8(32'h3ba1ea3a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7fe7a),
	.w1(32'hbbe9ea53),
	.w2(32'h3a54384c),
	.w3(32'h3b812f94),
	.w4(32'hbc4cb173),
	.w5(32'hb9ca5fdd),
	.w6(32'h3beb5a7d),
	.w7(32'hbb830997),
	.w8(32'hb9f2a9d0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11f411),
	.w1(32'hb93cacfb),
	.w2(32'h3bc79a48),
	.w3(32'hbb42ddc8),
	.w4(32'hbb6eee11),
	.w5(32'h3a70e620),
	.w6(32'hba91fa0f),
	.w7(32'hbad47613),
	.w8(32'h3b43cc7e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6da30),
	.w1(32'h3b22c8de),
	.w2(32'h3c2823bf),
	.w3(32'h3b9f1cdc),
	.w4(32'h3901977b),
	.w5(32'hbc0ae9c9),
	.w6(32'hbab7b8fa),
	.w7(32'hba173e45),
	.w8(32'h3ad491a2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64fc3b),
	.w1(32'h3ca32058),
	.w2(32'h3b956cff),
	.w3(32'h3bad0676),
	.w4(32'h3c4048b8),
	.w5(32'h3be94fd1),
	.w6(32'h3c4a10e1),
	.w7(32'h3c171cc8),
	.w8(32'h3b80abbb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0827f3),
	.w1(32'h3b1c2dd7),
	.w2(32'h3bb1a5e0),
	.w3(32'h39f10292),
	.w4(32'h3b5fe78d),
	.w5(32'hba4df55f),
	.w6(32'h3c115055),
	.w7(32'hbb52925a),
	.w8(32'h3b52e6ed),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04f91c),
	.w1(32'h3b59a6ad),
	.w2(32'h3aca3965),
	.w3(32'hbaaca93e),
	.w4(32'h3b4f60a0),
	.w5(32'h3b3c0f52),
	.w6(32'hbc07a7c8),
	.w7(32'h3baad0a3),
	.w8(32'h3bb1850b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ec62b),
	.w1(32'hbc39420f),
	.w2(32'h3b9cedce),
	.w3(32'hbc121b15),
	.w4(32'hbc925f4b),
	.w5(32'h3c490ca6),
	.w6(32'hbac8a67f),
	.w7(32'hbc1e6787),
	.w8(32'h3b5ede5e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb631e5),
	.w1(32'h3b98391b),
	.w2(32'hba8a3aac),
	.w3(32'h3b838dc3),
	.w4(32'h3c0f2704),
	.w5(32'h3bd007c8),
	.w6(32'h3bb6a4fe),
	.w7(32'h3be01c48),
	.w8(32'h3c0aafdc),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19eefc),
	.w1(32'hbc2c64cf),
	.w2(32'h3baa3b51),
	.w3(32'hbbe514c5),
	.w4(32'hbc614554),
	.w5(32'h3b935185),
	.w6(32'h3ac2ed48),
	.w7(32'hbbf06533),
	.w8(32'h3bb6d45c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30974f),
	.w1(32'h3cc0ac6c),
	.w2(32'h3d184e56),
	.w3(32'hbd127ea0),
	.w4(32'hbbafdd9e),
	.w5(32'h3c6fa631),
	.w6(32'h3bd97dda),
	.w7(32'h3c53420e),
	.w8(32'h3c27e2c9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52e6eb),
	.w1(32'hbb8b62bd),
	.w2(32'h3ba961da),
	.w3(32'h3c2bc97c),
	.w4(32'h3c1525af),
	.w5(32'h3c9313af),
	.w6(32'hbc9fb4d8),
	.w7(32'hbbc48376),
	.w8(32'hbb3a0634),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07f99),
	.w1(32'h3c128692),
	.w2(32'h3bd84298),
	.w3(32'h3b81d5ef),
	.w4(32'h3c853d7c),
	.w5(32'hba98441c),
	.w6(32'h3baf5b34),
	.w7(32'h3bb656e7),
	.w8(32'hbbc5fa04),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99fcb1),
	.w1(32'hbbdc9a80),
	.w2(32'hbcb930ce),
	.w3(32'hbc596bf5),
	.w4(32'hbbb05a73),
	.w5(32'hbca6be77),
	.w6(32'hbc78bcd6),
	.w7(32'hbbe3cdbe),
	.w8(32'hbbe22f1e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72990d),
	.w1(32'h3b320031),
	.w2(32'h3b7c604b),
	.w3(32'h3b25da61),
	.w4(32'h3be53159),
	.w5(32'h3c5b20a1),
	.w6(32'hb8b452f3),
	.w7(32'h3b847b68),
	.w8(32'h3c34566d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8e586),
	.w1(32'hbc190869),
	.w2(32'h3afc53d3),
	.w3(32'h3c1190ab),
	.w4(32'hbc9885d8),
	.w5(32'h3aa9359e),
	.w6(32'h3c32d7b1),
	.w7(32'hbc59a437),
	.w8(32'hbb548ad9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c367d),
	.w1(32'hbbe44eb3),
	.w2(32'h3c304d46),
	.w3(32'h3c7872b7),
	.w4(32'hbb3c5b60),
	.w5(32'h3c484ba9),
	.w6(32'h3c50f2c2),
	.w7(32'h384cd320),
	.w8(32'h3c938437),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82ddd3),
	.w1(32'hbb604f3e),
	.w2(32'h3c587627),
	.w3(32'hbb60f907),
	.w4(32'hbb49432f),
	.w5(32'h3c26d454),
	.w6(32'h3bc5f01d),
	.w7(32'h3bd8419b),
	.w8(32'h3c0283f3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04178c),
	.w1(32'h3be60f62),
	.w2(32'h3b5af750),
	.w3(32'hbb1f3857),
	.w4(32'h3bb0b890),
	.w5(32'h3beaafd5),
	.w6(32'h3952b3af),
	.w7(32'h3c0d939d),
	.w8(32'h3b8ed090),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97173e),
	.w1(32'h3c19e267),
	.w2(32'h3c45fe91),
	.w3(32'h3c3fb728),
	.w4(32'h3ba3a462),
	.w5(32'h3c2d941a),
	.w6(32'h3c124f3d),
	.w7(32'h3bac9302),
	.w8(32'h3c2617ff),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc106c18),
	.w1(32'h3b5b1de1),
	.w2(32'h3c5cda25),
	.w3(32'h3b26dd8a),
	.w4(32'hba78bc2b),
	.w5(32'h3c6367fb),
	.w6(32'hbb393fc2),
	.w7(32'h3c251ed5),
	.w8(32'hba42348f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef69d3),
	.w1(32'hbb6b154a),
	.w2(32'hbbcacf0b),
	.w3(32'hbaa9b163),
	.w4(32'hbba1f394),
	.w5(32'h3b335a1f),
	.w6(32'hba97665e),
	.w7(32'hbbf190d0),
	.w8(32'hbb9e0e17),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52b47b),
	.w1(32'hbbe54b96),
	.w2(32'h3be79bfe),
	.w3(32'h3ca1c955),
	.w4(32'hbc1d6325),
	.w5(32'h3b614748),
	.w6(32'h3c1bd17f),
	.w7(32'hbb3daefd),
	.w8(32'h3a451a07),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfbfd5),
	.w1(32'h3b945d5f),
	.w2(32'h3c26bc05),
	.w3(32'hbbd46500),
	.w4(32'hbaa36783),
	.w5(32'hbac86507),
	.w6(32'hb98ae68a),
	.w7(32'h3ba366c9),
	.w8(32'hbb1693eb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb5666),
	.w1(32'h3c1b60dd),
	.w2(32'h3b33194e),
	.w3(32'h3a6cfad7),
	.w4(32'h3c71bf66),
	.w5(32'h3bd6707d),
	.w6(32'h3b7b098d),
	.w7(32'h3bf59b39),
	.w8(32'h3ba77438),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb206782),
	.w1(32'h3bc4a0cd),
	.w2(32'h3c022c2b),
	.w3(32'hbb91d712),
	.w4(32'hbae46d4e),
	.w5(32'hbad83a1d),
	.w6(32'hbad67be5),
	.w7(32'hbb2f56fe),
	.w8(32'hbc0c7709),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6efbc),
	.w1(32'hba313f6b),
	.w2(32'hbb788e1e),
	.w3(32'h3a65c225),
	.w4(32'h3b0890b4),
	.w5(32'hba8f325d),
	.w6(32'h3b08a9ea),
	.w7(32'h3aa5d7aa),
	.w8(32'hba52272b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa25a4),
	.w1(32'hbbced4e8),
	.w2(32'hba408a41),
	.w3(32'h3c1c3723),
	.w4(32'h3ba49246),
	.w5(32'h3b35f322),
	.w6(32'hbadd5dad),
	.w7(32'h3b5fb706),
	.w8(32'hbb964310),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23c96e),
	.w1(32'hbbcf8d62),
	.w2(32'hbc3698e5),
	.w3(32'h3bf47882),
	.w4(32'hbb8e0051),
	.w5(32'h3bed3f65),
	.w6(32'hbb0bd8b6),
	.w7(32'hbbcc222e),
	.w8(32'h3c526f04),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8156d0),
	.w1(32'hbcd06c9a),
	.w2(32'h398112c8),
	.w3(32'hbb056959),
	.w4(32'hbcf28c2f),
	.w5(32'h3bbd29ad),
	.w6(32'hbb99c7fe),
	.w7(32'hbce88679),
	.w8(32'h3bb6195f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57b616),
	.w1(32'hbc36b079),
	.w2(32'hbbdb13e6),
	.w3(32'h390af0a8),
	.w4(32'hbc6cb568),
	.w5(32'hbb985124),
	.w6(32'h3b7f7498),
	.w7(32'hbc272278),
	.w8(32'h3a3b61ed),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf7fa3),
	.w1(32'hba883161),
	.w2(32'h3ab4f200),
	.w3(32'h3b3b610e),
	.w4(32'hb9a59de1),
	.w5(32'hba12b734),
	.w6(32'h3a9cc04a),
	.w7(32'h3a5904de),
	.w8(32'h3c0e9069),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb335a25),
	.w1(32'hbb715202),
	.w2(32'h3ba7f0a4),
	.w3(32'hba69411f),
	.w4(32'hbaa562b0),
	.w5(32'h3bf21720),
	.w6(32'hb6a9cbe6),
	.w7(32'hbb25d379),
	.w8(32'hbba89a10),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b6e99),
	.w1(32'h3c1a28a3),
	.w2(32'h3c9d0d48),
	.w3(32'h3b8b0f2e),
	.w4(32'h3b525672),
	.w5(32'h3c876446),
	.w6(32'hbb6d745b),
	.w7(32'hbb166e0c),
	.w8(32'hba503916),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca272f),
	.w1(32'h3c9237bc),
	.w2(32'h3ba8085d),
	.w3(32'hbc665924),
	.w4(32'h3b16c441),
	.w5(32'hbc03f469),
	.w6(32'h38d746fd),
	.w7(32'hbb0dacf1),
	.w8(32'hbbeb124c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb662b25),
	.w1(32'h3ab65659),
	.w2(32'h3cdef794),
	.w3(32'hbd253993),
	.w4(32'hbcdafb89),
	.w5(32'h3bab814f),
	.w6(32'hbc92036f),
	.w7(32'hbb9ac8a2),
	.w8(32'h3c7dd949),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2af456),
	.w1(32'h3b5a0d33),
	.w2(32'h3a7cab88),
	.w3(32'h38dad827),
	.w4(32'h3b6c97ca),
	.w5(32'hbb36a926),
	.w6(32'hba354558),
	.w7(32'hb9c83be4),
	.w8(32'hbb377a46),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c204e),
	.w1(32'h3c051396),
	.w2(32'h3c72ad03),
	.w3(32'hbc0fdb27),
	.w4(32'h3a48f6fb),
	.w5(32'h3c2735c0),
	.w6(32'hbaba03e4),
	.w7(32'h3b59ae87),
	.w8(32'h3c9039ef),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6d501),
	.w1(32'h3b09b129),
	.w2(32'h3aa6d08e),
	.w3(32'h3bbe96c9),
	.w4(32'h3b347a1c),
	.w5(32'hbc2b5c97),
	.w6(32'h3c535301),
	.w7(32'h3b8ab7fd),
	.w8(32'h3ae6b1d7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0247d),
	.w1(32'hbb9a0255),
	.w2(32'hbc8e4189),
	.w3(32'hbbdbbca2),
	.w4(32'h3ac3160c),
	.w5(32'hbc2bcf1c),
	.w6(32'h3c313b00),
	.w7(32'hbbf0b4f0),
	.w8(32'hbc65f2e2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39498ab7),
	.w1(32'hb9f9cf5e),
	.w2(32'hbb69a2ee),
	.w3(32'h3af94e4d),
	.w4(32'hbaf5cbd7),
	.w5(32'h3b3fef7e),
	.w6(32'hbbd979a4),
	.w7(32'hbaa94ed8),
	.w8(32'hbba8fab3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4c373),
	.w1(32'h3b7b19c0),
	.w2(32'h3c97936b),
	.w3(32'h3c68f831),
	.w4(32'h3c3810ba),
	.w5(32'h3c5721ab),
	.w6(32'hbbc33456),
	.w7(32'h3b8a6d03),
	.w8(32'hbb81cd65),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43865d),
	.w1(32'hba7f70ac),
	.w2(32'h3cda6fd6),
	.w3(32'hbcc95f30),
	.w4(32'hbc62b513),
	.w5(32'hbc44f910),
	.w6(32'hbc8c216b),
	.w7(32'hbc19681c),
	.w8(32'hbbae35b3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceec11b),
	.w1(32'hbbc7b734),
	.w2(32'hbb806487),
	.w3(32'h3b882646),
	.w4(32'h3c619c73),
	.w5(32'hbc855bcd),
	.w6(32'hbd077263),
	.w7(32'hbaac4dae),
	.w8(32'hbc830223),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18762d),
	.w1(32'hbb921f1d),
	.w2(32'hbcabb136),
	.w3(32'h3ae9d853),
	.w4(32'hbbb136fd),
	.w5(32'hbc442bc1),
	.w6(32'h3a553ca0),
	.w7(32'hbb9462fe),
	.w8(32'hbbba6649),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf946d),
	.w1(32'hb8bdd948),
	.w2(32'hbc825fa5),
	.w3(32'h3c4ef393),
	.w4(32'h3c2a2f83),
	.w5(32'hbbf0f650),
	.w6(32'h3a0a8166),
	.w7(32'h3b552ab1),
	.w8(32'h3aa040d7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb01bf4),
	.w1(32'hbbf148cf),
	.w2(32'h3c9788ac),
	.w3(32'hbb814820),
	.w4(32'hbca6027c),
	.w5(32'hbbbb3109),
	.w6(32'hbb0e8a69),
	.w7(32'hbc0347b7),
	.w8(32'h3aa7baba),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6fe6c),
	.w1(32'h39a0fc93),
	.w2(32'h3a6ac8bf),
	.w3(32'h3b83772e),
	.w4(32'h3943fd8c),
	.w5(32'h3c0590b0),
	.w6(32'h3b82bd7a),
	.w7(32'h3b8f06cf),
	.w8(32'h3bad2d10),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baba9fa),
	.w1(32'hbc8c837d),
	.w2(32'h3bc15f51),
	.w3(32'h3beb2543),
	.w4(32'hbc8004f0),
	.w5(32'hbcc8bc9d),
	.w6(32'hbcae3eea),
	.w7(32'hbc233cec),
	.w8(32'hbc96629e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7eb638),
	.w1(32'hbb185f93),
	.w2(32'h3c2b5b00),
	.w3(32'h3c262c3d),
	.w4(32'hbc0458f5),
	.w5(32'h3c74083c),
	.w6(32'h3befcaa3),
	.w7(32'hbc0f5a60),
	.w8(32'h3c518d4f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb013c41),
	.w1(32'hbbf3ce91),
	.w2(32'hbc48c986),
	.w3(32'h3be1f46c),
	.w4(32'hbc4b81b3),
	.w5(32'hbc4b88b1),
	.w6(32'h3c26d6f4),
	.w7(32'hbc0a7cc0),
	.w8(32'hbc826282),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeca969),
	.w1(32'h3b25f1b0),
	.w2(32'hbaa6db48),
	.w3(32'h3bb0c6c6),
	.w4(32'h3c3230a7),
	.w5(32'h3b570f8e),
	.w6(32'hbbf3a42e),
	.w7(32'hba7ed74a),
	.w8(32'hba5f60c1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc429977),
	.w1(32'hbb40f696),
	.w2(32'h3c01bc9e),
	.w3(32'hbbdd3126),
	.w4(32'hbba2bea9),
	.w5(32'h3c19a258),
	.w6(32'hbc17b7dd),
	.w7(32'hbbe406bb),
	.w8(32'hba8e33cd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f1b3c),
	.w1(32'h3b7cabf4),
	.w2(32'hba9f4c8f),
	.w3(32'hbadc78a6),
	.w4(32'h3b10704a),
	.w5(32'h3b6b9ce3),
	.w6(32'hbb914261),
	.w7(32'hbbe7b3ae),
	.w8(32'h3b05aaaf),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c31de),
	.w1(32'h3c205244),
	.w2(32'h3bd4ba21),
	.w3(32'h3b9c63a1),
	.w4(32'h3c6533cf),
	.w5(32'h3b1fd792),
	.w6(32'h3b302a73),
	.w7(32'h3c808555),
	.w8(32'hbb5fd1b1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b205d67),
	.w1(32'hbb0f73ba),
	.w2(32'hbb508f82),
	.w3(32'h3b83e590),
	.w4(32'hbb819aae),
	.w5(32'hba5694ff),
	.w6(32'h3bc211ad),
	.w7(32'hba9a76e2),
	.w8(32'h3c2a975f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27de65),
	.w1(32'hbc255d3f),
	.w2(32'hbc16b55a),
	.w3(32'h3af8364c),
	.w4(32'hbacd3004),
	.w5(32'hbbcda06d),
	.w6(32'hbc039d8c),
	.w7(32'hbbfcc7b5),
	.w8(32'hbc1e9156),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86c38d),
	.w1(32'h3be69b7e),
	.w2(32'h3c8f1e69),
	.w3(32'h3b17afc4),
	.w4(32'h3c75e925),
	.w5(32'hbbb58678),
	.w6(32'hbb88fe10),
	.w7(32'hbb4611b7),
	.w8(32'h3b72bb7c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ce69b8),
	.w1(32'hbbe1778e),
	.w2(32'hbbaa6ec8),
	.w3(32'hbc3a1c73),
	.w4(32'hbbe8b2e9),
	.w5(32'hbc17a59f),
	.w6(32'hbc22343b),
	.w7(32'hbc8484a6),
	.w8(32'hbc2d6008),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacf47f),
	.w1(32'h3a543e93),
	.w2(32'h3c13eb59),
	.w3(32'h3b438a80),
	.w4(32'h3ba8024b),
	.w5(32'h3c4f0f5b),
	.w6(32'hbbb9a9a8),
	.w7(32'h3b0307cf),
	.w8(32'h3b6e524c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5fc14),
	.w1(32'h3b44b5e3),
	.w2(32'hba01d605),
	.w3(32'h3c59b1de),
	.w4(32'h3b0e512a),
	.w5(32'h3893f98b),
	.w6(32'h3c52fa51),
	.w7(32'h391229d7),
	.w8(32'h3b942862),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a3ba9),
	.w1(32'h3a7cefc6),
	.w2(32'h3acb484f),
	.w3(32'h3b3395b6),
	.w4(32'h3b4cb783),
	.w5(32'hbafc68ef),
	.w6(32'h3b53dd9d),
	.w7(32'h3be867c7),
	.w8(32'hbad6a0e3),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af74a0b),
	.w1(32'hba996ff0),
	.w2(32'h3b9c57e9),
	.w3(32'h3b1c6f3d),
	.w4(32'h3a95b3ce),
	.w5(32'h3a7857d8),
	.w6(32'h3b2f3cb3),
	.w7(32'hbadac26e),
	.w8(32'h3b007b14),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2515b9),
	.w1(32'h3b9d2f4b),
	.w2(32'h39bfa8da),
	.w3(32'h3bf3d2f1),
	.w4(32'h3c1421d8),
	.w5(32'hbb80cc00),
	.w6(32'hbb9c8681),
	.w7(32'hbb820ce2),
	.w8(32'hba281f39),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c1af2),
	.w1(32'h3bb79d7b),
	.w2(32'hbadc472f),
	.w3(32'h3b323427),
	.w4(32'h3bdc4f9c),
	.w5(32'hb9a42538),
	.w6(32'hbb5f00ff),
	.w7(32'hb9fe33ac),
	.w8(32'hb9a8dd62),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf655dd),
	.w1(32'hbb9a8692),
	.w2(32'h3c0610b6),
	.w3(32'hbbde0cd3),
	.w4(32'hbc21e9cc),
	.w5(32'h3b97a3cf),
	.w6(32'hbb8a0ab4),
	.w7(32'hbb9ccf20),
	.w8(32'h3b7b8a28),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2e835),
	.w1(32'hbb5f31f3),
	.w2(32'hbbe870c2),
	.w3(32'h3c1e7ac0),
	.w4(32'h3b81abe4),
	.w5(32'h3c9f01ab),
	.w6(32'h3beded69),
	.w7(32'h3b64ed4a),
	.w8(32'h3cc008b6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c15b6d),
	.w1(32'hbb8e0508),
	.w2(32'h3bcfa780),
	.w3(32'h3ccc02e2),
	.w4(32'h3bfe559a),
	.w5(32'h3c219cec),
	.w6(32'h3cc12625),
	.w7(32'h3bc4b727),
	.w8(32'h3b90811f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6ea9e),
	.w1(32'hbbb80263),
	.w2(32'hba98d21d),
	.w3(32'h3ae0db06),
	.w4(32'hbc2face5),
	.w5(32'h3bdd41f6),
	.w6(32'hbb3c94bf),
	.w7(32'hbc366e4d),
	.w8(32'h3b5fc6eb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ef47),
	.w1(32'hbb7e7ec0),
	.w2(32'h3b0ca485),
	.w3(32'hbb6bf05a),
	.w4(32'hbb027de0),
	.w5(32'h3c2cd6d8),
	.w6(32'h3ae15f1a),
	.w7(32'hbc6d26bd),
	.w8(32'h3a52734f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b314fb3),
	.w1(32'h3b4696bd),
	.w2(32'h3b0e03e8),
	.w3(32'h3caf21a1),
	.w4(32'h3a2196aa),
	.w5(32'h3bcc6dac),
	.w6(32'h3c8b62a2),
	.w7(32'hbc59be75),
	.w8(32'h3930f99a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61b779),
	.w1(32'hbb59ecaf),
	.w2(32'h3c0c52b9),
	.w3(32'h3cca2ec7),
	.w4(32'h3c72806b),
	.w5(32'h3ca55e1b),
	.w6(32'hbaddc92a),
	.w7(32'h3bc8ea8d),
	.w8(32'h3aa53a15),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f378b),
	.w1(32'hbc5d9de9),
	.w2(32'h3c67bd4e),
	.w3(32'h3a4ffca2),
	.w4(32'hbc0f9f58),
	.w5(32'h3bdfa976),
	.w6(32'hb91fdbba),
	.w7(32'hbc01b049),
	.w8(32'hbc0aff03),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a590ed8),
	.w1(32'h3bdf4f9c),
	.w2(32'h3c17a23b),
	.w3(32'hbb59a39d),
	.w4(32'h3b088589),
	.w5(32'h3b5221a7),
	.w6(32'hbb1b52cd),
	.w7(32'hbc029868),
	.w8(32'h3c215b68),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19b1bb),
	.w1(32'hbc128d9c),
	.w2(32'h3af893c0),
	.w3(32'hbbd4ab39),
	.w4(32'h3998aaa4),
	.w5(32'h3b5b0108),
	.w6(32'hbbce62ae),
	.w7(32'h3c5b1913),
	.w8(32'hb982c4b6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b540f83),
	.w1(32'h3a5fd431),
	.w2(32'hbc17b484),
	.w3(32'h3bda6351),
	.w4(32'h3b6b6b6a),
	.w5(32'hbc0ac861),
	.w6(32'hba941b4a),
	.w7(32'hbb83cb7a),
	.w8(32'h3b17bb59),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b1e2c),
	.w1(32'hbba7dfcf),
	.w2(32'hbb1535ec),
	.w3(32'hbaaf7a39),
	.w4(32'hbbd2ea8c),
	.w5(32'h3beef5d5),
	.w6(32'h3af258cc),
	.w7(32'h3c1c6d4e),
	.w8(32'h3a5b26a0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d4760),
	.w1(32'h3bfacc24),
	.w2(32'h3a569e76),
	.w3(32'h3c93713e),
	.w4(32'h3c288363),
	.w5(32'hbb70f9e6),
	.w6(32'h3c441e52),
	.w7(32'h3bab81e8),
	.w8(32'h3a072003),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1270a8),
	.w1(32'h3c7ed2a9),
	.w2(32'h3d0f0330),
	.w3(32'hbc8ca8e3),
	.w4(32'hbb368554),
	.w5(32'h3c9f5790),
	.w6(32'hbc0b419b),
	.w7(32'h3acafaa1),
	.w8(32'h3c2421ee),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5aff76),
	.w1(32'hba8ed08e),
	.w2(32'hbc8869f0),
	.w3(32'h3c3ad99d),
	.w4(32'h3b1ed78d),
	.w5(32'hbafdaf4d),
	.w6(32'hbb801136),
	.w7(32'hbae1bd43),
	.w8(32'h3baa0a48),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc088ced),
	.w1(32'hbb9c198d),
	.w2(32'h3c94ef9f),
	.w3(32'hbbc947d2),
	.w4(32'hbc7059af),
	.w5(32'hbae605a6),
	.w6(32'hbc0c8e4c),
	.w7(32'hbc3f3ed4),
	.w8(32'hba924fe9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb30b14),
	.w1(32'h3be682ec),
	.w2(32'h3c887f19),
	.w3(32'hbcaa1e4d),
	.w4(32'hbc383f37),
	.w5(32'h3c1b4b6f),
	.w6(32'hbce3c86f),
	.w7(32'hbc2bbabf),
	.w8(32'h3afba407),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b1f8b),
	.w1(32'hbbcc2e22),
	.w2(32'hbaea0b25),
	.w3(32'h3a35f9a0),
	.w4(32'hbb7d0a9f),
	.w5(32'hbbd77f7a),
	.w6(32'hbb8b3acd),
	.w7(32'hbb968952),
	.w8(32'hbc128c62),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb402c14),
	.w1(32'h3a6a3cbc),
	.w2(32'h3c5d6d13),
	.w3(32'h3b514815),
	.w4(32'h3b2a3b0c),
	.w5(32'h3bf4b38d),
	.w6(32'h3b8e631a),
	.w7(32'h3bd94351),
	.w8(32'h3bc54bd5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc47d2),
	.w1(32'h3b869995),
	.w2(32'h3b998d5f),
	.w3(32'h3ba7ec6e),
	.w4(32'h3b9c240c),
	.w5(32'h3ba703a2),
	.w6(32'h3b798172),
	.w7(32'h3b906940),
	.w8(32'h3b8cad68),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9852f3),
	.w1(32'h3b8eedcb),
	.w2(32'hbc6f06ff),
	.w3(32'h3b784c4e),
	.w4(32'h3bf3e4ea),
	.w5(32'hbbbbc4ca),
	.w6(32'hbbaa6211),
	.w7(32'h3b511442),
	.w8(32'hb90c1354),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ce94f),
	.w1(32'h3a0d0cbb),
	.w2(32'hbbbd4c1d),
	.w3(32'hbc329e96),
	.w4(32'hbc0258bf),
	.w5(32'hbc7c9ed0),
	.w6(32'hbb95ef9d),
	.w7(32'hbc5a73ce),
	.w8(32'hbc1d5a2a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce3efa),
	.w1(32'h3aee4bbd),
	.w2(32'h3b31b338),
	.w3(32'hbc1258bf),
	.w4(32'h3b57ec9d),
	.w5(32'h3b0e5566),
	.w6(32'hbbdca88d),
	.w7(32'h3c16ec44),
	.w8(32'h3b2bb8b1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c7f45),
	.w1(32'hbae8d028),
	.w2(32'hbbaf76c9),
	.w3(32'h3b4a5c6e),
	.w4(32'hbb251585),
	.w5(32'hbc48b586),
	.w6(32'h3b5b0cf8),
	.w7(32'hbb168f22),
	.w8(32'hbc8cdbe1),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37461c),
	.w1(32'h3accc001),
	.w2(32'h3b07ba83),
	.w3(32'hbc873f73),
	.w4(32'hbbb07e79),
	.w5(32'hbb2ed3a9),
	.w6(32'hbca4b10f),
	.w7(32'hbc422673),
	.w8(32'hba46654b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe510c),
	.w1(32'hb95cec9d),
	.w2(32'hbc8bf20f),
	.w3(32'hbac6b13d),
	.w4(32'hbbe039c7),
	.w5(32'hbb90aabb),
	.w6(32'hb6d7234c),
	.w7(32'hbae78878),
	.w8(32'hbc3738ec),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccd1c4f),
	.w1(32'hbc86f9f2),
	.w2(32'h3c1b0345),
	.w3(32'hbb9fc928),
	.w4(32'hbc9a28ec),
	.w5(32'h3bcc3f25),
	.w6(32'hbc39b747),
	.w7(32'hbbcc8212),
	.w8(32'hbb5d364f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b800d7a),
	.w1(32'h3bd4fe86),
	.w2(32'h3ba12549),
	.w3(32'h3b6887e0),
	.w4(32'h3bc906fe),
	.w5(32'hba360907),
	.w6(32'hba3f89a4),
	.w7(32'h3afae356),
	.w8(32'h3aaec24d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8546de),
	.w1(32'h3aafd55e),
	.w2(32'h3b9effe7),
	.w3(32'hbb53388e),
	.w4(32'hb9fcb3bf),
	.w5(32'h3bed2475),
	.w6(32'hbb7830b7),
	.w7(32'h3ae8e0a7),
	.w8(32'h3b06fda5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb785a832),
	.w1(32'hbbacb597),
	.w2(32'h3afecd7f),
	.w3(32'h3c749bf1),
	.w4(32'h3bc9cbf3),
	.w5(32'h3b7fe1ef),
	.w6(32'h3b916e67),
	.w7(32'hbb0b7cec),
	.w8(32'h3b5f194d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe24615),
	.w1(32'h3b1c9439),
	.w2(32'h3c98175c),
	.w3(32'hbc81971a),
	.w4(32'hbc73cc3e),
	.w5(32'h3b09b950),
	.w6(32'hbb455022),
	.w7(32'hbbaed351),
	.w8(32'h3b9968ea),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becc715),
	.w1(32'h3cb6979d),
	.w2(32'h3bd9b975),
	.w3(32'hbb758915),
	.w4(32'h3bb073ef),
	.w5(32'h3c2ff709),
	.w6(32'h3c833bee),
	.w7(32'h3bebe4f7),
	.w8(32'h3c1c4797),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafc5a9),
	.w1(32'h3be1a6c8),
	.w2(32'hbc264f05),
	.w3(32'h3a9b5dde),
	.w4(32'h3c16a394),
	.w5(32'h3c18334c),
	.w6(32'hbbc5ac19),
	.w7(32'hbc1984e2),
	.w8(32'h3c0f026b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dfcf5),
	.w1(32'hbbae1a7d),
	.w2(32'hba6707ea),
	.w3(32'h3c1665e8),
	.w4(32'h3c341579),
	.w5(32'hbac78fad),
	.w6(32'h3bb3fa06),
	.w7(32'h3afb63c2),
	.w8(32'h395a512e),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0d974),
	.w1(32'hbb1d75f7),
	.w2(32'hbbbc18c3),
	.w3(32'h3a9c5d07),
	.w4(32'hbb3818e3),
	.w5(32'hbb4b5dcd),
	.w6(32'hbb0f17df),
	.w7(32'hbb1d3b06),
	.w8(32'hbc140ac0),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd01b75),
	.w1(32'h3a82dcac),
	.w2(32'h3c6a3c08),
	.w3(32'hbac03560),
	.w4(32'h3bdb0b80),
	.w5(32'hba8a86a1),
	.w6(32'hbc1974e9),
	.w7(32'hbc514970),
	.w8(32'hbcdf27d1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c823c68),
	.w1(32'h39f370ab),
	.w2(32'hbbe28147),
	.w3(32'h3c942b8e),
	.w4(32'h3b9b89ae),
	.w5(32'hbc0740ca),
	.w6(32'hbc7246ef),
	.w7(32'hbc1ecf09),
	.w8(32'hbbf091a9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9003bc),
	.w1(32'h3c153814),
	.w2(32'hbc16943a),
	.w3(32'hbb9005f2),
	.w4(32'h3a84455f),
	.w5(32'hbb55cfb8),
	.w6(32'hbb811738),
	.w7(32'h3ab5bc21),
	.w8(32'h3b25a0a6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81f56d),
	.w1(32'hbc15802c),
	.w2(32'hbbc03365),
	.w3(32'h3c9ac127),
	.w4(32'h3c43bd9b),
	.w5(32'hbbcc45e6),
	.w6(32'h3ce49219),
	.w7(32'h3c790925),
	.w8(32'h3b3149c4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc890048),
	.w1(32'hba0add2c),
	.w2(32'h3b96baca),
	.w3(32'hb8bfca26),
	.w4(32'h397f1ba7),
	.w5(32'h3b7cc903),
	.w6(32'h3c1f6bcf),
	.w7(32'h3c3167ac),
	.w8(32'h3bbda227),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17b4fd),
	.w1(32'hbb4f27b6),
	.w2(32'h3c04e40c),
	.w3(32'h3ac40348),
	.w4(32'h3b8095de),
	.w5(32'h3c5c3648),
	.w6(32'h3b757d39),
	.w7(32'h3b662c59),
	.w8(32'h3b378e99),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a824b),
	.w1(32'hbbb6f13d),
	.w2(32'hbc0ca4fb),
	.w3(32'h3c94d20b),
	.w4(32'hb93dccb4),
	.w5(32'hb996cee0),
	.w6(32'h3bedfb7f),
	.w7(32'h3ab9e64d),
	.w8(32'hbb1be0b2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3e019),
	.w1(32'hbbfbe16a),
	.w2(32'h3c6fc766),
	.w3(32'h3ba0e5d7),
	.w4(32'h3b85007f),
	.w5(32'h3bcf9ef9),
	.w6(32'h3b39489e),
	.w7(32'hba6c0039),
	.w8(32'hbbb4f00e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e7ba6),
	.w1(32'h3b0c56c6),
	.w2(32'hbbbc215f),
	.w3(32'hbc5474df),
	.w4(32'hbc013f46),
	.w5(32'h3b0e0906),
	.w6(32'hbce0f576),
	.w7(32'hbc435bf3),
	.w8(32'h3bae4020),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37600b),
	.w1(32'hbc13fda0),
	.w2(32'hbc1f3a7d),
	.w3(32'h3c24ed75),
	.w4(32'h3b890852),
	.w5(32'h3bc19d16),
	.w6(32'h39011c1b),
	.w7(32'hbbb2e059),
	.w8(32'h3c99aa59),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba465a66),
	.w1(32'hbb335864),
	.w2(32'h3c042f83),
	.w3(32'h3d0d0141),
	.w4(32'h3d04dbb1),
	.w5(32'hbbc9df0c),
	.w6(32'h3d0d62d5),
	.w7(32'h3d0a68cf),
	.w8(32'h3c30f4cf),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ca6d7),
	.w1(32'h3b981170),
	.w2(32'hb9eebede),
	.w3(32'hbc7122d0),
	.w4(32'hbc005542),
	.w5(32'h3bc77a83),
	.w6(32'h3ad88d28),
	.w7(32'hbbb434f5),
	.w8(32'h3c2e4021),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e27ae),
	.w1(32'hbbad2763),
	.w2(32'hb88fbd09),
	.w3(32'h3b1929ec),
	.w4(32'hb9cc4e4d),
	.w5(32'hbc467bf6),
	.w6(32'h3ba3d0cb),
	.w7(32'h3c025a1a),
	.w8(32'hb9aad3d0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47f66d),
	.w1(32'hbc165146),
	.w2(32'hbbd9cac6),
	.w3(32'hbc4e6b63),
	.w4(32'hbba94e2c),
	.w5(32'h3a56d8c6),
	.w6(32'h3ce9111d),
	.w7(32'h3ce99cd8),
	.w8(32'hbbae78f6),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb855bb7),
	.w1(32'hbc89d9a7),
	.w2(32'hbc70dbfc),
	.w3(32'h3c8922b5),
	.w4(32'h3c168016),
	.w5(32'hbb461439),
	.w6(32'h3b720f5a),
	.w7(32'h3a8a1eb2),
	.w8(32'hba37e3a4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc720e14),
	.w1(32'hbbcae719),
	.w2(32'h3c5ecb59),
	.w3(32'h3bbe6672),
	.w4(32'h3bd4e17e),
	.w5(32'hbb2ac5cb),
	.w6(32'h3c25904d),
	.w7(32'h3bdc9a55),
	.w8(32'hbc413bc9),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8bd2d6),
	.w1(32'h3c843809),
	.w2(32'h3c299158),
	.w3(32'hbc09e0df),
	.w4(32'h3c1ca407),
	.w5(32'h3b734402),
	.w6(32'h3b29402b),
	.w7(32'hba59cb6a),
	.w8(32'hbb83c326),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6870c8),
	.w1(32'h3ad8ad55),
	.w2(32'h3c2fb222),
	.w3(32'hbc433464),
	.w4(32'hbbb7bbb3),
	.w5(32'hbc0b0f35),
	.w6(32'hbb8291b0),
	.w7(32'hbbb2d43a),
	.w8(32'hbc430899),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd859c8),
	.w1(32'h3ba44efb),
	.w2(32'h3c7985e1),
	.w3(32'hbc6f4492),
	.w4(32'h3bf24205),
	.w5(32'h3c2c19dc),
	.w6(32'hbba76062),
	.w7(32'hbc1141bd),
	.w8(32'hbb46e51e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19ba6a),
	.w1(32'hb9e0c861),
	.w2(32'hbb46c3bf),
	.w3(32'hbbe2c359),
	.w4(32'hbc5bd0cf),
	.w5(32'h3b1da10a),
	.w6(32'hbbf24279),
	.w7(32'hbc1c55d6),
	.w8(32'hbb58ab3f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9ea53),
	.w1(32'hbb367f08),
	.w2(32'hba86bcc7),
	.w3(32'hb8c156ea),
	.w4(32'h3b9858ea),
	.w5(32'h3b2d9d09),
	.w6(32'hbae64cc6),
	.w7(32'hbaca5ff0),
	.w8(32'h3c6aca7e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fb732),
	.w1(32'hbc0e9608),
	.w2(32'h3b34f1c9),
	.w3(32'hbad89ac7),
	.w4(32'h3ba8a399),
	.w5(32'h3aa49847),
	.w6(32'h3ce97a31),
	.w7(32'h3c9cf9e9),
	.w8(32'hbbdda665),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba580e05),
	.w1(32'hbb89b15d),
	.w2(32'h39de09c4),
	.w3(32'h3c16fe54),
	.w4(32'h3b914f64),
	.w5(32'hbb9fdb99),
	.w6(32'h39e34438),
	.w7(32'h3c0eade6),
	.w8(32'hbc965ebf),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae008c4),
	.w1(32'hba8c51b2),
	.w2(32'hbb18b6e0),
	.w3(32'h3bb8b42d),
	.w4(32'hbbcb0c23),
	.w5(32'h3bc1ffdf),
	.w6(32'hbc59bfb2),
	.w7(32'h3a30f4f9),
	.w8(32'hbae910ef),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab431ee),
	.w1(32'h3a9e397e),
	.w2(32'h3bed7fd3),
	.w3(32'h3ba82b62),
	.w4(32'h3b17a04b),
	.w5(32'hbb30f3e9),
	.w6(32'h3bbddc56),
	.w7(32'hb9c4842a),
	.w8(32'hbb2cab78),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9d1f8),
	.w1(32'h3bd2ab65),
	.w2(32'hbbc4e671),
	.w3(32'h3be406a4),
	.w4(32'hbb29fb98),
	.w5(32'h3b7b6e2a),
	.w6(32'hbb33c764),
	.w7(32'hbc41fb84),
	.w8(32'hbc25f87d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1408a9),
	.w1(32'hbb9649c9),
	.w2(32'h39a4d608),
	.w3(32'h3c7c78c1),
	.w4(32'h3c75dfc3),
	.w5(32'hbbdfe73c),
	.w6(32'hb97b1376),
	.w7(32'hbb160853),
	.w8(32'h39e20a24),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c241ce6),
	.w1(32'h3bc4f281),
	.w2(32'hbc5af980),
	.w3(32'h3ba8f634),
	.w4(32'h3c0d5c55),
	.w5(32'hbbc50478),
	.w6(32'h3c76bdf3),
	.w7(32'h3c57d420),
	.w8(32'hbb06f791),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e9c9f),
	.w1(32'hbb93ba66),
	.w2(32'h3c550b2e),
	.w3(32'hbbd76c55),
	.w4(32'h39afcca3),
	.w5(32'hbc722503),
	.w6(32'h3b3b0991),
	.w7(32'hbb9e2138),
	.w8(32'hbc0eee1b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdd96c),
	.w1(32'hbc5152e6),
	.w2(32'hbc138665),
	.w3(32'hbc93b747),
	.w4(32'hbb8a1707),
	.w5(32'hbc5aa935),
	.w6(32'h39167380),
	.w7(32'h3ca40e6c),
	.w8(32'hbc9c8fc8),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb740c),
	.w1(32'hbb471434),
	.w2(32'hbc5b831f),
	.w3(32'hb9df62ac),
	.w4(32'hb9b4d545),
	.w5(32'hbc847553),
	.w6(32'hbc171909),
	.w7(32'hbb5bf0fe),
	.w8(32'h3b2649e7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcefdc49),
	.w1(32'hbbdb51df),
	.w2(32'h3d3450fc),
	.w3(32'hbcf68bca),
	.w4(32'hbc13634c),
	.w5(32'h3ca17f88),
	.w6(32'h3cb8dcad),
	.w7(32'h3cf08154),
	.w8(32'h3a22fd88),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c961a2b),
	.w1(32'h3cfbf1f8),
	.w2(32'hbab50ce6),
	.w3(32'hbd2eef74),
	.w4(32'hbcae39fc),
	.w5(32'h3a16e5b9),
	.w6(32'hba43dd38),
	.w7(32'hbc179a6d),
	.w8(32'h3b8b8397),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91d45b),
	.w1(32'hbb197a59),
	.w2(32'h3c1b71bf),
	.w3(32'h3b350f34),
	.w4(32'h3c52493e),
	.w5(32'h3bfca579),
	.w6(32'h3a76c273),
	.w7(32'h3c086d4b),
	.w8(32'h3b4aacdd),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4639bc),
	.w1(32'h3c088ae6),
	.w2(32'hbb982c5c),
	.w3(32'hbafd1e37),
	.w4(32'hba9f977d),
	.w5(32'hbc799420),
	.w6(32'hbb412720),
	.w7(32'hbc1a7247),
	.w8(32'h3b488758),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46502a),
	.w1(32'hbbc2f065),
	.w2(32'hb9fa6fe7),
	.w3(32'hbc79d4f4),
	.w4(32'hbc16e421),
	.w5(32'hbc24db18),
	.w6(32'h3c8498a0),
	.w7(32'h3cb88860),
	.w8(32'hb93314de),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba544319),
	.w1(32'h3b227a66),
	.w2(32'h3bbbd7af),
	.w3(32'hbc36708a),
	.w4(32'hbc3d1593),
	.w5(32'h3bd9c4d9),
	.w6(32'hbacee99a),
	.w7(32'h3bcfd28e),
	.w8(32'hbb424a4f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb490b9),
	.w1(32'h3b918dd6),
	.w2(32'h3b7dc77e),
	.w3(32'h3bea8e1d),
	.w4(32'h3b20db4a),
	.w5(32'h3ba17ff1),
	.w6(32'hbc03029c),
	.w7(32'hbb33cbbb),
	.w8(32'h3c0cfe88),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ef0c4),
	.w1(32'hbb9b6f7b),
	.w2(32'hbacac074),
	.w3(32'h3b2b96a0),
	.w4(32'h3b407926),
	.w5(32'h3b1e111b),
	.w6(32'hbb20a62f),
	.w7(32'h3b0dd932),
	.w8(32'hbb101f72),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfeb63b),
	.w1(32'hbba453ab),
	.w2(32'hbc0dd427),
	.w3(32'h3c4255ee),
	.w4(32'h3b0a144a),
	.w5(32'hbafbbb97),
	.w6(32'h3b736760),
	.w7(32'h3c0e9fe6),
	.w8(32'hbbcccac0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c027aac),
	.w1(32'hbbaa513a),
	.w2(32'hbb63bd7f),
	.w3(32'h3b9bbbf4),
	.w4(32'h3ae89d05),
	.w5(32'hbb8afae9),
	.w6(32'h390efb6c),
	.w7(32'h3b68c145),
	.w8(32'hbbc1ed9c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cd05d),
	.w1(32'hbb841184),
	.w2(32'hbaf03757),
	.w3(32'hbc1ee7e1),
	.w4(32'hbba88d72),
	.w5(32'h3c1895c6),
	.w6(32'hbc5dda7f),
	.w7(32'hbc1ba1b7),
	.w8(32'h3c1c8be3),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ffe02),
	.w1(32'hbbe48e1c),
	.w2(32'h3baa4d92),
	.w3(32'h3afedf59),
	.w4(32'hbc98dbfd),
	.w5(32'hba27b611),
	.w6(32'h3c41c24f),
	.w7(32'hbc0a0a11),
	.w8(32'hbb24b1de),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c139da7),
	.w1(32'h3bd39562),
	.w2(32'h3ade117a),
	.w3(32'h3b002f67),
	.w4(32'h3ba7ba1e),
	.w5(32'h3b5bd36c),
	.w6(32'hbc101860),
	.w7(32'hbb0a5071),
	.w8(32'hbb8543cc),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d1320),
	.w1(32'h3b9f25ac),
	.w2(32'hbbdd3438),
	.w3(32'h3c2dfb94),
	.w4(32'h3ad753e7),
	.w5(32'hbc68a99d),
	.w6(32'h3aa8824c),
	.w7(32'hbc142579),
	.w8(32'hbc8543d0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaebbbd),
	.w1(32'h3b9a4e40),
	.w2(32'h3ac7eede),
	.w3(32'h3abf955f),
	.w4(32'h3c0970e7),
	.w5(32'h3bd8dd1d),
	.w6(32'h3c2a3c88),
	.w7(32'h3c537285),
	.w8(32'h3a684507),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c9f95),
	.w1(32'h3b6a47b7),
	.w2(32'hbad69a64),
	.w3(32'h3be185c2),
	.w4(32'h3c4ccc3a),
	.w5(32'h3b76e812),
	.w6(32'hba959b82),
	.w7(32'h3b331269),
	.w8(32'h3b613c9c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb892829),
	.w1(32'hbbea467b),
	.w2(32'hbc29c782),
	.w3(32'h3c4f4caf),
	.w4(32'h3b4ad263),
	.w5(32'hbcae4c1f),
	.w6(32'h3ca218ce),
	.w7(32'h3c9a31c5),
	.w8(32'hbc70a6b0),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb855442),
	.w1(32'hbc114a48),
	.w2(32'hbb4dc3f9),
	.w3(32'hbc2802cd),
	.w4(32'hbb935ed3),
	.w5(32'hbc2019d3),
	.w6(32'hbbe25ed1),
	.w7(32'hbba03573),
	.w8(32'hbc8dcd98),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7a34e),
	.w1(32'hbc172ef0),
	.w2(32'h3a5dd929),
	.w3(32'hbb67ef38),
	.w4(32'hbb2cb313),
	.w5(32'hbb1e024c),
	.w6(32'hba8fb97b),
	.w7(32'h3c2721aa),
	.w8(32'h3b38e112),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cb97e),
	.w1(32'hbc87c750),
	.w2(32'hbc3cf8b5),
	.w3(32'hbb72b6ff),
	.w4(32'hbbd13b0f),
	.w5(32'hbb1a939a),
	.w6(32'hba8f7149),
	.w7(32'hbb840448),
	.w8(32'hbb9d81ee),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a42b6),
	.w1(32'h3b92a7a3),
	.w2(32'hbaf80171),
	.w3(32'h3c03a2be),
	.w4(32'h3becd690),
	.w5(32'h3ac51cc0),
	.w6(32'h3790e418),
	.w7(32'h3ac61fb1),
	.w8(32'hbba3975e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17b455),
	.w1(32'hbb9776dc),
	.w2(32'h3b89773f),
	.w3(32'hb9dcefc0),
	.w4(32'hbb6ab725),
	.w5(32'hba6c9094),
	.w6(32'hbbc47cbe),
	.w7(32'h39b07130),
	.w8(32'h3ac0ec24),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb895fe),
	.w1(32'hba432d69),
	.w2(32'hba3457b8),
	.w3(32'hbb60eb2d),
	.w4(32'hbae2b24a),
	.w5(32'h3c867dc5),
	.w6(32'hbb01714e),
	.w7(32'h3b28c2a9),
	.w8(32'h3c36fe17),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1517f1),
	.w1(32'h3bac4d13),
	.w2(32'hbbeff335),
	.w3(32'h3b903acb),
	.w4(32'hba8625db),
	.w5(32'h3b3d1e2a),
	.w6(32'h3be61afe),
	.w7(32'hb9a4e921),
	.w8(32'hbc07e5db),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51d74d),
	.w1(32'h3c2f1a32),
	.w2(32'h3c6a407d),
	.w3(32'h3c2f0b6b),
	.w4(32'h3c3c735a),
	.w5(32'h3c4806fc),
	.w6(32'hbcc0fb8c),
	.w7(32'hbac96bf2),
	.w8(32'hbb98bf29),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7f100),
	.w1(32'hba8ca72e),
	.w2(32'h3b886c28),
	.w3(32'h3bf7c5d2),
	.w4(32'h3c4664f4),
	.w5(32'h3b729ffb),
	.w6(32'hbbc7b8e7),
	.w7(32'h3adb51a4),
	.w8(32'h3c0356e1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe78558),
	.w1(32'hbbabab82),
	.w2(32'hbbbd694e),
	.w3(32'hbbc80e08),
	.w4(32'hbbce4854),
	.w5(32'hbbc6d592),
	.w6(32'h3ac2dc6e),
	.w7(32'hbbac233d),
	.w8(32'hbc4cc1c5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62ac09),
	.w1(32'hbb8068a9),
	.w2(32'h3ca1404a),
	.w3(32'hbcb08168),
	.w4(32'hbc9ae21c),
	.w5(32'hbba287c0),
	.w6(32'h3ba9d770),
	.w7(32'hbb35eea1),
	.w8(32'h3c203fb6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984afdd),
	.w1(32'h3ac917a2),
	.w2(32'h3aaea49d),
	.w3(32'h3b32541f),
	.w4(32'h3b8eb74e),
	.w5(32'hbb68b30b),
	.w6(32'h3bbf190a),
	.w7(32'h3c09725b),
	.w8(32'hbbf1223c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb975194),
	.w1(32'hbbbaf2eb),
	.w2(32'h3c99a77d),
	.w3(32'hbb39e1ce),
	.w4(32'hb96ce4c6),
	.w5(32'h3ca09d08),
	.w6(32'hb95a0fd3),
	.w7(32'hba58ee1e),
	.w8(32'hbc4c759f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d4c8f),
	.w1(32'h3b961b08),
	.w2(32'h3cbca509),
	.w3(32'h3d58ab01),
	.w4(32'h3cacae66),
	.w5(32'h3c0fcd27),
	.w6(32'hbb9b1848),
	.w7(32'hbc29316a),
	.w8(32'hbb467174),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82a828),
	.w1(32'h3c735d7b),
	.w2(32'h3d31e599),
	.w3(32'hba87ae38),
	.w4(32'hba69907e),
	.w5(32'h3ccd98ce),
	.w6(32'hbcb367b4),
	.w7(32'hbcb0779b),
	.w8(32'h3c2c2e3d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08cc55),
	.w1(32'h3aaa929a),
	.w2(32'h3c01f804),
	.w3(32'hbcbcf0eb),
	.w4(32'hbcce3d4a),
	.w5(32'h3b64e132),
	.w6(32'hbcefc892),
	.w7(32'hbca95da9),
	.w8(32'h3ac63cca),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c074a9f),
	.w1(32'h3b53a8ca),
	.w2(32'hbbbdfebc),
	.w3(32'h3c31bff0),
	.w4(32'h3c302400),
	.w5(32'hbbbe634e),
	.w6(32'h3c4e19a0),
	.w7(32'h3c472d3d),
	.w8(32'h39bd87b4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e9646),
	.w1(32'h3bdde14a),
	.w2(32'hbbdfc1ef),
	.w3(32'hbbb2d74d),
	.w4(32'h3a52800b),
	.w5(32'hbb8ab2f2),
	.w6(32'h3a8b75d2),
	.w7(32'h3bc27a34),
	.w8(32'hbb32d422),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a229652),
	.w1(32'hbbc16c6a),
	.w2(32'h3b28f463),
	.w3(32'h3bdbadf9),
	.w4(32'hbb02de0c),
	.w5(32'h3c73ed0c),
	.w6(32'h3b35b2e6),
	.w7(32'h3b6c21fc),
	.w8(32'h3c778301),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c1722),
	.w1(32'hbbd41e5c),
	.w2(32'hbc6f27ef),
	.w3(32'h3c4d31f8),
	.w4(32'h3bbe047a),
	.w5(32'h3bfe57bb),
	.w6(32'h3c10838f),
	.w7(32'h3b280ef6),
	.w8(32'h3c817532),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94cdcf),
	.w1(32'hbc24d7d8),
	.w2(32'hbb99f238),
	.w3(32'h3ca650c2),
	.w4(32'h3ca5f65c),
	.w5(32'h3b86ed49),
	.w6(32'h3c3a3ff6),
	.w7(32'h3c3989a4),
	.w8(32'h3bc92599),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f631f),
	.w1(32'h3b6f74e2),
	.w2(32'hbc7752f0),
	.w3(32'h3bab6da9),
	.w4(32'h3b5def09),
	.w5(32'hbc167ca5),
	.w6(32'h3b007623),
	.w7(32'hbb8bbdd5),
	.w8(32'hbc365676),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6dbb1e),
	.w1(32'hbc46c7d2),
	.w2(32'h3bc13d90),
	.w3(32'h3c706c2c),
	.w4(32'h3c54d039),
	.w5(32'h3cb56617),
	.w6(32'h3b2d3f10),
	.w7(32'h3cae22a9),
	.w8(32'h3c220ab9),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ef7e4),
	.w1(32'hbc67c73f),
	.w2(32'hbc60e2f7),
	.w3(32'h3b2444dc),
	.w4(32'hbb685e56),
	.w5(32'h3b500791),
	.w6(32'hbc3321f8),
	.w7(32'hbbfb9569),
	.w8(32'h3adea84d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8715a6),
	.w1(32'hbc483711),
	.w2(32'hbc1d2f71),
	.w3(32'h3baaef0d),
	.w4(32'hbad09b14),
	.w5(32'hbb8e3326),
	.w6(32'h3c368c16),
	.w7(32'h3bce156f),
	.w8(32'hbab33e5c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0bef5),
	.w1(32'hbbc099b4),
	.w2(32'hbc3dad9c),
	.w3(32'h3c11b90e),
	.w4(32'hba420403),
	.w5(32'hbc129474),
	.w6(32'h3c431b91),
	.w7(32'h3b2d738d),
	.w8(32'hbb94a8e7),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd026b9b),
	.w1(32'hbc072f9b),
	.w2(32'h3c855e5b),
	.w3(32'hbc52a973),
	.w4(32'hbbe4db49),
	.w5(32'h39433414),
	.w6(32'hbc7826af),
	.w7(32'h3b94c87e),
	.w8(32'hbc833edb),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af80e95),
	.w1(32'h3a20e729),
	.w2(32'h3c212fc3),
	.w3(32'h3bc31333),
	.w4(32'h37c35c07),
	.w5(32'h3c53b1b5),
	.w6(32'hbc176b32),
	.w7(32'hbc8066de),
	.w8(32'h3b6a27a8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68c827),
	.w1(32'hbc3362df),
	.w2(32'hbc01590a),
	.w3(32'hbb0df16d),
	.w4(32'hbb57d8c8),
	.w5(32'hbba3296e),
	.w6(32'hbc42e554),
	.w7(32'hbc60f58e),
	.w8(32'h3b658a92),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6bf4c3),
	.w1(32'hbc0390d9),
	.w2(32'h3c18d561),
	.w3(32'hbc39e42f),
	.w4(32'hbbe4bc84),
	.w5(32'h3c2c09b1),
	.w6(32'hba6e1744),
	.w7(32'hbb262135),
	.w8(32'h3c02f395),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a6244),
	.w1(32'hbbbd6fdb),
	.w2(32'hbc04e959),
	.w3(32'h3b2468af),
	.w4(32'hb8e998fd),
	.w5(32'hbb479304),
	.w6(32'h3c0330c3),
	.w7(32'hbacd8aa9),
	.w8(32'hbc05b853),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8218dc),
	.w1(32'hbc2b9287),
	.w2(32'hbc2ebc6f),
	.w3(32'hbb78d5b8),
	.w4(32'hbbc54dcb),
	.w5(32'h3b5db7df),
	.w6(32'h3b950db7),
	.w7(32'h3b305cec),
	.w8(32'hbbfb1144),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27d6e3),
	.w1(32'hbb71f667),
	.w2(32'hbc1f6529),
	.w3(32'h3b004161),
	.w4(32'hbab737a2),
	.w5(32'hbb5fd3f9),
	.w6(32'h3b56232a),
	.w7(32'hbaa43302),
	.w8(32'hbbb2da18),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29e390),
	.w1(32'hbbf39cd0),
	.w2(32'h3b69b514),
	.w3(32'h3c8c2ec8),
	.w4(32'h3cbb1006),
	.w5(32'h3bb3dc6f),
	.w6(32'h3c57f849),
	.w7(32'h3c4f5761),
	.w8(32'h397ff371),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bfd01),
	.w1(32'h3ba5ff59),
	.w2(32'hbc3fb0fc),
	.w3(32'h3c369c9e),
	.w4(32'h3c199531),
	.w5(32'h3b29ea78),
	.w6(32'hbb1045ff),
	.w7(32'hba0f6154),
	.w8(32'h3af745e0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf772b2),
	.w1(32'h3c90865d),
	.w2(32'h3c5c019c),
	.w3(32'hbc6a855b),
	.w4(32'hb9ed6d27),
	.w5(32'h3c18dd65),
	.w6(32'h3bb8f990),
	.w7(32'hba84bf59),
	.w8(32'h3c55be4a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6195cc),
	.w1(32'h391bafa4),
	.w2(32'h3b23600c),
	.w3(32'hbc7e64dc),
	.w4(32'hbb8d4fd4),
	.w5(32'h3b370076),
	.w6(32'hbae9ac8e),
	.w7(32'h3bb56654),
	.w8(32'hbc4d4d19),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39e0f3),
	.w1(32'hbafa8a9d),
	.w2(32'h3c54f9a1),
	.w3(32'h3c2d24f3),
	.w4(32'h3c56db1d),
	.w5(32'hbbca82f3),
	.w6(32'h3c9f9ad7),
	.w7(32'h3c1c757f),
	.w8(32'hbbdfec64),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1139a1),
	.w1(32'hbc12a83a),
	.w2(32'h39ce729b),
	.w3(32'hbd153781),
	.w4(32'hbd0c633b),
	.w5(32'h3b185a30),
	.w6(32'hbc24b931),
	.w7(32'hba5c022f),
	.w8(32'hb96d058d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c308d),
	.w1(32'hbb892e56),
	.w2(32'h3c647f86),
	.w3(32'hb99e7eb5),
	.w4(32'h3aa09e60),
	.w5(32'h3c42e7cd),
	.w6(32'hba103a9e),
	.w7(32'h3b971174),
	.w8(32'hba8eb0a4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf09d2b),
	.w1(32'h3cca5a15),
	.w2(32'hbc514755),
	.w3(32'h3c82ac97),
	.w4(32'h3c38c2f7),
	.w5(32'hbc3c7969),
	.w6(32'hbc97683e),
	.w7(32'hbcb11e52),
	.w8(32'hbb01fa10),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ba1a9),
	.w1(32'hbc69d3ff),
	.w2(32'hbc1bcb4a),
	.w3(32'hbc4ad323),
	.w4(32'hbc2c6dcc),
	.w5(32'h3b897aa2),
	.w6(32'h3c3e2afa),
	.w7(32'h3c537bd0),
	.w8(32'hb9eb3dc1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fbb87),
	.w1(32'hbb8487c2),
	.w2(32'h3b5d48eb),
	.w3(32'h3cb5c759),
	.w4(32'h3ca919ea),
	.w5(32'h3bd6a561),
	.w6(32'h3ccfe70e),
	.w7(32'h3cb92174),
	.w8(32'hbaf367ce),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ea682),
	.w1(32'hbbc23e80),
	.w2(32'hbb4fb7a8),
	.w3(32'hbb45fb8a),
	.w4(32'hbc08c9c5),
	.w5(32'h3947c16f),
	.w6(32'h3c218acb),
	.w7(32'h3b65efc8),
	.w8(32'h3b431101),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0f96f),
	.w1(32'h3b500e2a),
	.w2(32'h39810290),
	.w3(32'hbb11d50c),
	.w4(32'hbaedd0d8),
	.w5(32'hb9c2d807),
	.w6(32'h3b2763cc),
	.w7(32'hbc4fd1d4),
	.w8(32'hbb41afd0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcc7dc),
	.w1(32'h3b60b4fc),
	.w2(32'h3a3ecf27),
	.w3(32'h3b92f676),
	.w4(32'h3afe9892),
	.w5(32'hb889fe0e),
	.w6(32'h3bb100c3),
	.w7(32'h3a284074),
	.w8(32'hbaf07daf),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3aef7),
	.w1(32'h3b527b98),
	.w2(32'hbbb20332),
	.w3(32'hbb13a30b),
	.w4(32'h39b1120e),
	.w5(32'h3c0e13c6),
	.w6(32'h3b1cf5ed),
	.w7(32'h3b4be3fe),
	.w8(32'hbb67ba20),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84bc11),
	.w1(32'hbcee6dd5),
	.w2(32'hbbb8ece8),
	.w3(32'h3a879776),
	.w4(32'h3bae2171),
	.w5(32'hbbd4b080),
	.w6(32'hbaa5da47),
	.w7(32'h3c2a0025),
	.w8(32'hba93a5f1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd37c1b),
	.w1(32'hbbcaa3ba),
	.w2(32'hbc2137e5),
	.w3(32'hbb991b1b),
	.w4(32'hbbb3ae97),
	.w5(32'hbc4dc3a7),
	.w6(32'h3be849f6),
	.w7(32'hba1310dd),
	.w8(32'hbb91fefb),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75e30e),
	.w1(32'h3b4d2e08),
	.w2(32'h3cac65a9),
	.w3(32'hbcf5838a),
	.w4(32'h3b5c450f),
	.w5(32'h3c9d28e5),
	.w6(32'h3c80ee0f),
	.w7(32'h3ca086b1),
	.w8(32'h3be76b7d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba334be),
	.w1(32'hba3ab52a),
	.w2(32'h3bb714c5),
	.w3(32'h3bbbc55f),
	.w4(32'h3b25fe8b),
	.w5(32'h3c5b05a7),
	.w6(32'h3b4ef629),
	.w7(32'h3c1a6943),
	.w8(32'h3bb807ee),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d69444),
	.w1(32'hbc49ed4e),
	.w2(32'h3bbf86b0),
	.w3(32'h3ca3bacb),
	.w4(32'h3a6eecee),
	.w5(32'hbad75da7),
	.w6(32'h3c41a055),
	.w7(32'hbaf51015),
	.w8(32'hbbdd9121),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule