module layer_10_featuremap_230(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15c353),
	.w1(32'h3b43988d),
	.w2(32'h3acc394b),
	.w3(32'hbb14bf57),
	.w4(32'hbb979d13),
	.w5(32'h3d47bc5d),
	.w6(32'hbaf50974),
	.w7(32'h3b0fba6e),
	.w8(32'h3a8eb720),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe969dc),
	.w1(32'h3c57717c),
	.w2(32'h3b360162),
	.w3(32'hbc128051),
	.w4(32'h3bb35597),
	.w5(32'hba20b9fe),
	.w6(32'hbb7dd91a),
	.w7(32'h3c0a112e),
	.w8(32'hba0be5c5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a5592),
	.w1(32'hbaa01920),
	.w2(32'hbc992d23),
	.w3(32'h3b231a3c),
	.w4(32'h3cc5193a),
	.w5(32'hbb8850a8),
	.w6(32'hbb895a79),
	.w7(32'h39b8b73b),
	.w8(32'hbba6147c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc194079),
	.w1(32'hbbfda082),
	.w2(32'hbad2ac4f),
	.w3(32'hbbe674e7),
	.w4(32'hba84bdbd),
	.w5(32'hbc38e9fe),
	.w6(32'hbc368779),
	.w7(32'hba6397ee),
	.w8(32'h3b9edcb0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f35ee),
	.w1(32'hbbe48690),
	.w2(32'hbbb5341e),
	.w3(32'hbc1f3788),
	.w4(32'hbb7efd52),
	.w5(32'h3b9369f0),
	.w6(32'hba7c804d),
	.w7(32'hbb98cb45),
	.w8(32'hb892eca8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc087845),
	.w1(32'hbb41dde6),
	.w2(32'hbb739b9e),
	.w3(32'hbbc6ba58),
	.w4(32'hbb082dfc),
	.w5(32'h3c5ee21a),
	.w6(32'h3c42b8a9),
	.w7(32'hbbf99d57),
	.w8(32'hbb998778),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23b519),
	.w1(32'hbb875c0b),
	.w2(32'hb8284522),
	.w3(32'h3c1a5d13),
	.w4(32'h3b92bf9f),
	.w5(32'h3b98ebb2),
	.w6(32'h3c1eda01),
	.w7(32'hb9cc68d5),
	.w8(32'hbb2753e6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fb8cc),
	.w1(32'h3c53fb59),
	.w2(32'hbc2f3690),
	.w3(32'hbbf82fa2),
	.w4(32'h3bfe5389),
	.w5(32'h3a5b3816),
	.w6(32'hbc3b1ea6),
	.w7(32'h3b2072b8),
	.w8(32'hbbb068bf),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80baa6),
	.w1(32'hbb07b56b),
	.w2(32'h3a4de3fe),
	.w3(32'h3b5553d8),
	.w4(32'h3ad7a15a),
	.w5(32'hbb9850ce),
	.w6(32'h3b014b6d),
	.w7(32'h3acb4a36),
	.w8(32'hbafc3615),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85b57f),
	.w1(32'hb9bf1340),
	.w2(32'hbcd573ca),
	.w3(32'hbbf8c0d4),
	.w4(32'hba238203),
	.w5(32'hbb04e55e),
	.w6(32'h3b051c05),
	.w7(32'hbc2ded43),
	.w8(32'hbb77f59e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aead7f),
	.w1(32'hb9b941d6),
	.w2(32'hbc095934),
	.w3(32'h3bbf1296),
	.w4(32'hbbc887aa),
	.w5(32'h3b67458c),
	.w6(32'hbb35f8d3),
	.w7(32'hbc158443),
	.w8(32'hbbebf75c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7868c),
	.w1(32'h3b1da224),
	.w2(32'hbad0357c),
	.w3(32'hb89b0dce),
	.w4(32'h3be5ed26),
	.w5(32'hbb0bad22),
	.w6(32'h3acea396),
	.w7(32'hb94a841d),
	.w8(32'hbb899b73),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5ca35),
	.w1(32'hbc204178),
	.w2(32'h3c200cdf),
	.w3(32'hbaeb72bd),
	.w4(32'hbb5be566),
	.w5(32'h3c0936ac),
	.w6(32'h3c05fef3),
	.w7(32'h3bcb9228),
	.w8(32'hbb7ce118),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4694a),
	.w1(32'h3b833121),
	.w2(32'h3b84d139),
	.w3(32'h3b232a52),
	.w4(32'h3bbde439),
	.w5(32'hbbaaf963),
	.w6(32'hbabaed3b),
	.w7(32'h3bdea016),
	.w8(32'hba546a5a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47a044),
	.w1(32'hbbf76d82),
	.w2(32'hbbe07322),
	.w3(32'h3baa5701),
	.w4(32'hbc132cb5),
	.w5(32'h3c2e9b13),
	.w6(32'hbc70fc11),
	.w7(32'hbb0c9cfb),
	.w8(32'h3b565764),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ce671),
	.w1(32'hbc03c501),
	.w2(32'hbc58144a),
	.w3(32'h3bf19cce),
	.w4(32'hbb03bed4),
	.w5(32'hbb7ec589),
	.w6(32'h3ba97ad9),
	.w7(32'h3a6bb961),
	.w8(32'h3bad1b8b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4622c8),
	.w1(32'hbb22819c),
	.w2(32'h3ba816be),
	.w3(32'h3b2c433c),
	.w4(32'hb7aab733),
	.w5(32'h3b8c1ac2),
	.w6(32'h3b670af6),
	.w7(32'hbaa55c1f),
	.w8(32'h3b908fe3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf451c0),
	.w1(32'hbb47e2d0),
	.w2(32'hb9ad934b),
	.w3(32'hbc0133a8),
	.w4(32'hbbcfa962),
	.w5(32'hb8d387da),
	.w6(32'hbad5828b),
	.w7(32'h3c015937),
	.w8(32'h3b782a6d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b758999),
	.w1(32'hbc7d4c42),
	.w2(32'hbbb372f2),
	.w3(32'hbc5b18d2),
	.w4(32'hb9f6aa3e),
	.w5(32'hbb4ccef5),
	.w6(32'h3ad480bd),
	.w7(32'h3bd06ba4),
	.w8(32'h3b36d8fa),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62b4d8),
	.w1(32'hbb01c535),
	.w2(32'h3c1849fc),
	.w3(32'hbc34bf8c),
	.w4(32'hbbe4c429),
	.w5(32'hbbabfb9b),
	.w6(32'hbbb956a6),
	.w7(32'hbb070180),
	.w8(32'hbb540d63),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82ecb2),
	.w1(32'hbbffbdb4),
	.w2(32'h3c6a101f),
	.w3(32'h3b1e4a4d),
	.w4(32'h3abf1cfc),
	.w5(32'hbc8a5502),
	.w6(32'hbadf6df6),
	.w7(32'h3b7956a5),
	.w8(32'h3a8e6f51),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccbe4eb),
	.w1(32'h3b23c416),
	.w2(32'hb8e43461),
	.w3(32'hba7534b5),
	.w4(32'h3aba2c48),
	.w5(32'hba9e0781),
	.w6(32'h3aeb5b38),
	.w7(32'h39440eb4),
	.w8(32'hbb9678bb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b400c9c),
	.w1(32'hba811734),
	.w2(32'hb6f9984b),
	.w3(32'hbc39d4c8),
	.w4(32'hbb85b0c8),
	.w5(32'h3cbf8aa1),
	.w6(32'h3a8bba82),
	.w7(32'hbc2c12ba),
	.w8(32'hbb47bbb5),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3837bc),
	.w1(32'hbbd520a3),
	.w2(32'h3c04cdf8),
	.w3(32'hbbda9a24),
	.w4(32'hbb8112ce),
	.w5(32'hbc1f8d77),
	.w6(32'hbc3e86aa),
	.w7(32'hbb6cb530),
	.w8(32'h3b3ae764),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a992e58),
	.w1(32'h3bbe3944),
	.w2(32'hbbb01e1c),
	.w3(32'hbbb98b68),
	.w4(32'hbba3c610),
	.w5(32'hbb908b5e),
	.w6(32'hbc10dd3e),
	.w7(32'h3c3162b7),
	.w8(32'h3c2d7638),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b09a7),
	.w1(32'hbc6435b5),
	.w2(32'h3c33bd8b),
	.w3(32'hbbd24f07),
	.w4(32'h3cf5a9e7),
	.w5(32'hb9aeb8a9),
	.w6(32'h3bb97d6b),
	.w7(32'h3bc635bf),
	.w8(32'hb9ce6aa6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19ce38),
	.w1(32'hbb6f6f24),
	.w2(32'hbc47474b),
	.w3(32'h3b8442d1),
	.w4(32'h3b9575ce),
	.w5(32'hba5005e9),
	.w6(32'h3c13bacf),
	.w7(32'h3ba75cb7),
	.w8(32'h3bfe7818),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb17e67),
	.w1(32'hbc14579d),
	.w2(32'hba4e8b44),
	.w3(32'hbb6923d1),
	.w4(32'h3b060802),
	.w5(32'hbbffbf9b),
	.w6(32'h3a127aa6),
	.w7(32'h3cca385e),
	.w8(32'hbad6c5a9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd08787),
	.w1(32'h3bdf46b7),
	.w2(32'h3cb087b0),
	.w3(32'h3b2e8ab1),
	.w4(32'hbc1f5637),
	.w5(32'hbbafaccb),
	.w6(32'hbc2c42fd),
	.w7(32'h3bde51ee),
	.w8(32'hbc1cda31),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beca3e1),
	.w1(32'hba83ab5f),
	.w2(32'h3c557b9d),
	.w3(32'h3bf0ae79),
	.w4(32'h3c4293b5),
	.w5(32'hbbc2b045),
	.w6(32'h3c409628),
	.w7(32'hbc031817),
	.w8(32'hbc7c2cd8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68bc80),
	.w1(32'h3b997175),
	.w2(32'hbc98b798),
	.w3(32'hbc0b7f3f),
	.w4(32'h3830f4fb),
	.w5(32'h3c588aee),
	.w6(32'h3b35d44a),
	.w7(32'h3ad51b46),
	.w8(32'hbb6033d5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb282449),
	.w1(32'hbbc062bb),
	.w2(32'h3b94529c),
	.w3(32'hbbcf9f74),
	.w4(32'h3b57aacb),
	.w5(32'h3c881479),
	.w6(32'hba9f6ce3),
	.w7(32'hbb8014bc),
	.w8(32'h3b034dbb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6775c2),
	.w1(32'hbb18a278),
	.w2(32'hbcaf4419),
	.w3(32'h3c11bc55),
	.w4(32'hbb72ce7c),
	.w5(32'hbc8aa8fb),
	.w6(32'h3bfb41ef),
	.w7(32'hbcc5cb17),
	.w8(32'h3c632ff7),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8123c7),
	.w1(32'h3a4b201a),
	.w2(32'h3cb0dfcd),
	.w3(32'h3b8bcd89),
	.w4(32'h395ad104),
	.w5(32'h3bc4a51b),
	.w6(32'h390ca584),
	.w7(32'hbb926319),
	.w8(32'h3a490582),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc603796),
	.w1(32'hbb80f144),
	.w2(32'hbc20a86d),
	.w3(32'hbaea5777),
	.w4(32'hba5920d3),
	.w5(32'hbc35607a),
	.w6(32'h3b656629),
	.w7(32'hbc9efa9b),
	.w8(32'h3d2d55db),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb162c9c),
	.w1(32'hbba32b74),
	.w2(32'hbcd9c448),
	.w3(32'h3c0025ef),
	.w4(32'hbc9544ba),
	.w5(32'hbacd3ccd),
	.w6(32'hbcc00fb2),
	.w7(32'h3bd39611),
	.w8(32'hbb10ec51),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fd569),
	.w1(32'hbc119604),
	.w2(32'h3b4766cb),
	.w3(32'h3c1b67d4),
	.w4(32'h3c0b2647),
	.w5(32'hbd3c5a3f),
	.w6(32'hbb99d016),
	.w7(32'hbb01dc4f),
	.w8(32'hbc424763),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d7992),
	.w1(32'hbae6babc),
	.w2(32'h3c976925),
	.w3(32'hbc0df17f),
	.w4(32'hbcfe3edc),
	.w5(32'h38dd873c),
	.w6(32'h3ae9c387),
	.w7(32'h3bb3b57e),
	.w8(32'hbb9c7b8b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ba1d3),
	.w1(32'hbc27ac20),
	.w2(32'h3c6a16aa),
	.w3(32'h3d2477f7),
	.w4(32'hbbc60885),
	.w5(32'hbc12c141),
	.w6(32'hbc685104),
	.w7(32'h3a387ede),
	.w8(32'hbca6e692),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08f5ac),
	.w1(32'hbb5f7f2e),
	.w2(32'hba8f4b20),
	.w3(32'h3aa6e6b1),
	.w4(32'h3b30990b),
	.w5(32'hbbcd6fd1),
	.w6(32'h3a79f6ff),
	.w7(32'hbc4301e2),
	.w8(32'h3cabb5e9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aa1ac7),
	.w1(32'h3b50d835),
	.w2(32'hbc0e9174),
	.w3(32'h3c20bce6),
	.w4(32'hbc567e01),
	.w5(32'hbc2504e5),
	.w6(32'hbb55e85b),
	.w7(32'hbc3dabc6),
	.w8(32'hbab21e90),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37330b),
	.w1(32'hbb84ad66),
	.w2(32'hbada894e),
	.w3(32'hbba4d2b1),
	.w4(32'hbce68595),
	.w5(32'hbc040dec),
	.w6(32'h3bab1208),
	.w7(32'h3bb9c4cf),
	.w8(32'h3ce63069),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3feb2d),
	.w1(32'hbc095b3b),
	.w2(32'hbbbc12d4),
	.w3(32'hbc2af4f7),
	.w4(32'h3c7b4390),
	.w5(32'h39851181),
	.w6(32'hbabf3ec6),
	.w7(32'hbb01f25a),
	.w8(32'h3bc0745e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d7d84),
	.w1(32'hba9ac666),
	.w2(32'hbbe0386c),
	.w3(32'h3bb3a084),
	.w4(32'hbc07a5dd),
	.w5(32'hbbba6ece),
	.w6(32'hba9f83f8),
	.w7(32'hbac0c64d),
	.w8(32'hbb9a27dc),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc521a02),
	.w1(32'hbd52d2f7),
	.w2(32'hbb89dc1f),
	.w3(32'hbc026318),
	.w4(32'hbbe6ae27),
	.w5(32'hb964b099),
	.w6(32'h3baf7eec),
	.w7(32'hbb969847),
	.w8(32'h398f3cc6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f262bb),
	.w1(32'hbbdde1e1),
	.w2(32'h3c8d189a),
	.w3(32'hbc8c9d18),
	.w4(32'hbb65f354),
	.w5(32'h3c9d7e58),
	.w6(32'hba85a584),
	.w7(32'hbb37ac44),
	.w8(32'h3caa265c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f2697),
	.w1(32'h3ace2831),
	.w2(32'hbca61826),
	.w3(32'h3c4c842b),
	.w4(32'hbca387a6),
	.w5(32'h3a9adf82),
	.w6(32'h3a9457ff),
	.w7(32'hbc02d93f),
	.w8(32'hbc1b9b40),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1a4a8),
	.w1(32'h3bd9215b),
	.w2(32'hbbd1d526),
	.w3(32'h3bc4dfd3),
	.w4(32'hbc3b544d),
	.w5(32'hbc2d7fb1),
	.w6(32'hbb3373ad),
	.w7(32'hbbe1f68e),
	.w8(32'hbc614f17),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5bfde0),
	.w1(32'h3b91bb10),
	.w2(32'h3bc60702),
	.w3(32'h3a5101e1),
	.w4(32'h3bf95a6d),
	.w5(32'hbaf82bcc),
	.w6(32'hbc09e5d5),
	.w7(32'hbbd32be8),
	.w8(32'h3a874bed),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14071b),
	.w1(32'h3d0a1d91),
	.w2(32'hbbaa548e),
	.w3(32'hbcc305ed),
	.w4(32'h3c3b7d8e),
	.w5(32'h3a8e7e87),
	.w6(32'h3b71801b),
	.w7(32'h3a6dfd41),
	.w8(32'hba8589d3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9815dca),
	.w1(32'hbb04e0b3),
	.w2(32'h3a12846d),
	.w3(32'h3a872939),
	.w4(32'hba561829),
	.w5(32'hb88b7e08),
	.w6(32'hbbd689a7),
	.w7(32'hbc3cdaa0),
	.w8(32'hbb25846e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d23cc3),
	.w1(32'hb8970428),
	.w2(32'h3bae655f),
	.w3(32'hbd07f79c),
	.w4(32'hbc033734),
	.w5(32'h3b2b6b39),
	.w6(32'h3d0c720e),
	.w7(32'hbb699883),
	.w8(32'hbbad69d2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15bf38),
	.w1(32'hbb14a735),
	.w2(32'h3c306970),
	.w3(32'hba439a86),
	.w4(32'hbaefdcc5),
	.w5(32'hbc70f107),
	.w6(32'hbba10dbf),
	.w7(32'h3c279457),
	.w8(32'h3ce2f2bd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9efa27),
	.w1(32'h3d24ade5),
	.w2(32'hbbcd90dd),
	.w3(32'hbb4acad2),
	.w4(32'h3cad477f),
	.w5(32'hbcabab83),
	.w6(32'h3a50fffa),
	.w7(32'h3b05376c),
	.w8(32'h3b805f70),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ef0ed),
	.w1(32'h3c4bf7d8),
	.w2(32'hb9161829),
	.w3(32'hb8421476),
	.w4(32'hbc02b600),
	.w5(32'hbc3d576d),
	.w6(32'hbc4819e8),
	.w7(32'hbc26ed0d),
	.w8(32'hbc0fd438),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacdecd),
	.w1(32'h3baf9996),
	.w2(32'h3c2e8bf0),
	.w3(32'hbb5c889a),
	.w4(32'h3cab040c),
	.w5(32'hbb83633a),
	.w6(32'h3b67b315),
	.w7(32'hbbb75284),
	.w8(32'h3d338eb8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cae69),
	.w1(32'hba4f2dae),
	.w2(32'hbb379f58),
	.w3(32'hbb2675f1),
	.w4(32'h3b3a7606),
	.w5(32'hbba8649d),
	.w6(32'hbb361cb1),
	.w7(32'hba992979),
	.w8(32'h39e817ce),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19d11a),
	.w1(32'h3af197b2),
	.w2(32'hbbef2d58),
	.w3(32'h3af69ee0),
	.w4(32'hbae2e8ea),
	.w5(32'hbb5673bb),
	.w6(32'hbc9fa3c2),
	.w7(32'hbb69e6b4),
	.w8(32'h3c1c5dcf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bade12b),
	.w1(32'hbc094bb1),
	.w2(32'h3c457ab6),
	.w3(32'hbc01103b),
	.w4(32'hbb62f654),
	.w5(32'h3c9c2d1b),
	.w6(32'hbc0af1a0),
	.w7(32'h3aaa7e08),
	.w8(32'hbba70065),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9688798),
	.w1(32'h3bdd5978),
	.w2(32'h3c86679d),
	.w3(32'hbbc19a8f),
	.w4(32'hbc12f648),
	.w5(32'hbbcd2c12),
	.w6(32'h3a5b0624),
	.w7(32'hbbcf2d2f),
	.w8(32'h3ba3ed7f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3bcff),
	.w1(32'hbb316c24),
	.w2(32'h3bb308e0),
	.w3(32'h3af4b6dc),
	.w4(32'h3b0259ce),
	.w5(32'hbaa2bfb3),
	.w6(32'h39ff18ce),
	.w7(32'h3b24812c),
	.w8(32'h3b846271),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb9ecd),
	.w1(32'h3c23e683),
	.w2(32'hba37a114),
	.w3(32'hbb3047f0),
	.w4(32'hbbffdbbf),
	.w5(32'hbc05c738),
	.w6(32'hbc36a966),
	.w7(32'h3ba5d4be),
	.w8(32'hbb9225c7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81e171),
	.w1(32'hbac204f1),
	.w2(32'hbc9658c0),
	.w3(32'h3c0e128a),
	.w4(32'hbb81e524),
	.w5(32'h3c3eaa10),
	.w6(32'hbb665b31),
	.w7(32'h3b3da3f9),
	.w8(32'h3a21b7bd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc127875),
	.w1(32'h384eb526),
	.w2(32'h3a93cdf0),
	.w3(32'hba6eac07),
	.w4(32'hba0028ee),
	.w5(32'h3b9ed3c4),
	.w6(32'h3c7f59c1),
	.w7(32'hbbddbb76),
	.w8(32'h3b271b41),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2fc22),
	.w1(32'hbbbb81db),
	.w2(32'h3a1ab4f0),
	.w3(32'hbc50efaa),
	.w4(32'hbc356a15),
	.w5(32'h3c2515dd),
	.w6(32'hba4e895e),
	.w7(32'h3b1a40aa),
	.w8(32'h3b4c1b0f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c731195),
	.w1(32'hbc4210db),
	.w2(32'hba409c94),
	.w3(32'hbba62cfa),
	.w4(32'h3b3cceb2),
	.w5(32'h3ab216f0),
	.w6(32'h3ae4630d),
	.w7(32'hbaf79896),
	.w8(32'h3c4fce96),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c6414),
	.w1(32'hbb85fd87),
	.w2(32'h3c4ab148),
	.w3(32'hbc07f9ff),
	.w4(32'hbb5635e7),
	.w5(32'h3c6fa5ed),
	.w6(32'hb9b0fe19),
	.w7(32'h3c00d9a1),
	.w8(32'hbc874260),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d09b14a),
	.w1(32'h3bab12ae),
	.w2(32'h3b4c9c9e),
	.w3(32'hbb92a257),
	.w4(32'h3bb7f1c5),
	.w5(32'h3c09227b),
	.w6(32'hbaca402e),
	.w7(32'h3b970068),
	.w8(32'hbaf6b74c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84da53),
	.w1(32'h3ac52d60),
	.w2(32'h3b2cf71f),
	.w3(32'h3b88501c),
	.w4(32'hb94b5be9),
	.w5(32'hbcab87dd),
	.w6(32'hbba3cf81),
	.w7(32'h3ac724b0),
	.w8(32'h3bfa63b8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd62c5c),
	.w1(32'hbad0db5c),
	.w2(32'hba7ccfdb),
	.w3(32'hbbd35f6d),
	.w4(32'h3b8ff155),
	.w5(32'h3c1b71b1),
	.w6(32'h3bd8d6dc),
	.w7(32'hbc46f713),
	.w8(32'h3c0f2094),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49797a),
	.w1(32'hbbb95eb6),
	.w2(32'hbb78593c),
	.w3(32'hbba5e03e),
	.w4(32'hb98fc377),
	.w5(32'h3a2d4a08),
	.w6(32'h3be3266b),
	.w7(32'hbc90e447),
	.w8(32'h3c04bf0d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d00f3),
	.w1(32'h3ba8661e),
	.w2(32'h3b2141f0),
	.w3(32'h3b41654a),
	.w4(32'h3b2b3d94),
	.w5(32'hba97b754),
	.w6(32'hbc0528dd),
	.w7(32'h3c8edf3d),
	.w8(32'hbb8787dd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f0fd5),
	.w1(32'h3b0ae601),
	.w2(32'hbb7bb8f9),
	.w3(32'hbc09d500),
	.w4(32'hbb8b0b86),
	.w5(32'hbc0ca35e),
	.w6(32'h3a536b44),
	.w7(32'h3b9577c7),
	.w8(32'hbb472f61),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b826024),
	.w1(32'hb86d43a6),
	.w2(32'h3a7abe42),
	.w3(32'h3aafdcd7),
	.w4(32'hb906efa4),
	.w5(32'h3a21f300),
	.w6(32'hbbdeabf7),
	.w7(32'h3bdd0b0a),
	.w8(32'h3a95d144),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89e4eb),
	.w1(32'hbb58e3a2),
	.w2(32'h3a0d05b2),
	.w3(32'h3aeb2826),
	.w4(32'h395a5272),
	.w5(32'h3b693867),
	.w6(32'hbbcb28b6),
	.w7(32'hb91bf7c1),
	.w8(32'hbbdb6756),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc287089),
	.w1(32'h3b402881),
	.w2(32'hbb596048),
	.w3(32'hb9c62eec),
	.w4(32'hbb92ac51),
	.w5(32'hbb3553db),
	.w6(32'hbbf46ff4),
	.w7(32'hbbb1d028),
	.w8(32'h3c0d6107),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1971e9),
	.w1(32'h3b1b9939),
	.w2(32'h3add56dd),
	.w3(32'h3c93a899),
	.w4(32'h3bff099c),
	.w5(32'hbb90bbac),
	.w6(32'hbbf7dff1),
	.w7(32'h3b2f49a3),
	.w8(32'hbc85f59c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7c281),
	.w1(32'h3a86a74b),
	.w2(32'hba68cf8b),
	.w3(32'h39860632),
	.w4(32'hbb13bab3),
	.w5(32'hbbdb76f5),
	.w6(32'hbc01ff41),
	.w7(32'h3b25742c),
	.w8(32'h3b67644a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38326fab),
	.w1(32'h3be1adfb),
	.w2(32'hbb3c3f41),
	.w3(32'h3c3e10a2),
	.w4(32'h389246ad),
	.w5(32'h3a30550d),
	.w6(32'hbbb80b59),
	.w7(32'hbaccd000),
	.w8(32'h3b9a8d69),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9680d0),
	.w1(32'h3c21aad5),
	.w2(32'hbca42aba),
	.w3(32'hb9e9bedf),
	.w4(32'h3c12d649),
	.w5(32'h3b2432a8),
	.w6(32'h3a3d9353),
	.w7(32'hbc170d15),
	.w8(32'hbabd5485),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a4769),
	.w1(32'h3c22daf3),
	.w2(32'hbbd64528),
	.w3(32'h3bc800e8),
	.w4(32'hba62226d),
	.w5(32'h3b357a96),
	.w6(32'hbab44354),
	.w7(32'hbbf9be8f),
	.w8(32'h3ba9d291),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9aee9),
	.w1(32'hbb90aee7),
	.w2(32'hbac33c92),
	.w3(32'hbc5c2029),
	.w4(32'h3b3957ed),
	.w5(32'hbb09fd15),
	.w6(32'hbb928d62),
	.w7(32'h3c2d3ca7),
	.w8(32'hbc1e115c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c34df),
	.w1(32'hbcbb11ad),
	.w2(32'hbc0543c2),
	.w3(32'hb8faacf1),
	.w4(32'hbb932775),
	.w5(32'h3c0cb844),
	.w6(32'h3aa8135b),
	.w7(32'hbbd19a1d),
	.w8(32'hbc4f9ceb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0d7fa),
	.w1(32'h3bd323b3),
	.w2(32'hbb249a53),
	.w3(32'h3c1c75d8),
	.w4(32'hbba98c97),
	.w5(32'h3b3cbb14),
	.w6(32'hbb826de7),
	.w7(32'hbabf4227),
	.w8(32'hba0cb000),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67a7eb),
	.w1(32'hbc515e62),
	.w2(32'h3c8e992f),
	.w3(32'hbc1c962c),
	.w4(32'hbc80a2d2),
	.w5(32'hb85b3106),
	.w6(32'h3c60c814),
	.w7(32'hbc713d02),
	.w8(32'h3b40350a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e5eb9),
	.w1(32'hbc21cf6f),
	.w2(32'h3b69ad34),
	.w3(32'hbb1b518f),
	.w4(32'h3c313dd4),
	.w5(32'hbacfa41a),
	.w6(32'h3c12e5d5),
	.w7(32'hbcee200b),
	.w8(32'h39985385),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89a2596),
	.w1(32'h3ce82677),
	.w2(32'hbc9d7e3f),
	.w3(32'h3ca29106),
	.w4(32'hbb92e7eb),
	.w5(32'hbc120113),
	.w6(32'h3ae22ecb),
	.w7(32'h3b3c199a),
	.w8(32'h3afd4bcb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be198b4),
	.w1(32'hbb370d56),
	.w2(32'h3aa77aee),
	.w3(32'hbaae336c),
	.w4(32'h38999c0c),
	.w5(32'hbcba468c),
	.w6(32'h3bcabfa1),
	.w7(32'hbb3bb5a7),
	.w8(32'hbb6cac2f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57d751),
	.w1(32'hbb9df41a),
	.w2(32'h3c1f25fc),
	.w3(32'hbc35a513),
	.w4(32'hba859184),
	.w5(32'hbcbca531),
	.w6(32'hba5af517),
	.w7(32'hbc7ff78f),
	.w8(32'hbb4a40b7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe45c84),
	.w1(32'h3c1da688),
	.w2(32'h3b5d4cbd),
	.w3(32'h39b1443f),
	.w4(32'h3b3bcc75),
	.w5(32'hb8245143),
	.w6(32'hbc066422),
	.w7(32'hbbd80ff0),
	.w8(32'hbae9d0ef),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd3c99),
	.w1(32'h3bf4a8f6),
	.w2(32'h3c304735),
	.w3(32'h3a8a4dac),
	.w4(32'h3b4abad9),
	.w5(32'hb9e9b2c7),
	.w6(32'h3cc72ee5),
	.w7(32'h3ac5cbb4),
	.w8(32'hbacca8fd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b476d60),
	.w1(32'hbb508801),
	.w2(32'h3a8fe471),
	.w3(32'hb8dec1fd),
	.w4(32'h3b1003a9),
	.w5(32'hbbd9be39),
	.w6(32'hbc281a25),
	.w7(32'hbb4a13f7),
	.w8(32'h3b0934bb),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0ceea),
	.w1(32'hbba98802),
	.w2(32'hb9c6b75e),
	.w3(32'h3bcb61e6),
	.w4(32'h3c0ed2ac),
	.w5(32'h3be623c2),
	.w6(32'h3c8b493b),
	.w7(32'hbbf0a04b),
	.w8(32'hbbb9cfac),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd08df9),
	.w1(32'h3c40e3bc),
	.w2(32'hbc9e539c),
	.w3(32'h3a92c6ac),
	.w4(32'h3b002f6e),
	.w5(32'h3b7d678d),
	.w6(32'h3c102a33),
	.w7(32'h3aa9087c),
	.w8(32'h3c019757),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf4d6a8),
	.w1(32'h3c473a71),
	.w2(32'hb8dd97e4),
	.w3(32'hbaf14b9c),
	.w4(32'h3b4054a4),
	.w5(32'hbc08bab8),
	.w6(32'h3a848fdb),
	.w7(32'h3a9cebfe),
	.w8(32'hbba01e03),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07a3f4),
	.w1(32'hbba085fd),
	.w2(32'hbc04d6d5),
	.w3(32'hbba3d645),
	.w4(32'h39ca79d5),
	.w5(32'h3c0fe703),
	.w6(32'h3b93af23),
	.w7(32'h3b515421),
	.w8(32'h3b99ab61),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb752c4c),
	.w1(32'hbc27bd34),
	.w2(32'h3bb85b78),
	.w3(32'h3bcbe9be),
	.w4(32'h3b83495b),
	.w5(32'h3c8c811c),
	.w6(32'hbaf0dd58),
	.w7(32'h3b53098c),
	.w8(32'hb925fb3d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47b609),
	.w1(32'hbbe9f3e0),
	.w2(32'hbc2d9e35),
	.w3(32'hbab66d62),
	.w4(32'hb9c24fd0),
	.w5(32'hbc18ff78),
	.w6(32'hbb800cd5),
	.w7(32'hba6caaa9),
	.w8(32'h38502720),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42b3ad),
	.w1(32'hbd831c7b),
	.w2(32'h3a85d0fc),
	.w3(32'hbc7f92ae),
	.w4(32'h3b7b5c81),
	.w5(32'hbc895091),
	.w6(32'hbaad09eb),
	.w7(32'h3ccf2fd6),
	.w8(32'h3aea7cc8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5ba43),
	.w1(32'h3cb06466),
	.w2(32'hba83bed8),
	.w3(32'h3c79d919),
	.w4(32'hbb913d77),
	.w5(32'h3b51a81e),
	.w6(32'h3beff14f),
	.w7(32'hbb74fc10),
	.w8(32'hbb0f6fff),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad553f3),
	.w1(32'hbbf3ab49),
	.w2(32'hbb6b109e),
	.w3(32'hbbfb80aa),
	.w4(32'h3c6b3c64),
	.w5(32'hba0140e5),
	.w6(32'hb93bfe0b),
	.w7(32'hbbb944b0),
	.w8(32'hbb544381),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb962a3c),
	.w1(32'hbba783f1),
	.w2(32'h3c809221),
	.w3(32'hba83f92e),
	.w4(32'h3a380ced),
	.w5(32'h39a9ce26),
	.w6(32'hbd33239b),
	.w7(32'h3ba9c2a0),
	.w8(32'h39babcc1),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38ebd2),
	.w1(32'hb8f38fca),
	.w2(32'h3ce87a85),
	.w3(32'hbc2b2021),
	.w4(32'h3aaddec1),
	.w5(32'h3a840a2f),
	.w6(32'hbb1446cb),
	.w7(32'h3984d4d5),
	.w8(32'h3c8e4fc3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc2052a),
	.w1(32'h3b967af1),
	.w2(32'h3a0b946c),
	.w3(32'h39f34d12),
	.w4(32'h3ba7876b),
	.w5(32'h38a8927e),
	.w6(32'h380fe2a3),
	.w7(32'hbb8c8cda),
	.w8(32'h3b4f08e2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386ae5be),
	.w1(32'hbc5423fa),
	.w2(32'hb87d7c11),
	.w3(32'hbc51fdd0),
	.w4(32'h3be0da8c),
	.w5(32'hbbfb820d),
	.w6(32'h3bb5caee),
	.w7(32'hbafcb21c),
	.w8(32'hbc46a0df),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb917b),
	.w1(32'hbb33fcce),
	.w2(32'h3aeaf2d8),
	.w3(32'hbb7adea0),
	.w4(32'hbc12ee39),
	.w5(32'hbbbce48d),
	.w6(32'h3c6ad24a),
	.w7(32'h3ac5642f),
	.w8(32'h3ad4f5e5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce5383),
	.w1(32'h3b4d7f68),
	.w2(32'hbc9da878),
	.w3(32'hbb85c7f9),
	.w4(32'hb97958ef),
	.w5(32'h3ad0a5de),
	.w6(32'hbb7c3790),
	.w7(32'hbc676a64),
	.w8(32'hb96b666e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c231d0b),
	.w1(32'hbb334028),
	.w2(32'hb88a9106),
	.w3(32'hbb8eecfd),
	.w4(32'h3bc18023),
	.w5(32'h3ae2a814),
	.w6(32'hbbbbe677),
	.w7(32'h3a7a6afb),
	.w8(32'hb9d7026d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc69237),
	.w1(32'hbcba483e),
	.w2(32'hbc627889),
	.w3(32'hbbd5acac),
	.w4(32'h3b8a04d7),
	.w5(32'hba1ac173),
	.w6(32'h3d190e9f),
	.w7(32'hb9ad3077),
	.w8(32'hbcfa675d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba02e7b),
	.w1(32'hbbbeec48),
	.w2(32'h3b912f54),
	.w3(32'h3c3af9c9),
	.w4(32'h3af270b7),
	.w5(32'h3d61e1d1),
	.w6(32'hbad8513a),
	.w7(32'hbb5b54e1),
	.w8(32'h3ac14e99),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47032c),
	.w1(32'hbc0174c7),
	.w2(32'h3b405525),
	.w3(32'hbbbb0633),
	.w4(32'hbc01b950),
	.w5(32'hbc7264d9),
	.w6(32'h3c7c1de5),
	.w7(32'hbbc2c80b),
	.w8(32'hba32965b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c89b3),
	.w1(32'hbb731128),
	.w2(32'h3cdf82db),
	.w3(32'h3ac7dfdc),
	.w4(32'hbbf3797d),
	.w5(32'h3aea5fd3),
	.w6(32'h3b95bc26),
	.w7(32'hbc000ff2),
	.w8(32'h3adb567b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad85f84),
	.w1(32'hbb237542),
	.w2(32'hba70d3fa),
	.w3(32'hbaf9c8a5),
	.w4(32'hbc337868),
	.w5(32'hbb70627c),
	.w6(32'hbb6fb179),
	.w7(32'hb78e36d3),
	.w8(32'hbc96cd2d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cb41d),
	.w1(32'hbbae2c14),
	.w2(32'hbbfd704d),
	.w3(32'h3a489da3),
	.w4(32'h3c4a29d8),
	.w5(32'h3ab53bed),
	.w6(32'hbc0619f2),
	.w7(32'hbb3e567b),
	.w8(32'hbadd36db),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12e893),
	.w1(32'hbc442049),
	.w2(32'hbb939da8),
	.w3(32'h3bb12d58),
	.w4(32'hbc833002),
	.w5(32'hbb11e850),
	.w6(32'hbb27ab77),
	.w7(32'h3c3e9e9f),
	.w8(32'h3c47e718),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca274be),
	.w1(32'h3cd8d93d),
	.w2(32'hbbdea6bc),
	.w3(32'hba760bfe),
	.w4(32'hbaf88055),
	.w5(32'hbc02167f),
	.w6(32'h3a2fe298),
	.w7(32'h3b680707),
	.w8(32'h3be102d3),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc109910),
	.w1(32'h3a8e60c5),
	.w2(32'hbb869d42),
	.w3(32'hbc366428),
	.w4(32'h3c869207),
	.w5(32'h3b52728e),
	.w6(32'h3bbc3063),
	.w7(32'h358b13d4),
	.w8(32'hb96f5c8e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa9081),
	.w1(32'hbc898f28),
	.w2(32'h3b6a10e9),
	.w3(32'h3bdf9b0d),
	.w4(32'h3bb9edc7),
	.w5(32'h3c0711df),
	.w6(32'h3bb1ba9f),
	.w7(32'hbc209b92),
	.w8(32'hbb8be368),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18709b),
	.w1(32'h3bafb790),
	.w2(32'hbac780dc),
	.w3(32'h3cdc6b09),
	.w4(32'hba505e9d),
	.w5(32'hbc042181),
	.w6(32'hbabcc9b8),
	.w7(32'h3b2637c0),
	.w8(32'h3aa81a10),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd61d4),
	.w1(32'hbb9a87fc),
	.w2(32'h3a9f9c5d),
	.w3(32'hbc0b7219),
	.w4(32'hbba67791),
	.w5(32'hbae8ac64),
	.w6(32'h38e53a08),
	.w7(32'h3be501ae),
	.w8(32'h3c56b6f5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07868b),
	.w1(32'hbb683706),
	.w2(32'h3b311087),
	.w3(32'hb872a9b1),
	.w4(32'h3cfc42eb),
	.w5(32'hbb9b9ec3),
	.w6(32'hbcdeb0cf),
	.w7(32'h3bf97fb7),
	.w8(32'hbc3ded66),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f19c2),
	.w1(32'h3b899b17),
	.w2(32'h3c2cc6b2),
	.w3(32'hbaaaaa9b),
	.w4(32'h3bdbe8ed),
	.w5(32'h3b0f07da),
	.w6(32'h3c0ff395),
	.w7(32'h3b0d1ed2),
	.w8(32'h3bdecd5e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08e88c),
	.w1(32'hbb6090e3),
	.w2(32'hb8b61645),
	.w3(32'hbc257645),
	.w4(32'h3a58d1ad),
	.w5(32'h3b98b245),
	.w6(32'hbba04e12),
	.w7(32'h3a05db9a),
	.w8(32'hb9b598ac),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6f2b9),
	.w1(32'h3aa1355b),
	.w2(32'h3c3eefb7),
	.w3(32'hb84bbf3a),
	.w4(32'hbbe73f26),
	.w5(32'h3aca6be7),
	.w6(32'h3c89e58f),
	.w7(32'hbb35c5ca),
	.w8(32'hbb7e5abb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb23df),
	.w1(32'hbba45d78),
	.w2(32'hbb851bf0),
	.w3(32'hbad1fe27),
	.w4(32'h3b4923f6),
	.w5(32'hbbeaaf57),
	.w6(32'h3ba719cd),
	.w7(32'h3b61a7d6),
	.w8(32'hbac853c0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a08b7),
	.w1(32'hb5b6014e),
	.w2(32'h3c9fa940),
	.w3(32'hbb147f22),
	.w4(32'h38acb087),
	.w5(32'h3c8d0d01),
	.w6(32'h3a2db087),
	.w7(32'hbac97417),
	.w8(32'hbb1b9de9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abea8ea),
	.w1(32'hb8c67de9),
	.w2(32'hbb0e1ba3),
	.w3(32'hbc083202),
	.w4(32'h3c7b3bb8),
	.w5(32'hbc281aa0),
	.w6(32'hbbb6a8e6),
	.w7(32'hbce3b61d),
	.w8(32'hbc0c3626),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd3db07),
	.w1(32'hbb6e6cb7),
	.w2(32'hbb1e699c),
	.w3(32'h3c252a22),
	.w4(32'h3d160f9a),
	.w5(32'hbc045e9b),
	.w6(32'h3adeac06),
	.w7(32'h3cafbc78),
	.w8(32'hbc0423f3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb128435),
	.w1(32'h37aecc75),
	.w2(32'h38350eb7),
	.w3(32'h3c7235cc),
	.w4(32'hbadb6852),
	.w5(32'h3a030ee8),
	.w6(32'hbc03bb93),
	.w7(32'hbc2ac3ae),
	.w8(32'h3ac97202),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc09f3a),
	.w1(32'hba243e63),
	.w2(32'hbada4745),
	.w3(32'hbb49e155),
	.w4(32'h3c2c60d1),
	.w5(32'h3c07255a),
	.w6(32'hbbf2f4b6),
	.w7(32'hbc2f1e43),
	.w8(32'hbc285d3b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1392a1),
	.w1(32'hbbe4e375),
	.w2(32'hbbe3e127),
	.w3(32'hbbb3343d),
	.w4(32'hbb96a1e0),
	.w5(32'hbb1839dd),
	.w6(32'h38b71760),
	.w7(32'hbc603008),
	.w8(32'hbc38deb6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba550c),
	.w1(32'h3bcfd081),
	.w2(32'hbb4d169f),
	.w3(32'hbc03e362),
	.w4(32'hbbaa4112),
	.w5(32'h3c0a3c54),
	.w6(32'hbb3fbcfe),
	.w7(32'hb9ff874c),
	.w8(32'hbb63270b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47f629),
	.w1(32'h3be8f3ba),
	.w2(32'h3bbb8a20),
	.w3(32'hb9ca0c39),
	.w4(32'h3cbf7a43),
	.w5(32'h3b1f99ea),
	.w6(32'hbc60db35),
	.w7(32'h3ace5ee5),
	.w8(32'hb92807b4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54cb29),
	.w1(32'hbad8ceb8),
	.w2(32'hba2e7247),
	.w3(32'hbbd0e0e1),
	.w4(32'hbc4125e8),
	.w5(32'h3c8c3759),
	.w6(32'h3bb14a18),
	.w7(32'hbbd8e874),
	.w8(32'hbc2e3600),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc1222),
	.w1(32'hbc09753a),
	.w2(32'hbc889efd),
	.w3(32'hbc05e0d8),
	.w4(32'hbc8de786),
	.w5(32'h3c126e17),
	.w6(32'h3c09052c),
	.w7(32'hba0bc9e2),
	.w8(32'h39deb0a7),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a915c),
	.w1(32'h38cbbda1),
	.w2(32'h3af262b1),
	.w3(32'h3c255dff),
	.w4(32'hbbb1ae33),
	.w5(32'hbb272309),
	.w6(32'h3b758066),
	.w7(32'h38a1ba5f),
	.w8(32'hbc10e101),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e366a),
	.w1(32'hbbcb5ba1),
	.w2(32'hbc8434a5),
	.w3(32'hb95dbe76),
	.w4(32'h3bfd66c7),
	.w5(32'hbb0a5791),
	.w6(32'hbbebd5d1),
	.w7(32'h372594dd),
	.w8(32'h3a8e198f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe2c5f),
	.w1(32'hbaf25cff),
	.w2(32'hb9f7428a),
	.w3(32'h3c651904),
	.w4(32'h3a87ebd1),
	.w5(32'hbb359f43),
	.w6(32'hbbfb53e3),
	.w7(32'h38dcccb9),
	.w8(32'h3b56f651),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda7dfe),
	.w1(32'hbc36efda),
	.w2(32'h3c8e3f41),
	.w3(32'h3c5e2d48),
	.w4(32'hbacbebc6),
	.w5(32'h3c1d1944),
	.w6(32'h3bbffb53),
	.w7(32'h3b855f0d),
	.w8(32'hbbbecbc7),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba447311),
	.w1(32'h3c7bf7b0),
	.w2(32'hbc84f9ed),
	.w3(32'h3c07ac39),
	.w4(32'h3cc8cbe1),
	.w5(32'h3bc6fe8f),
	.w6(32'hbc9f29ad),
	.w7(32'h39194e94),
	.w8(32'h3b9db199),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04078c),
	.w1(32'h3cbb5894),
	.w2(32'h3a9e29dc),
	.w3(32'hbbd73d86),
	.w4(32'h3bb03048),
	.w5(32'hbb5d43ce),
	.w6(32'hbb2bf3eb),
	.w7(32'h3a451fe4),
	.w8(32'hbb904faf),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb932dcd),
	.w1(32'hba8eebef),
	.w2(32'h3acaa6e7),
	.w3(32'hbbb8f99e),
	.w4(32'h3961cf19),
	.w5(32'h3b9e4d3d),
	.w6(32'h3c0c9b3f),
	.w7(32'hbc9cce4c),
	.w8(32'h3a439553),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1164b1),
	.w1(32'hbb489677),
	.w2(32'h3a9412fa),
	.w3(32'hbbf2a9fd),
	.w4(32'h3b85d7c3),
	.w5(32'h3a8b3dce),
	.w6(32'h3bdab067),
	.w7(32'hbc5c7eea),
	.w8(32'hbb3fa446),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83f662),
	.w1(32'h3a3bc5ef),
	.w2(32'hb9f50276),
	.w3(32'hbb6fae49),
	.w4(32'hba89e51a),
	.w5(32'h3b91431f),
	.w6(32'h3caac365),
	.w7(32'h3bef7810),
	.w8(32'h3bc4cb00),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea767e),
	.w1(32'h3baa2091),
	.w2(32'hbbce45a3),
	.w3(32'hbc226058),
	.w4(32'hbcc6a694),
	.w5(32'h3b5cf696),
	.w6(32'h3ba852de),
	.w7(32'hbbdbbd77),
	.w8(32'hbc016317),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc155e),
	.w1(32'h3b8bdcd5),
	.w2(32'h3bee1a0d),
	.w3(32'hbc0221f1),
	.w4(32'hbaac598a),
	.w5(32'h3b915939),
	.w6(32'hba408d91),
	.w7(32'hb9923480),
	.w8(32'hbbcbfdbf),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b09da),
	.w1(32'hbabbc2e1),
	.w2(32'h3b2ef369),
	.w3(32'hbac98860),
	.w4(32'h3b28ac9e),
	.w5(32'hbc1176fe),
	.w6(32'hba0e34df),
	.w7(32'h3c424b08),
	.w8(32'hbabc7ead),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381874da),
	.w1(32'hbb63168a),
	.w2(32'h3b19622e),
	.w3(32'hbcfc5bf6),
	.w4(32'h3aa5526d),
	.w5(32'h3b57b32c),
	.w6(32'hbbf9fb2c),
	.w7(32'hbbcf7724),
	.w8(32'hbb924596),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd3a73),
	.w1(32'hbb80b262),
	.w2(32'h3c8f1347),
	.w3(32'h3b8541e7),
	.w4(32'h3be83afa),
	.w5(32'hbba45868),
	.w6(32'hb9ec3fef),
	.w7(32'h3b5742b1),
	.w8(32'h3b9c7786),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd77cb3),
	.w1(32'hb98df76c),
	.w2(32'hbb041f41),
	.w3(32'h3b11a22a),
	.w4(32'h3b24a3bd),
	.w5(32'hbbde5c10),
	.w6(32'h3b158ed9),
	.w7(32'hbc19813a),
	.w8(32'h3bd68696),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a534b70),
	.w1(32'hbb074fae),
	.w2(32'h3a20ce58),
	.w3(32'h3b714138),
	.w4(32'hbaa343a4),
	.w5(32'hbc0594d0),
	.w6(32'hbc07c32b),
	.w7(32'hbb859d55),
	.w8(32'hbb8a6d87),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87ef50),
	.w1(32'h3b97aa9f),
	.w2(32'h3bec9365),
	.w3(32'h3b4b94bc),
	.w4(32'h3b953209),
	.w5(32'hbc226e6d),
	.w6(32'h3d04afec),
	.w7(32'h392e0c0a),
	.w8(32'hbb69703d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12c317),
	.w1(32'h3ab5ad1b),
	.w2(32'h3c35cf1c),
	.w3(32'h3ab004fe),
	.w4(32'hb9014413),
	.w5(32'h3a3db831),
	.w6(32'h3bc46aa1),
	.w7(32'h3bd30a86),
	.w8(32'h3c3f1916),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1321ee),
	.w1(32'hbb03bfbe),
	.w2(32'h3ca79d59),
	.w3(32'hbb22aa58),
	.w4(32'h3aecb71e),
	.w5(32'hb824f89b),
	.w6(32'h3bd59755),
	.w7(32'hbb23f432),
	.w8(32'h3bab5c92),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ab329),
	.w1(32'h3b86f561),
	.w2(32'h3b04291a),
	.w3(32'hbbfc5bea),
	.w4(32'h3b0a151f),
	.w5(32'hb9a00516),
	.w6(32'hbae18944),
	.w7(32'h3a6dc9cb),
	.w8(32'h3b5defc4),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fcf57),
	.w1(32'hbb49ef0e),
	.w2(32'hbd0798f3),
	.w3(32'h3bc11e30),
	.w4(32'hbc3477f1),
	.w5(32'h3affcdf8),
	.w6(32'hbc851c0a),
	.w7(32'h3b8d9beb),
	.w8(32'hbb5f3087),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb4b41),
	.w1(32'h3bb63dd7),
	.w2(32'hbbe6df6c),
	.w3(32'h3aea8192),
	.w4(32'hbb78c505),
	.w5(32'hbbd09ccf),
	.w6(32'hbbe7d863),
	.w7(32'h3c0948c7),
	.w8(32'hbaf895f3),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6e6eb),
	.w1(32'hbb3de627),
	.w2(32'hbabbc051),
	.w3(32'h3a359367),
	.w4(32'hbb9d814e),
	.w5(32'h3b76f488),
	.w6(32'hbb71d0f1),
	.w7(32'h3b1d6392),
	.w8(32'h3b0192ec),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba21758),
	.w1(32'hbb8428db),
	.w2(32'hb8ad7ef4),
	.w3(32'h3c05aed2),
	.w4(32'h3acce982),
	.w5(32'hbc08f441),
	.w6(32'hbae8941f),
	.w7(32'hba2f82b7),
	.w8(32'hbbc4510b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f1962),
	.w1(32'h3bd7226f),
	.w2(32'h3805e7ec),
	.w3(32'hbabf27b0),
	.w4(32'h39f52766),
	.w5(32'hbcccb63f),
	.w6(32'h3a97859d),
	.w7(32'hbbd480ce),
	.w8(32'h3bad3a61),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba198066),
	.w1(32'h3abcfb5d),
	.w2(32'h3b354e39),
	.w3(32'hbb7c1c49),
	.w4(32'h3ae5acd2),
	.w5(32'hbb3fad6a),
	.w6(32'h3acdcb1b),
	.w7(32'h39f682e2),
	.w8(32'hbaf4ac8f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ae731),
	.w1(32'hbb022ae4),
	.w2(32'h3cb5e2cd),
	.w3(32'hbb80da46),
	.w4(32'hb9120750),
	.w5(32'hba9f6e85),
	.w6(32'hbbaa575d),
	.w7(32'hba99bbfe),
	.w8(32'h3b80e159),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2fa3f),
	.w1(32'h3b32809c),
	.w2(32'hba636d9e),
	.w3(32'hbc2581ac),
	.w4(32'h3bb45c73),
	.w5(32'h3b14f64e),
	.w6(32'hbb435390),
	.w7(32'hbc217821),
	.w8(32'h3cf5a749),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6f609),
	.w1(32'hbab5d9b2),
	.w2(32'hbb6020be),
	.w3(32'hbbbf28b8),
	.w4(32'h3b665eec),
	.w5(32'hb85e529a),
	.w6(32'h3ba65c51),
	.w7(32'h3a43c701),
	.w8(32'hbb935856),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d0625),
	.w1(32'hbb01ca40),
	.w2(32'h3ba3fbeb),
	.w3(32'h3b5981fe),
	.w4(32'hba8f42ad),
	.w5(32'hbc059b8a),
	.w6(32'hbc308e3a),
	.w7(32'h393f0836),
	.w8(32'hbd54c7d0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73844a),
	.w1(32'h3ac62c56),
	.w2(32'h3b7f0bd6),
	.w3(32'hbc82dd17),
	.w4(32'h395129b8),
	.w5(32'h3c4f8a08),
	.w6(32'h3bd9cfbf),
	.w7(32'h3c1615c2),
	.w8(32'hba993f86),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb903bb85),
	.w1(32'h3b13293b),
	.w2(32'hbcbc8b30),
	.w3(32'hbbffd4d2),
	.w4(32'h3b2918a2),
	.w5(32'hbb3dcb7d),
	.w6(32'h3abbdbfd),
	.w7(32'h3b61147a),
	.w8(32'h3b4c023a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5e31f),
	.w1(32'h3be05870),
	.w2(32'hbcaa8cfb),
	.w3(32'hbc1f70c2),
	.w4(32'hbadab8bf),
	.w5(32'hbabe31de),
	.w6(32'hbc85370d),
	.w7(32'hbb2f3a8b),
	.w8(32'h3c3bd585),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a791218),
	.w1(32'hb9ce218a),
	.w2(32'hbb7334c4),
	.w3(32'h3ba2f540),
	.w4(32'h3b387e87),
	.w5(32'hbb814549),
	.w6(32'hbbba6836),
	.w7(32'h3bcf1608),
	.w8(32'h3a8c3433),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71d75b),
	.w1(32'h3bb5bb4c),
	.w2(32'h3c4f55bc),
	.w3(32'h3b289737),
	.w4(32'h3b3946a6),
	.w5(32'h3a14f485),
	.w6(32'hbc72397a),
	.w7(32'hbb56cf9e),
	.w8(32'h3bcbcb7c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bf031),
	.w1(32'h3b00ceab),
	.w2(32'h3af29339),
	.w3(32'h3ba680d5),
	.w4(32'h3bac9960),
	.w5(32'hba8289a9),
	.w6(32'h3b3fff41),
	.w7(32'hbba551fd),
	.w8(32'hbb855bc8),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d8804),
	.w1(32'hbb0e0b94),
	.w2(32'h3bc79115),
	.w3(32'hbbfb594d),
	.w4(32'hbaf2793f),
	.w5(32'h3ab7de09),
	.w6(32'h3b53cd14),
	.w7(32'hbbad8138),
	.w8(32'h3c18bd13),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e230a),
	.w1(32'hbb8485a8),
	.w2(32'h3b4da5f1),
	.w3(32'hbc0789d7),
	.w4(32'hbba95444),
	.w5(32'h3a982afc),
	.w6(32'h39cd9f33),
	.w7(32'h3bcf5e44),
	.w8(32'h3cc4b43c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52c806),
	.w1(32'hbc60ab46),
	.w2(32'hbba44b54),
	.w3(32'hbbf68784),
	.w4(32'h3c1fbc99),
	.w5(32'h3b0da546),
	.w6(32'hbb7548cf),
	.w7(32'hbac8ff87),
	.w8(32'h3b323ff0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98db35),
	.w1(32'h3bad691a),
	.w2(32'hbba636e7),
	.w3(32'h3c811b3b),
	.w4(32'hbb57af38),
	.w5(32'h3b349dc4),
	.w6(32'h3bb96256),
	.w7(32'hbc23a35c),
	.w8(32'hbc331580),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05683b),
	.w1(32'hbb7a2558),
	.w2(32'hbb1870fd),
	.w3(32'h3bb27562),
	.w4(32'hb7f3cff2),
	.w5(32'hbbce0e21),
	.w6(32'h3916fe4d),
	.w7(32'h3cdaef32),
	.w8(32'h3c02c455),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a8e79),
	.w1(32'h3b35af62),
	.w2(32'hbab41fc5),
	.w3(32'hba82c0ba),
	.w4(32'hbb9e90c7),
	.w5(32'hbb27e6a4),
	.w6(32'hbb89cd75),
	.w7(32'hba3f03c1),
	.w8(32'h3be284a5),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4cf50),
	.w1(32'h3931fee9),
	.w2(32'h3b85b3f9),
	.w3(32'hbb2387e4),
	.w4(32'h3c9adb9d),
	.w5(32'hbabd17f5),
	.w6(32'hbc2d6623),
	.w7(32'hbc414f4a),
	.w8(32'h3b5ab4c1),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85636d),
	.w1(32'h3ba2a0d5),
	.w2(32'h3ab735d7),
	.w3(32'hbb324dbb),
	.w4(32'hbb07849d),
	.w5(32'h3c04d52f),
	.w6(32'hbc2a9ac0),
	.w7(32'hbbc4bd63),
	.w8(32'hbaf9c923),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc296818),
	.w1(32'hba7fc216),
	.w2(32'hbca9a5a9),
	.w3(32'h3a5be290),
	.w4(32'h3b559d12),
	.w5(32'h3c576a25),
	.w6(32'h3af949ee),
	.w7(32'hbad5e935),
	.w8(32'h3cdc3cba),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96bf51a),
	.w1(32'h3afe2f5d),
	.w2(32'h3a1ed40c),
	.w3(32'hbb670c45),
	.w4(32'h3b8a305c),
	.w5(32'h3ba6a491),
	.w6(32'h3c215e84),
	.w7(32'h3c735ffd),
	.w8(32'h3bee7848),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb441b0),
	.w1(32'hbbb67c9d),
	.w2(32'h3b4dc4f8),
	.w3(32'hbb986a7b),
	.w4(32'hbc8fe0af),
	.w5(32'hbb3cdf61),
	.w6(32'hbbb55c5c),
	.w7(32'hbb8df075),
	.w8(32'h3ae9f0a4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b070129),
	.w1(32'hbca4fc91),
	.w2(32'hbafc80ea),
	.w3(32'hbc8a04a4),
	.w4(32'h3a2926b1),
	.w5(32'hbbccb51c),
	.w6(32'h35f866c6),
	.w7(32'hb8f3618c),
	.w8(32'hbbfcec9f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae77915),
	.w1(32'h3b3fdc61),
	.w2(32'hbc858190),
	.w3(32'hbbc38e5e),
	.w4(32'h3c3e9f26),
	.w5(32'hbb81116e),
	.w6(32'h3ba9c9e3),
	.w7(32'h3b908147),
	.w8(32'hbcc16919),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc111fd1),
	.w1(32'hbb6fd4b3),
	.w2(32'h3883a361),
	.w3(32'h3ca3d8d5),
	.w4(32'hbb2e673b),
	.w5(32'hbbae350f),
	.w6(32'hbc0c7807),
	.w7(32'h3bdcc609),
	.w8(32'hbbae5a67),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be73b79),
	.w1(32'hbbb43451),
	.w2(32'hbbe05283),
	.w3(32'hbb8b4563),
	.w4(32'h3bf103d2),
	.w5(32'hbba4dd71),
	.w6(32'hb9d83575),
	.w7(32'h3b2c37ff),
	.w8(32'hbb1b6505),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15c3ba),
	.w1(32'hba32aba0),
	.w2(32'hba8c8531),
	.w3(32'hbb0245a9),
	.w4(32'h3b35a3e2),
	.w5(32'hbb22283d),
	.w6(32'h3b9f004d),
	.w7(32'h3cfa509e),
	.w8(32'h3aef8e5d),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a927521),
	.w1(32'h3b95b15d),
	.w2(32'hba71c7ef),
	.w3(32'h395f6e91),
	.w4(32'h3c654767),
	.w5(32'h3b43fe40),
	.w6(32'h39a00486),
	.w7(32'h3a2af3b9),
	.w8(32'h3c0c2ce0),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad02830),
	.w1(32'h3c90650f),
	.w2(32'h3a9c5aba),
	.w3(32'h3c06cab7),
	.w4(32'h3abeda70),
	.w5(32'h3ac50933),
	.w6(32'h3c883580),
	.w7(32'hbb6b6bf5),
	.w8(32'hba9d3fa0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddffbb),
	.w1(32'hbb8fe61f),
	.w2(32'h3b94456e),
	.w3(32'h3b43870b),
	.w4(32'h3cc95cf9),
	.w5(32'hbaaf8015),
	.w6(32'h3c41f8fb),
	.w7(32'hbbb7f2a3),
	.w8(32'hba8d8001),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3955f356),
	.w1(32'h3c1bb2c8),
	.w2(32'hbc59b2b4),
	.w3(32'hbcf82847),
	.w4(32'hbbce04a2),
	.w5(32'hbb49d06f),
	.w6(32'hbbc79a7a),
	.w7(32'hbad3abcf),
	.w8(32'h39683368),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b31d4),
	.w1(32'hbab2d8d5),
	.w2(32'h3bf0c1fc),
	.w3(32'h3b2df0f3),
	.w4(32'hbb92f534),
	.w5(32'hbb0b9dcd),
	.w6(32'h3c307eb3),
	.w7(32'hbc2cce08),
	.w8(32'hbbaeb242),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc771a2),
	.w1(32'hbb39e403),
	.w2(32'h3b4119b4),
	.w3(32'h3968f9a0),
	.w4(32'h3ad01e94),
	.w5(32'h3820550e),
	.w6(32'hb90bac70),
	.w7(32'h3bd0d777),
	.w8(32'hb855336c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9696c98),
	.w1(32'h3d3c135e),
	.w2(32'h3ca227ae),
	.w3(32'h3a6fd458),
	.w4(32'h3c52d46b),
	.w5(32'h3b0ab1f3),
	.w6(32'hbb9e1deb),
	.w7(32'hbc280bc3),
	.w8(32'hbbf19b0c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c266091),
	.w1(32'h39ef52f5),
	.w2(32'hbba65a7f),
	.w3(32'hbbaf422d),
	.w4(32'hbbe6047c),
	.w5(32'hbb4620aa),
	.w6(32'h3c8c3139),
	.w7(32'h3c0616e0),
	.w8(32'hbaa5c29e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bfd90),
	.w1(32'h3c3822e5),
	.w2(32'h3ab4481f),
	.w3(32'hbc4b51b9),
	.w4(32'h3b89a44c),
	.w5(32'h3bbde077),
	.w6(32'h3b063e25),
	.w7(32'h3c9480be),
	.w8(32'hbb068601),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cf7e9),
	.w1(32'h3bc0f050),
	.w2(32'h3b217620),
	.w3(32'h3a9aa306),
	.w4(32'hbbd55a89),
	.w5(32'hba60aa04),
	.w6(32'h3b36c3cd),
	.w7(32'h3bad85e3),
	.w8(32'h3c2bd670),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc49269),
	.w1(32'hbb94823e),
	.w2(32'hba8e5ea4),
	.w3(32'h3b420e69),
	.w4(32'h399c68fd),
	.w5(32'h3ac762fa),
	.w6(32'hbba445f3),
	.w7(32'hbb8d3225),
	.w8(32'hbbce9559),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d9e28),
	.w1(32'hbbd4f3f3),
	.w2(32'hbbfe6b03),
	.w3(32'h3c220032),
	.w4(32'hbcc634a7),
	.w5(32'hbb29b21b),
	.w6(32'hbc7f35e7),
	.w7(32'hbb7fe62e),
	.w8(32'hbb040444),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb999f11),
	.w1(32'hbc3bd3b2),
	.w2(32'hbba375bf),
	.w3(32'h3a15af40),
	.w4(32'h3b0f67da),
	.w5(32'hba788ca9),
	.w6(32'hbb88139b),
	.w7(32'hbb85764d),
	.w8(32'h361d30c5),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87add6),
	.w1(32'h3a6358a5),
	.w2(32'hbc4450a8),
	.w3(32'hbbc95157),
	.w4(32'hbb85703b),
	.w5(32'hbb3d7f60),
	.w6(32'h3a00a79b),
	.w7(32'h3bc3fb6a),
	.w8(32'hbb846667),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b91a7),
	.w1(32'hbb7741bd),
	.w2(32'hbab863b7),
	.w3(32'hbbc070b6),
	.w4(32'hbb68a91c),
	.w5(32'hbba5c258),
	.w6(32'h3b09b6b6),
	.w7(32'h3c52df45),
	.w8(32'hbafeacd9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc25b1c),
	.w1(32'hbb9a7618),
	.w2(32'hbab137dc),
	.w3(32'hbb550ad5),
	.w4(32'hbc79d4d6),
	.w5(32'hbbbcf220),
	.w6(32'hbc0fb00f),
	.w7(32'hbbb7dc40),
	.w8(32'hbbde9d7a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c111591),
	.w1(32'h3abfc61d),
	.w2(32'h3a3bb242),
	.w3(32'hbb0d9f6e),
	.w4(32'hbb92f48b),
	.w5(32'hbb042075),
	.w6(32'hbbab804a),
	.w7(32'h3aee43fe),
	.w8(32'hbaaf78d3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cff491d),
	.w1(32'h3c0dc293),
	.w2(32'h3b16f464),
	.w3(32'hbc23b61c),
	.w4(32'hbb595672),
	.w5(32'h3a5712b0),
	.w6(32'hbbb6a41d),
	.w7(32'hbaa6b0b5),
	.w8(32'h3bca00b3),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c3701),
	.w1(32'hbb7f008d),
	.w2(32'hbb23dafd),
	.w3(32'h39e40236),
	.w4(32'h3bbe09dc),
	.w5(32'h39ae991d),
	.w6(32'hbc4e2d35),
	.w7(32'hbcb610ab),
	.w8(32'hbcaaf5d7),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4ffb5),
	.w1(32'hbc24bfad),
	.w2(32'hbb95bd91),
	.w3(32'h3b5e97fd),
	.w4(32'hbc3927b4),
	.w5(32'h3c2d8954),
	.w6(32'hba85e0e1),
	.w7(32'hbb24f6b2),
	.w8(32'hbb9ef0e3),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20148a),
	.w1(32'hbc1891ef),
	.w2(32'hbbc7e5e2),
	.w3(32'h39b26a34),
	.w4(32'hbbbe4dbf),
	.w5(32'hbb9b8068),
	.w6(32'hbb768879),
	.w7(32'hba86431c),
	.w8(32'hbb8d21e2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a1f92),
	.w1(32'hbc42981e),
	.w2(32'h3b7a4fe1),
	.w3(32'hbca82a0d),
	.w4(32'h397e2340),
	.w5(32'hbb26359b),
	.w6(32'h3b71c710),
	.w7(32'hbbdac983),
	.w8(32'hbc22b20a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43f23d),
	.w1(32'h3b877854),
	.w2(32'hbb9e3712),
	.w3(32'hbaac1026),
	.w4(32'hba2b4663),
	.w5(32'h3b03c62d),
	.w6(32'hbbfd07b8),
	.w7(32'hbc4ddb6d),
	.w8(32'hb998dadf),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a6fc71),
	.w1(32'hbb3623bf),
	.w2(32'h362a61e3),
	.w3(32'h3bde75e9),
	.w4(32'h3ab532f1),
	.w5(32'hbbc0001f),
	.w6(32'hbba7c108),
	.w7(32'hbc27fafe),
	.w8(32'h39366a55),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8050cf),
	.w1(32'h3a6cccde),
	.w2(32'hbb76f31f),
	.w3(32'hbbe56783),
	.w4(32'hbbb935dc),
	.w5(32'h38f60e24),
	.w6(32'h3ae8c703),
	.w7(32'hbba269a9),
	.w8(32'h3ac072aa),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4013a),
	.w1(32'hbbbebef2),
	.w2(32'hbc388337),
	.w3(32'hbb7b5a75),
	.w4(32'hbc4dd72c),
	.w5(32'hb9209460),
	.w6(32'hbc577cd4),
	.w7(32'h3c42d3ce),
	.w8(32'hbc854c17),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8325d2),
	.w1(32'h3b8025c6),
	.w2(32'hbb920433),
	.w3(32'hbc71267c),
	.w4(32'h3a5362ab),
	.w5(32'hba9be867),
	.w6(32'h3a5c18fe),
	.w7(32'hbab410a9),
	.w8(32'hbb007ff2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df9995),
	.w1(32'h39919387),
	.w2(32'hbb0e03e3),
	.w3(32'hbb884d0d),
	.w4(32'hbbf208ce),
	.w5(32'h3b20fa5c),
	.w6(32'hbc92eeca),
	.w7(32'h39f0830a),
	.w8(32'hbbee31e7),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7c634),
	.w1(32'hba2d630a),
	.w2(32'hbc281ad8),
	.w3(32'hbb9cc5ee),
	.w4(32'hbbb1bbeb),
	.w5(32'hbb0b965e),
	.w6(32'hbb95da6a),
	.w7(32'h34a6d13a),
	.w8(32'hbb4c26c9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a2117),
	.w1(32'hbb97423b),
	.w2(32'h3cececca),
	.w3(32'hbbeeba87),
	.w4(32'hbc271ab2),
	.w5(32'h3c214e55),
	.w6(32'hba3883ce),
	.w7(32'hba9f7f5b),
	.w8(32'h39b01864),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d237e),
	.w1(32'hbb8f87f9),
	.w2(32'hb8d36b22),
	.w3(32'hb8530d55),
	.w4(32'hbb209906),
	.w5(32'hbbdd7609),
	.w6(32'hbbe91fbf),
	.w7(32'hba9d6269),
	.w8(32'hbb5935af),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6b3be),
	.w1(32'hba053b62),
	.w2(32'h3b004e22),
	.w3(32'hbc0551c0),
	.w4(32'hbb8319a8),
	.w5(32'hbb5c0c0d),
	.w6(32'hbb845df6),
	.w7(32'hbd47b6f0),
	.w8(32'hba7b9137),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07d0ae),
	.w1(32'hbbe76378),
	.w2(32'hbbca26cf),
	.w3(32'hb9b43358),
	.w4(32'hbc039ce9),
	.w5(32'hbd23fb47),
	.w6(32'hbb277f72),
	.w7(32'h3b69093f),
	.w8(32'hba837040),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f5e13),
	.w1(32'h3b841eea),
	.w2(32'hb8ca9b45),
	.w3(32'h3c668444),
	.w4(32'hba5da68f),
	.w5(32'h3acae549),
	.w6(32'h3a2a469f),
	.w7(32'hbacd53a4),
	.w8(32'hbaaaa471),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b509a39),
	.w1(32'hba0d5d64),
	.w2(32'h3a2cebd0),
	.w3(32'h3b8810c0),
	.w4(32'h38c6764c),
	.w5(32'h3be47637),
	.w6(32'hbb0a06c5),
	.w7(32'hbace168c),
	.w8(32'h3be5e27c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82486b),
	.w1(32'h3b89f5c4),
	.w2(32'hbca1ffd5),
	.w3(32'hbb039463),
	.w4(32'hbbd10fd1),
	.w5(32'hbb812ddf),
	.w6(32'h3b4d59b5),
	.w7(32'h3b63364e),
	.w8(32'h3b8df6d0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb904e18),
	.w1(32'h3ad82243),
	.w2(32'hbc0a93be),
	.w3(32'h3b14306d),
	.w4(32'hbc17b640),
	.w5(32'h3c06015e),
	.w6(32'h3aad479c),
	.w7(32'hbc5d08be),
	.w8(32'hba848273),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf3cd8c),
	.w1(32'hbb2daeea),
	.w2(32'hbab0c36f),
	.w3(32'hbba35d5d),
	.w4(32'h3b1e3d39),
	.w5(32'h39fc5354),
	.w6(32'hbb0024b0),
	.w7(32'h3ba4ce3f),
	.w8(32'hbbaa249a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba277a4),
	.w1(32'hbc44fabd),
	.w2(32'hbbb85f9a),
	.w3(32'h3b38bf59),
	.w4(32'hbbf54edb),
	.w5(32'hbb429c48),
	.w6(32'h3b535062),
	.w7(32'hba2f27ce),
	.w8(32'hbb240153),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb416355),
	.w1(32'hbb0582a3),
	.w2(32'h3b65d306),
	.w3(32'hbb8cc79c),
	.w4(32'h3c0dfb87),
	.w5(32'h3b8fc91a),
	.w6(32'h3958a75f),
	.w7(32'hbc78cd85),
	.w8(32'h3d05db7d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d9d02),
	.w1(32'h3b83f010),
	.w2(32'h3b1df489),
	.w3(32'h3b808e4c),
	.w4(32'hba281df5),
	.w5(32'h3c03e78f),
	.w6(32'h3ae9e813),
	.w7(32'h3b073764),
	.w8(32'hbbfee795),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b8ecd),
	.w1(32'h3c6c63a2),
	.w2(32'h3b503cea),
	.w3(32'hbc009f0b),
	.w4(32'h3a98f67d),
	.w5(32'h3beadef0),
	.w6(32'hbc076459),
	.w7(32'hbbb06ac9),
	.w8(32'hbc04bf6a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd46acd),
	.w1(32'hbb938325),
	.w2(32'hb91a3513),
	.w3(32'hb8cc19d8),
	.w4(32'h3c37ca8b),
	.w5(32'hba52f25d),
	.w6(32'hbab287e0),
	.w7(32'hbac26a49),
	.w8(32'hb9f3fe81),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bcf84),
	.w1(32'hbbef73ff),
	.w2(32'h3b84ebfb),
	.w3(32'hbb246597),
	.w4(32'h3aa4bb72),
	.w5(32'hbc2c6190),
	.w6(32'h3bc624f4),
	.w7(32'hbbaa8fd3),
	.w8(32'h3c846a47),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34311f),
	.w1(32'hbb0827fd),
	.w2(32'h3bb4c82f),
	.w3(32'hbc4e6cf1),
	.w4(32'h3c07f4c1),
	.w5(32'h3b0f92a3),
	.w6(32'hbb963451),
	.w7(32'h3b86af73),
	.w8(32'h3b3252e9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0de8e8),
	.w1(32'h3a95058d),
	.w2(32'h3bafaee2),
	.w3(32'h3b8d49ea),
	.w4(32'h3c3b66a4),
	.w5(32'hbb543626),
	.w6(32'h3b5158fb),
	.w7(32'hbb0cb091),
	.w8(32'h3acdb170),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9646662),
	.w1(32'hba144786),
	.w2(32'h3b8dee8a),
	.w3(32'h3b068bec),
	.w4(32'h3a56363b),
	.w5(32'h3c96912c),
	.w6(32'h3bbdb949),
	.w7(32'h3978ad88),
	.w8(32'hbc1894a1),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c684c1b),
	.w1(32'h3c0b08dd),
	.w2(32'h3b9f7d50),
	.w3(32'hbc1af745),
	.w4(32'h3c01c536),
	.w5(32'hbc6c07eb),
	.w6(32'h3d335bf9),
	.w7(32'hbb786492),
	.w8(32'h3b6e49dc),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c1da3),
	.w1(32'hba848996),
	.w2(32'h3b13da2a),
	.w3(32'hbbabda64),
	.w4(32'hbc3a023d),
	.w5(32'hbc2bc41b),
	.w6(32'hbb65c801),
	.w7(32'hbb3ae4e2),
	.w8(32'hbc465574),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4ee7c),
	.w1(32'h3b590460),
	.w2(32'h3c279552),
	.w3(32'h3c00d51e),
	.w4(32'h3a709635),
	.w5(32'h3c9f6792),
	.w6(32'h3c31517a),
	.w7(32'h3c819972),
	.w8(32'h389f7f86),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcfd87),
	.w1(32'h3ba380c1),
	.w2(32'hbaab459b),
	.w3(32'h3ba180f5),
	.w4(32'h3b8eeeee),
	.w5(32'h3c37d2af),
	.w6(32'hbca1d333),
	.w7(32'h3b3c14b9),
	.w8(32'hbaa23035),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b5f0b),
	.w1(32'hbc30b2c7),
	.w2(32'hbb86e232),
	.w3(32'hbad90753),
	.w4(32'hb8cae81f),
	.w5(32'hba817c8b),
	.w6(32'hbb9b44c1),
	.w7(32'hb94895c8),
	.w8(32'hbbb7c9ac),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba396747),
	.w1(32'hbb9345e2),
	.w2(32'hbb6e08cb),
	.w3(32'h38d32046),
	.w4(32'hbc37f150),
	.w5(32'h3a98ef19),
	.w6(32'hbb828aa3),
	.w7(32'h3c558d9b),
	.w8(32'hbc145286),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf96f8),
	.w1(32'hbc130728),
	.w2(32'hbc114299),
	.w3(32'h3bd6109a),
	.w4(32'hbad376d7),
	.w5(32'h3b9062c3),
	.w6(32'h3c22cb60),
	.w7(32'h3c177ff3),
	.w8(32'h3baa1a23),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8ea65),
	.w1(32'h3c835127),
	.w2(32'h3b90113f),
	.w3(32'hbb3da408),
	.w4(32'h3a96f02d),
	.w5(32'h3ba4b2d2),
	.w6(32'h3cff2dbf),
	.w7(32'h3ae19e05),
	.w8(32'h3b5009fc),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c8bc1),
	.w1(32'h3bb5fcbb),
	.w2(32'hbafec928),
	.w3(32'h3bc53687),
	.w4(32'hbb03202a),
	.w5(32'hbbafc8ef),
	.w6(32'hbb758dea),
	.w7(32'hbbce9a19),
	.w8(32'hbba417cb),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40d44e),
	.w1(32'h3b7af192),
	.w2(32'h3c31f87d),
	.w3(32'h3ba62127),
	.w4(32'h3c424ca9),
	.w5(32'h3c3a0c0f),
	.w6(32'h3b184f44),
	.w7(32'h3c3e661f),
	.w8(32'hba522199),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e54a9f),
	.w1(32'hbb9062cf),
	.w2(32'h3a47bb2b),
	.w3(32'h3a38887b),
	.w4(32'hbbe2dced),
	.w5(32'hbc92e30c),
	.w6(32'hba73b265),
	.w7(32'hbbc8ea6a),
	.w8(32'h3c893d11),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba09d56),
	.w1(32'hba308426),
	.w2(32'h3b5ffe52),
	.w3(32'h3c5bf888),
	.w4(32'h3bd3db01),
	.w5(32'hbb97f3ed),
	.w6(32'h3aa67577),
	.w7(32'h3bcac71c),
	.w8(32'hb92d2edc),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba473bda),
	.w1(32'h3975ba67),
	.w2(32'hbac5ee8b),
	.w3(32'h3c2bcb48),
	.w4(32'h3a3fd930),
	.w5(32'hbba22f50),
	.w6(32'h3c2f56db),
	.w7(32'hb9820d98),
	.w8(32'hbc302926),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cff6519),
	.w1(32'hba3c8b74),
	.w2(32'hbc08c843),
	.w3(32'h3b08b1ad),
	.w4(32'h3ca8f720),
	.w5(32'hbb9e8076),
	.w6(32'hbba70a7c),
	.w7(32'h3a8f3195),
	.w8(32'hba6fe1b3),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18381d),
	.w1(32'hbc359c48),
	.w2(32'hb9a6a8d7),
	.w3(32'hbc010bbc),
	.w4(32'hbc4674c0),
	.w5(32'h3cee2a99),
	.w6(32'h3d0deb83),
	.w7(32'h3c31d4a5),
	.w8(32'h3bec1691),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82c47f),
	.w1(32'hbacc8bcb),
	.w2(32'h3b98afbf),
	.w3(32'hb93a8dd8),
	.w4(32'hbb190278),
	.w5(32'h3a33d956),
	.w6(32'h3c16e154),
	.w7(32'hbb5b16b2),
	.w8(32'hb9a38b9b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98a47d),
	.w1(32'hbabebea9),
	.w2(32'hbbd6e7db),
	.w3(32'hbb990497),
	.w4(32'hbb4c2956),
	.w5(32'hbbd638a1),
	.w6(32'h3c8fd959),
	.w7(32'h3b8932b4),
	.w8(32'hbb36316b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63e6c1),
	.w1(32'hbb66d1d8),
	.w2(32'hbba78118),
	.w3(32'h3bd266ee),
	.w4(32'h3b8e227a),
	.w5(32'hbbcbc1b6),
	.w6(32'hbbff4294),
	.w7(32'hbb10a3cf),
	.w8(32'h3c477789),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bdfef),
	.w1(32'h391cb954),
	.w2(32'hbb841890),
	.w3(32'h3b2051ed),
	.w4(32'h3cdaac82),
	.w5(32'h3aa7db6e),
	.w6(32'h3957f585),
	.w7(32'hbc2fc677),
	.w8(32'h3bbc3749),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac08244),
	.w1(32'h3a845298),
	.w2(32'hbbfd814c),
	.w3(32'h3b90265c),
	.w4(32'h3c1cd0ed),
	.w5(32'hb936f512),
	.w6(32'hbbb61506),
	.w7(32'h3bfc3202),
	.w8(32'h3c5959ac),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12c65e),
	.w1(32'hbb7ecde6),
	.w2(32'hba7d7d1d),
	.w3(32'hba5959d6),
	.w4(32'hba5611ca),
	.w5(32'h3ada2168),
	.w6(32'hbb84e68e),
	.w7(32'hbb23d31f),
	.w8(32'hbaa71bae),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eb0fb5),
	.w1(32'hb9eb752a),
	.w2(32'h3baa7875),
	.w3(32'h3a4e875f),
	.w4(32'h3bbd69f6),
	.w5(32'hbc10b496),
	.w6(32'hbbac1cd6),
	.w7(32'h3be5b40f),
	.w8(32'h3c1a87b9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule