module layer_10_featuremap_414(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e2425),
	.w1(32'hb9613dbe),
	.w2(32'hbc4caa8e),
	.w3(32'hbbc4470d),
	.w4(32'h3a7c5f49),
	.w5(32'hbab94c6f),
	.w6(32'h3c2ed1bc),
	.w7(32'h3bbe3c5a),
	.w8(32'h3bf6b065),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12adaa),
	.w1(32'h3c01a637),
	.w2(32'h3c0e74dc),
	.w3(32'hbbb143ea),
	.w4(32'hbc4873d8),
	.w5(32'hbc15aafa),
	.w6(32'h3b31113c),
	.w7(32'hbc34f010),
	.w8(32'hbc89428a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09b641),
	.w1(32'h3ae064e0),
	.w2(32'hbb11ad68),
	.w3(32'hbc8cfe72),
	.w4(32'h3b0946d0),
	.w5(32'h3b9a9ce3),
	.w6(32'hbca134bb),
	.w7(32'hbc46e9b2),
	.w8(32'hbc42a847),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be257af),
	.w1(32'h3b1e4fe8),
	.w2(32'h3c1941a4),
	.w3(32'h3b076df0),
	.w4(32'hbaedd364),
	.w5(32'h3c0adf4e),
	.w6(32'hbc35f770),
	.w7(32'hbbee1c44),
	.w8(32'hbc26a2fe),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89c6bb),
	.w1(32'h3b837eac),
	.w2(32'hbb277fc0),
	.w3(32'h3c2b8c34),
	.w4(32'hbbaaf9de),
	.w5(32'hbb9e5766),
	.w6(32'hbc651577),
	.w7(32'hbbb08ae0),
	.w8(32'hbc621aed),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc010aab),
	.w1(32'h3ac1ed5b),
	.w2(32'h3c6d262f),
	.w3(32'hbc60d5cc),
	.w4(32'hbab37a01),
	.w5(32'h3bb585ab),
	.w6(32'hbc401246),
	.w7(32'h3c153109),
	.w8(32'h3a81dbc6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959b513),
	.w1(32'h3c45eea0),
	.w2(32'h3b97f953),
	.w3(32'hbb5db8b0),
	.w4(32'h3b9ca38d),
	.w5(32'h3ca200c3),
	.w6(32'hbbbc8996),
	.w7(32'h3b8b0ab8),
	.w8(32'h3bb1c2a1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7164ef),
	.w1(32'h3bdbd58d),
	.w2(32'hbbf04893),
	.w3(32'h3af8b97e),
	.w4(32'h3c5ad5bc),
	.w5(32'h3bb07f42),
	.w6(32'hbbed8b57),
	.w7(32'hbc31d9de),
	.w8(32'hbabdb83a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e6121),
	.w1(32'h3c5db2fc),
	.w2(32'h3b0239e7),
	.w3(32'hbb006cfd),
	.w4(32'hba77a875),
	.w5(32'hbc2e82cc),
	.w6(32'hbbae1af8),
	.w7(32'h3b20cce4),
	.w8(32'hbc38b97d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c145d),
	.w1(32'h3c30f0f8),
	.w2(32'h3c1de3ce),
	.w3(32'h3b856251),
	.w4(32'hbc325943),
	.w5(32'hbbc55518),
	.w6(32'hbbfc8069),
	.w7(32'hb9eeb172),
	.w8(32'hbb2fbe83),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25e942),
	.w1(32'h3c2b7800),
	.w2(32'h3bcd7195),
	.w3(32'hbbe02b14),
	.w4(32'hbb0bf71c),
	.w5(32'h3a7fefd1),
	.w6(32'hbbf78e19),
	.w7(32'h3bbb0c50),
	.w8(32'hbc0a49d3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba54663),
	.w1(32'hbb0be61f),
	.w2(32'hbc936031),
	.w3(32'hbc307a37),
	.w4(32'h3c1569fb),
	.w5(32'h3c1ddd4a),
	.w6(32'hbc5ddb8b),
	.w7(32'h3c2803ba),
	.w8(32'h3c8448ff),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62c6fb),
	.w1(32'h3c49a9e1),
	.w2(32'h3cb1374b),
	.w3(32'h3ba3c0d2),
	.w4(32'hbb27084a),
	.w5(32'hbc2b6a2c),
	.w6(32'h3c2e540c),
	.w7(32'hbc5832cd),
	.w8(32'hbca86553),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e6587),
	.w1(32'h3be8697c),
	.w2(32'hbc319e74),
	.w3(32'h3b5039ff),
	.w4(32'h3c4220a1),
	.w5(32'h3c4d13ff),
	.w6(32'hbbd43be4),
	.w7(32'hbc34e02e),
	.w8(32'hbc1aaf5f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8bb2a),
	.w1(32'h3c4b6c41),
	.w2(32'h3cd0f5ab),
	.w3(32'h3b2445ab),
	.w4(32'h3b42a7b2),
	.w5(32'hb949685c),
	.w6(32'hbbaf16f5),
	.w7(32'hbc472562),
	.w8(32'hbcb12c3a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbf8a9),
	.w1(32'h3c0edb9b),
	.w2(32'h3c1557eb),
	.w3(32'hbb7b7f5f),
	.w4(32'h3c2be86b),
	.w5(32'hb9df5f27),
	.w6(32'hbc21ae3f),
	.w7(32'h3b9f1a33),
	.w8(32'h3b8c45be),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc28d62),
	.w1(32'h3c0aeba5),
	.w2(32'h3b905e63),
	.w3(32'h3b95c26e),
	.w4(32'h3c3dd199),
	.w5(32'h3c74a15f),
	.w6(32'h3bf392db),
	.w7(32'h3c2da43f),
	.w8(32'h3b57c393),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62f651),
	.w1(32'hbbda6f5b),
	.w2(32'hbc78a3aa),
	.w3(32'h3c014ed8),
	.w4(32'h3ba18621),
	.w5(32'h3bd8e273),
	.w6(32'hbaf14366),
	.w7(32'h3a854810),
	.w8(32'hbb8c7306),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88b1ab),
	.w1(32'h3c3a0fd5),
	.w2(32'h3c3065a1),
	.w3(32'h3c49a3e6),
	.w4(32'hbbce807b),
	.w5(32'hbc004b39),
	.w6(32'h395a7176),
	.w7(32'hbb02b085),
	.w8(32'hbc3453d6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0dd586),
	.w1(32'h3b9077e2),
	.w2(32'h3c89dde0),
	.w3(32'hbc0af6bb),
	.w4(32'h3b003d56),
	.w5(32'h3aae54dc),
	.w6(32'hbc5d3302),
	.w7(32'h3c35e6d8),
	.w8(32'hbc3982b2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f4b61),
	.w1(32'hbc0ff0b1),
	.w2(32'hbc2dfd18),
	.w3(32'hbbd6a6f8),
	.w4(32'h3b82b016),
	.w5(32'h3ba24950),
	.w6(32'hbcad6ab7),
	.w7(32'h3c2579b8),
	.w8(32'h3bcdcadf),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeda122),
	.w1(32'h3a2be3c6),
	.w2(32'h3cad153f),
	.w3(32'h3b17be32),
	.w4(32'hbb6b3b18),
	.w5(32'hbbd8bc6d),
	.w6(32'h3ba3edb8),
	.w7(32'h3ae69c30),
	.w8(32'hbcb8d734),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70a72c),
	.w1(32'hbc391c71),
	.w2(32'h3ce51480),
	.w3(32'hbc1b5c47),
	.w4(32'hbc956536),
	.w5(32'hbc37b87e),
	.w6(32'hbbc37070),
	.w7(32'hbc433f01),
	.w8(32'hbbc83110),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d02a1),
	.w1(32'h3ba289ff),
	.w2(32'h3c9d9589),
	.w3(32'hbbd8b796),
	.w4(32'hbcce82a4),
	.w5(32'hbc8590e4),
	.w6(32'hbb1f54b8),
	.w7(32'h3ac93f74),
	.w8(32'h3c380267),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacedf3),
	.w1(32'hba726c4b),
	.w2(32'h3d08c3bb),
	.w3(32'hbcdbb6e6),
	.w4(32'hbbc9fbfa),
	.w5(32'hbc3a5523),
	.w6(32'h3c283a00),
	.w7(32'hbc8784ec),
	.w8(32'hbd02a1f6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb04bef),
	.w1(32'hb99961c1),
	.w2(32'h3967ac90),
	.w3(32'hbc974fa4),
	.w4(32'h3ada289b),
	.w5(32'hbc3b9ae7),
	.w6(32'hbc6b9d89),
	.w7(32'h3bd3cb6e),
	.w8(32'h3b2907a0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04d356),
	.w1(32'hbbc2c1ba),
	.w2(32'hbb681962),
	.w3(32'hbaee4428),
	.w4(32'hbb0e4eb8),
	.w5(32'h3c7d5ccd),
	.w6(32'h3bb95620),
	.w7(32'hbc1dcb48),
	.w8(32'hbc264eff),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18a007),
	.w1(32'h3b4401fa),
	.w2(32'h3c55a728),
	.w3(32'hb9e1fb68),
	.w4(32'h3b2c1ded),
	.w5(32'hbc2a5b34),
	.w6(32'hbc67294d),
	.w7(32'hbab41143),
	.w8(32'hbc88b537),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c398512),
	.w1(32'hbc056f88),
	.w2(32'h3c504488),
	.w3(32'hbc3dcc08),
	.w4(32'hbc62f61b),
	.w5(32'h3b61e18d),
	.w6(32'hbc88c361),
	.w7(32'hbc2282f9),
	.w8(32'hb8b37ef9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a6112),
	.w1(32'hbc801b76),
	.w2(32'hbc9b8bf1),
	.w3(32'h3b94df8f),
	.w4(32'h3bbd39b6),
	.w5(32'h3c3a69fb),
	.w6(32'h3ca67c16),
	.w7(32'h3c7afd88),
	.w8(32'h3ce7d989),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba067d8),
	.w1(32'h3b1c8053),
	.w2(32'hbab26e6a),
	.w3(32'h3b96edde),
	.w4(32'hbb0337b9),
	.w5(32'hbab79473),
	.w6(32'h3c27c5f9),
	.w7(32'h3baca550),
	.w8(32'h3bdc8a4a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48d38d),
	.w1(32'h3ba51058),
	.w2(32'hbb8c1e96),
	.w3(32'h3b12be34),
	.w4(32'h3a2d3882),
	.w5(32'hbb4dadad),
	.w6(32'h3ba2c9c2),
	.w7(32'hbb66fdc0),
	.w8(32'hbbc02000),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac78914),
	.w1(32'hba15746b),
	.w2(32'hbbfd8475),
	.w3(32'hbbfa82a4),
	.w4(32'h3b998604),
	.w5(32'h3cb11476),
	.w6(32'hbc16ac38),
	.w7(32'h3ab4af7b),
	.w8(32'hba5733f9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa87a95),
	.w1(32'hbbee3bcf),
	.w2(32'h3bab46c6),
	.w3(32'h3b9ba9c5),
	.w4(32'hbbbc763d),
	.w5(32'hbc42e5b7),
	.w6(32'h3b30083d),
	.w7(32'hb978cd12),
	.w8(32'h3b33819f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd65a8e),
	.w1(32'h3b79eb50),
	.w2(32'hbc296d27),
	.w3(32'hbbf6f041),
	.w4(32'h3c3c4dce),
	.w5(32'hbb386468),
	.w6(32'h3a1206a9),
	.w7(32'h3b51b091),
	.w8(32'h3c116316),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a928b2a),
	.w1(32'hbc3ab139),
	.w2(32'h3b938946),
	.w3(32'h3b17604f),
	.w4(32'hbac885e2),
	.w5(32'h3bb109a4),
	.w6(32'hbb511af9),
	.w7(32'h3c088813),
	.w8(32'h3c5170cf),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc344cc7),
	.w1(32'h3b192f59),
	.w2(32'h3c5a74c5),
	.w3(32'hbb6b245d),
	.w4(32'hbbca2ccb),
	.w5(32'h3ce1bd95),
	.w6(32'h3aaa6929),
	.w7(32'hb98d3443),
	.w8(32'h3b73d844),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c9da9),
	.w1(32'h3b7c49d0),
	.w2(32'h3bb374ba),
	.w3(32'hb931e976),
	.w4(32'h3a97d4a5),
	.w5(32'h3ae96dfd),
	.w6(32'h3ad3aa6c),
	.w7(32'h3be1b713),
	.w8(32'hbb0cb02a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4d4d4),
	.w1(32'h3a906636),
	.w2(32'h3b332401),
	.w3(32'hbab638c1),
	.w4(32'h3bab486e),
	.w5(32'hbc64a730),
	.w6(32'h3c236016),
	.w7(32'h3c3bfa9f),
	.w8(32'hbb771fc7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c091561),
	.w1(32'h3a92384b),
	.w2(32'h3be5a110),
	.w3(32'hbb5e354b),
	.w4(32'hbb08ffba),
	.w5(32'hbc05a70d),
	.w6(32'hbaa481ac),
	.w7(32'hbbf6cb98),
	.w8(32'hbbdc3158),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb45ce),
	.w1(32'h3b17c6d0),
	.w2(32'h3c412548),
	.w3(32'h3b8a53a6),
	.w4(32'h3bc50ae7),
	.w5(32'h3bea4802),
	.w6(32'hbb8603ff),
	.w7(32'h3adc39ae),
	.w8(32'hbbd5d6e2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdeb8c8),
	.w1(32'h3a92470d),
	.w2(32'h3c14beb9),
	.w3(32'h3bb450fc),
	.w4(32'hbbb8e170),
	.w5(32'hbb1a562b),
	.w6(32'hbc17cd37),
	.w7(32'hbbbad3a0),
	.w8(32'hbc5e2401),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b712077),
	.w1(32'h3ae0f079),
	.w2(32'h3b9ee8c4),
	.w3(32'hbb2a37f2),
	.w4(32'hbb968aa8),
	.w5(32'hbb14b976),
	.w6(32'hbb81d244),
	.w7(32'hbc03fc40),
	.w8(32'hbb917185),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8eca6),
	.w1(32'h3c47d958),
	.w2(32'hbb5ae313),
	.w3(32'h3b92930b),
	.w4(32'h3c7655b7),
	.w5(32'h3921f3ce),
	.w6(32'hbc151bba),
	.w7(32'h3bb2a61f),
	.w8(32'h3b1fd795),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb131978),
	.w1(32'h3bbb5292),
	.w2(32'hba8d994c),
	.w3(32'h3b8ab7be),
	.w4(32'hbac636ef),
	.w5(32'h3ba237f0),
	.w6(32'hbb0c7ece),
	.w7(32'h3b0cb01d),
	.w8(32'hbb8b235d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacca41),
	.w1(32'h3bff6d82),
	.w2(32'h3c51feaf),
	.w3(32'h3ba9e972),
	.w4(32'h3b8a0849),
	.w5(32'h3c1b9e63),
	.w6(32'h3b6dc671),
	.w7(32'hbb05ea46),
	.w8(32'h39bd6aac),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ffa24),
	.w1(32'hbb40cc93),
	.w2(32'h3a87dfca),
	.w3(32'h3b8d49a7),
	.w4(32'h394336d7),
	.w5(32'hbb575460),
	.w6(32'hba533c5e),
	.w7(32'hbc426008),
	.w8(32'hbca08e5d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab924d),
	.w1(32'h3c711a9c),
	.w2(32'h3c1b5ff0),
	.w3(32'h39a08c4c),
	.w4(32'hbb605bca),
	.w5(32'hbc2001f8),
	.w6(32'hbc3a8f9b),
	.w7(32'hbc3c975e),
	.w8(32'hbcbaae83),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7a323),
	.w1(32'hbb0ed053),
	.w2(32'hbc7907ce),
	.w3(32'hbaa3f70c),
	.w4(32'hbb9be7a7),
	.w5(32'h3c5bf70a),
	.w6(32'hbc4e3246),
	.w7(32'h3937c86f),
	.w8(32'h3c8fc790),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc156a14),
	.w1(32'hbb4b13ed),
	.w2(32'hbc60cd01),
	.w3(32'hbaeeb045),
	.w4(32'h3c113723),
	.w5(32'h3c3c6d6a),
	.w6(32'h3bb5972d),
	.w7(32'h3bf4cbb5),
	.w8(32'h3c9bb3bf),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00eb96),
	.w1(32'h3b67836c),
	.w2(32'h3c3be08d),
	.w3(32'h397082fd),
	.w4(32'hbc3fcd5c),
	.w5(32'hba5fb733),
	.w6(32'h3b6c4d0e),
	.w7(32'hbb838a05),
	.w8(32'hbc995a72),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ce629),
	.w1(32'h3c1541e0),
	.w2(32'h3cbd5cd3),
	.w3(32'hbbc22e16),
	.w4(32'hbc06ffbe),
	.w5(32'hbc214ccd),
	.w6(32'hbc19b782),
	.w7(32'h3a954dd6),
	.w8(32'hbbe1b59c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23a722),
	.w1(32'hbcac0fef),
	.w2(32'hbc93a998),
	.w3(32'hbc820d5c),
	.w4(32'h3b7d764c),
	.w5(32'h3c679a9e),
	.w6(32'hbc8a7d66),
	.w7(32'h3ba03478),
	.w8(32'h3c9932f1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55d809),
	.w1(32'h3b088edc),
	.w2(32'hbc79c57f),
	.w3(32'h3c48dd2c),
	.w4(32'h3c4da178),
	.w5(32'hbc321b2e),
	.w6(32'h3c57bb46),
	.w7(32'h3be2a199),
	.w8(32'h3c6ed286),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fa6cb),
	.w1(32'h3ca14106),
	.w2(32'h3c99eba2),
	.w3(32'h3b5485e6),
	.w4(32'hba99c0eb),
	.w5(32'hbc082d21),
	.w6(32'h3ba16a78),
	.w7(32'hbc3db400),
	.w8(32'hbc8eb822),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a178223),
	.w1(32'h3c246ee8),
	.w2(32'h3c0298c1),
	.w3(32'hbb037bf4),
	.w4(32'hba04476e),
	.w5(32'hbbc0f64b),
	.w6(32'hbb49c4a5),
	.w7(32'hbb07b970),
	.w8(32'hbb9e1a82),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2de504),
	.w1(32'hbb617c35),
	.w2(32'h3b00cabd),
	.w3(32'hbc36c42d),
	.w4(32'h38422e0d),
	.w5(32'hbb128dca),
	.w6(32'hbbf18bc6),
	.w7(32'hbbc52879),
	.w8(32'hbc49dfa6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac95528),
	.w1(32'h3c9ab491),
	.w2(32'h3cbe836b),
	.w3(32'hbbf1c56f),
	.w4(32'h39e8b274),
	.w5(32'hbb03ea13),
	.w6(32'hbc4cd4ec),
	.w7(32'hbc3b22bb),
	.w8(32'hbcaef1d1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeae5d5),
	.w1(32'h3b54587b),
	.w2(32'h3cc28fe5),
	.w3(32'h3b5ce7d1),
	.w4(32'hbb13b067),
	.w5(32'h3acc8610),
	.w6(32'hbb6446a5),
	.w7(32'hbb676808),
	.w8(32'hbc21b951),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d72d5),
	.w1(32'h3c97a062),
	.w2(32'h3cfeae59),
	.w3(32'h390e9fda),
	.w4(32'hbbfb8b75),
	.w5(32'hbc50c39f),
	.w6(32'hbb828463),
	.w7(32'hbc78ac65),
	.w8(32'hbcd79c9a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99edb5d),
	.w1(32'h3a427a43),
	.w2(32'h3c5a5022),
	.w3(32'hbbd561b4),
	.w4(32'h37a72641),
	.w5(32'hbc403fb5),
	.w6(32'hbcbec3d4),
	.w7(32'hbb64f943),
	.w8(32'hbc82e1b6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c09b6),
	.w1(32'h3a8185dc),
	.w2(32'hbb8cebd3),
	.w3(32'hbb681144),
	.w4(32'h3a65f7ee),
	.w5(32'hbc0c87f1),
	.w6(32'hbb8d4f4b),
	.w7(32'h3b4e7f33),
	.w8(32'hbc45c18b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e977d),
	.w1(32'h3c7ac6bb),
	.w2(32'h3ce6719b),
	.w3(32'hbb9a4518),
	.w4(32'hbbda6eac),
	.w5(32'hbbfd07b7),
	.w6(32'hbc28adad),
	.w7(32'hbc76cb04),
	.w8(32'hbc9ac0ad),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc77bcb),
	.w1(32'hba36343c),
	.w2(32'hbbb469fe),
	.w3(32'hbbd25510),
	.w4(32'hbb334aac),
	.w5(32'hbc236431),
	.w6(32'hbc63aa0b),
	.w7(32'h3b96df8a),
	.w8(32'h3b3500d2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a13f7),
	.w1(32'hbc732e54),
	.w2(32'hbd086336),
	.w3(32'hbba8a1e6),
	.w4(32'hba0d2ab2),
	.w5(32'h3b1ce335),
	.w6(32'hbb02a4a2),
	.w7(32'h3ca120dd),
	.w8(32'h3cfbc3b2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc979c35),
	.w1(32'hba6666b9),
	.w2(32'hbcb3949f),
	.w3(32'h3b12538c),
	.w4(32'h3b19d2b6),
	.w5(32'h3b27fd4f),
	.w6(32'h3c8cfd6a),
	.w7(32'h3b247979),
	.w8(32'h3c9471b6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f5bbe),
	.w1(32'h3c3148df),
	.w2(32'hbc1067d7),
	.w3(32'h3c8a4784),
	.w4(32'h3a17efd2),
	.w5(32'hbca376bc),
	.w6(32'h3c65dd48),
	.w7(32'hb9ee7be5),
	.w8(32'hbc2353cf),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab37aec),
	.w1(32'h3c90ea12),
	.w2(32'h3cfdfa2b),
	.w3(32'hbc03481d),
	.w4(32'hbc04a457),
	.w5(32'hbacda902),
	.w6(32'hbc47f695),
	.w7(32'hbcbd070a),
	.w8(32'hbcc104ab),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccf0624),
	.w1(32'h3c96d75e),
	.w2(32'h3caa0d87),
	.w3(32'hbc5fcea2),
	.w4(32'hbc7a9580),
	.w5(32'hbbf040b3),
	.w6(32'hbccc9865),
	.w7(32'hbc859792),
	.w8(32'hbca47f50),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c021ee6),
	.w1(32'hbc031474),
	.w2(32'h3c22aaf2),
	.w3(32'hbbf26a7f),
	.w4(32'hbc53a57b),
	.w5(32'h3c3b927d),
	.w6(32'h3b3ed9d5),
	.w7(32'hbb3f2735),
	.w8(32'h3c3bf219),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba71b51),
	.w1(32'h3cadbf75),
	.w2(32'h3ba55523),
	.w3(32'h3c4550a4),
	.w4(32'h3c37794c),
	.w5(32'hbc08d8c6),
	.w6(32'hbb9d77a6),
	.w7(32'hbb98aa88),
	.w8(32'hbb8726b9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72002f),
	.w1(32'h39f692c3),
	.w2(32'h3c5627ee),
	.w3(32'h3aff9150),
	.w4(32'h3afd9497),
	.w5(32'h3c860c0c),
	.w6(32'h3b1ec379),
	.w7(32'h3c45d008),
	.w8(32'hbac5c89d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb4b86),
	.w1(32'h3b208dcf),
	.w2(32'hbacd5fbb),
	.w3(32'h3ae169c9),
	.w4(32'h3a80a2ef),
	.w5(32'hbb0f3b9b),
	.w6(32'hbc4402b3),
	.w7(32'h3b6fe686),
	.w8(32'h3c535d99),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf574d),
	.w1(32'hbb1209ca),
	.w2(32'h3b365cf2),
	.w3(32'h3c2f5862),
	.w4(32'h3b42f8f0),
	.w5(32'h3ba51299),
	.w6(32'h3b9d7c35),
	.w7(32'h3b2d101d),
	.w8(32'h3b125013),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa86084),
	.w1(32'hbb53a70c),
	.w2(32'hbb2590c3),
	.w3(32'hbba4533b),
	.w4(32'hbc8eedac),
	.w5(32'h3c0566f6),
	.w6(32'hba256621),
	.w7(32'hbbca418d),
	.w8(32'hbb142bca),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83097b),
	.w1(32'h3a8c33b6),
	.w2(32'h3af0d1d2),
	.w3(32'hbb11848a),
	.w4(32'h3b24b840),
	.w5(32'h3c04eecf),
	.w6(32'hbc16007e),
	.w7(32'h398bd6d3),
	.w8(32'h3b0e185f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e72e3),
	.w1(32'h3c9b7bd9),
	.w2(32'h3cdcda5e),
	.w3(32'h3aa427d9),
	.w4(32'h3c5dc97d),
	.w5(32'h3c9d0397),
	.w6(32'hbb159724),
	.w7(32'h3c5625c6),
	.w8(32'h3d06208c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf13183),
	.w1(32'hbc2fff1f),
	.w2(32'hbb558fde),
	.w3(32'h3cd22552),
	.w4(32'h398af125),
	.w5(32'hbc291b14),
	.w6(32'h3d084464),
	.w7(32'h3c515ee8),
	.w8(32'hbb2ea733),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ee094),
	.w1(32'h3b5a9a82),
	.w2(32'h3a9d1ab3),
	.w3(32'h3c246d5c),
	.w4(32'h3af18ac3),
	.w5(32'hbafeb275),
	.w6(32'hbbff7194),
	.w7(32'h3bced92f),
	.w8(32'hbb060466),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc2a61),
	.w1(32'h3bbd29f0),
	.w2(32'hba60e8f8),
	.w3(32'h3c851006),
	.w4(32'h3c002dca),
	.w5(32'h3cbe1210),
	.w6(32'h3c3fa449),
	.w7(32'hbc1c87ad),
	.w8(32'h3c88b2e1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89db4b),
	.w1(32'h3b229ce4),
	.w2(32'h3b606f9f),
	.w3(32'h3bffa15d),
	.w4(32'hbc1abd88),
	.w5(32'hbbf71577),
	.w6(32'h3ca767de),
	.w7(32'h3b838513),
	.w8(32'h3aef4e1b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a91f0),
	.w1(32'h3b6339bb),
	.w2(32'hbb904dce),
	.w3(32'h3ba3935f),
	.w4(32'hba54418e),
	.w5(32'hbbed43ff),
	.w6(32'h3a8c3440),
	.w7(32'hbb2f650c),
	.w8(32'hbb9dea5d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6b617),
	.w1(32'hba0b5792),
	.w2(32'hbc08c8f7),
	.w3(32'hbaa29800),
	.w4(32'h39d2835a),
	.w5(32'hbc15703d),
	.w6(32'hbb16554b),
	.w7(32'h3b4d1d74),
	.w8(32'hbb671ff1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcad4e3),
	.w1(32'h3c313b8a),
	.w2(32'h3b7cc898),
	.w3(32'hbbeb3c15),
	.w4(32'h3c026666),
	.w5(32'hbc1276b7),
	.w6(32'hbba1f6aa),
	.w7(32'h3a818298),
	.w8(32'h3c3e2e38),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384be22a),
	.w1(32'h3a8e476c),
	.w2(32'h39d1136a),
	.w3(32'h3c9462bd),
	.w4(32'h3b493423),
	.w5(32'hbbd97570),
	.w6(32'h3bf52622),
	.w7(32'h3bea7bc2),
	.w8(32'hbacd0ddb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaeaf23),
	.w1(32'h3a157a63),
	.w2(32'hbb064ce3),
	.w3(32'h3aa6a285),
	.w4(32'h3b929ace),
	.w5(32'hbba38b7d),
	.w6(32'hbad03551),
	.w7(32'h3b831d55),
	.w8(32'hbc6128e2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86c5ec),
	.w1(32'hbae93ffc),
	.w2(32'h3bb4d34b),
	.w3(32'hbc3cbf74),
	.w4(32'hbb81cd12),
	.w5(32'h3c36a225),
	.w6(32'hbc12c118),
	.w7(32'hbc0353a4),
	.w8(32'h3be35cbc),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9cab2),
	.w1(32'hba8bd347),
	.w2(32'h3a750d5c),
	.w3(32'h3b0b808f),
	.w4(32'hbb7f2a1a),
	.w5(32'h3c1ce6bc),
	.w6(32'h3b863511),
	.w7(32'hbbfee491),
	.w8(32'hba04d236),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc043ceb),
	.w1(32'hbba1a4b9),
	.w2(32'h3c1866df),
	.w3(32'hbc36f0cf),
	.w4(32'hb89e24d1),
	.w5(32'hbc6530eb),
	.w6(32'hbb45f824),
	.w7(32'hbbf837c8),
	.w8(32'h3bb4e3db),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb3478),
	.w1(32'h3bab3189),
	.w2(32'hbb11b446),
	.w3(32'h3b6da691),
	.w4(32'h3b820b75),
	.w5(32'h3a033080),
	.w6(32'h3b46d118),
	.w7(32'hbb62f7ca),
	.w8(32'h3a6d49ea),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62b934),
	.w1(32'h3bb4dbea),
	.w2(32'h3b737fba),
	.w3(32'hbba42207),
	.w4(32'h3bdae2bb),
	.w5(32'hba7fc70f),
	.w6(32'hb91c3cbd),
	.w7(32'h3bdf5e77),
	.w8(32'h3b8454fa),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13eef2),
	.w1(32'h3c3d6684),
	.w2(32'hbab56b6b),
	.w3(32'hbb05b471),
	.w4(32'hbc817cd0),
	.w5(32'hbbf818dd),
	.w6(32'h3c222a5e),
	.w7(32'hb9a9a936),
	.w8(32'hbb6e65d2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a020a37),
	.w1(32'h3c1e0a39),
	.w2(32'h3ac8d9c8),
	.w3(32'hbbf27417),
	.w4(32'hbb6ee72c),
	.w5(32'h3bc89590),
	.w6(32'hba083574),
	.w7(32'h3baaa667),
	.w8(32'h3a777df5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40bb2d),
	.w1(32'h3c49862e),
	.w2(32'hba9baf4b),
	.w3(32'hbb4f558a),
	.w4(32'h3b8e7d89),
	.w5(32'hbaab99d5),
	.w6(32'hbbe68f82),
	.w7(32'h3bf81eff),
	.w8(32'h3be14a1c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38602c),
	.w1(32'h3b048d77),
	.w2(32'hbb8c0caa),
	.w3(32'hb63b99d4),
	.w4(32'h3c61a932),
	.w5(32'hbb7e32b9),
	.w6(32'h3b883605),
	.w7(32'hbc43d9d4),
	.w8(32'h3b1784aa),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba964738),
	.w1(32'hba3e1f13),
	.w2(32'h3bf74410),
	.w3(32'h3b39832a),
	.w4(32'h3afc8ea1),
	.w5(32'h3c8813ec),
	.w6(32'h3c57ed29),
	.w7(32'h3c4763c5),
	.w8(32'h3b20bdb1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77c06f),
	.w1(32'h3b866d91),
	.w2(32'h3a3d1d7b),
	.w3(32'h39a0a199),
	.w4(32'hb997b1ed),
	.w5(32'hbbef0dfc),
	.w6(32'hbbeef68e),
	.w7(32'hbbbb6b8b),
	.w8(32'hbc5a89f0),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81423c),
	.w1(32'h3bc4b2b6),
	.w2(32'h3b6ea3a5),
	.w3(32'hbc199506),
	.w4(32'h3c7ada10),
	.w5(32'hbb32aa12),
	.w6(32'hbc0b8436),
	.w7(32'h3ab957ae),
	.w8(32'h3b4930c2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63b266),
	.w1(32'hbb4f9533),
	.w2(32'hba84ada8),
	.w3(32'hbb9a3d58),
	.w4(32'h3b56f084),
	.w5(32'hbc1a04fd),
	.w6(32'hbab8c9f7),
	.w7(32'h39a572f2),
	.w8(32'h3b18ddd4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5012d),
	.w1(32'h3b6dbe43),
	.w2(32'h3ca9a80b),
	.w3(32'h3aa1c705),
	.w4(32'hbc831158),
	.w5(32'h3ae34ba3),
	.w6(32'h3cac0506),
	.w7(32'hbc4d95f8),
	.w8(32'hbc1676e0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d582b),
	.w1(32'hbc086a14),
	.w2(32'h3b3001b7),
	.w3(32'hbc07c58b),
	.w4(32'hbb570c29),
	.w5(32'hbac2e0eb),
	.w6(32'h3c230623),
	.w7(32'hbb9f4141),
	.w8(32'h3b9615d4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba85f2a),
	.w1(32'hbbe7ced8),
	.w2(32'hbbda62a9),
	.w3(32'hbbaa13a7),
	.w4(32'hbc03fed8),
	.w5(32'h3a80015d),
	.w6(32'h3c1092c1),
	.w7(32'h3b5dde61),
	.w8(32'hba41e65d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c6d79),
	.w1(32'hbb577bb5),
	.w2(32'h3bac9611),
	.w3(32'hbc75c64f),
	.w4(32'hbc14cfaa),
	.w5(32'h3c711f38),
	.w6(32'hbc859403),
	.w7(32'h3c203c00),
	.w8(32'h3a0ecc28),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90b99f),
	.w1(32'hbb3ad296),
	.w2(32'hba46a0b4),
	.w3(32'h3a8ee5e6),
	.w4(32'hba59b029),
	.w5(32'hbb783fd3),
	.w6(32'hbb8cdc77),
	.w7(32'h3bb46be9),
	.w8(32'hba906a7f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb127d9),
	.w1(32'h3c3fb3a3),
	.w2(32'h3c0f83b8),
	.w3(32'h3a24a724),
	.w4(32'h3adaf60c),
	.w5(32'hbc15cf39),
	.w6(32'hbb13c1fc),
	.w7(32'hbc248622),
	.w8(32'h3c48aa72),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e27472),
	.w1(32'h3c06c921),
	.w2(32'h3b859036),
	.w3(32'h3ae3531b),
	.w4(32'h3bf441db),
	.w5(32'h3b41a250),
	.w6(32'h3bf4e4f1),
	.w7(32'h3c2af531),
	.w8(32'h3c46ac52),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae911c2),
	.w1(32'h3a29cdf4),
	.w2(32'hbba18d2e),
	.w3(32'h3a37c308),
	.w4(32'hb9b2bc63),
	.w5(32'hbbacd400),
	.w6(32'hb9103a85),
	.w7(32'hbb4202c7),
	.w8(32'hbb4d340e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2218c4),
	.w1(32'hbb88a989),
	.w2(32'hbc66f76b),
	.w3(32'hbb5f68c2),
	.w4(32'hbc333b3d),
	.w5(32'hbc0c7ca6),
	.w6(32'h3ab1c587),
	.w7(32'hbba7126b),
	.w8(32'hbc08d6c9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52485a),
	.w1(32'h3bf228df),
	.w2(32'h3baa7b4b),
	.w3(32'hbb5a1b1d),
	.w4(32'hb7d8b5e5),
	.w5(32'hbb9c6081),
	.w6(32'hbbba2351),
	.w7(32'hbb07748f),
	.w8(32'hba929b09),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfae503),
	.w1(32'h3c7771f1),
	.w2(32'h3ba5e720),
	.w3(32'hbb9f783b),
	.w4(32'h3c03deca),
	.w5(32'h3bfd4c34),
	.w6(32'h3ac5af56),
	.w7(32'hbbbc9feb),
	.w8(32'h3c45feae),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0720a6),
	.w1(32'h3ab5017f),
	.w2(32'hbbf8c22f),
	.w3(32'h3b601f0d),
	.w4(32'h3bbe059f),
	.w5(32'hbbf6068d),
	.w6(32'h3c0dc3ac),
	.w7(32'h3b6e1bcb),
	.w8(32'hbb2b3911),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9faccb),
	.w1(32'hbbfdca2e),
	.w2(32'hbbb7df56),
	.w3(32'hba367623),
	.w4(32'h3ba5d17c),
	.w5(32'hbcba7c30),
	.w6(32'hbac3c5c7),
	.w7(32'h3c0768b4),
	.w8(32'hbbd3cda4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdacd1),
	.w1(32'hbaff354a),
	.w2(32'h3c0df728),
	.w3(32'hbbb03c7b),
	.w4(32'hbbe7aa1d),
	.w5(32'h3c331510),
	.w6(32'hbbf52ed5),
	.w7(32'hbb89e92a),
	.w8(32'hbbc78c12),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d966c),
	.w1(32'h3b3563fe),
	.w2(32'h3a6d3807),
	.w3(32'hbc729c44),
	.w4(32'h3b9a8055),
	.w5(32'h3c28b9b3),
	.w6(32'hbac28b94),
	.w7(32'h3ad1c76b),
	.w8(32'h3aa404f1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd175db),
	.w1(32'h3ae9d0d7),
	.w2(32'hbb456e18),
	.w3(32'h3b8a067f),
	.w4(32'h3bd3dc54),
	.w5(32'hbb29d7a6),
	.w6(32'h3b8574b1),
	.w7(32'h3aa4f15e),
	.w8(32'h3a9aedeb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20ef86),
	.w1(32'h3c2cccf4),
	.w2(32'hbb8b961e),
	.w3(32'hbc5c908b),
	.w4(32'h394ac321),
	.w5(32'hbbce4bba),
	.w6(32'hbb531e43),
	.w7(32'h3b516dab),
	.w8(32'h3ae4fabc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f38459),
	.w1(32'h3c1ae2f1),
	.w2(32'hba83255f),
	.w3(32'h3c629162),
	.w4(32'h3c857d80),
	.w5(32'h3bf029de),
	.w6(32'h3b63d50c),
	.w7(32'h3afd78d0),
	.w8(32'h3bd3381b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09282b),
	.w1(32'h3bfef631),
	.w2(32'h3aba71a3),
	.w3(32'hbc3aa16e),
	.w4(32'h3c1a5ead),
	.w5(32'hbbb61664),
	.w6(32'hb995419b),
	.w7(32'h3b6fea43),
	.w8(32'h3ae0e8d7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d51e9),
	.w1(32'hbc89e909),
	.w2(32'h3b37b1e8),
	.w3(32'hbbbeab27),
	.w4(32'hbc5fd1b4),
	.w5(32'h3bca7a23),
	.w6(32'h3bb4ec2e),
	.w7(32'hbb5ff255),
	.w8(32'hba2887e8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971098e),
	.w1(32'hbba531cf),
	.w2(32'h3b895adb),
	.w3(32'hbb302c23),
	.w4(32'h3a4804b0),
	.w5(32'h3c884852),
	.w6(32'hba1b1ed4),
	.w7(32'h36658bf0),
	.w8(32'h3bdceb70),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ac0be),
	.w1(32'h3bb90e8c),
	.w2(32'h3b962dd5),
	.w3(32'hbbf8cb4a),
	.w4(32'h3b496155),
	.w5(32'hbc64910c),
	.w6(32'h3a8b2c23),
	.w7(32'hbb60ec30),
	.w8(32'h3c1c733e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ffe52),
	.w1(32'h3b85beb1),
	.w2(32'h3b0f6f8c),
	.w3(32'h3cc54606),
	.w4(32'hbc40efcf),
	.w5(32'h3c01d103),
	.w6(32'h3c8dff2a),
	.w7(32'hba853605),
	.w8(32'hbbb0ee0d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4de0e1),
	.w1(32'hbb5d29d4),
	.w2(32'hbb328f35),
	.w3(32'hbbb33f05),
	.w4(32'hbae29407),
	.w5(32'hbc23c6a9),
	.w6(32'hbb287b45),
	.w7(32'h3a86b1b2),
	.w8(32'hbb80ac3e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6ee2d),
	.w1(32'hbbb720d2),
	.w2(32'hbc039f0a),
	.w3(32'h39e3f5af),
	.w4(32'hbc3c2c61),
	.w5(32'hbb0de2d9),
	.w6(32'hbb82e5e8),
	.w7(32'hbb5fec9d),
	.w8(32'hbbdc5279),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa04af),
	.w1(32'hbbd8ce25),
	.w2(32'h3b0f1e93),
	.w3(32'hbc2483c1),
	.w4(32'hbc04f1f5),
	.w5(32'h3b49038a),
	.w6(32'hbc173f32),
	.w7(32'h3aa7adb3),
	.w8(32'hbb9c2ec0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaddee),
	.w1(32'h3bbd1f92),
	.w2(32'hbb93cdb3),
	.w3(32'hbaa2b15d),
	.w4(32'h3bec1636),
	.w5(32'hbbac07ab),
	.w6(32'hbc063a7e),
	.w7(32'hbaa89f11),
	.w8(32'hbb8d55bc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62538c),
	.w1(32'hbbc50a2e),
	.w2(32'hbbb243ba),
	.w3(32'h3b1f94f8),
	.w4(32'h3b8baec4),
	.w5(32'hbc36a780),
	.w6(32'hbbe0ee80),
	.w7(32'hba9b8051),
	.w8(32'hbc08c6b4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80f53b),
	.w1(32'h3ba6d3c3),
	.w2(32'h3c4ccfae),
	.w3(32'hbbadc5d9),
	.w4(32'hbb38a0e2),
	.w5(32'h3c055c0d),
	.w6(32'hbb8cd611),
	.w7(32'hbc1629cd),
	.w8(32'hbc6e0c65),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e02bf),
	.w1(32'h38d86e07),
	.w2(32'hbb8200b2),
	.w3(32'hbc0ced1c),
	.w4(32'h3c12350c),
	.w5(32'hbc3fdb5b),
	.w6(32'hbc504e02),
	.w7(32'hba0cc71b),
	.w8(32'hb8915acc),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c804ffa),
	.w1(32'hbb240080),
	.w2(32'h3aaabe7e),
	.w3(32'h3c3995d7),
	.w4(32'hba75ee92),
	.w5(32'h3b9b1ea9),
	.w6(32'h3c4676c6),
	.w7(32'hbb8274da),
	.w8(32'hbb0ede9d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc108ce9),
	.w1(32'h3ae496c1),
	.w2(32'hbaf24fa2),
	.w3(32'hbbd00132),
	.w4(32'h3c1be91b),
	.w5(32'hbb4ebfa0),
	.w6(32'hbbb394e5),
	.w7(32'hbb905dce),
	.w8(32'h3c0f4a32),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb592c),
	.w1(32'hbc3aab9c),
	.w2(32'hba6ec22a),
	.w3(32'hbb933b1d),
	.w4(32'hbb957e1e),
	.w5(32'h3c80a7b3),
	.w6(32'h3bd850d8),
	.w7(32'h3ba66fd2),
	.w8(32'hbb505032),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a558426),
	.w1(32'h3b94142c),
	.w2(32'hbbbb5fa9),
	.w3(32'hb9e652fe),
	.w4(32'h3b303b9e),
	.w5(32'hbb893be2),
	.w6(32'hbba7626e),
	.w7(32'h3b2c66a6),
	.w8(32'hbb91ec9f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae9bc6),
	.w1(32'h3b7284b5),
	.w2(32'h3a85c69a),
	.w3(32'hbb022aea),
	.w4(32'hb92ce9d8),
	.w5(32'hbbbb0b56),
	.w6(32'h3a4bf87b),
	.w7(32'hb99c854b),
	.w8(32'hbc36877c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f7324),
	.w1(32'hbbabb29a),
	.w2(32'h3c0fa471),
	.w3(32'hbc367b80),
	.w4(32'h3ba88dbc),
	.w5(32'h3bc8b4bd),
	.w6(32'hbc103d5c),
	.w7(32'h3c181fc2),
	.w8(32'hbbaaee62),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c032eb9),
	.w1(32'hba97baa9),
	.w2(32'hbb060a41),
	.w3(32'h3bb5b9b9),
	.w4(32'h3bc7c3b4),
	.w5(32'hbbd1ee58),
	.w6(32'hbae43d64),
	.w7(32'h3b8a4fee),
	.w8(32'hbc0854a5),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c031867),
	.w1(32'h3b4a1320),
	.w2(32'h3bcde108),
	.w3(32'hba9e95c6),
	.w4(32'hbae59ae7),
	.w5(32'h3bf50879),
	.w6(32'h3b6e4ab7),
	.w7(32'h3bc5ea13),
	.w8(32'h3c0eb262),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9a741),
	.w1(32'hbb8371b0),
	.w2(32'hba93da2a),
	.w3(32'h39ed417a),
	.w4(32'hbbef48e4),
	.w5(32'hbc6c05e1),
	.w6(32'h3b05580a),
	.w7(32'hbc6d214f),
	.w8(32'hbc942cf1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c9069),
	.w1(32'hbb877e84),
	.w2(32'h3b967dc0),
	.w3(32'hbc5b9c04),
	.w4(32'hbc16731f),
	.w5(32'hba0fca96),
	.w6(32'hbba8eeab),
	.w7(32'hbc55d990),
	.w8(32'hbb923308),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1058ee),
	.w1(32'h3bf76bf9),
	.w2(32'h3b3aaae8),
	.w3(32'hbbc0bd7e),
	.w4(32'hbbae2453),
	.w5(32'h3bf40bbd),
	.w6(32'hbb63d819),
	.w7(32'h3c3c43c6),
	.w8(32'h3c17251b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99daa9),
	.w1(32'h3bb9b213),
	.w2(32'hbb92f164),
	.w3(32'h3cf4cf3c),
	.w4(32'h3bc2774a),
	.w5(32'hbc7acfc4),
	.w6(32'h3c8f4a6a),
	.w7(32'h39d31ff6),
	.w8(32'hbbc063f1),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b8c54),
	.w1(32'h3a9af9a1),
	.w2(32'hbc5491e9),
	.w3(32'h3bbc31e9),
	.w4(32'h3c1abc62),
	.w5(32'hbc0d2f9a),
	.w6(32'h3b460ddf),
	.w7(32'h3c0d415b),
	.w8(32'h3acd83b8),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc322a4b),
	.w1(32'hbab4a7e6),
	.w2(32'hbc33f6cb),
	.w3(32'hbb147f56),
	.w4(32'hbaa194aa),
	.w5(32'hbc288893),
	.w6(32'hbb007283),
	.w7(32'h3b23a531),
	.w8(32'hb9fb5348),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc039f3d),
	.w1(32'h3b565c1f),
	.w2(32'h3b0a70ad),
	.w3(32'h3acf0a40),
	.w4(32'hbc413ff9),
	.w5(32'hbb87a994),
	.w6(32'hbaceb9a7),
	.w7(32'hb956423c),
	.w8(32'h3bd3d46e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a4285),
	.w1(32'hba78af2a),
	.w2(32'h3978aba8),
	.w3(32'h3cdc52c0),
	.w4(32'h3ba0be00),
	.w5(32'hbb59ab1e),
	.w6(32'h3c04ccdb),
	.w7(32'h3ba4b7c5),
	.w8(32'hbb0ca114),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88ef80),
	.w1(32'h3af07b07),
	.w2(32'h3c11c904),
	.w3(32'h3a93f88c),
	.w4(32'h3c544ec2),
	.w5(32'hbc3e0114),
	.w6(32'h3b6396b4),
	.w7(32'h3bf55652),
	.w8(32'hbb19c1c7),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb402aad),
	.w1(32'hbc0df5f3),
	.w2(32'hbb295af1),
	.w3(32'hbbc97617),
	.w4(32'hbb8d0023),
	.w5(32'hbc03a301),
	.w6(32'h3c3ac139),
	.w7(32'h39ab53b8),
	.w8(32'hba0bec8d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac44829),
	.w1(32'h3c13a350),
	.w2(32'h3c12170d),
	.w3(32'h3bb2d809),
	.w4(32'h3b91bdb2),
	.w5(32'hbc86929d),
	.w6(32'hbb140c2f),
	.w7(32'hbc07a7ba),
	.w8(32'hbb999829),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3783f2),
	.w1(32'hbb68b734),
	.w2(32'hbbb6ffbf),
	.w3(32'hbbb68320),
	.w4(32'hbb909bcb),
	.w5(32'h3b979877),
	.w6(32'h3b085b27),
	.w7(32'hbb1fa4bf),
	.w8(32'hbb3d4c45),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea74af),
	.w1(32'h38433026),
	.w2(32'hbc848f89),
	.w3(32'hbc267f12),
	.w4(32'h3ba38472),
	.w5(32'hbbc6e6f3),
	.w6(32'hbc3e16b2),
	.w7(32'h3a47f70f),
	.w8(32'hbbe8569c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a718e),
	.w1(32'h3b705c4a),
	.w2(32'h3b7eafce),
	.w3(32'hbc1cd47d),
	.w4(32'hb9e93a9b),
	.w5(32'h3c0a006b),
	.w6(32'hbc78ae23),
	.w7(32'h3b800aa5),
	.w8(32'hbbf86410),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3b6aa),
	.w1(32'h3baa7bc6),
	.w2(32'h3bdf17ed),
	.w3(32'h3a923685),
	.w4(32'hbab0ac45),
	.w5(32'h3a0c3899),
	.w6(32'hbc2a4c5d),
	.w7(32'hbb5e5cf1),
	.w8(32'hbb9985d1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88e20e),
	.w1(32'hbb04fa67),
	.w2(32'hbc751d99),
	.w3(32'hb9549445),
	.w4(32'h3ca06ad5),
	.w5(32'hbbd6bb97),
	.w6(32'hbbc46662),
	.w7(32'h3bb4dd01),
	.w8(32'hbbf3dea6),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4f016),
	.w1(32'h3baa06c0),
	.w2(32'h3b543645),
	.w3(32'hbc777a4d),
	.w4(32'h3b7653ac),
	.w5(32'h3cd064bc),
	.w6(32'hbbdbe6b9),
	.w7(32'h3b5d500a),
	.w8(32'hbba40b95),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11d897),
	.w1(32'hbc5586d2),
	.w2(32'h39d98db7),
	.w3(32'hbc8e1be0),
	.w4(32'hbc71aa1f),
	.w5(32'h3c236f66),
	.w6(32'hbbd19b5e),
	.w7(32'hbb9b9071),
	.w8(32'hbc02c415),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49a1bc),
	.w1(32'hbb9365fe),
	.w2(32'h3ad37f3d),
	.w3(32'hbbae3461),
	.w4(32'hbb092ae5),
	.w5(32'hbc44ab93),
	.w6(32'hbc185924),
	.w7(32'hba5cc3ce),
	.w8(32'hbc2a51ab),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f227e),
	.w1(32'hbc323d49),
	.w2(32'h3ca29e80),
	.w3(32'hbcbca708),
	.w4(32'h3cd19615),
	.w5(32'h3d0fde7a),
	.w6(32'hbc2d504e),
	.w7(32'h3cd4a997),
	.w8(32'hbaa5a969),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d2ed3),
	.w1(32'hbb8df083),
	.w2(32'hbba31a21),
	.w3(32'h3c7945e9),
	.w4(32'hbb6af0b2),
	.w5(32'hbbd87967),
	.w6(32'hbc19e408),
	.w7(32'h3a620545),
	.w8(32'hbc0f70ad),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e268d),
	.w1(32'hbb165ad0),
	.w2(32'h3c736e96),
	.w3(32'hbb8ab328),
	.w4(32'h3abd1a63),
	.w5(32'hbaaa8534),
	.w6(32'hbc06dbf1),
	.w7(32'h3977dad8),
	.w8(32'hbb8b857b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10662b),
	.w1(32'hba084738),
	.w2(32'hbb0c8fb4),
	.w3(32'h3c5972b0),
	.w4(32'h3804baa1),
	.w5(32'hbb7ab69a),
	.w6(32'h3bca1655),
	.w7(32'h37b493f5),
	.w8(32'h3a93cfd3),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba48ff9),
	.w1(32'h3bdabf6c),
	.w2(32'h3a796282),
	.w3(32'hbb686193),
	.w4(32'h3b95e446),
	.w5(32'hbbdc601c),
	.w6(32'hbc12c457),
	.w7(32'hbb8cc6f6),
	.w8(32'h3b496e85),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9cf9d),
	.w1(32'h3bb236df),
	.w2(32'h3c0b8586),
	.w3(32'hbb5f2e40),
	.w4(32'h3c0aefab),
	.w5(32'hbae4e675),
	.w6(32'hbbbb6f80),
	.w7(32'h3b8f8de5),
	.w8(32'hbb7d5b56),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba357b39),
	.w1(32'h3bb45b99),
	.w2(32'h3b085291),
	.w3(32'hbb27822d),
	.w4(32'h3bd66340),
	.w5(32'hbb9988d1),
	.w6(32'hbb8fb397),
	.w7(32'h3c7fb42e),
	.w8(32'hbbaedc58),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2effb0),
	.w1(32'hbb89c2e9),
	.w2(32'h3bfc1db7),
	.w3(32'hbb07a794),
	.w4(32'hbb87ad2b),
	.w5(32'h3c53bab2),
	.w6(32'hbb6c6dec),
	.w7(32'h3bae2c04),
	.w8(32'h3b9d1904),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc303a1),
	.w1(32'hbc12dced),
	.w2(32'hbc0e2671),
	.w3(32'h3b67b06c),
	.w4(32'hbc0f409f),
	.w5(32'h3be6baad),
	.w6(32'h3bb805ea),
	.w7(32'hbb80ff0f),
	.w8(32'hba84c6b4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0be135),
	.w1(32'hbc462d54),
	.w2(32'hbbfa2414),
	.w3(32'hba13b58d),
	.w4(32'hbbee61e2),
	.w5(32'hbc1e16ce),
	.w6(32'h3c07a2da),
	.w7(32'hbc164f9e),
	.w8(32'hbbabfa81),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c1fb3),
	.w1(32'h3bdd1178),
	.w2(32'hbbb4baa5),
	.w3(32'hbb78df5a),
	.w4(32'h3a91711f),
	.w5(32'hbb754ffd),
	.w6(32'hbb89727d),
	.w7(32'hbba6cebd),
	.w8(32'h3bd73692),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3c4d9),
	.w1(32'hbbf52ff8),
	.w2(32'hbb03ee47),
	.w3(32'h3bbef474),
	.w4(32'h3b7a8363),
	.w5(32'h3abef1fb),
	.w6(32'h3c519f41),
	.w7(32'hbbc57ca7),
	.w8(32'hbb7ebd79),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc788aa4),
	.w1(32'h3b6ffb1a),
	.w2(32'h3b858656),
	.w3(32'hbc37e7f4),
	.w4(32'hba959a51),
	.w5(32'h3d00a3fa),
	.w6(32'hbc436494),
	.w7(32'hbabef005),
	.w8(32'h3b0e7d7a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5daa35),
	.w1(32'hbbb15dbe),
	.w2(32'hbb550a49),
	.w3(32'h3c16d4e5),
	.w4(32'hbb88897d),
	.w5(32'h3c1e9088),
	.w6(32'hbb6a455c),
	.w7(32'hb9d1829d),
	.w8(32'hbb123c30),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03ea08),
	.w1(32'h3b449f5a),
	.w2(32'h3b1a3f2a),
	.w3(32'h3ae97072),
	.w4(32'h3b7b7bd8),
	.w5(32'h3c2dff50),
	.w6(32'h379edd15),
	.w7(32'h3b55c0bb),
	.w8(32'hbb2d92f5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7aee8),
	.w1(32'h3b780626),
	.w2(32'h3b83ef44),
	.w3(32'h3a2e221b),
	.w4(32'h39a83f2d),
	.w5(32'h3989c208),
	.w6(32'hbb1b4cc4),
	.w7(32'hbadbebed),
	.w8(32'h3bbbbdef),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c660a8a),
	.w1(32'h3c21e782),
	.w2(32'hbb5db1f9),
	.w3(32'h3b8549e9),
	.w4(32'h3b979659),
	.w5(32'hbbd736e7),
	.w6(32'hbae3219e),
	.w7(32'h3bd56165),
	.w8(32'hbb07f870),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b560f),
	.w1(32'h3c6cc66d),
	.w2(32'h3c59a7a0),
	.w3(32'h3bda63bd),
	.w4(32'hbc5b70be),
	.w5(32'h3ce931d1),
	.w6(32'hb96c8724),
	.w7(32'h3b9312b1),
	.w8(32'h3c9d2608),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4810d3),
	.w1(32'hba76f835),
	.w2(32'hbba3d7af),
	.w3(32'h3d1348f7),
	.w4(32'hbbdb5e59),
	.w5(32'hbbb2729c),
	.w6(32'h3c4fd0d7),
	.w7(32'hbbf0a0f9),
	.w8(32'h3b6b1870),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc036cd7),
	.w1(32'h3af19516),
	.w2(32'h3c3b37d6),
	.w3(32'hbbdc06d4),
	.w4(32'hba4856d1),
	.w5(32'h3c10dca9),
	.w6(32'hbc151ed0),
	.w7(32'h3a31a5de),
	.w8(32'h3c4cd682),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c426393),
	.w1(32'hb88afec4),
	.w2(32'h3b7344ec),
	.w3(32'h3c367fef),
	.w4(32'hbada9165),
	.w5(32'h3b21d70b),
	.w6(32'h3bbddfa5),
	.w7(32'hbab5df4f),
	.w8(32'hba01ebf8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0effa),
	.w1(32'hbac085ed),
	.w2(32'hbb57a256),
	.w3(32'h395f118b),
	.w4(32'hb9dc4722),
	.w5(32'h3c01147e),
	.w6(32'hbb691226),
	.w7(32'h3aa4bf18),
	.w8(32'hba5c1c58),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4a886),
	.w1(32'h37b77d36),
	.w2(32'h3b5c184f),
	.w3(32'h3a74f0d2),
	.w4(32'h3c336517),
	.w5(32'hbaa2ea22),
	.w6(32'hbafc23a6),
	.w7(32'hbbe088ba),
	.w8(32'hbbe256d8),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2f907),
	.w1(32'h3be7680b),
	.w2(32'h3c8ace4c),
	.w3(32'hbc68d8ad),
	.w4(32'hbc08ecca),
	.w5(32'h3cfe9182),
	.w6(32'hbc173856),
	.w7(32'hbb23941b),
	.w8(32'h3cb93da8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24f673),
	.w1(32'h3a3d9f0d),
	.w2(32'h3a04cbcb),
	.w3(32'h3c446f26),
	.w4(32'h3bcd3d67),
	.w5(32'hba5bd64b),
	.w6(32'h3c27515f),
	.w7(32'h3bd11035),
	.w8(32'hbb27a1c2),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a120d),
	.w1(32'hbad0dcc6),
	.w2(32'hbb529a4e),
	.w3(32'hbba96eb1),
	.w4(32'h3bc3c9ad),
	.w5(32'h3a4a4a5a),
	.w6(32'h3b5b8c23),
	.w7(32'h3b0d9e32),
	.w8(32'hbb069585),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89a20d),
	.w1(32'hbb8df65f),
	.w2(32'hbc255c6a),
	.w3(32'hbbea90d5),
	.w4(32'hba1d919c),
	.w5(32'hbc97832c),
	.w6(32'h3bc556ff),
	.w7(32'hbb8a9bd7),
	.w8(32'hbc122a3f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f8ceb),
	.w1(32'hbb7c95af),
	.w2(32'hbad6ed40),
	.w3(32'hbb474e62),
	.w4(32'h3bfd8639),
	.w5(32'hbb466630),
	.w6(32'h3a8f8498),
	.w7(32'h3bb637b6),
	.w8(32'hbb8b24fb),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd34b8),
	.w1(32'hbb93e0ce),
	.w2(32'h3adce17e),
	.w3(32'h3b9b32b0),
	.w4(32'hbc11d44b),
	.w5(32'h3ba38cb9),
	.w6(32'hba2cec1b),
	.w7(32'hbc0e0298),
	.w8(32'h3a7704fa),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b1c28),
	.w1(32'h3b71a0ed),
	.w2(32'hbb9b0ae9),
	.w3(32'hbb85b729),
	.w4(32'hbaf6360b),
	.w5(32'hbb62cf0e),
	.w6(32'hbab5b7a0),
	.w7(32'h3a8c00bb),
	.w8(32'hba75e110),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae83516),
	.w1(32'h3a3b0af5),
	.w2(32'hbc0befa2),
	.w3(32'hbbd29fe3),
	.w4(32'hbc3e4773),
	.w5(32'hbad07631),
	.w6(32'hbbdb2443),
	.w7(32'hbc19a930),
	.w8(32'hbb6502de),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6097b0),
	.w1(32'hba5141bf),
	.w2(32'hbc13b996),
	.w3(32'h3b8b50b0),
	.w4(32'h3b0bce56),
	.w5(32'hbb14e843),
	.w6(32'hbc3d5dd9),
	.w7(32'hbc4f4a55),
	.w8(32'hbbfe6dba),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d397b),
	.w1(32'h386dfef0),
	.w2(32'hbc06e56f),
	.w3(32'h3a292a57),
	.w4(32'h39c0028b),
	.w5(32'hbbe9bc75),
	.w6(32'hbb665d46),
	.w7(32'h3bf101c1),
	.w8(32'hbad0ce0d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc15621),
	.w1(32'h3b4fa179),
	.w2(32'h3c27f8b9),
	.w3(32'hbc3d7cd1),
	.w4(32'h3b6e5f63),
	.w5(32'h3c073a47),
	.w6(32'hbbaa703f),
	.w7(32'h3c083b70),
	.w8(32'h3c01a143),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47986c),
	.w1(32'hbc6b3772),
	.w2(32'hbba830de),
	.w3(32'hbb30c66e),
	.w4(32'hbc2f5a73),
	.w5(32'h3c8380d3),
	.w6(32'h3aaab9a9),
	.w7(32'hbc5a4a19),
	.w8(32'hbbe789a2),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb83402),
	.w1(32'h3b3d2fbf),
	.w2(32'hb9c1bf79),
	.w3(32'hbc4a080b),
	.w4(32'hbb3f2526),
	.w5(32'hbc457bd2),
	.w6(32'hbc373abe),
	.w7(32'hba818f38),
	.w8(32'h3b8cbab5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e4eaa),
	.w1(32'hbbee6a11),
	.w2(32'hbb35db56),
	.w3(32'h3c985c31),
	.w4(32'hbbf577a4),
	.w5(32'hbc057268),
	.w6(32'h3c7a5df2),
	.w7(32'hbbd452cf),
	.w8(32'hbba11f5c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ebb9b),
	.w1(32'h390cefe3),
	.w2(32'h3b3aeebc),
	.w3(32'hba04da08),
	.w4(32'hbc1b3d1f),
	.w5(32'h3cebc396),
	.w6(32'h397e81ff),
	.w7(32'hba8ea757),
	.w8(32'h3b9f9d59),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97b091),
	.w1(32'hb9ada008),
	.w2(32'h3bcac64b),
	.w3(32'hbbf391e2),
	.w4(32'h3b491e6c),
	.w5(32'h3ad0e84e),
	.w6(32'hbaf78ae1),
	.w7(32'hbadcb7d5),
	.w8(32'hba4f817c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe4421),
	.w1(32'h3a0be26c),
	.w2(32'h3c4df04d),
	.w3(32'hbc3b610c),
	.w4(32'h3c26d363),
	.w5(32'h3bc22ed3),
	.w6(32'hbb8961b4),
	.w7(32'h3baabae8),
	.w8(32'h3c432e85),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60650c),
	.w1(32'h3b90d3c5),
	.w2(32'h3c45b1c3),
	.w3(32'hbc5758ff),
	.w4(32'h3ce2be0c),
	.w5(32'hba0c07dd),
	.w6(32'hba71fb3d),
	.w7(32'h3b995ce2),
	.w8(32'h39c59467),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc085f7),
	.w1(32'hbb858795),
	.w2(32'h3c0572d9),
	.w3(32'hba1d7dc8),
	.w4(32'hbbc91112),
	.w5(32'h3cacc143),
	.w6(32'h3aa30690),
	.w7(32'hbbb5fcb5),
	.w8(32'hbc104057),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2075d5),
	.w1(32'h3b1190f9),
	.w2(32'h3c11312c),
	.w3(32'hbc48f7fe),
	.w4(32'hbb081df8),
	.w5(32'h3b2cab61),
	.w6(32'hbbf9d2df),
	.w7(32'hbb2c28d5),
	.w8(32'hbae19bf4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7af32d),
	.w1(32'h3ab1f17d),
	.w2(32'h3aeb4e6e),
	.w3(32'hbb930012),
	.w4(32'h395c0d9b),
	.w5(32'h3a9ab659),
	.w6(32'h3aa07923),
	.w7(32'hbb81a5bf),
	.w8(32'hbadd90b0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6faea6),
	.w1(32'h3c1fbafc),
	.w2(32'h3a5aa59b),
	.w3(32'h3be042d4),
	.w4(32'hb986c320),
	.w5(32'h3b94b62f),
	.w6(32'hbba64808),
	.w7(32'h3ad32850),
	.w8(32'h3ad76ec4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fede8),
	.w1(32'hba0a0ff8),
	.w2(32'h3af7fcd6),
	.w3(32'h3c093254),
	.w4(32'h3ad24f5c),
	.w5(32'hbb7197bf),
	.w6(32'h3c3203ed),
	.w7(32'h3b529cac),
	.w8(32'hb8e7252d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a6df9),
	.w1(32'hba925569),
	.w2(32'h3b49a88d),
	.w3(32'h3b43b569),
	.w4(32'hbb1bf82b),
	.w5(32'h3b17d381),
	.w6(32'h3af703ad),
	.w7(32'hbb38ba4e),
	.w8(32'h3a2a7ede),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95bc90),
	.w1(32'h3aa306e0),
	.w2(32'h3a23fe47),
	.w3(32'h3ac8fb1a),
	.w4(32'h3b10ff13),
	.w5(32'hbc557cf4),
	.w6(32'h3ad976bf),
	.w7(32'h3bb27556),
	.w8(32'hbaa53c7f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49d5f6),
	.w1(32'hbaa33423),
	.w2(32'hbb475d92),
	.w3(32'hbc1afde9),
	.w4(32'hbbd8dab1),
	.w5(32'hb98e6f5b),
	.w6(32'hb9911564),
	.w7(32'h3c086d52),
	.w8(32'h3ae485ef),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77bd9c),
	.w1(32'hbbb96938),
	.w2(32'hbbf742f3),
	.w3(32'h3c967831),
	.w4(32'h3bb22572),
	.w5(32'hbb99fea7),
	.w6(32'h3c814779),
	.w7(32'h3b850168),
	.w8(32'h3c0bf234),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b023a87),
	.w1(32'h3b94a723),
	.w2(32'h3ba0db2d),
	.w3(32'hbb223d41),
	.w4(32'hbb1814aa),
	.w5(32'h3bd94639),
	.w6(32'h3aa951d4),
	.w7(32'hbb3b14d5),
	.w8(32'h3bdc87b1),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25fd66),
	.w1(32'h3b7759a2),
	.w2(32'hbbca5b19),
	.w3(32'h3c1c8ab5),
	.w4(32'hbb66cf21),
	.w5(32'hb962ce2f),
	.w6(32'h398b4d79),
	.w7(32'h3c12862f),
	.w8(32'hbb38abf5),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19485f),
	.w1(32'h3afe626e),
	.w2(32'h3a0ada7f),
	.w3(32'h3c0b8658),
	.w4(32'hbb40bbeb),
	.w5(32'hbc86e4dc),
	.w6(32'h3a2f03a6),
	.w7(32'h3be91fb3),
	.w8(32'h3c9a0c97),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4a3b1),
	.w1(32'hbb9fb6b1),
	.w2(32'hbbb646e5),
	.w3(32'h3c53fd15),
	.w4(32'h3b332bf7),
	.w5(32'hbb3c2cdb),
	.w6(32'h3c422274),
	.w7(32'h3b9b24ae),
	.w8(32'h3bb0c9e5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba146c1c),
	.w1(32'h3b145aa6),
	.w2(32'h39d0adcd),
	.w3(32'hbba1c127),
	.w4(32'h3ba95aea),
	.w5(32'h3aeb3895),
	.w6(32'h3b03e2d6),
	.w7(32'h3b6bd7d9),
	.w8(32'h3a61f45c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88e851),
	.w1(32'h3c1a91df),
	.w2(32'h3c31b1a1),
	.w3(32'hbb437f82),
	.w4(32'h3c14113e),
	.w5(32'h3bd7dd83),
	.w6(32'hbb5a5e3c),
	.w7(32'h3b30eb07),
	.w8(32'hbb2c486b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc05849),
	.w1(32'h39ef1150),
	.w2(32'h3b12fa5c),
	.w3(32'hbabdfe2d),
	.w4(32'hbaf98575),
	.w5(32'h3c14c69e),
	.w6(32'h3b62127f),
	.w7(32'hbb01e1a0),
	.w8(32'h3b4f3928),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc37492),
	.w1(32'hbba0d5ce),
	.w2(32'hbab2e92d),
	.w3(32'hbb27b2f1),
	.w4(32'hbbf7c203),
	.w5(32'hbba582ed),
	.w6(32'h3b1a929b),
	.w7(32'hbc3d79ac),
	.w8(32'hbc3a4b6c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92cc5d),
	.w1(32'hbb827ba3),
	.w2(32'hbb70734f),
	.w3(32'hbc31354a),
	.w4(32'hbbaa3fd2),
	.w5(32'h3ab3d570),
	.w6(32'hbc5bcb8e),
	.w7(32'h3beb5184),
	.w8(32'h3b75c1f0),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc329ab2),
	.w1(32'hbb624d5d),
	.w2(32'h3b142b6f),
	.w3(32'hbbc27db4),
	.w4(32'hbb7b2bb0),
	.w5(32'hbc15ac76),
	.w6(32'hba8f0916),
	.w7(32'h3b355234),
	.w8(32'hba8503c7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba64e7b),
	.w1(32'h3b9afe46),
	.w2(32'h3a86348f),
	.w3(32'hbb6625a9),
	.w4(32'h3a7495fc),
	.w5(32'hbb00e0d7),
	.w6(32'hbba5e349),
	.w7(32'hbb8e4f7e),
	.w8(32'hbb947e90),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb62b1b),
	.w1(32'h3b945282),
	.w2(32'h3c1e947b),
	.w3(32'h3b9e935c),
	.w4(32'h3c18a53f),
	.w5(32'h3c203cc1),
	.w6(32'hbb472753),
	.w7(32'h3bc0402c),
	.w8(32'h39b83146),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee14be),
	.w1(32'hbb7af93d),
	.w2(32'hb9bae830),
	.w3(32'h39f7b17b),
	.w4(32'h3b2e990a),
	.w5(32'h3c24565a),
	.w6(32'hbbe567e5),
	.w7(32'hbb79ef55),
	.w8(32'hbb7666b8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addfc30),
	.w1(32'h3bf4c629),
	.w2(32'h3c33a465),
	.w3(32'hba611b22),
	.w4(32'hbb9d3e80),
	.w5(32'hbba471d4),
	.w6(32'hbb09e6c6),
	.w7(32'hbc51e9ac),
	.w8(32'hbbe23c83),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb994548),
	.w1(32'hbb6a1a7a),
	.w2(32'hbb0b4a00),
	.w3(32'hbb11cdcd),
	.w4(32'hbac168f6),
	.w5(32'h3b6705e9),
	.w6(32'h392e0d90),
	.w7(32'hb9b28929),
	.w8(32'h3be6598c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5ea1c),
	.w1(32'hbb1a336c),
	.w2(32'h3bc6ac74),
	.w3(32'h3b2ffbf9),
	.w4(32'hbb6b6187),
	.w5(32'hbabb8800),
	.w6(32'h3c13f101),
	.w7(32'h3bd754f8),
	.w8(32'h3bf84f5e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a8989),
	.w1(32'h3bc4f6d1),
	.w2(32'hbb993d2b),
	.w3(32'hbb56d7f0),
	.w4(32'h3a06a548),
	.w5(32'hba4aac5d),
	.w6(32'h3a55ef2b),
	.w7(32'hbbb2a810),
	.w8(32'hbb5af925),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa5481),
	.w1(32'h3ba73e4f),
	.w2(32'h3a5a6ac1),
	.w3(32'h3ac15e2c),
	.w4(32'hbc02bb04),
	.w5(32'h3c4c72a5),
	.w6(32'hbb10316c),
	.w7(32'hb9c1dbd6),
	.w8(32'hbc213da2),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc059df6),
	.w1(32'hbb73845d),
	.w2(32'h3b024186),
	.w3(32'hba3375b9),
	.w4(32'h3b16cf5b),
	.w5(32'hbbce7df9),
	.w6(32'hbb95f5d2),
	.w7(32'hba8f73c7),
	.w8(32'hbb8a8d27),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd4235),
	.w1(32'hbb9fd113),
	.w2(32'hbc09f93e),
	.w3(32'hbbdc34e5),
	.w4(32'hbc1e0c42),
	.w5(32'hbbaa8002),
	.w6(32'hbb77e3b8),
	.w7(32'h3a4424c4),
	.w8(32'hbb782e3c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3239a6),
	.w1(32'h3b0e463b),
	.w2(32'h3c18af57),
	.w3(32'h3ae77a01),
	.w4(32'h3b8563b8),
	.w5(32'h3c7f06da),
	.w6(32'hbb5733cf),
	.w7(32'hbb973343),
	.w8(32'h3aaaa73f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaef45f),
	.w1(32'hbb5de813),
	.w2(32'hbb8f9164),
	.w3(32'h3b486ed2),
	.w4(32'h3a837a73),
	.w5(32'hbaa7a8a0),
	.w6(32'hba3d553b),
	.w7(32'hbb16d63b),
	.w8(32'h3a0ee450),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ddfa1),
	.w1(32'hbb235fa1),
	.w2(32'h3bedafc9),
	.w3(32'hbb8332d5),
	.w4(32'hbb6a6441),
	.w5(32'hba9b75c5),
	.w6(32'hbc2d3b2c),
	.w7(32'h3b7d6bf7),
	.w8(32'h3b36d31e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a703de6),
	.w1(32'h3a3b28f0),
	.w2(32'hbb91625d),
	.w3(32'h3b843154),
	.w4(32'h3b6f7445),
	.w5(32'h38a88871),
	.w6(32'h3bf68398),
	.w7(32'hbbac141e),
	.w8(32'hbbaa6b19),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6db3d),
	.w1(32'h3c2e1e08),
	.w2(32'h3bfd7bcf),
	.w3(32'hbbd554cc),
	.w4(32'h3b651e7d),
	.w5(32'h3af4a2dd),
	.w6(32'hbbe10777),
	.w7(32'hbb424532),
	.w8(32'h39e4016f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74db44),
	.w1(32'h3b1addf3),
	.w2(32'h3a7cde67),
	.w3(32'h3b251924),
	.w4(32'h3b546152),
	.w5(32'h3ba14481),
	.w6(32'hbb8d828a),
	.w7(32'h3997ee7e),
	.w8(32'h3bc8cb78),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915acde),
	.w1(32'hba35a438),
	.w2(32'hbb110b4d),
	.w3(32'h3aa60dcd),
	.w4(32'h3be1c20a),
	.w5(32'hbba8b636),
	.w6(32'h3931e44f),
	.w7(32'hbae88a9e),
	.w8(32'h3bcdea8a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80efc3),
	.w1(32'h3c3c98fd),
	.w2(32'h3af1e677),
	.w3(32'h3ac58b6f),
	.w4(32'h3bc1e652),
	.w5(32'hbbd98329),
	.w6(32'h3b9dd44e),
	.w7(32'h3b54360d),
	.w8(32'h3b15a1fd),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0af775),
	.w1(32'hbbc7cf22),
	.w2(32'hbc1b9801),
	.w3(32'hbb8c0d5e),
	.w4(32'hbba0df11),
	.w5(32'hbb915651),
	.w6(32'hbb795bfc),
	.w7(32'h3a45f1da),
	.w8(32'hbb63feca),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42ebc0),
	.w1(32'hbbd5180a),
	.w2(32'h3bc120ed),
	.w3(32'hbc1de3bc),
	.w4(32'hbb8c19a4),
	.w5(32'h3b8c84da),
	.w6(32'hbbca9f26),
	.w7(32'hbbf41026),
	.w8(32'hba61aa16),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf61dd9),
	.w1(32'hbb9aea3f),
	.w2(32'hbaa4e311),
	.w3(32'h394e3fc5),
	.w4(32'hbac16036),
	.w5(32'hbb2319a4),
	.w6(32'hbb9bff5a),
	.w7(32'hbb7590ec),
	.w8(32'h3981b2e2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02ba80),
	.w1(32'h3be30c67),
	.w2(32'h3baa2966),
	.w3(32'hbbf5c908),
	.w4(32'hba5a2b7f),
	.w5(32'hbc426b5d),
	.w6(32'hbb7c15f2),
	.w7(32'h3b8ff733),
	.w8(32'h3b0152f7),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb60a9d),
	.w1(32'hbb8f5b05),
	.w2(32'h3b242df5),
	.w3(32'h3baccbcf),
	.w4(32'hbc233f4c),
	.w5(32'hbc22701d),
	.w6(32'h3b2d9375),
	.w7(32'hbc199998),
	.w8(32'hbbd8c804),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb029af1),
	.w1(32'h3b42cb03),
	.w2(32'hbc706807),
	.w3(32'hbbd1dde6),
	.w4(32'h3cdec09b),
	.w5(32'hbc2754cc),
	.w6(32'hbbf48cb2),
	.w7(32'h3bd20d11),
	.w8(32'hba10f081),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb515ed7),
	.w1(32'h3b954761),
	.w2(32'hba896068),
	.w3(32'hbbfacdea),
	.w4(32'h3bb00675),
	.w5(32'h3a3be7b9),
	.w6(32'hbc1b3f57),
	.w7(32'h3b6e983f),
	.w8(32'hba134a04),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc266ca),
	.w1(32'h3b051527),
	.w2(32'hbb4ad0e9),
	.w3(32'h3b70ea30),
	.w4(32'hba81ec23),
	.w5(32'hbc020997),
	.w6(32'h3baefa3b),
	.w7(32'h3c0a0f60),
	.w8(32'h3a44ded1),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78ce7e),
	.w1(32'hbbc8a3da),
	.w2(32'h3c14e5eb),
	.w3(32'h3a159c9b),
	.w4(32'hbc09ed61),
	.w5(32'h3c8e057c),
	.w6(32'hbc2a934e),
	.w7(32'hbbe34427),
	.w8(32'h3b70bff1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba949ef0),
	.w1(32'h3c0f6cb2),
	.w2(32'h3a68d89f),
	.w3(32'hbbce0276),
	.w4(32'h3c7901d3),
	.w5(32'hbbc922ff),
	.w6(32'hba6970c7),
	.w7(32'h39f62f62),
	.w8(32'h3b07f76f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bc00b),
	.w1(32'h3ba66713),
	.w2(32'hbb49bae0),
	.w3(32'hbad88317),
	.w4(32'h3bc5afd0),
	.w5(32'h3cb8c20d),
	.w6(32'h3a39bd3d),
	.w7(32'hba7f22e0),
	.w8(32'hbb8c2be4),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80e7ac),
	.w1(32'hbbe669f8),
	.w2(32'hbb7b2ad7),
	.w3(32'hbc2d1d17),
	.w4(32'hbae40d92),
	.w5(32'h3aceba5f),
	.w6(32'hbb8dad8e),
	.w7(32'hbb24d06d),
	.w8(32'hbb1e0ba7),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cce1ad),
	.w1(32'hb9667082),
	.w2(32'hbbf525b7),
	.w3(32'hba774144),
	.w4(32'h3bce73c4),
	.w5(32'hbb88af3f),
	.w6(32'hb7ff5cc0),
	.w7(32'hb74d8d6c),
	.w8(32'h398d38a9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b007ee1),
	.w1(32'h3c05d2d7),
	.w2(32'hbb096d82),
	.w3(32'h3b0f445b),
	.w4(32'h3bc350ef),
	.w5(32'h3c0d669d),
	.w6(32'h3b86984f),
	.w7(32'h3b9f1680),
	.w8(32'h3acb30cb),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3b622),
	.w1(32'h3aef1f65),
	.w2(32'h3b82bfbe),
	.w3(32'hb97d2adf),
	.w4(32'hbbc4e8e3),
	.w5(32'hbbeffc70),
	.w6(32'hbab606f1),
	.w7(32'h3b960936),
	.w8(32'h3b6df2ff),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c864a06),
	.w1(32'h3aaf76a5),
	.w2(32'hbba5f9f8),
	.w3(32'h3c3b1dc3),
	.w4(32'hbbd11d13),
	.w5(32'h3a346748),
	.w6(32'h3c73b366),
	.w7(32'hbbbb8393),
	.w8(32'hba91756f),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ec145),
	.w1(32'hbc1e77ff),
	.w2(32'h3a886792),
	.w3(32'hbc33c12d),
	.w4(32'h3a253b75),
	.w5(32'hbbdbaaae),
	.w6(32'hbc2ca380),
	.w7(32'hbaae43e2),
	.w8(32'hbb87df29),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7bd10),
	.w1(32'h3b440109),
	.w2(32'hbc472b93),
	.w3(32'hbbc10d3e),
	.w4(32'h3c448e1f),
	.w5(32'hbc937613),
	.w6(32'hbb5d1136),
	.w7(32'h3b757dac),
	.w8(32'hbbdb6e82),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99f4ce),
	.w1(32'hbbb76391),
	.w2(32'hbc375df0),
	.w3(32'hbc34d14c),
	.w4(32'h3c641499),
	.w5(32'hbafd76b7),
	.w6(32'hbc2663dc),
	.w7(32'h3b823860),
	.w8(32'h3c128b53),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c610882),
	.w1(32'h3b20920f),
	.w2(32'hbbcd9926),
	.w3(32'hbb4762cc),
	.w4(32'h3b556e28),
	.w5(32'hbbe9bd6b),
	.w6(32'hbb8e7fa9),
	.w7(32'h3b08bf7b),
	.w8(32'hbb9e8a7a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baac2f5),
	.w1(32'hbb664298),
	.w2(32'hbb1cfc06),
	.w3(32'h3b205666),
	.w4(32'hbbb3e27e),
	.w5(32'h3bd6a49f),
	.w6(32'h39dce13e),
	.w7(32'hbbc46a10),
	.w8(32'hbc466094),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36c9da),
	.w1(32'h3b646d71),
	.w2(32'h39e524c2),
	.w3(32'hbc96b29f),
	.w4(32'hbbbd42ef),
	.w5(32'hbb30c0d6),
	.w6(32'hbc6908ab),
	.w7(32'hbb8c0097),
	.w8(32'hbc4d4421),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule