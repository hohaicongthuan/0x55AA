module layer_8_featuremap_184(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d7ff8),
	.w1(32'h3c992db1),
	.w2(32'h3c480e83),
	.w3(32'h3a483afd),
	.w4(32'h3bf6bc28),
	.w5(32'h3c862563),
	.w6(32'h3ba4df85),
	.w7(32'hbc065936),
	.w8(32'hbb2b6657),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be09352),
	.w1(32'hbb562627),
	.w2(32'hbbe89a29),
	.w3(32'h3c7b6a93),
	.w4(32'hbb94d6a2),
	.w5(32'hbb686902),
	.w6(32'hba72b09e),
	.w7(32'hbb327067),
	.w8(32'hb91736e1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6646e),
	.w1(32'hbccc7ecd),
	.w2(32'hbd23aebd),
	.w3(32'hbb698c4f),
	.w4(32'hbcbce064),
	.w5(32'hbd1518be),
	.w6(32'hbc95df75),
	.w7(32'hbcadfd05),
	.w8(32'hbc8ab613),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf19201),
	.w1(32'h3bb8262c),
	.w2(32'hbbe4c876),
	.w3(32'hbce4cf52),
	.w4(32'hba80cc1d),
	.w5(32'hba4b140f),
	.w6(32'hbc469cee),
	.w7(32'hbc177c9a),
	.w8(32'h3b9517e6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc838e8d),
	.w1(32'hbb71cb14),
	.w2(32'h3b0ae0f4),
	.w3(32'hbc1dc980),
	.w4(32'hbb0d5dbc),
	.w5(32'h3b03717c),
	.w6(32'h3aa93606),
	.w7(32'h3b910072),
	.w8(32'h3ba9652f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c7a53),
	.w1(32'h3c803c98),
	.w2(32'h3d12e4e6),
	.w3(32'hba5b2a4e),
	.w4(32'h3c932710),
	.w5(32'h3ce545dd),
	.w6(32'hbb2a84ca),
	.w7(32'h3c8fd4c9),
	.w8(32'h3d136b09),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b175c25),
	.w1(32'h3bc6349e),
	.w2(32'h3c08e08e),
	.w3(32'hbbc7e565),
	.w4(32'h3bb0937d),
	.w5(32'h3c085e8c),
	.w6(32'h3b32b2bd),
	.w7(32'h3bbd2bf4),
	.w8(32'h3c01770f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ea6ac),
	.w1(32'hbac34629),
	.w2(32'h3c66e0a8),
	.w3(32'h3b39868b),
	.w4(32'hbbb42af5),
	.w5(32'h3c89eb9e),
	.w6(32'hbc89e971),
	.w7(32'hbca99234),
	.w8(32'hbbd2f520),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b720483),
	.w1(32'hbc6f2f13),
	.w2(32'hbc60f967),
	.w3(32'h3b3520ca),
	.w4(32'hbc8cd07c),
	.w5(32'hbc55e67c),
	.w6(32'hbc28411d),
	.w7(32'hbc147b5f),
	.w8(32'hbbea3de8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4aa81),
	.w1(32'hbbff259c),
	.w2(32'hbc71132c),
	.w3(32'h39f98c20),
	.w4(32'hbc2a8071),
	.w5(32'hbb72a963),
	.w6(32'hbaae74aa),
	.w7(32'hbc82af76),
	.w8(32'hbae4e74b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18794c),
	.w1(32'h3bbe033b),
	.w2(32'h3c34ca0b),
	.w3(32'hbc4afa5b),
	.w4(32'h3bba31ef),
	.w5(32'h3c3b4076),
	.w6(32'h3c0bd6b9),
	.w7(32'hbabdedac),
	.w8(32'h3b9314d2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6db674),
	.w1(32'h3c16f5c2),
	.w2(32'h3bdbfffa),
	.w3(32'h3c278515),
	.w4(32'hbab32c0c),
	.w5(32'h3ab857fc),
	.w6(32'hba207dcc),
	.w7(32'hbb9374d7),
	.w8(32'h3c2b1fc0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d6656),
	.w1(32'h3c10b87f),
	.w2(32'h3ade7edf),
	.w3(32'h3b10564d),
	.w4(32'h3bcd19b1),
	.w5(32'h3c8015d7),
	.w6(32'hbb8a4a99),
	.w7(32'hbb6fdd18),
	.w8(32'h3b2903c8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82466b),
	.w1(32'hbc6b426a),
	.w2(32'hbce8fc5e),
	.w3(32'h3bc6c9d3),
	.w4(32'hbc67b38b),
	.w5(32'hbce22a87),
	.w6(32'hbc94e228),
	.w7(32'hbca6685a),
	.w8(32'hbb822854),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc808b59),
	.w1(32'h3be6f6f4),
	.w2(32'h3bb3ff3c),
	.w3(32'hbcbf557e),
	.w4(32'h3b8cdc2c),
	.w5(32'h3b6f909f),
	.w6(32'h3a68c683),
	.w7(32'h3b549715),
	.w8(32'h3b3a653d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b180403),
	.w1(32'h3c6a4440),
	.w2(32'h3aedef21),
	.w3(32'h3a89d12f),
	.w4(32'h3c52c6c5),
	.w5(32'h3b91098a),
	.w6(32'h398ba864),
	.w7(32'h3ba75982),
	.w8(32'h3c110246),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8320f9),
	.w1(32'h3cb26a0f),
	.w2(32'h3c9ddb54),
	.w3(32'h3beeba4c),
	.w4(32'h3c1234d9),
	.w5(32'h3cc56e91),
	.w6(32'h3c2629fa),
	.w7(32'h3c3507c6),
	.w8(32'h3c059d1d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c524120),
	.w1(32'hbb03e835),
	.w2(32'hbc97d59f),
	.w3(32'h3b16fa84),
	.w4(32'hbbec2b0a),
	.w5(32'hbb081953),
	.w6(32'hbc72c28c),
	.w7(32'hbbdad80b),
	.w8(32'hbb357f83),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb866402),
	.w1(32'h3ca10ae3),
	.w2(32'h3c5acd2c),
	.w3(32'hbc4c8711),
	.w4(32'h3cd356cb),
	.w5(32'h3c96c0c7),
	.w6(32'h3b9e77d3),
	.w7(32'hbd2c8743),
	.w8(32'h39f920ef),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8611b),
	.w1(32'h3af709df),
	.w2(32'h3bd78839),
	.w3(32'hbc7c1e37),
	.w4(32'hbc5d16c7),
	.w5(32'hbaa46227),
	.w6(32'hbbda2ec1),
	.w7(32'hba02ac2b),
	.w8(32'h3b9ea374),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b427fdf),
	.w1(32'h3b96c812),
	.w2(32'h3ca39c93),
	.w3(32'hbaec5e8d),
	.w4(32'h3c2aac53),
	.w5(32'h3c81db29),
	.w6(32'h3c5d587d),
	.w7(32'h3cc679f5),
	.w8(32'h3c31ca92),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafa788),
	.w1(32'h3c38d3e6),
	.w2(32'h3d211717),
	.w3(32'h3b914240),
	.w4(32'h3c6605d8),
	.w5(32'h3ce84448),
	.w6(32'h3c1ffdfd),
	.w7(32'h3c3054aa),
	.w8(32'h3beec8a8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed0e51),
	.w1(32'hbd0261d2),
	.w2(32'hbd11fd4b),
	.w3(32'hbb403dc1),
	.w4(32'hbcc5aedb),
	.w5(32'hbc85c90c),
	.w6(32'hbc85f87f),
	.w7(32'hbd2e6be0),
	.w8(32'hbccf71f2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994b438),
	.w1(32'h3ca887bc),
	.w2(32'h3d3c7193),
	.w3(32'hbbff14b7),
	.w4(32'h3c433c63),
	.w5(32'h3d06ad1f),
	.w6(32'h3c126091),
	.w7(32'h3d017e78),
	.w8(32'h3cbecb46),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd75b59),
	.w1(32'h389d0b4f),
	.w2(32'h3b8af9ff),
	.w3(32'h3c827a9e),
	.w4(32'hbb5aa2ec),
	.w5(32'hb94c52ee),
	.w6(32'hba2a8219),
	.w7(32'h3bd6eb78),
	.w8(32'h3bea3b5d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa43ccd),
	.w1(32'hbb5ad216),
	.w2(32'hba5097b4),
	.w3(32'hbc5bb6ca),
	.w4(32'hbb82077c),
	.w5(32'h3c2188f1),
	.w6(32'hbb48d42e),
	.w7(32'hbc80ad56),
	.w8(32'hbca43ed7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b2fdc),
	.w1(32'hbbb557bd),
	.w2(32'hbc3c6e31),
	.w3(32'h3c779af4),
	.w4(32'hba29e2e8),
	.w5(32'hbc8aefc9),
	.w6(32'hbbe2bb53),
	.w7(32'hbc0603e9),
	.w8(32'h3b87b94b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc862bcd),
	.w1(32'hbcca8fc8),
	.w2(32'h3d794140),
	.w3(32'hbda208ff),
	.w4(32'h3c342ad8),
	.w5(32'h3e1681b3),
	.w6(32'h3dd99692),
	.w7(32'h3ccce68d),
	.w8(32'hbbade2ab),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08ff09),
	.w1(32'h3b907286),
	.w2(32'h3c690a84),
	.w3(32'h3b263e6b),
	.w4(32'hbbedb083),
	.w5(32'h3a6e1ce4),
	.w6(32'hbbdab236),
	.w7(32'hbb46c723),
	.w8(32'h3956664d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9153ad),
	.w1(32'h3b1041ff),
	.w2(32'h3c2d9d5a),
	.w3(32'h3aa427d8),
	.w4(32'h3b7b5263),
	.w5(32'h3c40e898),
	.w6(32'h3af629d2),
	.w7(32'h3bf50131),
	.w8(32'h3c6d15ba),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ba644),
	.w1(32'hbb2c8484),
	.w2(32'h3b57053f),
	.w3(32'h3c6e30c5),
	.w4(32'h39fe7ee8),
	.w5(32'h3ae183f7),
	.w6(32'hbba05b33),
	.w7(32'h3b1316cf),
	.w8(32'hbba7b53f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3aef77),
	.w1(32'hbb80a329),
	.w2(32'h3a669db2),
	.w3(32'hbbbe6b7a),
	.w4(32'h3c2da49b),
	.w5(32'h3bb8d528),
	.w6(32'hbaa8b074),
	.w7(32'h3baa20ef),
	.w8(32'h3c42144f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cb970),
	.w1(32'hbb66912f),
	.w2(32'hbc249b66),
	.w3(32'hba84b6d3),
	.w4(32'hbafae861),
	.w5(32'hbc00fa37),
	.w6(32'h3b6c6008),
	.w7(32'hbb45cee5),
	.w8(32'h3c07d70e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3392a6),
	.w1(32'h3c4e9364),
	.w2(32'h3d2362ff),
	.w3(32'hbbdc50f9),
	.w4(32'h3b72cca0),
	.w5(32'h3ca8ee46),
	.w6(32'h3ca69861),
	.w7(32'h3c8f766e),
	.w8(32'hbb0111a8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc9551e),
	.w1(32'h39cfad1d),
	.w2(32'hbb506482),
	.w3(32'h3d09ddd6),
	.w4(32'h3bb3e449),
	.w5(32'hbb1be8cc),
	.w6(32'h3b1f8c8d),
	.w7(32'h3b3e84e2),
	.w8(32'h3c107a57),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b3b58),
	.w1(32'h3b9582a9),
	.w2(32'hbc468bed),
	.w3(32'hbc3f924d),
	.w4(32'hbb1880bc),
	.w5(32'hbbd66166),
	.w6(32'h3b3132f6),
	.w7(32'h3ba0805f),
	.w8(32'h3c07a129),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84a6ce),
	.w1(32'hbb6280ba),
	.w2(32'hbaee9da8),
	.w3(32'hbc6bc0b4),
	.w4(32'hba4ce554),
	.w5(32'hb9b3c51e),
	.w6(32'hbba1deb6),
	.w7(32'hbbadc868),
	.w8(32'hbb4cb788),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bb349),
	.w1(32'hbaf954e5),
	.w2(32'hbbb661a3),
	.w3(32'hbaf86e51),
	.w4(32'hbbb29e94),
	.w5(32'hbbbce385),
	.w6(32'hbb7377a8),
	.w7(32'hbbbd59c6),
	.w8(32'hbb8656e9),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb935ef08),
	.w1(32'h3bda2a34),
	.w2(32'hbbe80551),
	.w3(32'hbb284c8d),
	.w4(32'h3b9e8c4f),
	.w5(32'h3b6c8793),
	.w6(32'h3bc8d131),
	.w7(32'h3acf203d),
	.w8(32'h3acf4402),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae5926),
	.w1(32'h3c2d7ae2),
	.w2(32'h3cfcf184),
	.w3(32'h3bc863cc),
	.w4(32'h3c311176),
	.w5(32'h3ca9c0db),
	.w6(32'h3ba3578f),
	.w7(32'h3c4459ba),
	.w8(32'h3c89fa92),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d02a3f2),
	.w1(32'h3aae304c),
	.w2(32'h3c875988),
	.w3(32'h3a2e4ac9),
	.w4(32'hbcefb990),
	.w5(32'h3b8d58b0),
	.w6(32'hbcb7369e),
	.w7(32'hbcb880bd),
	.w8(32'h3c044e58),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b3aa8),
	.w1(32'h3be9c55e),
	.w2(32'h3b2d48be),
	.w3(32'hbc222520),
	.w4(32'h3c795bd2),
	.w5(32'h3bca4011),
	.w6(32'h3ba3c5cd),
	.w7(32'h3a63c7de),
	.w8(32'h3b841a64),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c147883),
	.w1(32'hba77a6d8),
	.w2(32'h3bfdb267),
	.w3(32'h3bc5ed86),
	.w4(32'hbaf084b2),
	.w5(32'h3b91e20d),
	.w6(32'h3b936a8f),
	.w7(32'h3bc0f58a),
	.w8(32'h3c0b3fac),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8aa358),
	.w1(32'hbb6f5606),
	.w2(32'hbcdd2569),
	.w3(32'hbb1d855c),
	.w4(32'h3b1d964e),
	.w5(32'hbbf21326),
	.w6(32'hbc7135a3),
	.w7(32'hbc88365e),
	.w8(32'hbc0c541e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf675e),
	.w1(32'h3c73a925),
	.w2(32'h3c31da55),
	.w3(32'hbcecf765),
	.w4(32'h3c9895c1),
	.w5(32'h3c27f2fb),
	.w6(32'h3c1c3b6c),
	.w7(32'hbc2a0afa),
	.w8(32'h3ac3465a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9913f5e),
	.w1(32'h3ad86411),
	.w2(32'h3b94f9ee),
	.w3(32'h3b1b42f0),
	.w4(32'h3b30509d),
	.w5(32'h3ba6d7b6),
	.w6(32'hbbc7061f),
	.w7(32'hbb6a3ea8),
	.w8(32'h3b3624c3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f969a),
	.w1(32'h3c935924),
	.w2(32'h3cec37b6),
	.w3(32'hbab75e39),
	.w4(32'h3c868c52),
	.w5(32'h3cce9ed4),
	.w6(32'h3c3cfead),
	.w7(32'h3cbc5336),
	.w8(32'h3cbc696c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caeb4f1),
	.w1(32'h3a12cf06),
	.w2(32'h3a789f16),
	.w3(32'h3c8b4a7f),
	.w4(32'h3c224f85),
	.w5(32'h3c06dbf5),
	.w6(32'h3b28e312),
	.w7(32'hbbfbfc4e),
	.w8(32'hbbb2b50d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d275b),
	.w1(32'hbb220870),
	.w2(32'hbc3a64f2),
	.w3(32'h3bc5e685),
	.w4(32'hbbb2751c),
	.w5(32'hbbb58d09),
	.w6(32'hbbf79b77),
	.w7(32'hbbfa737c),
	.w8(32'hbb607b38),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7eafa1),
	.w1(32'h3c173cc1),
	.w2(32'h3cb8624b),
	.w3(32'hbb310fbf),
	.w4(32'h3bda4fa8),
	.w5(32'h3c8a112c),
	.w6(32'h3b550680),
	.w7(32'h3a8b1a1f),
	.w8(32'h383e6cc2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c5751),
	.w1(32'h3c74ef48),
	.w2(32'h3c5f3f79),
	.w3(32'h3ca17f23),
	.w4(32'h3c20d9d5),
	.w5(32'h3c5d532f),
	.w6(32'hbb849f38),
	.w7(32'h3b45b1ff),
	.w8(32'h3c99090d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9629c6),
	.w1(32'h3c11cb50),
	.w2(32'h3cbccfae),
	.w3(32'hba6d881c),
	.w4(32'h3c63cb01),
	.w5(32'h3cb7d5f6),
	.w6(32'hbc85b0f5),
	.w7(32'hbcc3f6da),
	.w8(32'h3c214d21),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b4dde),
	.w1(32'hbbd9a518),
	.w2(32'hbaeb4c22),
	.w3(32'hbc052b7a),
	.w4(32'hbc070486),
	.w5(32'hba95fac4),
	.w6(32'hbbcbee48),
	.w7(32'hbb7175ff),
	.w8(32'h3af97393),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68504a),
	.w1(32'h3bf09550),
	.w2(32'hbbb296ab),
	.w3(32'hbb489aa7),
	.w4(32'hbc78c450),
	.w5(32'hbc227930),
	.w6(32'hbbbd69da),
	.w7(32'hbc2f8119),
	.w8(32'hbc4886ee),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb085a9),
	.w1(32'h3ab53a24),
	.w2(32'h3b05bef4),
	.w3(32'h3b88344b),
	.w4(32'hbbaeaa9e),
	.w5(32'hbbdc70f2),
	.w6(32'hbb8f7a8b),
	.w7(32'hba147f35),
	.w8(32'h3bf5bf53),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28f8aa),
	.w1(32'h3c8698e5),
	.w2(32'h3c80c857),
	.w3(32'hbb890b00),
	.w4(32'h3bee9075),
	.w5(32'h3cb3fe6c),
	.w6(32'h3bcb4185),
	.w7(32'hbba601e2),
	.w8(32'hbb3d3fc5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17a194),
	.w1(32'h3be93a2b),
	.w2(32'h3beb2188),
	.w3(32'h3c54ec19),
	.w4(32'h3c61213e),
	.w5(32'h3ba45e4c),
	.w6(32'h3b871127),
	.w7(32'h3bd8e615),
	.w8(32'h3c496e92),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43c6b4),
	.w1(32'h3aa8baa3),
	.w2(32'h3c620ec3),
	.w3(32'hbb842c87),
	.w4(32'h3c0c07ad),
	.w5(32'h3c341b98),
	.w6(32'hbc0b7431),
	.w7(32'hbbdb74ad),
	.w8(32'h3c0da6ca),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86c40fa),
	.w1(32'hbb796e9d),
	.w2(32'hbab5dd95),
	.w3(32'h3aab5adb),
	.w4(32'h3b2f7cba),
	.w5(32'h3b413880),
	.w6(32'h3b254e2a),
	.w7(32'hb7189bf0),
	.w8(32'hbbb05698),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11c5f8),
	.w1(32'h3cb2ef0a),
	.w2(32'h3d217bcb),
	.w3(32'h3bf64ff5),
	.w4(32'h3cc1adb1),
	.w5(32'h3d193d78),
	.w6(32'h3c9bd103),
	.w7(32'h3cbebdba),
	.w8(32'h3bfbd613),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cbe1f),
	.w1(32'hbbfc56e2),
	.w2(32'hbbac7079),
	.w3(32'h3c6bd08c),
	.w4(32'hbab71f25),
	.w5(32'hbbc63198),
	.w6(32'h3b40b123),
	.w7(32'h3c0c243b),
	.w8(32'h3b967c7f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b9afb),
	.w1(32'h3afd098f),
	.w2(32'h3c4be6fb),
	.w3(32'hbafff0ad),
	.w4(32'h3b8f7908),
	.w5(32'h3c7be76f),
	.w6(32'hbbc6a91e),
	.w7(32'hba441fd7),
	.w8(32'hbaadf5c1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fec13),
	.w1(32'h3c0230ac),
	.w2(32'h3c3f8dc1),
	.w3(32'h3b8bcf54),
	.w4(32'hbcbc103c),
	.w5(32'hbbb1c7d0),
	.w6(32'hbc3d8ddc),
	.w7(32'hbc5b6725),
	.w8(32'hbb0a9706),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1639a1),
	.w1(32'h3b9c5583),
	.w2(32'h3bc2dbac),
	.w3(32'hbb291a8c),
	.w4(32'h3b83f693),
	.w5(32'h3b884a3a),
	.w6(32'h3be199f1),
	.w7(32'h3b2bcd8a),
	.w8(32'h3bce300e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b173b46),
	.w1(32'h3af8a910),
	.w2(32'h3a16fa16),
	.w3(32'h3af1b249),
	.w4(32'h3ac205c5),
	.w5(32'hba76927f),
	.w6(32'hb995022d),
	.w7(32'hb9957094),
	.w8(32'hbac6f487),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf1c65),
	.w1(32'h3b9bd614),
	.w2(32'h3cbb5251),
	.w3(32'hbb3a9052),
	.w4(32'h3c21571d),
	.w5(32'h3d0e6b11),
	.w6(32'h3b004732),
	.w7(32'h3c024e3a),
	.w8(32'h3bb96426),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f2595),
	.w1(32'h3c955aae),
	.w2(32'h3c234d16),
	.w3(32'h3c2fabf8),
	.w4(32'hbb6206ee),
	.w5(32'h3b8475cb),
	.w6(32'h3b77cf5e),
	.w7(32'h3b85a663),
	.w8(32'h3b619c13),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b8643c),
	.w1(32'h3c94891c),
	.w2(32'h3cb50488),
	.w3(32'hbaa17104),
	.w4(32'h3c164905),
	.w5(32'h3cb0b752),
	.w6(32'h3b68d9b8),
	.w7(32'h3c6470e6),
	.w8(32'h3c93512d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e97e6),
	.w1(32'h3cf48627),
	.w2(32'h3d602aa3),
	.w3(32'h3c06a546),
	.w4(32'h3ca57857),
	.w5(32'h3d2058a2),
	.w6(32'h3cb849c1),
	.w7(32'h3ce4df5b),
	.w8(32'h3c44d1bb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc43500),
	.w1(32'hbd1ac64b),
	.w2(32'hbd00cdef),
	.w3(32'h3ce5c4be),
	.w4(32'h3bd49098),
	.w5(32'h38513bc5),
	.w6(32'h3bcf1e1b),
	.w7(32'hbc99dceb),
	.w8(32'hbd22bccb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc51114),
	.w1(32'h3b8a83db),
	.w2(32'h3c25d2ae),
	.w3(32'hbcaf128d),
	.w4(32'hbaa524f8),
	.w5(32'h3b95dfe6),
	.w6(32'hb84c255e),
	.w7(32'h3c1cb1e9),
	.w8(32'hba8ddd62),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd371ca),
	.w1(32'hbcc9da93),
	.w2(32'hbd395465),
	.w3(32'hbbdc336f),
	.w4(32'hbcda5a31),
	.w5(32'hbd2a3ff9),
	.w6(32'hbc5dc92b),
	.w7(32'hbc9c5683),
	.w8(32'hba8c1ae5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd07a6a4),
	.w1(32'hbc701e42),
	.w2(32'hbd28cd1e),
	.w3(32'hbd0d5372),
	.w4(32'hbcaa09f3),
	.w5(32'hbd1ad657),
	.w6(32'hbc65fec3),
	.w7(32'hbc623494),
	.w8(32'hbb32cc08),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd8e00b),
	.w1(32'hbc0ae603),
	.w2(32'hbb5b6489),
	.w3(32'hbcde4c2d),
	.w4(32'hbbe844d6),
	.w5(32'h3b86f345),
	.w6(32'hbc40e2f2),
	.w7(32'hbba9c4f3),
	.w8(32'hbb0db957),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1ee99),
	.w1(32'hbb37df4c),
	.w2(32'hbb953040),
	.w3(32'hbb4d5100),
	.w4(32'hbb86362c),
	.w5(32'hbb7b51b0),
	.w6(32'hbb469a3e),
	.w7(32'hb9b404b8),
	.w8(32'h3b63420c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e82c9),
	.w1(32'hbc2da712),
	.w2(32'hbc2c0338),
	.w3(32'hbb805033),
	.w4(32'hbc0f2084),
	.w5(32'hbbdfabb1),
	.w6(32'hbac72d92),
	.w7(32'hbba90f8c),
	.w8(32'h3b8a9540),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7cd98),
	.w1(32'hbb6fa3dd),
	.w2(32'h3b1f1025),
	.w3(32'hbc31c7dd),
	.w4(32'h3ab9d946),
	.w5(32'hb915e191),
	.w6(32'hbac05ad0),
	.w7(32'h3acf6686),
	.w8(32'h3c325b1a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44962d),
	.w1(32'h3b969691),
	.w2(32'h3c179afd),
	.w3(32'hbbe84921),
	.w4(32'h3c1fd7d5),
	.w5(32'h3c44f28c),
	.w6(32'h3bc124f0),
	.w7(32'hbc18ca81),
	.w8(32'h3ab18302),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c389fc9),
	.w1(32'h3c3aa711),
	.w2(32'h3bf729aa),
	.w3(32'h3bf5cbdd),
	.w4(32'h3bd1c14e),
	.w5(32'h3b3bfb3c),
	.w6(32'h3b61a851),
	.w7(32'h3b41c9d9),
	.w8(32'hbb321223),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b612eb3),
	.w1(32'h3a8e3e00),
	.w2(32'h3c05d438),
	.w3(32'hbafcef04),
	.w4(32'h3b705a80),
	.w5(32'h3bb503af),
	.w6(32'hb9bc9ce4),
	.w7(32'h3b6eb6a0),
	.w8(32'h3bc415f2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef1822),
	.w1(32'hbc24aa3d),
	.w2(32'hbd18642d),
	.w3(32'h3b2c4dcc),
	.w4(32'hbc3edb9d),
	.w5(32'hbcfea4cd),
	.w6(32'hbbf19b4c),
	.w7(32'hbc72e2d6),
	.w8(32'hbb952408),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc62074),
	.w1(32'h3c43b0da),
	.w2(32'h3cd09b68),
	.w3(32'hbc80e7f9),
	.w4(32'h3c888b01),
	.w5(32'h3cbe73c0),
	.w6(32'h3c878b6c),
	.w7(32'h3ce6a088),
	.w8(32'h3c1224ac),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4c446),
	.w1(32'hbbbb23b6),
	.w2(32'hbbfc71fb),
	.w3(32'h3c528e16),
	.w4(32'hbb513bcb),
	.w5(32'hba25e375),
	.w6(32'hbbb15372),
	.w7(32'hbc68342a),
	.w8(32'hbbb5c5c2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a59ea),
	.w1(32'h3d249bdc),
	.w2(32'h3d4f870d),
	.w3(32'hbb127fcf),
	.w4(32'h3cd82ffc),
	.w5(32'h3c534918),
	.w6(32'hbcc1ed16),
	.w7(32'h36423520),
	.w8(32'h3d4b8c2a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c8558),
	.w1(32'hbc813df7),
	.w2(32'hbc471d24),
	.w3(32'hbc8f1dba),
	.w4(32'hbcba3b67),
	.w5(32'hbc6025d0),
	.w6(32'hbc4bd0b0),
	.w7(32'hbce66917),
	.w8(32'hbc1e68bf),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa567a3),
	.w1(32'hbbc15966),
	.w2(32'hbc080000),
	.w3(32'hbc6dffa9),
	.w4(32'hbae0c391),
	.w5(32'hbc171a44),
	.w6(32'h3b0936ac),
	.w7(32'hbb8dfc7d),
	.w8(32'h3ba5eb43),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd6c13),
	.w1(32'hbba90ee4),
	.w2(32'hba1cf9da),
	.w3(32'hbb9d4df0),
	.w4(32'hbb89fcfc),
	.w5(32'hbbabe226),
	.w6(32'hb94f896e),
	.w7(32'hbadb2309),
	.w8(32'hba8d8e7e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b4223),
	.w1(32'hbb0584f2),
	.w2(32'h3b8d3bdd),
	.w3(32'hbb5fc443),
	.w4(32'hbbb18698),
	.w5(32'h3b532a4d),
	.w6(32'hba05e5d6),
	.w7(32'h3b2c26ba),
	.w8(32'hb9f2121c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968c3a2),
	.w1(32'hbbb0f6e8),
	.w2(32'hbad2e282),
	.w3(32'h3abf43a1),
	.w4(32'h3ad5d49d),
	.w5(32'hbb57bde5),
	.w6(32'hbb1257d6),
	.w7(32'hbb0602c5),
	.w8(32'hbaa6d022),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03ddcd),
	.w1(32'hbc863470),
	.w2(32'hbcfc1a20),
	.w3(32'hba15913b),
	.w4(32'hbb8c70ef),
	.w5(32'hbcdf6ee1),
	.w6(32'hbc5d6c4f),
	.w7(32'hbca1ca26),
	.w8(32'hbc6f4c4c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc58069),
	.w1(32'hbc51d7e6),
	.w2(32'hbd1c51ac),
	.w3(32'hbcb99b28),
	.w4(32'hbc81c3a1),
	.w5(32'hbd0e5a26),
	.w6(32'h3adcbb34),
	.w7(32'hba9c7a9a),
	.w8(32'h3c2165d0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce39ff0),
	.w1(32'h3c130b40),
	.w2(32'h3cd8cccf),
	.w3(32'hbd04a394),
	.w4(32'h3bb66b1e),
	.w5(32'h3c3456de),
	.w6(32'h3c612764),
	.w7(32'h3c4fc007),
	.w8(32'h3c06805c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c758b8f),
	.w1(32'hbadf7495),
	.w2(32'h3bd962ac),
	.w3(32'h3ca3e77c),
	.w4(32'h3aaf0310),
	.w5(32'h3b6d76e5),
	.w6(32'hbb5d6fab),
	.w7(32'h39af8a68),
	.w8(32'h3b91a409),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88c900),
	.w1(32'h3b247dc5),
	.w2(32'h3c10bcb9),
	.w3(32'hbb46344d),
	.w4(32'hbb09af23),
	.w5(32'h3baf7dfb),
	.w6(32'hbb966320),
	.w7(32'hba178f94),
	.w8(32'h3b323d5b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c290372),
	.w1(32'h3bc08bf2),
	.w2(32'h3bc07645),
	.w3(32'h3c054359),
	.w4(32'h3c156ce2),
	.w5(32'h3c187d86),
	.w6(32'h3b756291),
	.w7(32'h3abdd130),
	.w8(32'h3c142639),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ccc83),
	.w1(32'h3bd661fb),
	.w2(32'h3c2c0bda),
	.w3(32'h3c10f53b),
	.w4(32'h3bc81a5a),
	.w5(32'h3ba14953),
	.w6(32'h3a9b7e2e),
	.w7(32'h3a861e01),
	.w8(32'h3bc773c0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c0e15),
	.w1(32'hbbda79bd),
	.w2(32'hbc1e8450),
	.w3(32'hbc312ddd),
	.w4(32'hbca0d2b2),
	.w5(32'hbc3e2565),
	.w6(32'hbca6b1c1),
	.w7(32'hbc7de0ec),
	.w8(32'h3b82b046),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f03cd),
	.w1(32'hbbe02d99),
	.w2(32'hbd15399e),
	.w3(32'hbbc63dc6),
	.w4(32'h3bb8e7ef),
	.w5(32'hbc82ad01),
	.w6(32'hbbab444e),
	.w7(32'hbc9acdfe),
	.w8(32'hb9f3eb54),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ed1e3),
	.w1(32'h3bac82d6),
	.w2(32'hbcb47497),
	.w3(32'hbc18a696),
	.w4(32'h3bb06c54),
	.w5(32'hbbeb1ec7),
	.w6(32'h3b3c59a9),
	.w7(32'hbb32f6d0),
	.w8(32'h3b8e72e1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76c86d5),
	.w1(32'hbb0d5987),
	.w2(32'h3b61c188),
	.w3(32'hbb574468),
	.w4(32'hbb2e64fa),
	.w5(32'h3a46169d),
	.w6(32'h3a9a063d),
	.w7(32'h3bd75bb7),
	.w8(32'hba0acfd3),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc09df9),
	.w1(32'h3bddd3fe),
	.w2(32'h39f32d68),
	.w3(32'h3aa29235),
	.w4(32'hbc3ef98a),
	.w5(32'hbbc8623a),
	.w6(32'h3c1f8054),
	.w7(32'h3c277dfe),
	.w8(32'h3b8f380a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a0c9c),
	.w1(32'hbc43259f),
	.w2(32'hbc91f999),
	.w3(32'h3bf6b75c),
	.w4(32'hbaf83367),
	.w5(32'hbc156f3b),
	.w6(32'hbc10b23d),
	.w7(32'hbc776fc8),
	.w8(32'hbb739aac),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00f0d9),
	.w1(32'hbbdf551c),
	.w2(32'hbc533660),
	.w3(32'hbb919fd1),
	.w4(32'hbb7a3e2c),
	.w5(32'hbc67c3f2),
	.w6(32'h3940b04e),
	.w7(32'hbaff5289),
	.w8(32'hbab802a2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc331adb),
	.w1(32'hbc991a8a),
	.w2(32'hbc285e5b),
	.w3(32'hbca39977),
	.w4(32'hbc1875d5),
	.w5(32'hbb21e10b),
	.w6(32'hbc11563e),
	.w7(32'h39acd207),
	.w8(32'h3b354ac4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ae6cb),
	.w1(32'hbacda779),
	.w2(32'hbba5798f),
	.w3(32'hbbad0abc),
	.w4(32'h3c47ffbc),
	.w5(32'h3aedf56c),
	.w6(32'h3c272dc1),
	.w7(32'h3bdf201f),
	.w8(32'h3bc20664),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea8db9),
	.w1(32'hbc484487),
	.w2(32'hb9fbff2d),
	.w3(32'hbc193e96),
	.w4(32'hbaabe21d),
	.w5(32'h3c2bd62c),
	.w6(32'hbab0634b),
	.w7(32'hbbf7ce9f),
	.w8(32'hbc5796e3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0557a9),
	.w1(32'hbbc69fce),
	.w2(32'hb9cbff07),
	.w3(32'hbc0277cd),
	.w4(32'hbb9d472b),
	.w5(32'hbbb46105),
	.w6(32'hbb3f2077),
	.w7(32'hbb248f50),
	.w8(32'h3a610811),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d3697),
	.w1(32'hbc54e9c5),
	.w2(32'hbadaca55),
	.w3(32'hbaa4e01f),
	.w4(32'hbc04353d),
	.w5(32'hbbf16e29),
	.w6(32'hbbddbe9b),
	.w7(32'hba246320),
	.w8(32'hba58793e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc54dc1),
	.w1(32'hbb3c84b8),
	.w2(32'h3c2192d1),
	.w3(32'hbbaad8b9),
	.w4(32'hbc1ca943),
	.w5(32'hbac60f37),
	.w6(32'hbb217609),
	.w7(32'h3b8015ae),
	.w8(32'h3b022bfb),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba56739),
	.w1(32'hbbe57e52),
	.w2(32'hbb896351),
	.w3(32'hbaf4668f),
	.w4(32'hbbe0e489),
	.w5(32'hbb61ba41),
	.w6(32'hbb402231),
	.w7(32'hbb3fce42),
	.w8(32'hbba881da),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1705d8),
	.w1(32'h3b196380),
	.w2(32'h3b459a3b),
	.w3(32'h3aec3085),
	.w4(32'hbc48611f),
	.w5(32'hbbae0797),
	.w6(32'h398ebb4c),
	.w7(32'h3a9e2fc6),
	.w8(32'h3c3f165f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc16937),
	.w1(32'h3c0a121a),
	.w2(32'h3c8a21b1),
	.w3(32'hbc34b44a),
	.w4(32'h3b998ad2),
	.w5(32'h3c429ebc),
	.w6(32'h3b5d7cde),
	.w7(32'h3bc2808c),
	.w8(32'h3c39c7ff),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a02cd),
	.w1(32'hb9a72d28),
	.w2(32'h3ae71ab2),
	.w3(32'h39fef9e0),
	.w4(32'h3c0a758b),
	.w5(32'h3b04884d),
	.w6(32'h3c35ba45),
	.w7(32'h3b386a3f),
	.w8(32'h3bcc4c5f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97acfc),
	.w1(32'hbc14edc1),
	.w2(32'hbcf41147),
	.w3(32'h3bc5a20d),
	.w4(32'hbb84ccd7),
	.w5(32'hbc73e982),
	.w6(32'hbbfaff3f),
	.w7(32'hbc32a679),
	.w8(32'hbc6b018d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52030a),
	.w1(32'hbbb108b3),
	.w2(32'hbb8b45be),
	.w3(32'hbc617afc),
	.w4(32'h3b0cb7cb),
	.w5(32'hbc143081),
	.w6(32'hbbd9df37),
	.w7(32'hbbadf86e),
	.w8(32'hbb140fe7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb052f60),
	.w1(32'hbb8aa298),
	.w2(32'hbb3fd4d8),
	.w3(32'hbba34e49),
	.w4(32'hbb4a473f),
	.w5(32'hba411b27),
	.w6(32'hb9ca0671),
	.w7(32'hbaf1fea7),
	.w8(32'hb9f0e41f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab63921),
	.w1(32'hbb932621),
	.w2(32'hbba08040),
	.w3(32'hbb47fd5f),
	.w4(32'hbc348935),
	.w5(32'hbc219407),
	.w6(32'hbc35309c),
	.w7(32'hbbe1f621),
	.w8(32'hbb59dfa1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb882ed7),
	.w1(32'h3c0435f5),
	.w2(32'h3c6cce0a),
	.w3(32'hbc1e8a55),
	.w4(32'h3be52883),
	.w5(32'h3c4a6f59),
	.w6(32'h3c189430),
	.w7(32'hbba40c66),
	.w8(32'hb8cf52bc),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba647f),
	.w1(32'hbb63d2f2),
	.w2(32'h3b5220a6),
	.w3(32'h3b948680),
	.w4(32'hbaab826e),
	.w5(32'hbacabbaa),
	.w6(32'hbc4abc82),
	.w7(32'hbc3a2700),
	.w8(32'hbc7941d7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19c18d),
	.w1(32'h3b2ca6ca),
	.w2(32'hbb215c74),
	.w3(32'hbb1749eb),
	.w4(32'h3a11482e),
	.w5(32'hbad0ec2a),
	.w6(32'hbbb334bd),
	.w7(32'hba881921),
	.w8(32'h3ba2466c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57f0fd),
	.w1(32'h3d152e14),
	.w2(32'h3d847673),
	.w3(32'h3c2b7e8f),
	.w4(32'h3c82502f),
	.w5(32'h3d3b5a28),
	.w6(32'h3ce06763),
	.w7(32'h3d2e0aae),
	.w8(32'h3cb9608a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2709de),
	.w1(32'hbb5a42e7),
	.w2(32'h3b8273f9),
	.w3(32'h3cff929e),
	.w4(32'hbae1d0b3),
	.w5(32'hb9e45f59),
	.w6(32'hbb9d127f),
	.w7(32'h3ac79e8b),
	.w8(32'h3a301151),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1658d8),
	.w1(32'h3a460f45),
	.w2(32'h3ad0856d),
	.w3(32'hbb81d448),
	.w4(32'hb8f33d30),
	.w5(32'h3b3919fb),
	.w6(32'h3b7b65f2),
	.w7(32'h3b3a84c8),
	.w8(32'h3aa923b2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27e3e5),
	.w1(32'h3c3ae3a6),
	.w2(32'h3bf8ce93),
	.w3(32'hb9f3698b),
	.w4(32'h3c8bc7b6),
	.w5(32'h3c0d58ce),
	.w6(32'h3c12f147),
	.w7(32'h3b78f099),
	.w8(32'h3c409b07),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a9f58),
	.w1(32'hbc06cf61),
	.w2(32'hbc0d527a),
	.w3(32'h3b8295ff),
	.w4(32'hbbdd80bc),
	.w5(32'hbbb02bde),
	.w6(32'hbb5ed949),
	.w7(32'hbc137b51),
	.w8(32'hbc0221e9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc084a70),
	.w1(32'h3b9fd2e6),
	.w2(32'h3c7cf663),
	.w3(32'hbc46cdfa),
	.w4(32'h3c25aa22),
	.w5(32'h3c3ef38c),
	.w6(32'h3b223118),
	.w7(32'h3bbb32de),
	.w8(32'h3b2306c9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad6cf2),
	.w1(32'h3a97d166),
	.w2(32'h3b3d3632),
	.w3(32'h39b03f26),
	.w4(32'hbb22b013),
	.w5(32'h3b491172),
	.w6(32'hbb1d90b9),
	.w7(32'h3abcf447),
	.w8(32'h3b8e7309),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c44e3),
	.w1(32'h3ca5effb),
	.w2(32'h3c154b48),
	.w3(32'h3b0d1146),
	.w4(32'h3ce41432),
	.w5(32'h3a188662),
	.w6(32'h3bb1956d),
	.w7(32'hb81a285c),
	.w8(32'hbc541fe8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule