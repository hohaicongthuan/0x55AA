module layer_10_featuremap_157(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361fbf3d),
	.w1(32'h35ffdf07),
	.w2(32'h36d14f05),
	.w3(32'h36625700),
	.w4(32'hb347f086),
	.w5(32'hb59a223b),
	.w6(32'hb585308c),
	.w7(32'h358c0227),
	.w8(32'h36070159),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9482036),
	.w1(32'hb76b71a6),
	.w2(32'h3845b015),
	.w3(32'hb9399486),
	.w4(32'hb8c5767a),
	.w5(32'hb8f5d8d6),
	.w6(32'hb96c0be0),
	.w7(32'hb8d4bc23),
	.w8(32'hb92e9c06),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ca3109),
	.w1(32'hb52156b5),
	.w2(32'h369632ec),
	.w3(32'h3565de2b),
	.w4(32'hb5901cf4),
	.w5(32'h366244a4),
	.w6(32'hb59db6c7),
	.w7(32'h35c58521),
	.w8(32'h365c0f65),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb47dd483),
	.w1(32'hb6f6ebcf),
	.w2(32'h36a0e3ff),
	.w3(32'hb63f3aa8),
	.w4(32'hb645d8e1),
	.w5(32'h373b3bb6),
	.w6(32'hb6ac62ae),
	.w7(32'h35b476dd),
	.w8(32'h370eae1e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b81466),
	.w1(32'h36b24925),
	.w2(32'hb5fcfc97),
	.w3(32'h36df9d1f),
	.w4(32'h36577fce),
	.w5(32'h31e18c6f),
	.w6(32'h376d93ef),
	.w7(32'h3693f633),
	.w8(32'h35c7d976),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363fb1e3),
	.w1(32'h3617f296),
	.w2(32'h34170417),
	.w3(32'h361518ef),
	.w4(32'h355591fb),
	.w5(32'h3383232f),
	.w6(32'h36f9534e),
	.w7(32'h35fec2ec),
	.w8(32'h361aca27),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b009a4),
	.w1(32'h380b4c02),
	.w2(32'hb8c322fc),
	.w3(32'h367abb57),
	.w4(32'h38f87588),
	.w5(32'hb715be74),
	.w6(32'h38a8637d),
	.w7(32'h38d3c8fa),
	.w8(32'h3891810b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aae74d),
	.w1(32'h375ff275),
	.w2(32'hb9de811e),
	.w3(32'h39965c7d),
	.w4(32'h37808d80),
	.w5(32'h370d189e),
	.w6(32'h39b6161d),
	.w7(32'h3947fc26),
	.w8(32'h3910dbfe),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aba954),
	.w1(32'h38d83cfb),
	.w2(32'hb7de0e86),
	.w3(32'h38158f3c),
	.w4(32'h38d31ed8),
	.w5(32'h368d89fa),
	.w6(32'h373817df),
	.w7(32'h389d7664),
	.w8(32'h379072ae),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382fd401),
	.w1(32'h388a94d5),
	.w2(32'hba8920f4),
	.w3(32'h3a0ff3b6),
	.w4(32'h3a4831ea),
	.w5(32'hb8aab8b0),
	.w6(32'h3a46eb59),
	.w7(32'h3a7fff41),
	.w8(32'h39fd1469),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373f31cc),
	.w1(32'h38af81ec),
	.w2(32'h389d681e),
	.w3(32'h383c852d),
	.w4(32'h38a8dd12),
	.w5(32'h3884c374),
	.w6(32'h380d0cd9),
	.w7(32'h38a0414f),
	.w8(32'h3798dc98),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f3bdf),
	.w1(32'h390117b3),
	.w2(32'h397f465c),
	.w3(32'hba45445a),
	.w4(32'h39bf80a2),
	.w5(32'h3a253272),
	.w6(32'hba528eba),
	.w7(32'h399226ac),
	.w8(32'h39e74ba9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945f866),
	.w1(32'h390211ee),
	.w2(32'hba8beea1),
	.w3(32'h3a44c957),
	.w4(32'h3a816e91),
	.w5(32'h38ea69d9),
	.w6(32'h3a7fb8a7),
	.w7(32'h3aa45912),
	.w8(32'h3a4eabd2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374518f3),
	.w1(32'h382c1b67),
	.w2(32'h38446457),
	.w3(32'hb8401a0a),
	.w4(32'hb74f817e),
	.w5(32'h3518cde2),
	.w6(32'hb7cc228d),
	.w7(32'h3783f99c),
	.w8(32'hb6150102),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3484a4f8),
	.w1(32'h38760d3e),
	.w2(32'hb9be091d),
	.w3(32'h3912d8ae),
	.w4(32'h39918fa7),
	.w5(32'hb70015c5),
	.w6(32'h38f65679),
	.w7(32'h399385fb),
	.w8(32'hb760cbe3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3808cacb),
	.w1(32'hb944bc0a),
	.w2(32'hba6b8edb),
	.w3(32'h39cceec5),
	.w4(32'h39c86e2b),
	.w5(32'hb9dcbd82),
	.w6(32'h3a107762),
	.w7(32'h3a077441),
	.w8(32'hb69f27e8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e5a7fc),
	.w1(32'h37fd89ab),
	.w2(32'h38088e09),
	.w3(32'h3802ffb9),
	.w4(32'h383e7d0c),
	.w5(32'hb52561a5),
	.w6(32'h381708ce),
	.w7(32'h382d42ed),
	.w8(32'hb796e1aa),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367cbafb),
	.w1(32'hb9512b0a),
	.w2(32'hba930698),
	.w3(32'h39a5200d),
	.w4(32'h3986e16c),
	.w5(32'hb9bb7b05),
	.w6(32'h3a1a2cae),
	.w7(32'h39ed1879),
	.w8(32'h39059afa),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb487d8a1),
	.w1(32'hb8099fa9),
	.w2(32'hba00563e),
	.w3(32'h3948fee8),
	.w4(32'h398817c7),
	.w5(32'h375be4e9),
	.w6(32'h39966616),
	.w7(32'h39ce4721),
	.w8(32'h399c7c79),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363fb7f9),
	.w1(32'hb594e3e3),
	.w2(32'hb494057b),
	.w3(32'h36b146e7),
	.w4(32'hb60e8130),
	.w5(32'hb608e07f),
	.w6(32'h36d0dd5e),
	.w7(32'h32fb8c54),
	.w8(32'h359f4f35),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360fa61a),
	.w1(32'hb705bdd3),
	.w2(32'hb5965ee7),
	.w3(32'h363d353b),
	.w4(32'hb729da9a),
	.w5(32'hb6e3d2e6),
	.w6(32'h34ac5fde),
	.w7(32'hb61a1ff2),
	.w8(32'hb6c8c4cb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86761f7),
	.w1(32'h38788466),
	.w2(32'h383105cb),
	.w3(32'hb890a799),
	.w4(32'h388966f5),
	.w5(32'h3838070c),
	.w6(32'hb8d279ab),
	.w7(32'h384c6c47),
	.w8(32'h381eb143),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba628f59),
	.w1(32'hba49891f),
	.w2(32'hbacab612),
	.w3(32'hba289b93),
	.w4(32'hb9509d78),
	.w5(32'hbaa69e02),
	.w6(32'hba2c7750),
	.w7(32'hb994aa3b),
	.w8(32'hbaaa2a35),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b452cd),
	.w1(32'h3900c2d6),
	.w2(32'hba87113d),
	.w3(32'h39fe4c69),
	.w4(32'h3a2ede3f),
	.w5(32'hb98c96cd),
	.w6(32'h3a172739),
	.w7(32'h3a542ec9),
	.w8(32'h3924fd53),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c98f7),
	.w1(32'hb90b20c6),
	.w2(32'hba31e11b),
	.w3(32'hb9198329),
	.w4(32'h39961aa2),
	.w5(32'hb93ed976),
	.w6(32'hb881498d),
	.w7(32'h39c18bd3),
	.w8(32'hb7cc6a45),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3828a45a),
	.w1(32'h3867ad18),
	.w2(32'h37ccf17d),
	.w3(32'h37c4c3ac),
	.w4(32'h37a9f831),
	.w5(32'h3744e09d),
	.w6(32'h3804639b),
	.w7(32'h371ccc75),
	.w8(32'h371b2dd2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6166d8c),
	.w1(32'hb6722cf1),
	.w2(32'h37336c0f),
	.w3(32'hb69b753b),
	.w4(32'hb7481c84),
	.w5(32'h36052c3e),
	.w6(32'hb61248c7),
	.w7(32'hb704ac15),
	.w8(32'h35989ee4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3cb3d),
	.w1(32'h38d92547),
	.w2(32'h380f36b0),
	.w3(32'hb8f50c3e),
	.w4(32'h396487cf),
	.w5(32'h39b95253),
	.w6(32'hb8b61151),
	.w7(32'h39404ddc),
	.w8(32'h39c0f912),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba224614),
	.w1(32'hb9aa5451),
	.w2(32'h38dbb3ac),
	.w3(32'hba13f048),
	.w4(32'hb99ef6a0),
	.w5(32'h3844aa26),
	.w6(32'hba249cf0),
	.w7(32'hb9c255e7),
	.w8(32'hb7c1313c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3827f34c),
	.w1(32'h392fb42f),
	.w2(32'hb9a86ea9),
	.w3(32'h38d17437),
	.w4(32'h39ab3fda),
	.w5(32'hb7d9b2fe),
	.w6(32'h38b1bb79),
	.w7(32'h399fbd8c),
	.w8(32'h38b17f01),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62dbaa2),
	.w1(32'hb59eb41d),
	.w2(32'h35ad8b15),
	.w3(32'hb608fcd2),
	.w4(32'h34a66411),
	.w5(32'h363c22c4),
	.w6(32'hb6ba3bde),
	.w7(32'hb5d72027),
	.w8(32'h34eb0dd6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e3970a),
	.w1(32'h380b48aa),
	.w2(32'h37d7228f),
	.w3(32'h3702af78),
	.w4(32'h3822d041),
	.w5(32'h3832c702),
	.w6(32'h374a6d12),
	.w7(32'h38030f95),
	.w8(32'h380a5da2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392eaf40),
	.w1(32'h383b5801),
	.w2(32'hba14b911),
	.w3(32'h39b803c7),
	.w4(32'h399d5e77),
	.w5(32'hb96fee35),
	.w6(32'h39cacc23),
	.w7(32'h39bbcf1f),
	.w8(32'hb86210df),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb890b609),
	.w1(32'h38d09dd7),
	.w2(32'hb845c6cd),
	.w3(32'hb83c059f),
	.w4(32'h38c0daad),
	.w5(32'hb80f0de5),
	.w6(32'hb893ad8f),
	.w7(32'h37d21dec),
	.w8(32'hb91c9256),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369c82b9),
	.w1(32'hb61558ad),
	.w2(32'h370cb3fc),
	.w3(32'h37063d62),
	.w4(32'hb58f2a72),
	.w5(32'h3796f881),
	.w6(32'hb64dbe77),
	.w7(32'h355b0d9a),
	.w8(32'h35cfa90a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38383a53),
	.w1(32'hb79e1213),
	.w2(32'hb95d6d4d),
	.w3(32'h39143b51),
	.w4(32'h39373af7),
	.w5(32'h38843590),
	.w6(32'h39300fac),
	.w7(32'h395f5cda),
	.w8(32'h391cb002),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a317d79),
	.w1(32'hb8914db8),
	.w2(32'hba5d51ac),
	.w3(32'h3a497d0f),
	.w4(32'h398fd9c7),
	.w5(32'hba189715),
	.w6(32'h3a338c38),
	.w7(32'h3a0e6639),
	.w8(32'hb9f696ea),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae597be),
	.w1(32'hba5e292e),
	.w2(32'h3a066c06),
	.w3(32'hbaf619fd),
	.w4(32'hba8f8959),
	.w5(32'hb9db3b42),
	.w6(32'hbb003c1f),
	.w7(32'hba8f7d2f),
	.w8(32'hba01b241),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6bc29),
	.w1(32'hba14f589),
	.w2(32'hb8e5a0a8),
	.w3(32'hbadadc7b),
	.w4(32'hba507a57),
	.w5(32'hba236f3b),
	.w6(32'hbafebed5),
	.w7(32'hba966765),
	.w8(32'hba8a21a8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9826043),
	.w1(32'hb8e3a786),
	.w2(32'h38b51846),
	.w3(32'hb972c18e),
	.w4(32'hb8d77e4c),
	.w5(32'h383692b3),
	.w6(32'hb98e4d0c),
	.w7(32'hb90e45fc),
	.w8(32'hb81ee96c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3827e1df),
	.w1(32'h38a21c22),
	.w2(32'h38c2fe31),
	.w3(32'h3843b0da),
	.w4(32'h389568f7),
	.w5(32'h388a1c9d),
	.w6(32'h382d55c1),
	.w7(32'h38397721),
	.w8(32'h38543629),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3663603c),
	.w1(32'hb817a65f),
	.w2(32'h3798b720),
	.w3(32'hb807c1f5),
	.w4(32'hb85205d6),
	.w5(32'h370a5c8f),
	.w6(32'hb82e1dcf),
	.w7(32'hb82e5d4f),
	.w8(32'hb62eb584),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77f475),
	.w1(32'hb91af957),
	.w2(32'h396eaf9c),
	.w3(32'hba800c4e),
	.w4(32'hb913e502),
	.w5(32'h39504abe),
	.w6(32'hba8c467b),
	.w7(32'hb9614330),
	.w8(32'h3942d080),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896577f),
	.w1(32'hb9bc916e),
	.w2(32'hba25472d),
	.w3(32'h397d5b62),
	.w4(32'h392228be),
	.w5(32'hb887916a),
	.w6(32'h39e57d86),
	.w7(32'h39e079a6),
	.w8(32'h39d055a1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38332129),
	.w1(32'h38708e35),
	.w2(32'hba4b3dd8),
	.w3(32'h39a1058f),
	.w4(32'h39f663cd),
	.w5(32'hb9409cf1),
	.w6(32'h39ba92cb),
	.w7(32'h3a0a9a3b),
	.w8(32'h389bb73e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908dd20),
	.w1(32'h3903c0da),
	.w2(32'hba9e2903),
	.w3(32'h3a14254e),
	.w4(32'h3a482e7c),
	.w5(32'hb9c1c61f),
	.w6(32'h3a2ddcef),
	.w7(32'h3a8147d1),
	.w8(32'h394b27df),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e687e),
	.w1(32'hb887a799),
	.w2(32'hb9a6d474),
	.w3(32'hb8cf6105),
	.w4(32'h38ac4a55),
	.w5(32'hb90a66d9),
	.w6(32'hb9723cbf),
	.w7(32'hb7ed3dd5),
	.w8(32'hb919b9c6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e10396),
	.w1(32'h38a73ae9),
	.w2(32'hba2067b0),
	.w3(32'h39c5dff4),
	.w4(32'h3a025cc1),
	.w5(32'hb47c4e62),
	.w6(32'h3a1baf7e),
	.w7(32'h3a3b87ac),
	.w8(32'h3a035120),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d33287),
	.w1(32'h385abbe0),
	.w2(32'h390e7025),
	.w3(32'h384de45c),
	.w4(32'h3539efac),
	.w5(32'h38ce17d9),
	.w6(32'h37be33e3),
	.w7(32'h37a1a530),
	.w8(32'h3881e803),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390594e9),
	.w1(32'h3972e3e2),
	.w2(32'h39516aef),
	.w3(32'h376d9f68),
	.w4(32'h3941e843),
	.w5(32'h392c6f05),
	.w6(32'hb7b2628c),
	.w7(32'h38bf2d1c),
	.w8(32'h38e85ebd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e68960),
	.w1(32'h37c9c22c),
	.w2(32'hb7947da8),
	.w3(32'h37c8fde5),
	.w4(32'h38220d28),
	.w5(32'hb64d9bd9),
	.w6(32'hb7153b0a),
	.w7(32'h3856abdc),
	.w8(32'h3898818e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a8550e),
	.w1(32'h3944bf5a),
	.w2(32'hba1cc99a),
	.w3(32'h39d46b80),
	.w4(32'h3a0b6faa),
	.w5(32'hb89b4e0c),
	.w6(32'h3a06535c),
	.w7(32'h3a30a8b9),
	.w8(32'h398f487f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76ff825),
	.w1(32'h37e38a9d),
	.w2(32'hb96db67c),
	.w3(32'h3831ec87),
	.w4(32'h38ca64fc),
	.w5(32'hb930833b),
	.w6(32'h37964dfd),
	.w7(32'h38a02331),
	.w8(32'hb8906052),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76ae2d5),
	.w1(32'hb97b5427),
	.w2(32'hba9ebb2f),
	.w3(32'h39cc7a36),
	.w4(32'h39ad508b),
	.w5(32'hb9e8a5b8),
	.w6(32'h3a26e1dd),
	.w7(32'h3a15a583),
	.w8(32'h3967b63d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9061a9c),
	.w1(32'hb88325c2),
	.w2(32'hb82629cc),
	.w3(32'hb8d68aa2),
	.w4(32'hb88759e4),
	.w5(32'hb7d3bc07),
	.w6(32'hb8cf1b56),
	.w7(32'hb8a505d4),
	.w8(32'hb82e75ed),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367e04eb),
	.w1(32'h3685463b),
	.w2(32'h36df84a0),
	.w3(32'h35874c6a),
	.w4(32'h36008319),
	.w5(32'h36a11cbc),
	.w6(32'hb60259d0),
	.w7(32'h3552db59),
	.w8(32'hb49266fd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3691b946),
	.w1(32'hb360d89d),
	.w2(32'h36b53116),
	.w3(32'h36043758),
	.w4(32'hb61cb551),
	.w5(32'h3680861e),
	.w6(32'hb5ca9580),
	.w7(32'hb4535a14),
	.w8(32'h35e8601a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb672e0f7),
	.w1(32'h368bbc13),
	.w2(32'h37403d71),
	.w3(32'hb720bcab),
	.w4(32'hb6e77f01),
	.w5(32'h3713a0d1),
	.w6(32'hb609f5a2),
	.w7(32'hb61bf2da),
	.w8(32'h371f2dc9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c76c3),
	.w1(32'hb8a589a2),
	.w2(32'h3852a078),
	.w3(32'hb99c9a78),
	.w4(32'hb8e90184),
	.w5(32'h35c31426),
	.w6(32'hb9b6ee4d),
	.w7(32'hb93b900c),
	.w8(32'hb8bad770),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38768795),
	.w1(32'h353e60ed),
	.w2(32'hb6d80920),
	.w3(32'h3852ca64),
	.w4(32'h3809532d),
	.w5(32'h3700693f),
	.w6(32'h3775535c),
	.w7(32'h3833eb86),
	.w8(32'h37a5f883),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e9945),
	.w1(32'hb885faf4),
	.w2(32'hb9f1a601),
	.w3(32'h39937d80),
	.w4(32'h3998ac85),
	.w5(32'h38472d54),
	.w6(32'h39cb44d5),
	.w7(32'h39ebc098),
	.w8(32'h399d0036),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a5b0d9),
	.w1(32'hb8fd5262),
	.w2(32'hb9629640),
	.w3(32'hb8515835),
	.w4(32'hb866ffea),
	.w5(32'hb961bd9d),
	.w6(32'h3767dec2),
	.w7(32'hb8dfb173),
	.w8(32'hb93f94f6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c1d723),
	.w1(32'h3837efe6),
	.w2(32'h37e44f23),
	.w3(32'h3764be24),
	.w4(32'h37eb4985),
	.w5(32'h3798eb90),
	.w6(32'h3736ede3),
	.w7(32'h37a6cf68),
	.w8(32'h379725b5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a04d88),
	.w1(32'h36a88f64),
	.w2(32'h36bff7cd),
	.w3(32'h363bfacd),
	.w4(32'h36a8b1bb),
	.w5(32'h36a0d757),
	.w6(32'h36c4b257),
	.w7(32'h367ed80c),
	.w8(32'h36973f6d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f65bd1),
	.w1(32'h36af05c7),
	.w2(32'h37840b8c),
	.w3(32'hb50716f0),
	.w4(32'hb5724f2d),
	.w5(32'h36c6dcf3),
	.w6(32'hb7204b99),
	.w7(32'hb71ab7f6),
	.w8(32'h3710b363),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36342cab),
	.w1(32'hb603db71),
	.w2(32'h36b9fc29),
	.w3(32'h36361887),
	.w4(32'hb6e1f624),
	.w5(32'hb4d9e948),
	.w6(32'hb5934672),
	.w7(32'hb63d0aa8),
	.w8(32'h35490a0f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8019f4d),
	.w1(32'hb932afc5),
	.w2(32'hb9b98491),
	.w3(32'h38d5eaae),
	.w4(32'hb7a7d06b),
	.w5(32'hb96a5063),
	.w6(32'h3942198a),
	.w7(32'h37c81510),
	.w8(32'hb8e57c71),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3858662f),
	.w1(32'h35a765d8),
	.w2(32'hba9389ae),
	.w3(32'h3a134ad8),
	.w4(32'h3a0f6251),
	.w5(32'hba085a38),
	.w6(32'h3a187984),
	.w7(32'h3a5927cf),
	.w8(32'h37702090),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a937b9),
	.w1(32'hb8ef2088),
	.w2(32'hba670632),
	.w3(32'h3926d6c9),
	.w4(32'h39708eaa),
	.w5(32'hb9fc9842),
	.w6(32'h38ce9aa1),
	.w7(32'h390cd8f7),
	.w8(32'hb9d7aa1a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc0b98),
	.w1(32'h3a20a77b),
	.w2(32'hb925792b),
	.w3(32'h399ca708),
	.w4(32'h3a9e6cdb),
	.w5(32'h3a52379b),
	.w6(32'h393524ae),
	.w7(32'h3a8b2829),
	.w8(32'h39fcec28),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374d04d5),
	.w1(32'h36817947),
	.w2(32'h36d31828),
	.w3(32'h3733774f),
	.w4(32'h361ac3e1),
	.w5(32'h36c1e9b3),
	.w6(32'h36e22a2d),
	.w7(32'h36947d00),
	.w8(32'h36e612db),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37352274),
	.w1(32'h36dc8610),
	.w2(32'h375e4bd9),
	.w3(32'h36da5517),
	.w4(32'h356f35df),
	.w5(32'h36f7a6f6),
	.w6(32'h37548bac),
	.w7(32'h362ce32e),
	.w8(32'h370cae1b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37821a40),
	.w1(32'h33db1661),
	.w2(32'h372a2299),
	.w3(32'h371ac5fd),
	.w4(32'hb5c1b5ff),
	.w5(32'h36b699ca),
	.w6(32'h371a277e),
	.w7(32'h35e4dafd),
	.w8(32'h370cdfdd),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8049c9e),
	.w1(32'hb89bb355),
	.w2(32'hb95caa22),
	.w3(32'h3824c4f7),
	.w4(32'h37cb0cd7),
	.w5(32'hb842d89d),
	.w6(32'h38869ad8),
	.w7(32'h387f6ddb),
	.w8(32'h382c1f22),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3761702d),
	.w1(32'h35053469),
	.w2(32'h38157c59),
	.w3(32'hb738b118),
	.w4(32'hb7bec3eb),
	.w5(32'h37f16be1),
	.w6(32'hb6eabefb),
	.w7(32'hb775bf47),
	.w8(32'h37d4ffb6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d6dc1e),
	.w1(32'hb8ee83fd),
	.w2(32'hb998ca74),
	.w3(32'hb81bf281),
	.w4(32'hb8dcba5d),
	.w5(32'hb8987cb3),
	.w6(32'h38bc1af6),
	.w7(32'h38728cdd),
	.w8(32'h38363220),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a08e19),
	.w1(32'hb98537b5),
	.w2(32'hb9d5f0ec),
	.w3(32'h398a8f3c),
	.w4(32'h390e7988),
	.w5(32'hb7b2ba97),
	.w6(32'h39cf2498),
	.w7(32'h39cf74e4),
	.w8(32'h38aa31ef),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cb341f),
	.w1(32'h38a40276),
	.w2(32'hba1dc20a),
	.w3(32'h39cb4122),
	.w4(32'h3a1d0f26),
	.w5(32'h3920124c),
	.w6(32'h39f4080a),
	.w7(32'h3a36f2db),
	.w8(32'h39d258d6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3814a386),
	.w1(32'hb9262e8f),
	.w2(32'hba27f173),
	.w3(32'h396fb66a),
	.w4(32'h38c84159),
	.w5(32'hb9a37bc1),
	.w6(32'h39a94f26),
	.w7(32'h394214ea),
	.w8(32'hb9040422),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ffde4e),
	.w1(32'h3858b4d4),
	.w2(32'hb9d838b6),
	.w3(32'h397c6530),
	.w4(32'h398e6706),
	.w5(32'hb88ee9c5),
	.w6(32'h397d96a3),
	.w7(32'h39b9eeb4),
	.w8(32'h393a40da),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386a0351),
	.w1(32'h388881db),
	.w2(32'hb9c1df74),
	.w3(32'h394b19c0),
	.w4(32'h397502f7),
	.w5(32'hb91fdc39),
	.w6(32'h397b45d3),
	.w7(32'h3983e35d),
	.w8(32'hb8043d67),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d44cc9),
	.w1(32'h36b3cf71),
	.w2(32'hba295e0f),
	.w3(32'h3956bcf5),
	.w4(32'h397885ea),
	.w5(32'hb99ca152),
	.w6(32'h39a81d55),
	.w7(32'h39ade4c4),
	.w8(32'h37274617),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb541fe39),
	.w1(32'hb5848c71),
	.w2(32'h34429deb),
	.w3(32'hb61d803d),
	.w4(32'hb5f05a87),
	.w5(32'hb5a975fd),
	.w6(32'hb5307d59),
	.w7(32'hb5a6e1cf),
	.w8(32'hb4a729e4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362948f2),
	.w1(32'h364721b5),
	.w2(32'h3690826f),
	.w3(32'h36018786),
	.w4(32'h35a7c4e6),
	.w5(32'h3619e2d7),
	.w6(32'hb2de934e),
	.w7(32'h344cb693),
	.w8(32'h35bf6abe),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3721b098),
	.w1(32'h35fd3d34),
	.w2(32'h371d8bbb),
	.w3(32'h372b697c),
	.w4(32'h368d0c02),
	.w5(32'h3738456c),
	.w6(32'hb40c4082),
	.w7(32'h370b2702),
	.w8(32'h371c2b67),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e7dbbf),
	.w1(32'hb5bf4700),
	.w2(32'h37150188),
	.w3(32'hb6c11e79),
	.w4(32'h3653b921),
	.w5(32'h3784f361),
	.w6(32'hb76a65a0),
	.w7(32'hb667cee4),
	.w8(32'h3761905c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de7da3),
	.w1(32'hb9301a27),
	.w2(32'h381d9d76),
	.w3(32'hb9d7704c),
	.w4(32'hb965ffee),
	.w5(32'hb9106412),
	.w6(32'hb9d93edc),
	.w7(32'hb98ea1db),
	.w8(32'hb98380da),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63b1541),
	.w1(32'h38b3f34b),
	.w2(32'h382c236f),
	.w3(32'h37b0c942),
	.w4(32'h390d1495),
	.w5(32'h3897ac30),
	.w6(32'hb83572cb),
	.w7(32'h38939a85),
	.w8(32'h374745f7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79e326e),
	.w1(32'h3787ff89),
	.w2(32'hba211934),
	.w3(32'h39341185),
	.w4(32'h3984f5fc),
	.w5(32'hb9c90b81),
	.w6(32'h3987c688),
	.w7(32'h39de39c9),
	.w8(32'hb75e0b35),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4327e8),
	.w1(32'hba4889de),
	.w2(32'hba97d8d3),
	.w3(32'hba375eb4),
	.w4(32'hba5f2810),
	.w5(32'hba980cfb),
	.w6(32'hb9fb2671),
	.w7(32'hba33fcc8),
	.w8(32'hbaa0ada5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c9ada),
	.w1(32'hb989064f),
	.w2(32'h3787dd41),
	.w3(32'hba32f216),
	.w4(32'hb98438d1),
	.w5(32'hb8b087a1),
	.w6(32'hba62433b),
	.w7(32'hb9fdfea9),
	.w8(32'hb9998af4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a8cb5f),
	.w1(32'hb8ab0368),
	.w2(32'hba08376b),
	.w3(32'h38e617df),
	.w4(32'h386ba0cd),
	.w5(32'hb9c7fe40),
	.w6(32'h38f7345e),
	.w7(32'h396b16a7),
	.w8(32'hb9b08c46),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39778e88),
	.w1(32'h3993e425),
	.w2(32'hb7865cd4),
	.w3(32'h39e9ceb6),
	.w4(32'h3a0aa200),
	.w5(32'h399253f3),
	.w6(32'h39bb5c2e),
	.w7(32'h3a257f5c),
	.w8(32'h39fe7207),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfdc54),
	.w1(32'hb951a253),
	.w2(32'hba15f299),
	.w3(32'hb985f972),
	.w4(32'hb9098e8b),
	.w5(32'hba068085),
	.w6(32'hb9589c9d),
	.w7(32'hb92c652f),
	.w8(32'hba16014d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d59d24),
	.w1(32'h38dce7d8),
	.w2(32'hb9c3772e),
	.w3(32'hb77db740),
	.w4(32'h3950c821),
	.w5(32'hb95e2232),
	.w6(32'h385a464c),
	.w7(32'h39785285),
	.w8(32'hb9786144),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be7cc4),
	.w1(32'hb81a1181),
	.w2(32'hb834c69d),
	.w3(32'hb98ae622),
	.w4(32'h39098b00),
	.w5(32'h379897a7),
	.w6(32'hb9b5344d),
	.w7(32'h38503ef2),
	.w8(32'h389a25c6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386f632b),
	.w1(32'h393dcb51),
	.w2(32'h38a049f0),
	.w3(32'h37955362),
	.w4(32'h3935c809),
	.w5(32'h38dc878a),
	.w6(32'h36935268),
	.w7(32'h39434778),
	.w8(32'h38e1ee1e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39249de1),
	.w1(32'h39579a42),
	.w2(32'hba41b99b),
	.w3(32'h39b09569),
	.w4(32'h3a447d6a),
	.w5(32'hb61d0114),
	.w6(32'h39b24d94),
	.w7(32'h3a531dbe),
	.w8(32'h39a45d77),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a71c04),
	.w1(32'h38876e69),
	.w2(32'hba38c171),
	.w3(32'h39da3708),
	.w4(32'h39c9674d),
	.w5(32'hb9410ac4),
	.w6(32'h39d3dc77),
	.w7(32'h39c5953f),
	.w8(32'hb9a828cb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1046ab),
	.w1(32'h381274d1),
	.w2(32'hba980ce0),
	.w3(32'h3a487f3f),
	.w4(32'h39b83ae3),
	.w5(32'hba4615cc),
	.w6(32'h3a58614d),
	.w7(32'h3a303a9c),
	.w8(32'hb9feeeaa),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09763b),
	.w1(32'hba965d63),
	.w2(32'h3a48bbbf),
	.w3(32'hbb1aeb23),
	.w4(32'hbac6786b),
	.w5(32'hb9d7090c),
	.w6(32'hbb379f9c),
	.w7(32'hbb003301),
	.w8(32'hba76b2f4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb55f719c),
	.w1(32'h3a034e22),
	.w2(32'hba3c4161),
	.w3(32'h39acf4d1),
	.w4(32'h3a5c82be),
	.w5(32'hb8e56fdd),
	.w6(32'h3a047e1c),
	.w7(32'h3a80f8ce),
	.w8(32'h39b36235),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3976bbdd),
	.w1(32'hb885170c),
	.w2(32'hb9498d08),
	.w3(32'h39843bb3),
	.w4(32'h3938033f),
	.w5(32'h388a8cef),
	.w6(32'h394d595a),
	.w7(32'h39703316),
	.w8(32'h385b05fc),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d10b7),
	.w1(32'h39037524),
	.w2(32'h38cab1fa),
	.w3(32'h38ae5a73),
	.w4(32'h39276faf),
	.w5(32'h3959432f),
	.w6(32'hb71ba6cb),
	.w7(32'h38e8ac97),
	.w8(32'h38dc5254),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39088a4c),
	.w1(32'hb78e4ef3),
	.w2(32'hbaa71483),
	.w3(32'h3a199abe),
	.w4(32'h395e0911),
	.w5(32'hba04d2e5),
	.w6(32'h3a43996b),
	.w7(32'h3a1fafd1),
	.w8(32'h380bef11),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e4183),
	.w1(32'h39bab713),
	.w2(32'h392dc69b),
	.w3(32'h38a05d3a),
	.w4(32'h3a0d4141),
	.w5(32'h3a11ac94),
	.w6(32'h38b2351a),
	.w7(32'h3a2e9299),
	.w8(32'h3a1169e6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6993e17),
	.w1(32'hb70b5f2c),
	.w2(32'hb63a1053),
	.w3(32'hb63aebae),
	.w4(32'h35f8da23),
	.w5(32'h36e9ae81),
	.w6(32'hb694e9e8),
	.w7(32'h359cec71),
	.w8(32'hb596fd37),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8285867),
	.w1(32'h38470f3c),
	.w2(32'hb8464fc3),
	.w3(32'hb80320a8),
	.w4(32'h38956365),
	.w5(32'hb8bc3700),
	.w6(32'hb89c23e3),
	.w7(32'h370aaa62),
	.w8(32'hb8f97a81),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986a00b),
	.w1(32'hb9407596),
	.w2(32'hb93e6e29),
	.w3(32'hb888adb1),
	.w4(32'h3910afce),
	.w5(32'h3908e314),
	.w6(32'h360a2cb3),
	.w7(32'h395d2fdd),
	.w8(32'h397087fb),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7ca13),
	.w1(32'h39cb36d8),
	.w2(32'hb98b9351),
	.w3(32'h39f84a7a),
	.w4(32'h3a2911f6),
	.w5(32'h3964c785),
	.w6(32'h39e848f6),
	.w7(32'h3a3a1309),
	.w8(32'h39e81a22),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9c670),
	.w1(32'hb9a7d828),
	.w2(32'hb9aad22f),
	.w3(32'hb9a5573e),
	.w4(32'hb9a9191e),
	.w5(32'hb9c21b22),
	.w6(32'hb9e5d8bd),
	.w7(32'hb9ee5620),
	.w8(32'hb9dabd26),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3895b58b),
	.w1(32'h39708bf6),
	.w2(32'hb9600d94),
	.w3(32'h396c60b8),
	.w4(32'h39b30d9b),
	.w5(32'hb7879959),
	.w6(32'h38ffe379),
	.w7(32'h3983dd77),
	.w8(32'hb9027145),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9896872),
	.w1(32'hb8bf47b9),
	.w2(32'h382a15d4),
	.w3(32'hb91b58ee),
	.w4(32'hb8cbee5a),
	.w5(32'h384b1555),
	.w6(32'hb7e8ddf1),
	.w7(32'h3858b344),
	.w8(32'h38dfadd3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dfcb2e),
	.w1(32'hb53d3d92),
	.w2(32'hb9fecc40),
	.w3(32'h39a700d3),
	.w4(32'h393bc813),
	.w5(32'hb9caac74),
	.w6(32'h39d56db7),
	.w7(32'h39b92828),
	.w8(32'hb926b12d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8539756),
	.w1(32'h376440d9),
	.w2(32'hb9acffe3),
	.w3(32'h38c1228e),
	.w4(32'h394211ae),
	.w5(32'hb8c42128),
	.w6(32'h38d9f69d),
	.w7(32'h39721144),
	.w8(32'h37b9ede2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb610f498),
	.w1(32'hb571941f),
	.w2(32'hb62a4268),
	.w3(32'hb6acdefd),
	.w4(32'hb688f99a),
	.w5(32'hb5fb50d8),
	.w6(32'h35471ea4),
	.w7(32'hb687a2ef),
	.w8(32'hb627ad57),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3726b52d),
	.w1(32'h37a93dbf),
	.w2(32'h370af9dc),
	.w3(32'h3765a2ef),
	.w4(32'h3616af25),
	.w5(32'hb5613ca3),
	.w6(32'h3798b501),
	.w7(32'h370f3478),
	.w8(32'hb607cfec),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3661c21e),
	.w1(32'hb39eb92d),
	.w2(32'h362df62f),
	.w3(32'h366f883a),
	.w4(32'hb543c3d2),
	.w5(32'h3517c5cf),
	.w6(32'h366f0e00),
	.w7(32'h34bef342),
	.w8(32'h36b85050),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369dc747),
	.w1(32'hb69c099b),
	.w2(32'hb5d9cbde),
	.w3(32'h36aa0b72),
	.w4(32'hb58212bf),
	.w5(32'h34d0266c),
	.w6(32'h369dcc9e),
	.w7(32'h36165b5d),
	.w8(32'h361bbdca),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74f0305),
	.w1(32'h3710450b),
	.w2(32'hba22aeed),
	.w3(32'h397e25ae),
	.w4(32'h39b0ea66),
	.w5(32'hb8fdcfe9),
	.w6(32'h39a3c0f2),
	.w7(32'h39fb8eaa),
	.w8(32'h3927ad4b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38211706),
	.w1(32'h3722c014),
	.w2(32'h35b481f0),
	.w3(32'h37db779b),
	.w4(32'h36f2ba68),
	.w5(32'h36dfc94e),
	.w6(32'h37f90dc2),
	.w7(32'h373b07e5),
	.w8(32'h36ebd87a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37553a9e),
	.w1(32'h37b7a004),
	.w2(32'hb94a61a6),
	.w3(32'h3911cdd9),
	.w4(32'h39395d3b),
	.w5(32'h38801660),
	.w6(32'h39506692),
	.w7(32'h396e61b9),
	.w8(32'h3921adbb),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995d47e),
	.w1(32'hb8c698a3),
	.w2(32'hb8e76f0c),
	.w3(32'hb96ede55),
	.w4(32'hb8ce8d40),
	.w5(32'hb9b0a987),
	.w6(32'hb9a8af2c),
	.w7(32'hb981b515),
	.w8(32'hba197571),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379dda42),
	.w1(32'h379b8c51),
	.w2(32'hb7a525bf),
	.w3(32'h37afa654),
	.w4(32'h374aeac2),
	.w5(32'hb70af501),
	.w6(32'h37b480e8),
	.w7(32'h3739c730),
	.w8(32'hb7210d2f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378cc6fb),
	.w1(32'h37405796),
	.w2(32'h36f64885),
	.w3(32'h37a6aa45),
	.w4(32'h3767f6d6),
	.w5(32'h36b72648),
	.w6(32'h371b50cb),
	.w7(32'h375a3bdb),
	.w8(32'h375d26d5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69a0f4e),
	.w1(32'hb6c9b51c),
	.w2(32'hb5a8a240),
	.w3(32'hb6ceac5c),
	.w4(32'hb65e00bc),
	.w5(32'h35503b09),
	.w6(32'hb7247df6),
	.w7(32'hb6dcadbc),
	.w8(32'hb5c16829),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9248398),
	.w1(32'hb8aaa503),
	.w2(32'hb871a4d1),
	.w3(32'hb919ebdf),
	.w4(32'hb8f54d82),
	.w5(32'hb908eb19),
	.w6(32'hb926ecc8),
	.w7(32'hb90ad795),
	.w8(32'hb92e8e48),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399bda6a),
	.w1(32'h39344b4c),
	.w2(32'hb9cc2a7d),
	.w3(32'h39b2e341),
	.w4(32'h396e5955),
	.w5(32'hb9be46b9),
	.w6(32'h3a0e3d35),
	.w7(32'h39f3795c),
	.w8(32'hb8079028),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f46e7),
	.w1(32'hb833069c),
	.w2(32'hba6c996d),
	.w3(32'h3a027317),
	.w4(32'h39e41d42),
	.w5(32'hb969f945),
	.w6(32'h3a22f9e8),
	.w7(32'h3a0f4799),
	.w8(32'h391ad119),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368bdc37),
	.w1(32'hb7689b9f),
	.w2(32'hb7024a04),
	.w3(32'hb724e74b),
	.w4(32'hb7a6ee9c),
	.w5(32'hb816374b),
	.w6(32'h35795f13),
	.w7(32'hb7b83935),
	.w8(32'hb7db686e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c7190),
	.w1(32'h37066d63),
	.w2(32'hb7953348),
	.w3(32'hb774158e),
	.w4(32'h378aecc5),
	.w5(32'h381089cf),
	.w6(32'hb76b7637),
	.w7(32'h3844420a),
	.w8(32'h37db6a12),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9935fe6),
	.w1(32'hb8c88e4b),
	.w2(32'hb965ca2c),
	.w3(32'hb942a13a),
	.w4(32'hb7df06d2),
	.w5(32'hb956968c),
	.w6(32'hb95d5e2a),
	.w7(32'hb814ec4c),
	.w8(32'hb8ad7928),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb849c1de),
	.w1(32'h3696b9c6),
	.w2(32'hb976ed5a),
	.w3(32'h3869614f),
	.w4(32'h391617ea),
	.w5(32'hb8c96fb9),
	.w6(32'h38a7e277),
	.w7(32'h39256e3d),
	.w8(32'h370b76b0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bea899),
	.w1(32'h39154c7a),
	.w2(32'hb98561a3),
	.w3(32'h385725be),
	.w4(32'h3921680e),
	.w5(32'hb9d96ca3),
	.w6(32'h39441a30),
	.w7(32'h3913bc2b),
	.w8(32'hb989d23c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb2e16),
	.w1(32'hb86737a5),
	.w2(32'hba7447a1),
	.w3(32'h39b4adef),
	.w4(32'h39a13543),
	.w5(32'hb9a565aa),
	.w6(32'h3a0739e5),
	.w7(32'h3a115d4e),
	.w8(32'h3899ae03),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997bcde),
	.w1(32'hb86fa75b),
	.w2(32'hb8df2967),
	.w3(32'hb980f752),
	.w4(32'hb50c5c0e),
	.w5(32'hb84df810),
	.w6(32'hb99f45b3),
	.w7(32'hb88fbddd),
	.w8(32'hb91b0920),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3867411e),
	.w1(32'hb83fc294),
	.w2(32'hba02067b),
	.w3(32'h39b18582),
	.w4(32'h39a95aad),
	.w5(32'hb906d466),
	.w6(32'h3998c089),
	.w7(32'h396baefe),
	.w8(32'hb7b79703),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92efc71),
	.w1(32'hb993214f),
	.w2(32'hba64c6e7),
	.w3(32'hb850a4aa),
	.w4(32'h38983d01),
	.w5(32'hba094994),
	.w6(32'h391a7be4),
	.w7(32'h39544a1a),
	.w8(32'hb9597bde),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98733a3),
	.w1(32'hb8c4250a),
	.w2(32'hb914023a),
	.w3(32'hb928621d),
	.w4(32'hb880c496),
	.w5(32'hb91de806),
	.w6(32'hb93dbd10),
	.w7(32'hb88b6985),
	.w8(32'hb92cedc4),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb890b208),
	.w1(32'hb7a77a97),
	.w2(32'hb968d6e4),
	.w3(32'h3828b788),
	.w4(32'h390120c2),
	.w5(32'hb808a58d),
	.w6(32'h373f4952),
	.w7(32'h38f71c6c),
	.w8(32'hb809d34c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38607823),
	.w1(32'h377b6471),
	.w2(32'hb9826de7),
	.w3(32'h391d77a0),
	.w4(32'h392158d0),
	.w5(32'hb840a403),
	.w6(32'h394951a5),
	.w7(32'h39526d34),
	.w8(32'h3862f04f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8638f),
	.w1(32'hb883d311),
	.w2(32'hb92c7262),
	.w3(32'hb96162a2),
	.w4(32'h388771bd),
	.w5(32'hb8de90f0),
	.w6(32'hb9d3a4dd),
	.w7(32'hb92facc7),
	.w8(32'hb9c9e9a5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94da0cc),
	.w1(32'hb8f45f37),
	.w2(32'hb93644df),
	.w3(32'hb91ce14e),
	.w4(32'hb8cf2d12),
	.w5(32'hb928ee94),
	.w6(32'hb9205b04),
	.w7(32'hb902174d),
	.w8(32'hb94de89d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h356474bd),
	.w1(32'h364d7a8f),
	.w2(32'h3657e1c3),
	.w3(32'h366e9095),
	.w4(32'h36531fb5),
	.w5(32'h36834742),
	.w6(32'h3656cff4),
	.w7(32'h365113ae),
	.w8(32'h367fe35a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5be10af),
	.w1(32'h3437122c),
	.w2(32'hb56a2e85),
	.w3(32'h35cc43e5),
	.w4(32'h35eda8db),
	.w5(32'hb62bb29a),
	.w6(32'h349b52e3),
	.w7(32'h3591046d),
	.w8(32'hb594116c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f7e29),
	.w1(32'h38a69d95),
	.w2(32'hb7bd8872),
	.w3(32'hb82c44f4),
	.w4(32'h38ee2164),
	.w5(32'h38d9d02b),
	.w6(32'hb83749f4),
	.w7(32'h3915c319),
	.w8(32'h38dc50ef),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a858eb),
	.w1(32'hb807c7b7),
	.w2(32'hb923ba89),
	.w3(32'hb974d982),
	.w4(32'h36441084),
	.w5(32'hb8f5d728),
	.w6(32'hb9bc54d8),
	.w7(32'hb8910363),
	.w8(32'hb90a28e8),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f19c76),
	.w1(32'hb75e8e23),
	.w2(32'hba90716d),
	.w3(32'h3a32605b),
	.w4(32'h3a3ddcb5),
	.w5(32'h37ac081c),
	.w6(32'h3a56b7d4),
	.w7(32'h3a7dd881),
	.w8(32'h3a05984c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b6a10a),
	.w1(32'h378dcf77),
	.w2(32'h35f47bc6),
	.w3(32'h361bf15d),
	.w4(32'h375cc881),
	.w5(32'h362e9f7e),
	.w6(32'h368cdc56),
	.w7(32'h37308d01),
	.w8(32'h36c0ca96),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38932887),
	.w1(32'hb8807507),
	.w2(32'hba55d43b),
	.w3(32'h39b5f068),
	.w4(32'h39c9afb1),
	.w5(32'hb9210cae),
	.w6(32'h39efc1b0),
	.w7(32'h39fb0cba),
	.w8(32'h39010f73),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d26a92),
	.w1(32'h38ccb5c7),
	.w2(32'hb9c91d3b),
	.w3(32'h383d66db),
	.w4(32'h39ac8eeb),
	.w5(32'hb8b005c8),
	.w6(32'h38dfc926),
	.w7(32'h39c5eb2c),
	.w8(32'h3895f7ce),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aaa44e),
	.w1(32'hb84a2504),
	.w2(32'hb99fa961),
	.w3(32'h3975fa69),
	.w4(32'h397f5d7d),
	.w5(32'h387e5ffc),
	.w6(32'h39c17bbe),
	.w7(32'h39b7ac7a),
	.w8(32'h3990da12),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c40332),
	.w1(32'h39de5a6e),
	.w2(32'hb9c1b461),
	.w3(32'h3a4067e1),
	.w4(32'h3a53982e),
	.w5(32'h39ada34e),
	.w6(32'h3a4c424b),
	.w7(32'h3a7b11b0),
	.w8(32'h3a177cb7),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05f205),
	.w1(32'hb9a88e51),
	.w2(32'hb88ff1c7),
	.w3(32'hba25cd59),
	.w4(32'hb9d75f5d),
	.w5(32'hb99f5aec),
	.w6(32'hba33edba),
	.w7(32'hba00c816),
	.w8(32'hb9c16967),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392cae73),
	.w1(32'h38d99c3a),
	.w2(32'h38349801),
	.w3(32'h38d5a8fa),
	.w4(32'h39284bf3),
	.w5(32'h381b7a4c),
	.w6(32'h38059fd4),
	.w7(32'h38bc53bf),
	.w8(32'hb7656753),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991cf49),
	.w1(32'h38ec8ea3),
	.w2(32'h38931651),
	.w3(32'hb9c2fb30),
	.w4(32'h38d57975),
	.w5(32'h38492494),
	.w6(32'hba14d85d),
	.w7(32'hb9237a6f),
	.w8(32'hb93b40e1),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51c6a1),
	.w1(32'hb9f290e1),
	.w2(32'hb95e067b),
	.w3(32'hba5f219d),
	.w4(32'hba205981),
	.w5(32'hba1a201d),
	.w6(32'hba6dcadd),
	.w7(32'hba39c9ad),
	.w8(32'hba24c3cb),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9958068),
	.w1(32'h3743d772),
	.w2(32'h394ecc08),
	.w3(32'hb99ac092),
	.w4(32'hb79d4c8b),
	.w5(32'h38c73c22),
	.w6(32'hb9ca73a3),
	.w7(32'hb8e60f44),
	.w8(32'hb7b46748),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79179a9),
	.w1(32'hb81807dc),
	.w2(32'hb9251967),
	.w3(32'h37e075f3),
	.w4(32'hb74ee0a5),
	.w5(32'hb8d37910),
	.w6(32'h385022b5),
	.w7(32'h3882ee27),
	.w8(32'hb81ab27b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82b05ea),
	.w1(32'hb8135e24),
	.w2(32'hb84cd065),
	.w3(32'hb871da4e),
	.w4(32'hb8697a29),
	.w5(32'hb8a308c5),
	.w6(32'hb881eb22),
	.w7(32'hb88da777),
	.w8(32'hb8ca124b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d0c10d),
	.w1(32'hb81d4671),
	.w2(32'hb9901fd1),
	.w3(32'hb7aa2f13),
	.w4(32'h38dc4ebf),
	.w5(32'hb8e036f8),
	.w6(32'h37bed9d7),
	.w7(32'h392e1d93),
	.w8(32'hb632d202),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ed564e),
	.w1(32'h37299c12),
	.w2(32'h374211d0),
	.w3(32'h379250b3),
	.w4(32'h36b8cd87),
	.w5(32'h37e2ebd1),
	.w6(32'h37419bbb),
	.w7(32'h3724e07b),
	.w8(32'h37516bf7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ce869d),
	.w1(32'h38ceccfb),
	.w2(32'hb9086e2b),
	.w3(32'h38c07eec),
	.w4(32'h3974a4b2),
	.w5(32'h38dc9d7f),
	.w6(32'h390d6230),
	.w7(32'h39895d2c),
	.w8(32'h396bff3c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3782ed39),
	.w1(32'hb7895b4c),
	.w2(32'h379c969c),
	.w3(32'h379226d2),
	.w4(32'h36b3a8f0),
	.w5(32'h377f2716),
	.w6(32'h37e7e4df),
	.w7(32'h37a48cc3),
	.w8(32'h37196172),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39189135),
	.w1(32'h391d54e9),
	.w2(32'hb8d6e9b1),
	.w3(32'h39a331f4),
	.w4(32'h39d0a8c4),
	.w5(32'h39a15192),
	.w6(32'h39800056),
	.w7(32'h39c8775a),
	.w8(32'h39a9b884),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3782c172),
	.w1(32'h35ac9a9b),
	.w2(32'h3802b348),
	.w3(32'h36f42a8a),
	.w4(32'h374b356c),
	.w5(32'h384533bf),
	.w6(32'hb61dcdf4),
	.w7(32'h371c28c7),
	.w8(32'h38389290),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ecdb75),
	.w1(32'hb441cd13),
	.w2(32'hb7312399),
	.w3(32'hb5e6c320),
	.w4(32'h37db8e69),
	.w5(32'hb730bae8),
	.w6(32'h36f3c3d4),
	.w7(32'h380edb28),
	.w8(32'hb6c90935),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3c614),
	.w1(32'hb94d3bb3),
	.w2(32'hb7b3cca0),
	.w3(32'hb9fa673c),
	.w4(32'hb989847d),
	.w5(32'hb96b343c),
	.w6(32'hba163852),
	.w7(32'hb9b79d7f),
	.w8(32'hb9a86a84),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9226856),
	.w1(32'hba0880cc),
	.w2(32'hbab654de),
	.w3(32'h39155a88),
	.w4(32'hb919e7b5),
	.w5(32'hbaba4ca2),
	.w6(32'h390fdeda),
	.w7(32'h3933daed),
	.w8(32'hba2f89e0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b83110),
	.w1(32'hb8c36ab3),
	.w2(32'h382ec905),
	.w3(32'hb9b67200),
	.w4(32'hb8caefdf),
	.w5(32'h379469ad),
	.w6(32'hb9d2fc65),
	.w7(32'hb939cd2f),
	.w8(32'hb886374c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9599dc7),
	.w1(32'hb8447743),
	.w2(32'hb9c74970),
	.w3(32'h380be13d),
	.w4(32'h39670bbe),
	.w5(32'hb70724fa),
	.w6(32'h37b7ead0),
	.w7(32'h3982feb7),
	.w8(32'h388b153b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9146d5d),
	.w1(32'hb841fda7),
	.w2(32'hb7d3e16d),
	.w3(32'hb8c65208),
	.w4(32'hb6c9a767),
	.w5(32'hb5e3d976),
	.w6(32'hb8f75702),
	.w7(32'hb861ddbd),
	.w8(32'hb7ab9837),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c45fa5),
	.w1(32'hb90ec229),
	.w2(32'hba85736a),
	.w3(32'h39fe9171),
	.w4(32'h3a333127),
	.w5(32'h36989e5f),
	.w6(32'h3a434cd5),
	.w7(32'h3a633497),
	.w8(32'h3a216d19),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953a055),
	.w1(32'h3853fc91),
	.w2(32'hb9e1a9aa),
	.w3(32'hb83fee33),
	.w4(32'h39965d30),
	.w5(32'hb910482b),
	.w6(32'h37e40b3c),
	.w7(32'h39948319),
	.w8(32'hb83971c4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec9dc4),
	.w1(32'h38af03f7),
	.w2(32'hba9bf229),
	.w3(32'h3a396bde),
	.w4(32'h3a159da3),
	.w5(32'hba1af8af),
	.w6(32'h3a451710),
	.w7(32'h3a24b7f2),
	.w8(32'hb852c095),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384a88f5),
	.w1(32'hb659340a),
	.w2(32'h384ea2be),
	.w3(32'h3839d126),
	.w4(32'hb780860d),
	.w5(32'h384e8b66),
	.w6(32'h37d0ca68),
	.w7(32'hb7db7850),
	.w8(32'h37fd01a8),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39494e42),
	.w1(32'hb7ebc4a9),
	.w2(32'hb9ec7c7d),
	.w3(32'h39a63579),
	.w4(32'h39203927),
	.w5(32'hb9a7a1fe),
	.w6(32'h39b07105),
	.w7(32'h3951178f),
	.w8(32'hb90ee2e8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a8f6f2),
	.w1(32'h360e6e7f),
	.w2(32'h366e72a3),
	.w3(32'h368fbd48),
	.w4(32'h3642ca6c),
	.w5(32'h36a8f836),
	.w6(32'h3691346f),
	.w7(32'h36905af2),
	.w8(32'h36a138b9),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39815f44),
	.w1(32'h38b3f5f6),
	.w2(32'hb98a005c),
	.w3(32'h39a852ab),
	.w4(32'h39245c7f),
	.w5(32'hb949db00),
	.w6(32'h39a4e6da),
	.w7(32'h395532fa),
	.w8(32'hb9066c75),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9757330),
	.w1(32'h38ae533a),
	.w2(32'h3895b3b2),
	.w3(32'hb973074e),
	.w4(32'h38613e1e),
	.w5(32'h38177276),
	.w6(32'hb984562c),
	.w7(32'h387407d1),
	.w8(32'h380c0b9e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88d7ce4),
	.w1(32'hb8752c29),
	.w2(32'hb99b8f01),
	.w3(32'h38ba8552),
	.w4(32'h3911b334),
	.w5(32'hb8abca9f),
	.w6(32'h392b0bab),
	.w7(32'h3930bb77),
	.w8(32'h380cfd72),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b5f30c),
	.w1(32'h34b11082),
	.w2(32'h33f6dbfd),
	.w3(32'h367fa8be),
	.w4(32'hb5cf104f),
	.w5(32'h358e4fab),
	.w6(32'h367a01aa),
	.w7(32'h3633e842),
	.w8(32'h3603cb22),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f8d136),
	.w1(32'h3845ad79),
	.w2(32'h38381471),
	.w3(32'h3720019c),
	.w4(32'h37e11b9f),
	.w5(32'h37edd511),
	.w6(32'hb67caf3d),
	.w7(32'h3773a39a),
	.w8(32'h3797f272),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b405b),
	.w1(32'hb875fc46),
	.w2(32'h380dc29d),
	.w3(32'hb95cc280),
	.w4(32'hb88382ea),
	.w5(32'h38617a15),
	.w6(32'hb951a0d0),
	.w7(32'hb8bf6435),
	.w8(32'hb7d8bb5f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8af72e7),
	.w1(32'hb7c08efa),
	.w2(32'hb9a03ec7),
	.w3(32'hb84e60eb),
	.w4(32'h38a740f6),
	.w5(32'hb93df4d5),
	.w6(32'hb83faa41),
	.w7(32'h37c50cf0),
	.w8(32'hb96fa222),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3836ec81),
	.w1(32'hb83267f9),
	.w2(32'hb7f9f3bb),
	.w3(32'h38655e51),
	.w4(32'hb8945b50),
	.w5(32'hb6f12570),
	.w6(32'h371b077c),
	.w7(32'h37cd0841),
	.w8(32'hb7a151cd),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80210a2),
	.w1(32'hb836cf87),
	.w2(32'hb8c72636),
	.w3(32'hb785e642),
	.w4(32'h36b9e431),
	.w5(32'hb862fe31),
	.w6(32'hb76fe61a),
	.w7(32'h37a69816),
	.w8(32'hb81602f4),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399dc7b7),
	.w1(32'hb93ffdf4),
	.w2(32'hba9c144a),
	.w3(32'h3a86015a),
	.w4(32'h3a8d3a32),
	.w5(32'h3a368a37),
	.w6(32'h3a969122),
	.w7(32'h3ab3726c),
	.w8(32'h3aa8c45c),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a7988),
	.w1(32'hb9b8816f),
	.w2(32'hb9ca0433),
	.w3(32'hba5cf67d),
	.w4(32'hb9f34a75),
	.w5(32'hba22419e),
	.w6(32'hba5d8c86),
	.w7(32'hba0e09ef),
	.w8(32'hba23743f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38633dcf),
	.w1(32'h37498512),
	.w2(32'h3839e2b1),
	.w3(32'h3865aef7),
	.w4(32'h36c7e4d5),
	.w5(32'h3886cd5e),
	.w6(32'h3807d530),
	.w7(32'h3806c651),
	.w8(32'h383f25be),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3722d0f1),
	.w1(32'h37050499),
	.w2(32'hb5c0cd18),
	.w3(32'h36ee8dbd),
	.w4(32'h36dba00e),
	.w5(32'hb6f98229),
	.w6(32'h366dbef0),
	.w7(32'hb5e326dc),
	.w8(32'hb6ad6e05),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c7e0a4),
	.w1(32'h39290868),
	.w2(32'h389b875c),
	.w3(32'h371d3191),
	.w4(32'h38a29fbd),
	.w5(32'hb6972ddd),
	.w6(32'hb8629f21),
	.w7(32'hb5dc3016),
	.w8(32'hb8183d94),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f21a58),
	.w1(32'hb3dd4ccf),
	.w2(32'h3605b234),
	.w3(32'h363fa44c),
	.w4(32'hb5e1a621),
	.w5(32'h3537a6cb),
	.w6(32'h3622c67b),
	.w7(32'hb5a0f9be),
	.w8(32'h361ed905),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d5b669),
	.w1(32'hb8395aac),
	.w2(32'hb81c72db),
	.w3(32'hb80ee4ef),
	.w4(32'hb8868e80),
	.w5(32'hb89ad7ae),
	.w6(32'hb83349b2),
	.w7(32'hb87b56b6),
	.w8(32'hb8adf209),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f7dad),
	.w1(32'hb8414a38),
	.w2(32'hba415499),
	.w3(32'h386f003c),
	.w4(32'h3940f372),
	.w5(32'hba0496cf),
	.w6(32'hb6cff8b6),
	.w7(32'h394a6594),
	.w8(32'hb99aecfd),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382216cf),
	.w1(32'hb8b02cf3),
	.w2(32'hba2869ea),
	.w3(32'h39a96399),
	.w4(32'h39c779b2),
	.w5(32'hb81274c6),
	.w6(32'h39cd5cc4),
	.w7(32'h3a142fed),
	.w8(32'h39905a26),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb891f8a9),
	.w1(32'hb75ab46a),
	.w2(32'h379d8cf3),
	.w3(32'hb81f5795),
	.w4(32'h37443a51),
	.w5(32'h37e69488),
	.w6(32'hb87fb745),
	.w7(32'hb6895fac),
	.w8(32'hb474d75c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a1378a),
	.w1(32'hb8b34f7a),
	.w2(32'hba095b7a),
	.w3(32'h39816b4f),
	.w4(32'h39d94d8a),
	.w5(32'h389352c3),
	.w6(32'h39b37096),
	.w7(32'h3a19f3d9),
	.w8(32'h39d87c25),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a721d),
	.w1(32'h39241b13),
	.w2(32'h36d61137),
	.w3(32'h39a3012f),
	.w4(32'h39a9803b),
	.w5(32'h39ae7b37),
	.w6(32'h39acb6c1),
	.w7(32'h39cf8b85),
	.w8(32'h39d47636),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f8c788),
	.w1(32'h363322dd),
	.w2(32'h36c207c4),
	.w3(32'h36d0e1b8),
	.w4(32'h355997e1),
	.w5(32'h369cf5f1),
	.w6(32'h36ee47bf),
	.w7(32'h361ea883),
	.w8(32'h36985739),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e990e0),
	.w1(32'h374e64ec),
	.w2(32'hb85a577c),
	.w3(32'hb5b0dc90),
	.w4(32'h3719ed97),
	.w5(32'hb87a2cf0),
	.w6(32'h385fcdad),
	.w7(32'h37aeebbe),
	.w8(32'hb7d0e5cf),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37684f72),
	.w1(32'h36ab953d),
	.w2(32'h3752d4aa),
	.w3(32'h37294c8a),
	.w4(32'h357663c6),
	.w5(32'h36ca238b),
	.w6(32'h373ae5b6),
	.w7(32'h3629da2c),
	.w8(32'h36d3c777),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ccd7b6),
	.w1(32'h3994428d),
	.w2(32'hb8c74c78),
	.w3(32'h39693158),
	.w4(32'h39f713b4),
	.w5(32'h39aa8f4e),
	.w6(32'h3961c748),
	.w7(32'h3a27d0e6),
	.w8(32'h39ec8e05),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1735b1),
	.w1(32'hb95a3ac5),
	.w2(32'hb90fc864),
	.w3(32'hba182608),
	.w4(32'hb99e10c7),
	.w5(32'hb9d18042),
	.w6(32'hba1f99a9),
	.w7(32'hb9c79c08),
	.w8(32'hb9fcabdd),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4588f),
	.w1(32'hb83a0637),
	.w2(32'hb95d13fd),
	.w3(32'hb94c9da0),
	.w4(32'h3897766f),
	.w5(32'hb8c06507),
	.w6(32'hb968ccaa),
	.w7(32'h384b67e2),
	.w8(32'hb8d7d252),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0e466),
	.w1(32'hb974f892),
	.w2(32'h38af4983),
	.w3(32'hb9bf5e82),
	.w4(32'hb9986f17),
	.w5(32'hb852cde7),
	.w6(32'hb9d8dc7d),
	.w7(32'hb9b685bc),
	.w8(32'hb94c4cfb),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b4a3b),
	.w1(32'hb9341db8),
	.w2(32'hb95cdabd),
	.w3(32'hb9d8a5a7),
	.w4(32'hb89e2788),
	.w5(32'hb91b0144),
	.w6(32'hb9eb86c0),
	.w7(32'hb8f9e96d),
	.w8(32'hb94ab1c0),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902828a),
	.w1(32'h38c122fd),
	.w2(32'hb9adfef5),
	.w3(32'h39792174),
	.w4(32'h3992a3d1),
	.w5(32'h366c7f7c),
	.w6(32'h39a16a88),
	.w7(32'h39c7ca36),
	.w8(32'h395252bf),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c39d98),
	.w1(32'h37f57152),
	.w2(32'hba913c89),
	.w3(32'h3a8188bb),
	.w4(32'h3a83a641),
	.w5(32'h3921748c),
	.w6(32'h3a97b498),
	.w7(32'h3aae04dd),
	.w8(32'h3a515e3f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d594e0),
	.w1(32'h37435df2),
	.w2(32'hb6dd2b07),
	.w3(32'h368a7f21),
	.w4(32'h3798ef50),
	.w5(32'h3546e78a),
	.w6(32'hb5fd8d1d),
	.w7(32'h37867c34),
	.w8(32'h36541350),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57949d7),
	.w1(32'hb6b9a118),
	.w2(32'hb63c801b),
	.w3(32'h34dbd3d5),
	.w4(32'hb5fc8ae6),
	.w5(32'hb6eb2183),
	.w6(32'h36b01e32),
	.w7(32'h35ee497b),
	.w8(32'hb69f2fb8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bcab9e),
	.w1(32'h3885875b),
	.w2(32'hb9f7d4ab),
	.w3(32'h38eb81ab),
	.w4(32'h399aee29),
	.w5(32'hb94293c7),
	.w6(32'h39074975),
	.w7(32'h39dbd416),
	.w8(32'hb73b7a1a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a75270),
	.w1(32'h39434628),
	.w2(32'hbab4be41),
	.w3(32'h39fafca9),
	.w4(32'h3a149072),
	.w5(32'hba755285),
	.w6(32'h39f2912b),
	.w7(32'h3a2d097f),
	.w8(32'hb9dde1a0),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3605bdef),
	.w1(32'hb70521e4),
	.w2(32'hba2d0a93),
	.w3(32'h39a340b5),
	.w4(32'h39c7c7b3),
	.w5(32'hb90e3598),
	.w6(32'h39ba8a68),
	.w7(32'h39f5c272),
	.w8(32'h388747cf),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38502f40),
	.w1(32'hb84eb203),
	.w2(32'hb717227f),
	.w3(32'h383121db),
	.w4(32'hb8234883),
	.w5(32'h3750f4e4),
	.w6(32'h383b8f2d),
	.w7(32'hb6ea36be),
	.w8(32'hb8b43915),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b7d9e7),
	.w1(32'hb5f1c1c7),
	.w2(32'h36d7ed09),
	.w3(32'h36ee3d2b),
	.w4(32'h367c897e),
	.w5(32'h369db125),
	.w6(32'h3738df0c),
	.w7(32'h36089c17),
	.w8(32'h3746cf15),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e233d5),
	.w1(32'h382abdbe),
	.w2(32'h381a3b39),
	.w3(32'h380563e7),
	.w4(32'h3825a52e),
	.w5(32'h379421f4),
	.w6(32'h3828464a),
	.w7(32'h38496f28),
	.w8(32'h37a3a10d),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394427ef),
	.w1(32'hb78b9166),
	.w2(32'h38351d6e),
	.w3(32'h3939f5e1),
	.w4(32'h3863cf7e),
	.w5(32'h38b01084),
	.w6(32'h38c1f799),
	.w7(32'h39134e8e),
	.w8(32'h38d41105),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e16a28),
	.w1(32'hb911834b),
	.w2(32'hba1eae8c),
	.w3(32'h3a08808d),
	.w4(32'h3a14f3a3),
	.w5(32'h39e9eef4),
	.w6(32'h3a4753be),
	.w7(32'h3a554c55),
	.w8(32'h3a4e7f60),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3743ca82),
	.w1(32'hb8ae5a7e),
	.w2(32'hb8dfeea7),
	.w3(32'h380c5c63),
	.w4(32'hb86bf46f),
	.w5(32'hb8f54b1a),
	.w6(32'h38dd69a0),
	.w7(32'h37ea9eed),
	.w8(32'hb8821642),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c37b80),
	.w1(32'hb8f2e11b),
	.w2(32'hb82b1aca),
	.w3(32'hb9a625b3),
	.w4(32'hb8acc4d0),
	.w5(32'hb8464f3c),
	.w6(32'hb9c8c5a4),
	.w7(32'hb93d4b04),
	.w8(32'hb9422f16),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382f4bc5),
	.w1(32'hb91e7cd6),
	.w2(32'hba1d48b8),
	.w3(32'h3916ae7a),
	.w4(32'hb83562d5),
	.w5(32'hba148cf5),
	.w6(32'h3841320e),
	.w7(32'hb91b7d0b),
	.w8(32'hba30561c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35910701),
	.w1(32'hb58115d9),
	.w2(32'h3583c545),
	.w3(32'h357efbba),
	.w4(32'hb50b2703),
	.w5(32'h35781f63),
	.w6(32'h359b397c),
	.w7(32'h35a2d0e8),
	.w8(32'h365bd315),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3640e4e3),
	.w1(32'hb4b01018),
	.w2(32'h36905a2e),
	.w3(32'h35a28d79),
	.w4(32'hb5ffe8d0),
	.w5(32'h36258f89),
	.w6(32'hb46c876a),
	.w7(32'hb51aacf6),
	.w8(32'h3666cc5b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a68599),
	.w1(32'h36c60627),
	.w2(32'h37b86b50),
	.w3(32'hb7a56aac),
	.w4(32'hb75ef86c),
	.w5(32'h36d4f8b8),
	.w6(32'h3788550c),
	.w7(32'h369c9534),
	.w8(32'h36ac74a6),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f8b836),
	.w1(32'hb5a98810),
	.w2(32'h369b48ee),
	.w3(32'h36b3b90f),
	.w4(32'h33c65ec1),
	.w5(32'h36bca08d),
	.w6(32'h36940a7e),
	.w7(32'h35893b10),
	.w8(32'h36d3a002),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85655fe),
	.w1(32'h36bc622e),
	.w2(32'h383edb36),
	.w3(32'hb876a2e2),
	.w4(32'hb70d4f33),
	.w5(32'h38869150),
	.w6(32'hb868ccc3),
	.w7(32'hb7c31986),
	.w8(32'h380a2472),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c6e402),
	.w1(32'h38a447b8),
	.w2(32'hba08f457),
	.w3(32'h39866acd),
	.w4(32'h398ce539),
	.w5(32'hb9c822fa),
	.w6(32'h39ab79ae),
	.w7(32'h39a337a4),
	.w8(32'hb92e4cae),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa10af),
	.w1(32'hb8d783ee),
	.w2(32'hb9299cc6),
	.w3(32'hb93cf36b),
	.w4(32'h388f0857),
	.w5(32'h377ec6a8),
	.w6(32'hb98488e2),
	.w7(32'hb813f9d6),
	.w8(32'hb874ea28),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370adaf1),
	.w1(32'hb585666e),
	.w2(32'h35dd3b88),
	.w3(32'h36ec59c1),
	.w4(32'hb673e653),
	.w5(32'h3516d136),
	.w6(32'h36497ae1),
	.w7(32'h365a2b12),
	.w8(32'h36a0ee19),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39907b12),
	.w1(32'h38b2010e),
	.w2(32'hba02054a),
	.w3(32'h39dadee3),
	.w4(32'h39d9dca9),
	.w5(32'hb85031dc),
	.w6(32'h3a2128ed),
	.w7(32'h3a1451bd),
	.w8(32'h39560283),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39132388),
	.w1(32'h3865d36c),
	.w2(32'hb9ce07c6),
	.w3(32'h3995f2ce),
	.w4(32'h398ff9f4),
	.w5(32'hb8c227d3),
	.w6(32'h39c0e194),
	.w7(32'h39d713a1),
	.w8(32'h38f6d25d),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36973ae6),
	.w1(32'hb6c156ed),
	.w2(32'h361dd319),
	.w3(32'h3621e805),
	.w4(32'hb6fe24e7),
	.w5(32'hb4fe25e4),
	.w6(32'h3672795c),
	.w7(32'hb6ac3a82),
	.w8(32'hb4f3b97e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f22182),
	.w1(32'hb893d352),
	.w2(32'hb9407aeb),
	.w3(32'h387e08ff),
	.w4(32'h382ef2c5),
	.w5(32'hb61bed3f),
	.w6(32'h3912285c),
	.w7(32'h391c7b67),
	.w8(32'h38fc8cfd),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370c5a1f),
	.w1(32'hb78385a6),
	.w2(32'hb7bd5d54),
	.w3(32'hb6d4b582),
	.w4(32'hb7df5a21),
	.w5(32'hb8011092),
	.w6(32'hb70efe37),
	.w7(32'hb7528923),
	.w8(32'hb7d56355),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e7631d),
	.w1(32'h3607b5ec),
	.w2(32'h37479c91),
	.w3(32'h37d8ef4b),
	.w4(32'h37ba0dc0),
	.w5(32'h37f73ab5),
	.w6(32'h36d7b936),
	.w7(32'h378a85d3),
	.w8(32'h37eef017),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a61d3a),
	.w1(32'h36a0c652),
	.w2(32'h368768e7),
	.w3(32'h3688f905),
	.w4(32'h36e65374),
	.w5(32'h368c4c53),
	.w6(32'h36b7122f),
	.w7(32'h3725e445),
	.w8(32'h36d66b2f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4a707ed),
	.w1(32'hb69ff504),
	.w2(32'hb61072ea),
	.w3(32'h3293919e),
	.w4(32'hb653e9a6),
	.w5(32'hb629912c),
	.w6(32'hb61fac85),
	.w7(32'hb50ce118),
	.w8(32'h36311300),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f95f6b),
	.w1(32'hb88a76be),
	.w2(32'h38196c65),
	.w3(32'hb8c72e9d),
	.w4(32'hb79f8830),
	.w5(32'h388e6001),
	.w6(32'hb8e54609),
	.w7(32'hb81e581e),
	.w8(32'h37efa29e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39854fe2),
	.w1(32'h3753e486),
	.w2(32'hba8cfc5d),
	.w3(32'h3a086ed4),
	.w4(32'h3a064c6a),
	.w5(32'hba047d30),
	.w6(32'h3a319e92),
	.w7(32'h3a28bdf1),
	.w8(32'hb85ef658),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c78a97),
	.w1(32'hb84f418d),
	.w2(32'hb9df538c),
	.w3(32'h39663816),
	.w4(32'h398572ae),
	.w5(32'h37a7aa63),
	.w6(32'h39a6780e),
	.w7(32'h39c110e0),
	.w8(32'h396b5fed),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c81d51),
	.w1(32'hb921004f),
	.w2(32'hba389045),
	.w3(32'h38fbc77b),
	.w4(32'h39568c2f),
	.w5(32'hb94d50fb),
	.w6(32'h39a1f635),
	.w7(32'h39f61955),
	.w8(32'h39619e42),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368d03cd),
	.w1(32'h36932490),
	.w2(32'h3617721a),
	.w3(32'h36a82004),
	.w4(32'h371a508d),
	.w5(32'h3685314c),
	.w6(32'h36a42cd3),
	.w7(32'h370c11c8),
	.w8(32'h35efd13c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d186e5),
	.w1(32'h369fffde),
	.w2(32'h37151c3a),
	.w3(32'h36897b0f),
	.w4(32'hb67758db),
	.w5(32'hb3ff7970),
	.w6(32'h36c5449c),
	.w7(32'hb5885c03),
	.w8(32'hb62e5d0d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e0cece),
	.w1(32'h379ed3a4),
	.w2(32'hb55af577),
	.w3(32'hb5008954),
	.w4(32'h378ce625),
	.w5(32'h36afee81),
	.w6(32'h36191adf),
	.w7(32'h375f52d9),
	.w8(32'h36039bbd),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3577822b),
	.w1(32'hb481b9a1),
	.w2(32'h3638f70f),
	.w3(32'h35a8074c),
	.w4(32'hb5d2acf9),
	.w5(32'h364149b1),
	.w6(32'h342e1ba7),
	.w7(32'hb612f0f0),
	.w8(32'h3532fe94),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8430fe9),
	.w1(32'hb795d9c3),
	.w2(32'hb9bb356c),
	.w3(32'h38b032ea),
	.w4(32'h390273f0),
	.w5(32'hb93a8349),
	.w6(32'h39117677),
	.w7(32'h3923228e),
	.w8(32'hb86066dc),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d0cc70),
	.w1(32'h38d19824),
	.w2(32'h37f35d35),
	.w3(32'h389a2aed),
	.w4(32'h389de245),
	.w5(32'h37b7dea1),
	.w6(32'h3791adba),
	.w7(32'h37e98d36),
	.w8(32'h375c6011),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb963d899),
	.w1(32'hb8a1ba9a),
	.w2(32'h3619f7e9),
	.w3(32'hb9679c8f),
	.w4(32'hb8e65577),
	.w5(32'hb85ffabf),
	.w6(32'hb9850f02),
	.w7(32'hb9276b5d),
	.w8(32'hb903d8be),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8307149),
	.w1(32'hb80b0ca9),
	.w2(32'hb7a340d8),
	.w3(32'hb84d90ce),
	.w4(32'hb841808e),
	.w5(32'hb8537263),
	.w6(32'hb882cde8),
	.w7(32'hb882eb76),
	.w8(32'hb86cebce),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b5b67a),
	.w1(32'h38395218),
	.w2(32'h36710067),
	.w3(32'hb5feb90b),
	.w4(32'h3783214a),
	.w5(32'hb64dcdf6),
	.w6(32'hb7c302ec),
	.w7(32'hb7c0bd4d),
	.w8(32'hb797860a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb791f73d),
	.w1(32'hb7ba2c8b),
	.w2(32'hb93ebd87),
	.w3(32'h389515c4),
	.w4(32'h38d7d14b),
	.w5(32'h360ab8df),
	.w6(32'h38b4c763),
	.w7(32'h39259cfd),
	.w8(32'h38e0fbbb),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379ebec0),
	.w1(32'h375c351d),
	.w2(32'h370f7365),
	.w3(32'h375089ea),
	.w4(32'h370860fa),
	.w5(32'h363fdb51),
	.w6(32'h36b307d6),
	.w7(32'hb4585216),
	.w8(32'hb5b5f12f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952e7a5),
	.w1(32'hb954b0e9),
	.w2(32'hb9ed41cd),
	.w3(32'hb8d84fdb),
	.w4(32'h37218d96),
	.w5(32'hb9b08fd6),
	.w6(32'h383a33af),
	.w7(32'h349d7a34),
	.w8(32'hb99d1170),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c41c77),
	.w1(32'hba9b0419),
	.w2(32'hbab7cb9f),
	.w3(32'h36ad70ee),
	.w4(32'hba87a5a2),
	.w5(32'hbacb3c50),
	.w6(32'hbaa73f8b),
	.w7(32'hbaa4c5ca),
	.w8(32'hb9c14c05),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99b69a),
	.w1(32'hba866211),
	.w2(32'hb9fd8817),
	.w3(32'hba8902fa),
	.w4(32'hba61484b),
	.w5(32'hb9384ea8),
	.w6(32'hbab49126),
	.w7(32'hba888e15),
	.w8(32'hb9d5a703),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule