module layer_10_featuremap_207(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2a690),
	.w1(32'h3a9b8675),
	.w2(32'h3d1bb0b1),
	.w3(32'hbb3f8b48),
	.w4(32'hbcb6527c),
	.w5(32'h39de9b1f),
	.w6(32'h3a9142e0),
	.w7(32'h3c6252cf),
	.w8(32'h3bef3164),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d0797),
	.w1(32'hb82c15cd),
	.w2(32'hb9d5293d),
	.w3(32'h3c23f2bb),
	.w4(32'hbaa6dc88),
	.w5(32'hbb9704c4),
	.w6(32'h3b6d1280),
	.w7(32'h3bc5cd8c),
	.w8(32'h3b2e8f5d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b407651),
	.w1(32'hb86d9b37),
	.w2(32'hbb86e00c),
	.w3(32'h3aa334fc),
	.w4(32'h3b870dfa),
	.w5(32'h3b47569b),
	.w6(32'hb944d6bc),
	.w7(32'hbb792171),
	.w8(32'hbb5257b9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7584d),
	.w1(32'hbb182438),
	.w2(32'h3b8f1391),
	.w3(32'h3b2c3e8d),
	.w4(32'hbc22f1d7),
	.w5(32'hbc9b39c8),
	.w6(32'h3afdb3a2),
	.w7(32'h3a7a8016),
	.w8(32'h3aaac9b8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab41d1e),
	.w1(32'hbc55cd86),
	.w2(32'hbc7e9f32),
	.w3(32'hbc8a535b),
	.w4(32'hbbec99b2),
	.w5(32'hbc914a4f),
	.w6(32'hbc042093),
	.w7(32'hbb21b714),
	.w8(32'h3be06663),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f4a04a),
	.w1(32'h3b7f33b2),
	.w2(32'h3b3565c9),
	.w3(32'hbc4fccbf),
	.w4(32'hbba6201e),
	.w5(32'hbc163c94),
	.w6(32'h3c160727),
	.w7(32'h3c115ea3),
	.w8(32'h3bdbd36a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd3502),
	.w1(32'hbae48075),
	.w2(32'hbbbb5f98),
	.w3(32'hbbbfbe94),
	.w4(32'h3b270694),
	.w5(32'hbb6d48ee),
	.w6(32'hba5dbb94),
	.w7(32'hb93b38a8),
	.w8(32'hbab7bbce),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6733c),
	.w1(32'hba8f4da9),
	.w2(32'hbb65fd81),
	.w3(32'hba781313),
	.w4(32'h3aca9e75),
	.w5(32'h39d0f3b8),
	.w6(32'hb940efa4),
	.w7(32'hbbdee46a),
	.w8(32'hbb994c14),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb859fe0),
	.w1(32'hbb029778),
	.w2(32'hba09da10),
	.w3(32'hbb41a4f8),
	.w4(32'hbba56468),
	.w5(32'hbb59e4e1),
	.w6(32'hbaa0e4c8),
	.w7(32'h3ae00ce9),
	.w8(32'hbaebda2f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37bce3),
	.w1(32'h3a813b52),
	.w2(32'hba4df627),
	.w3(32'hbaa8c086),
	.w4(32'hbaf93f23),
	.w5(32'hbb59c58b),
	.w6(32'h3ad74741),
	.w7(32'h3bc6b3a5),
	.w8(32'h3a9098a7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39490197),
	.w1(32'hba8c0d8d),
	.w2(32'h39b3dde6),
	.w3(32'h3b1290db),
	.w4(32'h3bc6a329),
	.w5(32'h3c65ba82),
	.w6(32'h3bd8e6aa),
	.w7(32'h3bd9d3bc),
	.w8(32'h3b03b4e5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8b3f8),
	.w1(32'hbc9ffd36),
	.w2(32'hbc950340),
	.w3(32'h3c03e757),
	.w4(32'hbc9702ac),
	.w5(32'hbcda8ce3),
	.w6(32'hbc57c919),
	.w7(32'hbc26c24c),
	.w8(32'hbc1feae4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc844022),
	.w1(32'hbb293cf4),
	.w2(32'hbb49db44),
	.w3(32'hbc91b693),
	.w4(32'h3b1c89d5),
	.w5(32'h3ad3ad0f),
	.w6(32'hb97fd0cf),
	.w7(32'hbb840c3e),
	.w8(32'h39f39e5c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d9a6c),
	.w1(32'h3acba8c9),
	.w2(32'hbb63889d),
	.w3(32'hb8b9068c),
	.w4(32'h3bdf8c09),
	.w5(32'h3c4b9838),
	.w6(32'hb9f29816),
	.w7(32'hbc326a3e),
	.w8(32'hbc61126b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe9143),
	.w1(32'hbca5f323),
	.w2(32'hbc389af6),
	.w3(32'h3bad631d),
	.w4(32'hbbd07aae),
	.w5(32'hbc9d6339),
	.w6(32'hbc04e081),
	.w7(32'hbaa5e708),
	.w8(32'h3b1303d6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b6382),
	.w1(32'hbaf91cc5),
	.w2(32'hba835ea7),
	.w3(32'hbc0a9a8d),
	.w4(32'hbc001259),
	.w5(32'hbbdfb195),
	.w6(32'h394923ab),
	.w7(32'h3b7a7383),
	.w8(32'h3a22fe7e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6dfde),
	.w1(32'hbabd89eb),
	.w2(32'h3a7000d6),
	.w3(32'hbb5207dc),
	.w4(32'h3a09f50f),
	.w5(32'h3bdff517),
	.w6(32'hbb9aeaf2),
	.w7(32'hbb69cf94),
	.w8(32'h3ac9582f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baec6e4),
	.w1(32'hbb618f96),
	.w2(32'hbbc66682),
	.w3(32'h3addb943),
	.w4(32'h371c97a8),
	.w5(32'hbb3a2f2e),
	.w6(32'hbb8ce53c),
	.w7(32'hbadc30f6),
	.w8(32'hbbb2a5de),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9f0fc),
	.w1(32'hbb152d88),
	.w2(32'hba80b753),
	.w3(32'hbb6dffb0),
	.w4(32'h3a062ba2),
	.w5(32'hbae01a86),
	.w6(32'hba8b2646),
	.w7(32'hbb04fd67),
	.w8(32'hb9feca92),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5920b1),
	.w1(32'h387bbc2a),
	.w2(32'hbab1eb8f),
	.w3(32'hba6e1667),
	.w4(32'hbb6072cb),
	.w5(32'hbad4a07a),
	.w6(32'hba1d7cbd),
	.w7(32'h39a5d757),
	.w8(32'hbb25b3f3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60ff43),
	.w1(32'hbb3183ba),
	.w2(32'hbc01d2c6),
	.w3(32'h3955950d),
	.w4(32'hba60de22),
	.w5(32'hbadd6d88),
	.w6(32'h39830ad8),
	.w7(32'hbb6a8bad),
	.w8(32'hbb56bf60),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb06396),
	.w1(32'hbc80f533),
	.w2(32'hbb81d53b),
	.w3(32'h391ce0f6),
	.w4(32'h38e174ba),
	.w5(32'hbc221219),
	.w6(32'hbba1d439),
	.w7(32'hbc1f4c4d),
	.w8(32'hba8fc714),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f8e32),
	.w1(32'h3b46b640),
	.w2(32'hbb683d62),
	.w3(32'hbc1beadb),
	.w4(32'hbb6ee0b4),
	.w5(32'hbb8a3a36),
	.w6(32'h3bc3aacf),
	.w7(32'hba83e8c6),
	.w8(32'hbaa2508a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25e3d0),
	.w1(32'h3b02abdf),
	.w2(32'h3ab6c7eb),
	.w3(32'hbb84d8dc),
	.w4(32'h3afb87cd),
	.w5(32'h3b59337d),
	.w6(32'h3b34c78d),
	.w7(32'hbb3777bc),
	.w8(32'hbb2f6323),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a51f7),
	.w1(32'hbbe96c64),
	.w2(32'hbae7d4c3),
	.w3(32'h3aa89211),
	.w4(32'hbc17c0e7),
	.w5(32'hbc270053),
	.w6(32'h3b8152b6),
	.w7(32'h3c2844b0),
	.w8(32'h3bf1554a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f2a0e),
	.w1(32'hbbdc64e1),
	.w2(32'hbb9910e8),
	.w3(32'h39620394),
	.w4(32'hba3c4c29),
	.w5(32'hbb474083),
	.w6(32'hbbdff166),
	.w7(32'hbbecf02f),
	.w8(32'hbbc6c3a6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c6417),
	.w1(32'h3a596a28),
	.w2(32'hbade0cd3),
	.w3(32'hbc111db8),
	.w4(32'hbafe4e43),
	.w5(32'hba91a5bc),
	.w6(32'hb9594e87),
	.w7(32'h39dff886),
	.w8(32'hba4ab7a5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb085cd1),
	.w1(32'hbc1e80fe),
	.w2(32'hbba409e3),
	.w3(32'hba277dd7),
	.w4(32'hbc2c5b65),
	.w5(32'hbc5eb966),
	.w6(32'hba57bf81),
	.w7(32'h3c33fb88),
	.w8(32'h3a5600c3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0a51a),
	.w1(32'hb969d4e9),
	.w2(32'hbc14a4cf),
	.w3(32'hbbab5bc9),
	.w4(32'hba025b92),
	.w5(32'hbadb37f5),
	.w6(32'h3bc2b73d),
	.w7(32'hbae0decd),
	.w8(32'h3b12d570),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eea96),
	.w1(32'hbb523a6f),
	.w2(32'hbb0afed0),
	.w3(32'hbb021fbe),
	.w4(32'hb92e72c0),
	.w5(32'h3b830d6e),
	.w6(32'hba9ab292),
	.w7(32'hba1ef659),
	.w8(32'h3b3e7d41),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb351d47),
	.w1(32'h392a753c),
	.w2(32'hbb393fff),
	.w3(32'h3ba0404f),
	.w4(32'h3b0b70c5),
	.w5(32'h3b1b243f),
	.w6(32'h3b0cd861),
	.w7(32'h390e8f6c),
	.w8(32'h3a778f30),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d178d),
	.w1(32'h38ddd699),
	.w2(32'h390976aa),
	.w3(32'h3b140194),
	.w4(32'hba2dd212),
	.w5(32'hba18b1c2),
	.w6(32'h3b605732),
	.w7(32'h3a93fe15),
	.w8(32'h3ace1eda),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378f13df),
	.w1(32'hb9d1bd60),
	.w2(32'h3b88ea1b),
	.w3(32'h39e69456),
	.w4(32'hbb3550bb),
	.w5(32'h3bac7494),
	.w6(32'h3b94fec9),
	.w7(32'h3b29434e),
	.w8(32'hbbf01410),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2875e2),
	.w1(32'hbba63139),
	.w2(32'hbc6a8a97),
	.w3(32'hbac2a583),
	.w4(32'hbc004323),
	.w5(32'hbc45dfcc),
	.w6(32'hbc515796),
	.w7(32'hbc637c88),
	.w8(32'h3ba53fbf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfd10b),
	.w1(32'hbb8cf8f4),
	.w2(32'hbb993943),
	.w3(32'hbc5106f0),
	.w4(32'hbbc151cb),
	.w5(32'hbc1ed1f1),
	.w6(32'h3a982ec5),
	.w7(32'h3c147dea),
	.w8(32'h3bd7ffcb),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b398272),
	.w1(32'hbb217f03),
	.w2(32'hba7d66ec),
	.w3(32'hbb054b8a),
	.w4(32'hbada2526),
	.w5(32'hb9db38f5),
	.w6(32'h3abb1e6e),
	.w7(32'h38efb257),
	.w8(32'hba529fc1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75cb73),
	.w1(32'hbbed0244),
	.w2(32'hbbd6d760),
	.w3(32'hbac927d6),
	.w4(32'hbb92aed3),
	.w5(32'hbc78a4a6),
	.w6(32'hbb5c81cd),
	.w7(32'h3b8e0906),
	.w8(32'h3b739c2d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a678e3),
	.w1(32'hbaa6d7c4),
	.w2(32'hbb5d784e),
	.w3(32'hbc33f38d),
	.w4(32'h3a1be832),
	.w5(32'hbad51cc0),
	.w6(32'h3a8a7474),
	.w7(32'h3b21fac2),
	.w8(32'h3ab7a32e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99957a0),
	.w1(32'h3ab6db7a),
	.w2(32'h3af32b78),
	.w3(32'h39b0f921),
	.w4(32'hba6bbef5),
	.w5(32'h3a9a63bb),
	.w6(32'h3b56d81c),
	.w7(32'h39d4fe0b),
	.w8(32'hba234837),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a7335),
	.w1(32'hbaec3522),
	.w2(32'hbb7cf9eb),
	.w3(32'h3a12f7fe),
	.w4(32'hba4f2b2c),
	.w5(32'hbbaf30bc),
	.w6(32'hba06db35),
	.w7(32'h3adbf9e7),
	.w8(32'h3ae11257),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ebf9fb),
	.w1(32'hbb942092),
	.w2(32'hbbd6f91b),
	.w3(32'hbb3526df),
	.w4(32'hbb20a6bc),
	.w5(32'hbaf3a4f2),
	.w6(32'hbaa2a0e8),
	.w7(32'hba6a328e),
	.w8(32'h3bb86b3d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fc569),
	.w1(32'h3aa00eab),
	.w2(32'hbb1003e5),
	.w3(32'hba09429a),
	.w4(32'h3af1a67d),
	.w5(32'h39e2168c),
	.w6(32'h3b23a4dc),
	.w7(32'h3a9920d3),
	.w8(32'hbb51c566),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacc8a6),
	.w1(32'h3a8b79c7),
	.w2(32'h3b950744),
	.w3(32'h3b80154c),
	.w4(32'hba815a39),
	.w5(32'h3ad02d09),
	.w6(32'h3b3acc55),
	.w7(32'h3b217cfa),
	.w8(32'h3a233708),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80913c),
	.w1(32'hba403668),
	.w2(32'hbb48fd22),
	.w3(32'hba80bdbd),
	.w4(32'h3b070667),
	.w5(32'hbb9f05ce),
	.w6(32'hbbb05966),
	.w7(32'hbaaca018),
	.w8(32'h388f65a9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba714989),
	.w1(32'h3bff1730),
	.w2(32'h3c910d4f),
	.w3(32'hbb04ada6),
	.w4(32'h3bf78c27),
	.w5(32'h3cca0f9e),
	.w6(32'h3ac27bde),
	.w7(32'hbb98b000),
	.w8(32'hbc29f6af),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd2410),
	.w1(32'h3aa13f07),
	.w2(32'hba82c85b),
	.w3(32'h3c8467c9),
	.w4(32'h3c5e31ab),
	.w5(32'h3c3333e0),
	.w6(32'hba223dea),
	.w7(32'hbbccbbe0),
	.w8(32'hb9b6f168),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5ef3c),
	.w1(32'hbc9f3868),
	.w2(32'hbc5b42a4),
	.w3(32'h3bc22f3b),
	.w4(32'hbc215f91),
	.w5(32'hbcbb7f96),
	.w6(32'hbbf0cbb1),
	.w7(32'h3a87d873),
	.w8(32'h3b427baf),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43e624),
	.w1(32'hbb13a6a5),
	.w2(32'hbb9f37fb),
	.w3(32'hbc315d71),
	.w4(32'hbbe7ee29),
	.w5(32'h3a2dc605),
	.w6(32'h3b66c42a),
	.w7(32'h3a5be27f),
	.w8(32'h3a852667),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb740ec5),
	.w1(32'hb99898a0),
	.w2(32'h3b1dd5ca),
	.w3(32'hbabe65bc),
	.w4(32'hbb16260c),
	.w5(32'hb97c9a30),
	.w6(32'h3ab24890),
	.w7(32'h3b5719dd),
	.w8(32'h3b287ba0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a174112),
	.w1(32'h3b07b215),
	.w2(32'h3a2fcc00),
	.w3(32'h37df5fd4),
	.w4(32'h3b7195d6),
	.w5(32'h3bc2864d),
	.w6(32'h3b444ded),
	.w7(32'hbb6f5b96),
	.w8(32'hbb6d4e75),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ac8bc),
	.w1(32'hbacee841),
	.w2(32'hbc2edb36),
	.w3(32'h3ac56093),
	.w4(32'h3bcdd8f9),
	.w5(32'h3ba9513a),
	.w6(32'hbbf9936d),
	.w7(32'hbc6af6ca),
	.w8(32'hbc06b10e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05f6dd),
	.w1(32'hbc342e87),
	.w2(32'hbbddd681),
	.w3(32'h3a3309e4),
	.w4(32'hbccebb90),
	.w5(32'hbcdfa230),
	.w6(32'h3b8ded5b),
	.w7(32'h3cadece6),
	.w8(32'hba1c3e73),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00f183),
	.w1(32'hbb357ca0),
	.w2(32'hbb10f009),
	.w3(32'h3a0c21b0),
	.w4(32'hbc358332),
	.w5(32'hbc6636a2),
	.w6(32'h3bda761d),
	.w7(32'h3c19f2f9),
	.w8(32'h3c06819c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ea01d),
	.w1(32'hbc32a4d8),
	.w2(32'hbc614a4b),
	.w3(32'hbbeba3f7),
	.w4(32'hbb9b911e),
	.w5(32'hbcb116f3),
	.w6(32'hbb11f04a),
	.w7(32'hbb3dd9a0),
	.w8(32'h3c0aa05b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20c8b6),
	.w1(32'hbb2745f2),
	.w2(32'h3a9cbd3c),
	.w3(32'hbc7376b8),
	.w4(32'hbba88633),
	.w5(32'hbb10e154),
	.w6(32'hba9725b5),
	.w7(32'h3b7de968),
	.w8(32'h3b40420a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3897640d),
	.w1(32'hbbc63846),
	.w2(32'hbbe72445),
	.w3(32'h3b17adc9),
	.w4(32'hbb09b2a7),
	.w5(32'hbb44e6b9),
	.w6(32'h3a64f8bc),
	.w7(32'h3a5f78ba),
	.w8(32'h3bb9a493),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd69db),
	.w1(32'hbad9a646),
	.w2(32'hbbe25b3a),
	.w3(32'hbb032331),
	.w4(32'h39b2cead),
	.w5(32'h3b73bfb2),
	.w6(32'h3a6acd2c),
	.w7(32'hbb8dcc3b),
	.w8(32'h3af32901),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3268ef),
	.w1(32'hbc996dad),
	.w2(32'hbcba407b),
	.w3(32'h3bb55df1),
	.w4(32'hbb6d3382),
	.w5(32'hbcc3df9d),
	.w6(32'hbc88801e),
	.w7(32'hbca3aa12),
	.w8(32'hb933b0a7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86a874),
	.w1(32'h3946d989),
	.w2(32'h3b4f1604),
	.w3(32'hbc18b235),
	.w4(32'hbb84d782),
	.w5(32'hbb82e6f2),
	.w6(32'h3b4fed8c),
	.w7(32'h3ba29efa),
	.w8(32'h3a98e4c2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10174e),
	.w1(32'h3a81f6aa),
	.w2(32'h3aa14bf6),
	.w3(32'h3b30355f),
	.w4(32'h378657c9),
	.w5(32'h3aec41ed),
	.w6(32'h3b187a03),
	.w7(32'hba9ac7f7),
	.w8(32'hbb443147),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffc239),
	.w1(32'hb9c162eb),
	.w2(32'hbab9aeef),
	.w3(32'h39cb1a2e),
	.w4(32'hbacc30f4),
	.w5(32'hba484b98),
	.w6(32'hbb2d7c93),
	.w7(32'hbaee05dc),
	.w8(32'hbb89c918),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf50409),
	.w1(32'h3b3c798a),
	.w2(32'h3c0bd282),
	.w3(32'h3a8a31db),
	.w4(32'h3bdf46ba),
	.w5(32'h3c18118f),
	.w6(32'h3aebf102),
	.w7(32'hb9e971f6),
	.w8(32'hb902df7f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62ff10),
	.w1(32'hbc6236c6),
	.w2(32'hbc3ca2c7),
	.w3(32'h3b423d21),
	.w4(32'hbbc1b418),
	.w5(32'hba1b03d6),
	.w6(32'hbc289a5a),
	.w7(32'hbc0fc3ab),
	.w8(32'hbc1750df),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe29ef),
	.w1(32'hba5182ee),
	.w2(32'hbacc143d),
	.w3(32'hbc2fea37),
	.w4(32'hb81a84eb),
	.w5(32'hbb98e65a),
	.w6(32'hbb4786a0),
	.w7(32'h3a706011),
	.w8(32'h3a303d6d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5688c),
	.w1(32'h3aeda9f6),
	.w2(32'h3bae714c),
	.w3(32'hbace5a8d),
	.w4(32'h3aff2902),
	.w5(32'h3bddcac9),
	.w6(32'hb90d1da2),
	.w7(32'h3b12e035),
	.w8(32'hbb62b0c6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dc418),
	.w1(32'hbb673735),
	.w2(32'hbc42dbf4),
	.w3(32'h3b1aade9),
	.w4(32'h3c5bfb87),
	.w5(32'hbc15fb09),
	.w6(32'hbc30a08b),
	.w7(32'hbc96feb9),
	.w8(32'h3bcdb6cf),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd0ab0),
	.w1(32'hbba80a25),
	.w2(32'hbb94ae64),
	.w3(32'hbc03e8f5),
	.w4(32'h3b0b83eb),
	.w5(32'h3ab1c82b),
	.w6(32'h3b035c42),
	.w7(32'h3b8c80c9),
	.w8(32'h3bfad2a8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf97366),
	.w1(32'hbb6bcef8),
	.w2(32'hbc316a43),
	.w3(32'h3b9d6588),
	.w4(32'hbb17f01a),
	.w5(32'hbbf812a2),
	.w6(32'h3b3d7583),
	.w7(32'hbb29e947),
	.w8(32'hba01d5ff),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9b3ae),
	.w1(32'hb9622a68),
	.w2(32'hba783561),
	.w3(32'hbbac285b),
	.w4(32'hbb777028),
	.w5(32'hbbb04a7c),
	.w6(32'h3b3d1b72),
	.w7(32'h3b65700c),
	.w8(32'hba4ca566),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcc33b),
	.w1(32'hbbcf0ec4),
	.w2(32'hbc9a5ee2),
	.w3(32'hbb3a6d8b),
	.w4(32'h3c75b5c8),
	.w5(32'h3c277ad4),
	.w6(32'hbc8ca7ee),
	.w7(32'hbd0008b0),
	.w8(32'hbc83465d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d83da),
	.w1(32'h39309337),
	.w2(32'hb9b62db9),
	.w3(32'hbb8aca7e),
	.w4(32'h3aaba5c1),
	.w5(32'hb9232da3),
	.w6(32'h398b1cc0),
	.w7(32'h3ad4eb7e),
	.w8(32'h3a082560),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabd917),
	.w1(32'h393d36e5),
	.w2(32'hbb2bd088),
	.w3(32'h3b4a68c6),
	.w4(32'h3acb9c89),
	.w5(32'h39f154e0),
	.w6(32'hb9df6fd8),
	.w7(32'hbb91da68),
	.w8(32'hbb0a59dc),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae3a5f),
	.w1(32'h3a9bf833),
	.w2(32'h3ab8b2c9),
	.w3(32'hba928427),
	.w4(32'hb9a0a481),
	.w5(32'h3a8617ca),
	.w6(32'h3b2f184c),
	.w7(32'h39d3c22d),
	.w8(32'hbac1b639),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba806fd3),
	.w1(32'hb9a454ac),
	.w2(32'hb942a7c2),
	.w3(32'h39d05930),
	.w4(32'hbb11f75c),
	.w5(32'h39e919c0),
	.w6(32'h3b622de4),
	.w7(32'h3a8faf97),
	.w8(32'hba82da2b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f86aa),
	.w1(32'hbb494e55),
	.w2(32'hb9ab610a),
	.w3(32'h39fe1be6),
	.w4(32'hbbc37e78),
	.w5(32'hbc01aa69),
	.w6(32'h3a4deccf),
	.w7(32'h3bde3e5a),
	.w8(32'h3aa76876),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d64607),
	.w1(32'hbc0ac2e1),
	.w2(32'hbc6efeea),
	.w3(32'h3a3db420),
	.w4(32'h3b0dd419),
	.w5(32'hbb756af3),
	.w6(32'h3ba5cc4a),
	.w7(32'h3bbc5468),
	.w8(32'hbbf50650),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98570b),
	.w1(32'hb95f29d4),
	.w2(32'hba543b32),
	.w3(32'h3bf5dcc6),
	.w4(32'h3b873667),
	.w5(32'h3bb6fe9e),
	.w6(32'h38b1caf5),
	.w7(32'hbbcffef2),
	.w8(32'hbb99fc45),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb861cbe),
	.w1(32'hba940f0d),
	.w2(32'h3b2d542f),
	.w3(32'hb9c8ef97),
	.w4(32'hbb11c3ca),
	.w5(32'h3b063de3),
	.w6(32'hbaea01bc),
	.w7(32'hbb887dda),
	.w8(32'hbbdbc5a5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dec37),
	.w1(32'hba4a8ce8),
	.w2(32'h3c17ea84),
	.w3(32'h3b5c6f4b),
	.w4(32'hbc014b7c),
	.w5(32'hba5e1c0f),
	.w6(32'h3a105993),
	.w7(32'h3a18a6e9),
	.w8(32'hbb89490b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ee196),
	.w1(32'h3a984e39),
	.w2(32'hbb470a15),
	.w3(32'h39d72085),
	.w4(32'h3a660526),
	.w5(32'h3a8071cd),
	.w6(32'h3b60524e),
	.w7(32'h39cf9c6b),
	.w8(32'h3b04bf98),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ade66),
	.w1(32'hbb7bf834),
	.w2(32'hbc23495f),
	.w3(32'h3b32ef7e),
	.w4(32'hba34724b),
	.w5(32'hbbc3cac4),
	.w6(32'h3b8e1c4b),
	.w7(32'h3a690f6f),
	.w8(32'h3bb6f1eb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92f03c),
	.w1(32'h3ba3a7f1),
	.w2(32'hbb0b632f),
	.w3(32'hbb19b596),
	.w4(32'h3ac643aa),
	.w5(32'hba8fc9f9),
	.w6(32'h3b6a5748),
	.w7(32'h3b3c4de9),
	.w8(32'hbac97ebb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94384eb),
	.w1(32'hbb44be01),
	.w2(32'hbaa174f2),
	.w3(32'hba86507d),
	.w4(32'hbb885fc4),
	.w5(32'hbb41caf6),
	.w6(32'h3abd1852),
	.w7(32'h3b6bfe39),
	.w8(32'h3b67a54a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac02898),
	.w1(32'h3a007d0e),
	.w2(32'h3bb47179),
	.w3(32'h3af91da4),
	.w4(32'hbb68dc75),
	.w5(32'hbb0fd1ad),
	.w6(32'h3ab72e63),
	.w7(32'h3b7ab0ff),
	.w8(32'h3ac6f903),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b357366),
	.w1(32'h3c448377),
	.w2(32'h39330b17),
	.w3(32'h3b7f85ba),
	.w4(32'h3a3c58f5),
	.w5(32'h3b420828),
	.w6(32'h3c0b6ce5),
	.w7(32'h3bf5edc9),
	.w8(32'h3c0c493b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c007593),
	.w1(32'h3a72f368),
	.w2(32'hbb93d914),
	.w3(32'h3a89a500),
	.w4(32'h3b9b3645),
	.w5(32'h3b9a24e0),
	.w6(32'h3a75c727),
	.w7(32'hbb23517e),
	.w8(32'hb9e587de),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bc69d),
	.w1(32'h3955b407),
	.w2(32'hbc0f21cb),
	.w3(32'h3b710cca),
	.w4(32'h39b974c5),
	.w5(32'hbbb3290e),
	.w6(32'hbbd437e5),
	.w7(32'hbc04aa43),
	.w8(32'hbbd01f6c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18cb66),
	.w1(32'h38a7e2e9),
	.w2(32'hbb0e6539),
	.w3(32'h3a50c60a),
	.w4(32'h3aaca119),
	.w5(32'h3b220de3),
	.w6(32'h3b0889a2),
	.w7(32'h3a61a2ee),
	.w8(32'h3a821c5f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e572ce),
	.w1(32'hb9108053),
	.w2(32'h3b3b3273),
	.w3(32'h3b27415d),
	.w4(32'hbb9b69a4),
	.w5(32'hbb79510d),
	.w6(32'h3b5f7d7e),
	.w7(32'h3c20aa01),
	.w8(32'h3beed94a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b962753),
	.w1(32'h3965983f),
	.w2(32'hbb0bc8e0),
	.w3(32'h3b23c24a),
	.w4(32'h3a870c7b),
	.w5(32'h39c4ccb0),
	.w6(32'h3b1ceb2b),
	.w7(32'h3a044cd5),
	.w8(32'h3ade55d4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7861fb),
	.w1(32'h3ad8ff2b),
	.w2(32'h3a1423a8),
	.w3(32'h3ad89035),
	.w4(32'h3ab1d201),
	.w5(32'h3b0e7f44),
	.w6(32'h3b8465b3),
	.w7(32'h3b2b04e0),
	.w8(32'h3a78bd38),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12c1fd),
	.w1(32'h3b848059),
	.w2(32'hbad52c91),
	.w3(32'h3aacc1ed),
	.w4(32'h3bf7b914),
	.w5(32'h3be07a6d),
	.w6(32'hba35c198),
	.w7(32'hba923cdd),
	.w8(32'hbaeec6df),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7401f8),
	.w1(32'h3a811727),
	.w2(32'h3bf3c38d),
	.w3(32'h3bd19a19),
	.w4(32'hbbab71d9),
	.w5(32'hbb95fd02),
	.w6(32'h3be173ee),
	.w7(32'h3c59e7d3),
	.w8(32'h3c1a9d92),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f36b0),
	.w1(32'hbba214bf),
	.w2(32'hbc28e8f2),
	.w3(32'h3b97d2de),
	.w4(32'hbb4f3cd1),
	.w5(32'hbbd15213),
	.w6(32'h3b4a0787),
	.w7(32'hb9afb35f),
	.w8(32'h3b80b020),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba84256),
	.w1(32'h393c886b),
	.w2(32'hbb1993f9),
	.w3(32'hbadb61e5),
	.w4(32'h3b0eb06b),
	.w5(32'hbaf39ebc),
	.w6(32'hba119dac),
	.w7(32'hbb0cf392),
	.w8(32'hbb50d3eb),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e7310),
	.w1(32'h3b43647c),
	.w2(32'h3bda0fe2),
	.w3(32'h3a37ab06),
	.w4(32'h3ad9d41d),
	.w5(32'hbc585a45),
	.w6(32'h3bce4952),
	.w7(32'h38bd9e92),
	.w8(32'h3bcc42b3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc21047),
	.w1(32'h3b8f027a),
	.w2(32'hbb933049),
	.w3(32'hbbc4b8ac),
	.w4(32'hb937d6db),
	.w5(32'hbb33ac39),
	.w6(32'h3b66f621),
	.w7(32'hbb6b1e99),
	.w8(32'hbb4f93eb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac15453),
	.w1(32'hbbf36e5f),
	.w2(32'h3b21a4b3),
	.w3(32'hbba3d384),
	.w4(32'hbc13f6db),
	.w5(32'hbbad3eec),
	.w6(32'h3aad201c),
	.w7(32'h3b5c85f3),
	.w8(32'hbc2a7010),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c9bbb),
	.w1(32'h3b1606ea),
	.w2(32'hbb939d80),
	.w3(32'hbbc38e85),
	.w4(32'h3a6aeaaf),
	.w5(32'hbb815195),
	.w6(32'h3ad6d8fc),
	.w7(32'hba2691a2),
	.w8(32'hbb843d98),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38185c37),
	.w1(32'hbbf75cb0),
	.w2(32'hbbde7a92),
	.w3(32'hbb6ca3f4),
	.w4(32'hbc4850d2),
	.w5(32'hbc846ccb),
	.w6(32'h3bb3d175),
	.w7(32'h3bf4c255),
	.w8(32'h3be03e42),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39721370),
	.w1(32'hbae532b3),
	.w2(32'hbc590d45),
	.w3(32'hbb862f42),
	.w4(32'h3c87e700),
	.w5(32'hbc470fbf),
	.w6(32'hbbbdfe44),
	.w7(32'hbc526c63),
	.w8(32'h3ba5c0ab),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8d5cf),
	.w1(32'hbb8c3732),
	.w2(32'hbc3e0c30),
	.w3(32'hbb86facb),
	.w4(32'h3c9b7c00),
	.w5(32'hbc4ae347),
	.w6(32'hbaccb159),
	.w7(32'hbc05b7d3),
	.w8(32'h3a79e4d9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbc426),
	.w1(32'hba2ad767),
	.w2(32'hbaf9e4bd),
	.w3(32'hbc15e903),
	.w4(32'h3bdabd04),
	.w5(32'h3c0a1773),
	.w6(32'hb99704cf),
	.w7(32'hbc2a48c5),
	.w8(32'hbbf089b5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2499b),
	.w1(32'hb7d5289f),
	.w2(32'hbb2941a6),
	.w3(32'hba5d2e3e),
	.w4(32'hb9731c47),
	.w5(32'hbae7690e),
	.w6(32'h3ae60e3d),
	.w7(32'hba3ab123),
	.w8(32'h3ac7c53c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca7911),
	.w1(32'hb8809300),
	.w2(32'hb902688b),
	.w3(32'hbadd556d),
	.w4(32'h3b2a2a1e),
	.w5(32'h3b7c3a46),
	.w6(32'h39c4fd11),
	.w7(32'hbb837b80),
	.w8(32'hbb66f72b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aadfd),
	.w1(32'h3ad1738b),
	.w2(32'hb9c34be8),
	.w3(32'hb9e6fc87),
	.w4(32'hbb03fe35),
	.w5(32'hba47e477),
	.w6(32'h3af0e3eb),
	.w7(32'h3ad4cb76),
	.w8(32'hbb0b0485),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43cb25),
	.w1(32'hbaae4730),
	.w2(32'hbb627a6e),
	.w3(32'hbafe0a15),
	.w4(32'h3a805a3e),
	.w5(32'hb9fc659b),
	.w6(32'h3a8b72ce),
	.w7(32'hb94e4db3),
	.w8(32'hbb323a0a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80fdcd),
	.w1(32'h3a2a4fc6),
	.w2(32'hbb348eaf),
	.w3(32'h3a8c35e7),
	.w4(32'h3b618c20),
	.w5(32'h3b93ade4),
	.w6(32'h3b28532a),
	.w7(32'h3a8e8691),
	.w8(32'hbae6d80d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dc9c3),
	.w1(32'hb99a59ed),
	.w2(32'hbaa16ccc),
	.w3(32'h3b82fa51),
	.w4(32'h3b84170e),
	.w5(32'h3b9fb91e),
	.w6(32'hb987125f),
	.w7(32'hbbc6db4e),
	.w8(32'hbb83e6ee),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e5178),
	.w1(32'h3b2c61d8),
	.w2(32'h3a5a7d65),
	.w3(32'hb9835b02),
	.w4(32'h3b817bb8),
	.w5(32'h3c3b20ca),
	.w6(32'hb9f8db09),
	.w7(32'hbbbc3cdb),
	.w8(32'hbc333d4c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79bf97),
	.w1(32'hbb1fa84d),
	.w2(32'hb824cf91),
	.w3(32'h3c446f8d),
	.w4(32'hbc078f2d),
	.w5(32'hbbd91145),
	.w6(32'h3b86d9b8),
	.w7(32'h3bdda00d),
	.w8(32'hbada0478),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91ade5),
	.w1(32'hba3e7939),
	.w2(32'h3cb4da6a),
	.w3(32'hba9ab060),
	.w4(32'hbc77c9b9),
	.w5(32'h3a05eef6),
	.w6(32'h3abcfddf),
	.w7(32'h3c329ace),
	.w8(32'hbb76b2b0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09b5d4),
	.w1(32'hbbbbe0f8),
	.w2(32'hbb2d638d),
	.w3(32'h3c3a820e),
	.w4(32'hbc317b49),
	.w5(32'hbc2cbb21),
	.w6(32'h3b964416),
	.w7(32'h3c00ffb4),
	.w8(32'h3b2c5ceb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00fa5c),
	.w1(32'h3b1ab283),
	.w2(32'hbbc77313),
	.w3(32'hbbb57894),
	.w4(32'h3b7a5d99),
	.w5(32'h3988ab1f),
	.w6(32'hba8e880c),
	.w7(32'hbb686881),
	.w8(32'hbb2fc9d0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56c8ff),
	.w1(32'h3b2231c6),
	.w2(32'h3b724a61),
	.w3(32'h3b722a8d),
	.w4(32'hba3af647),
	.w5(32'h3b204ea0),
	.w6(32'h3bd76916),
	.w7(32'h3a28c99a),
	.w8(32'h39ae03eb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2808c2),
	.w1(32'hb96e9b67),
	.w2(32'hba6cca6c),
	.w3(32'h3b814a43),
	.w4(32'h3b9978f0),
	.w5(32'h3bcfc41d),
	.w6(32'h38dcb391),
	.w7(32'hbbeb5117),
	.w8(32'hbbaedfa1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97d586),
	.w1(32'h3b64c6c6),
	.w2(32'h3adfa701),
	.w3(32'hb9e68bdb),
	.w4(32'h3b9a3eff),
	.w5(32'h3bc90b7a),
	.w6(32'h3b174a6f),
	.w7(32'hbb544ca2),
	.w8(32'hbb7f3fb7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397c88b7),
	.w1(32'h3b35eb25),
	.w2(32'h3ac1ef1c),
	.w3(32'h3acc7f11),
	.w4(32'h3b3b2abb),
	.w5(32'h3b80c905),
	.w6(32'h3b5bd0ed),
	.w7(32'hb9f935a6),
	.w8(32'hbb488ae4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20fbf0),
	.w1(32'h3b2b96b1),
	.w2(32'h3c97bbb0),
	.w3(32'hba48ff8e),
	.w4(32'h3c00cb9e),
	.w5(32'h3c74a45f),
	.w6(32'h3c01e3b1),
	.w7(32'hba27f486),
	.w8(32'hbb56c1f8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb931f8),
	.w1(32'hbb48951c),
	.w2(32'hbbd7bb52),
	.w3(32'h3be6f75d),
	.w4(32'h3c1cbc2a),
	.w5(32'hbb0ddab8),
	.w6(32'hbb9a434b),
	.w7(32'hbbf22367),
	.w8(32'h38328190),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a2f73d),
	.w1(32'h38578ddc),
	.w2(32'hbbb76a3a),
	.w3(32'hbb13529a),
	.w4(32'hbba2cfea),
	.w5(32'hbc21b133),
	.w6(32'h3b426965),
	.w7(32'hb996911a),
	.w8(32'h392c9872),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c2e7a),
	.w1(32'h39f96a40),
	.w2(32'hbb63cdc7),
	.w3(32'hbbc6fc23),
	.w4(32'hbbaff005),
	.w5(32'hbbd08f6b),
	.w6(32'h3aee1b7e),
	.w7(32'h3b61fb7a),
	.w8(32'hb81b2e17),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb786aa0),
	.w1(32'h3a9f67b7),
	.w2(32'h3adf4b83),
	.w3(32'hba679797),
	.w4(32'h3acf9eb5),
	.w5(32'h3b579331),
	.w6(32'h3b2a5854),
	.w7(32'hbb2e7142),
	.w8(32'hbb336f20),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54c157),
	.w1(32'h3c0c5ed0),
	.w2(32'h3ccdaf72),
	.w3(32'h3a9f5354),
	.w4(32'h3bdf598a),
	.w5(32'h3c066a65),
	.w6(32'h3c708946),
	.w7(32'h3c1a9d9a),
	.w8(32'h3c4d6aca),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21cc0c),
	.w1(32'h3a7d5371),
	.w2(32'hba404238),
	.w3(32'h3bdd01b9),
	.w4(32'hbc22da6e),
	.w5(32'hbc794fbd),
	.w6(32'h3c25fa60),
	.w7(32'h3c584ac0),
	.w8(32'h3c80e91b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbc952),
	.w1(32'hba722fb1),
	.w2(32'hbb524907),
	.w3(32'hbc17482e),
	.w4(32'h3a3b17ed),
	.w5(32'h3b74bca5),
	.w6(32'h3b493057),
	.w7(32'h3b238fbe),
	.w8(32'h39fa2974),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb119c05),
	.w1(32'hb5fa4680),
	.w2(32'hb5981fcf),
	.w3(32'h3b308a2d),
	.w4(32'hb5264272),
	.w5(32'hb4d3166d),
	.w6(32'hb6476b00),
	.w7(32'hb5ec26cc),
	.w8(32'hb6277aa2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f596c1),
	.w1(32'h36ac713a),
	.w2(32'h372dd6de),
	.w3(32'hb6a016ec),
	.w4(32'h36acb5b6),
	.w5(32'h373fdd51),
	.w6(32'hb69c7aa5),
	.w7(32'hb6584f4d),
	.w8(32'hb49f8181),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb764f745),
	.w1(32'hb727f228),
	.w2(32'h355e78c8),
	.w3(32'hb6e42329),
	.w4(32'h353f4ee0),
	.w5(32'h3688306c),
	.w6(32'hb735e435),
	.w7(32'hb77a3e6a),
	.w8(32'hb7381578),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3598beee),
	.w1(32'h35200dd6),
	.w2(32'h35a97eab),
	.w3(32'hb65de49f),
	.w4(32'h35fcd547),
	.w5(32'h3546b84d),
	.w6(32'hb52b6055),
	.w7(32'hb57f464f),
	.w8(32'hb5ac12ea),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6800f4e),
	.w1(32'hb6017811),
	.w2(32'h35b4389f),
	.w3(32'hb55162ad),
	.w4(32'hb617b967),
	.w5(32'h3610e442),
	.w6(32'hb66ba40b),
	.w7(32'hb50937e5),
	.w8(32'hb625b9a1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6efad33),
	.w1(32'hb70542cd),
	.w2(32'hb6db6187),
	.w3(32'hb6898886),
	.w4(32'hb6bb3620),
	.w5(32'h3676a25f),
	.w6(32'h3595b2d6),
	.w7(32'hb6bbad9a),
	.w8(32'hb6dbdad2),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb782aee8),
	.w1(32'h35947198),
	.w2(32'h37411770),
	.w3(32'hb70e1ce3),
	.w4(32'hb6c34018),
	.w5(32'h3689f97d),
	.w6(32'h3647adda),
	.w7(32'h362cc318),
	.w8(32'hb6288aa7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb520a748),
	.w1(32'hb6fe2f29),
	.w2(32'hb690c09a),
	.w3(32'h3630745f),
	.w4(32'hb6ce3412),
	.w5(32'hb6a1a001),
	.w6(32'hb630d5d1),
	.w7(32'hb69319bc),
	.w8(32'hb7098736),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76c6b1f),
	.w1(32'hb787df70),
	.w2(32'hb6155be3),
	.w3(32'h35a0692c),
	.w4(32'h368817a1),
	.w5(32'h36919985),
	.w6(32'hb72c213a),
	.w7(32'hb79a9176),
	.w8(32'hb773f036),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361abaa4),
	.w1(32'h36418f7c),
	.w2(32'h36a344d9),
	.w3(32'h3641d989),
	.w4(32'hb63ae9cc),
	.w5(32'hb4d9c4f2),
	.w6(32'h3643ce11),
	.w7(32'h368f2a1b),
	.w8(32'h34c1a82f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76235ef),
	.w1(32'hb69a29a9),
	.w2(32'h37038aa4),
	.w3(32'hb72943cb),
	.w4(32'hb5f69f20),
	.w5(32'h36fb0bb5),
	.w6(32'hb70d32e0),
	.w7(32'hb6a0c440),
	.w8(32'hb654606b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76a32fb),
	.w1(32'hb72c8661),
	.w2(32'h34a85e62),
	.w3(32'hb7811189),
	.w4(32'hb70fe956),
	.w5(32'h3619c445),
	.w6(32'hb7e4b4bc),
	.w7(32'hb7c1ed06),
	.w8(32'hb742d4a3),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7048f9c),
	.w1(32'hb66e070d),
	.w2(32'hb6684846),
	.w3(32'hb638e847),
	.w4(32'hb5196ff9),
	.w5(32'h368876e4),
	.w6(32'hb5fa030d),
	.w7(32'hb61a5962),
	.w8(32'h36efa2bd),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365bd892),
	.w1(32'h371c405a),
	.w2(32'h35f0b1c1),
	.w3(32'h371e7d2d),
	.w4(32'h36ec9c27),
	.w5(32'h369aeb39),
	.w6(32'h3760eee1),
	.w7(32'h35c596c4),
	.w8(32'hb72960ad),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a3978b),
	.w1(32'hb54246c5),
	.w2(32'hb60ebed4),
	.w3(32'h367e0b92),
	.w4(32'hb610eb99),
	.w5(32'hb613d69c),
	.w6(32'h3632be91),
	.w7(32'hb457a269),
	.w8(32'hb5b279d4),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c9804f),
	.w1(32'h3747e9f3),
	.w2(32'h361f49f6),
	.w3(32'h375765db),
	.w4(32'h3726e4d0),
	.w5(32'hb5e2ecfe),
	.w6(32'h3756736e),
	.w7(32'h3745a666),
	.w8(32'h365e4b57),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d2a62c),
	.w1(32'hb6892477),
	.w2(32'h35f20877),
	.w3(32'hb5b58b9c),
	.w4(32'hb69ecf84),
	.w5(32'h3657d64e),
	.w6(32'h36917b82),
	.w7(32'hb6cc3dff),
	.w8(32'hb74d8e3f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7085c5e),
	.w1(32'hb5bd7513),
	.w2(32'h35a315d7),
	.w3(32'h36ce27ef),
	.w4(32'hb60b6601),
	.w5(32'hb4854154),
	.w6(32'h350579ad),
	.w7(32'h35810375),
	.w8(32'h351a3472),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h350ba57e),
	.w1(32'hb6c8e364),
	.w2(32'h357cac1c),
	.w3(32'h33d20dad),
	.w4(32'hb71c176b),
	.w5(32'hb56a2f8f),
	.w6(32'hb6802054),
	.w7(32'h368e160a),
	.w8(32'h34736f64),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb628ca55),
	.w1(32'h363f5f72),
	.w2(32'h35814d14),
	.w3(32'hb584987e),
	.w4(32'h3526c737),
	.w5(32'hb3733c26),
	.w6(32'h363ee15d),
	.w7(32'h36a810e4),
	.w8(32'h3576082e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6015866),
	.w1(32'hb43254a0),
	.w2(32'h358dfae6),
	.w3(32'h365e3e3d),
	.w4(32'hb6775f38),
	.w5(32'hb70890c0),
	.w6(32'hb60845fd),
	.w7(32'hb3a2d246),
	.w8(32'hb6a304be),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c6e7dc),
	.w1(32'hb77ebfb0),
	.w2(32'hb6abae8e),
	.w3(32'hb6c7aa48),
	.w4(32'hb7060dc9),
	.w5(32'hb6bbb73d),
	.w6(32'h377be912),
	.w7(32'h36c5d17c),
	.w8(32'h36881050),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d8a1c2),
	.w1(32'hb5776e7e),
	.w2(32'hb57f7589),
	.w3(32'h3547c1ff),
	.w4(32'hb5a8a69c),
	.w5(32'hb5507488),
	.w6(32'h344f3eaf),
	.w7(32'hb5a690d5),
	.w8(32'hb636f24b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e88658),
	.w1(32'h3629bc9c),
	.w2(32'hb7099a39),
	.w3(32'hb6931649),
	.w4(32'h35bceb02),
	.w5(32'hb66fbb02),
	.w6(32'h369666f5),
	.w7(32'hb67b9960),
	.w8(32'hb6eed9cf),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb506609e),
	.w1(32'h372ff792),
	.w2(32'hb6dc3b49),
	.w3(32'hb6a991de),
	.w4(32'h36d329b0),
	.w5(32'hb6b4302f),
	.w6(32'h36cb0770),
	.w7(32'h3524bf55),
	.w8(32'hb5497156),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75b75a8),
	.w1(32'hb7013af4),
	.w2(32'hb5abf9ad),
	.w3(32'hb6a4dfa2),
	.w4(32'hb62e4483),
	.w5(32'h3540144a),
	.w6(32'hb49cfe83),
	.w7(32'hb72f17ad),
	.w8(32'hb708d042),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37175112),
	.w1(32'h359a463f),
	.w2(32'h35a0ba76),
	.w3(32'h37894165),
	.w4(32'h372452b0),
	.w5(32'h3636fea3),
	.w6(32'h37b35add),
	.w7(32'h36f185d1),
	.w8(32'h35f43419),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6820fe3),
	.w1(32'h36ac5fae),
	.w2(32'h36f81c09),
	.w3(32'hb6bd9faf),
	.w4(32'hb5aa3cf8),
	.w5(32'h3643e02e),
	.w6(32'hb5688ab7),
	.w7(32'h365f4a88),
	.w8(32'h3617f741),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb673be64),
	.w1(32'hb68bbd60),
	.w2(32'hb4ca412b),
	.w3(32'hb6eac895),
	.w4(32'hb69fc478),
	.w5(32'hb66e6fc9),
	.w6(32'hb50efcf2),
	.w7(32'hb5cd05ba),
	.w8(32'hb5dafb27),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3763782b),
	.w1(32'h377c0161),
	.w2(32'h36f257f7),
	.w3(32'h371faa74),
	.w4(32'h37376cfe),
	.w5(32'h357c5804),
	.w6(32'h36f3f7c6),
	.w7(32'h37539238),
	.w8(32'h36cd82c2),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb667f761),
	.w1(32'h3725c74d),
	.w2(32'h3778cef8),
	.w3(32'hb706933e),
	.w4(32'hb3a22db3),
	.w5(32'h36acfc4b),
	.w6(32'hb6fbd49a),
	.w7(32'hb6f7e589),
	.w8(32'h361dd40b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b7e970),
	.w1(32'h368b86a9),
	.w2(32'h3683716a),
	.w3(32'hb60a63ff),
	.w4(32'hb3541c8e),
	.w5(32'h35fe6406),
	.w6(32'h369f9d08),
	.w7(32'h3586b85d),
	.w8(32'h367ad5fe),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d16e42),
	.w1(32'hb6719f39),
	.w2(32'hb4d75329),
	.w3(32'hb6b1a43e),
	.w4(32'hb5b2bcfa),
	.w5(32'hb45c94bf),
	.w6(32'hb63d0d36),
	.w7(32'hb6b572f1),
	.w8(32'hb6584ffe),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3525611d),
	.w1(32'h35aaf228),
	.w2(32'h35873c84),
	.w3(32'h3510795f),
	.w4(32'h3574ab9e),
	.w5(32'hb2130f87),
	.w6(32'h35c86620),
	.w7(32'h34a27bcc),
	.w8(32'h3519dec0),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61fd3ca),
	.w1(32'hb6a9d522),
	.w2(32'hb69406f5),
	.w3(32'h3630b566),
	.w4(32'hb5c76905),
	.w5(32'hb58814b4),
	.w6(32'hb63c09e0),
	.w7(32'hb7050899),
	.w8(32'hb704dbfd),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c4fbd2),
	.w1(32'h35e07f98),
	.w2(32'h36732731),
	.w3(32'hb6dd8357),
	.w4(32'h36e24856),
	.w5(32'h347d62e9),
	.w6(32'h36274ac2),
	.w7(32'h35a98e68),
	.w8(32'hb549e43b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36460fbf),
	.w1(32'h370903ad),
	.w2(32'h35afed3d),
	.w3(32'hb580b979),
	.w4(32'h36c0af42),
	.w5(32'h35535481),
	.w6(32'h367b8e3d),
	.w7(32'h365413e0),
	.w8(32'hb6705b6a),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5157684),
	.w1(32'h34abcda4),
	.w2(32'h36043b02),
	.w3(32'h358c19d1),
	.w4(32'h351bbb3d),
	.w5(32'h362bf42e),
	.w6(32'h35a4fb75),
	.w7(32'h35759599),
	.w8(32'h35a34676),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37daf114),
	.w1(32'h36afabc0),
	.w2(32'h36a2adfa),
	.w3(32'h37c19a9c),
	.w4(32'h3665d6d2),
	.w5(32'hb5123cd6),
	.w6(32'h37d7e3dd),
	.w7(32'h36cc09ef),
	.w8(32'hb6502b09),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h357259e3),
	.w1(32'hb39feb54),
	.w2(32'h35d63b11),
	.w3(32'h35ae1efe),
	.w4(32'h34d8af94),
	.w5(32'h34339ded),
	.w6(32'h34375f90),
	.w7(32'h35d78a0a),
	.w8(32'h35e4dd83),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365b2557),
	.w1(32'hb610ac63),
	.w2(32'h344a8b81),
	.w3(32'h36009ec0),
	.w4(32'hb68f6159),
	.w5(32'hb5fcada7),
	.w6(32'hb627dbb3),
	.w7(32'hb60ac150),
	.w8(32'h341d8e34),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37765ebe),
	.w1(32'h37313a3b),
	.w2(32'h35d5d47d),
	.w3(32'h370100b9),
	.w4(32'h3620ac3a),
	.w5(32'h367c284f),
	.w6(32'hb638f242),
	.w7(32'hb65667d3),
	.w8(32'h362fc4b5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35efcb83),
	.w1(32'h371e9bb3),
	.w2(32'hb6088b4d),
	.w3(32'h36b35118),
	.w4(32'h37822ac5),
	.w5(32'hb74476e5),
	.w6(32'hb72fcd34),
	.w7(32'hb7ad81c0),
	.w8(32'hb795ab8b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368b52a1),
	.w1(32'hb6512485),
	.w2(32'hb64b8a59),
	.w3(32'hb64d2bcc),
	.w4(32'hb5c72562),
	.w5(32'hb5e4d2cf),
	.w6(32'h36115a2e),
	.w7(32'hb619c4c1),
	.w8(32'hb5f48ded),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7353a51),
	.w1(32'h3694065c),
	.w2(32'h367d4b32),
	.w3(32'hb68c75d8),
	.w4(32'h35d255dd),
	.w5(32'hb49fc50b),
	.w6(32'h36ce96f7),
	.w7(32'h36a0fae2),
	.w8(32'hb4adcc5a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360808ed),
	.w1(32'h332e91ce),
	.w2(32'h33143498),
	.w3(32'h36454ec4),
	.w4(32'h35f6aa7b),
	.w5(32'h35bc3cc2),
	.w6(32'hb6e7d067),
	.w7(32'hb59bcdbc),
	.w8(32'h34d90650),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e1ec97),
	.w1(32'hb7476c4c),
	.w2(32'h3755bc9e),
	.w3(32'hb5a1b0e0),
	.w4(32'h3736a0a0),
	.w5(32'h37827f9c),
	.w6(32'h3781ad45),
	.w7(32'hb5f56008),
	.w8(32'h37b925bc),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a7b9ac),
	.w1(32'hb7050b81),
	.w2(32'hb6594827),
	.w3(32'hb66d858b),
	.w4(32'hb599987c),
	.w5(32'hb49fec46),
	.w6(32'hb7050517),
	.w7(32'hb6cc2992),
	.w8(32'hb655d7e7),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb703d872),
	.w1(32'hb7303d42),
	.w2(32'hb7333ad3),
	.w3(32'hb6896ba3),
	.w4(32'h352e489b),
	.w5(32'hb677212a),
	.w6(32'h3747826a),
	.w7(32'hb686d6ec),
	.w8(32'hb79a1091),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6573f1e),
	.w1(32'h36266e6e),
	.w2(32'h3598ab9b),
	.w3(32'h36abc679),
	.w4(32'hb60691b5),
	.w5(32'hb6bf92a8),
	.w6(32'h35ff2f0b),
	.w7(32'h33d82d8a),
	.w8(32'hb6499840),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366df046),
	.w1(32'h36148874),
	.w2(32'h34c53b07),
	.w3(32'hb69dacbe),
	.w4(32'h368e869e),
	.w5(32'hb66ed54f),
	.w6(32'hb5cde7bf),
	.w7(32'hb68b5062),
	.w8(32'hb70b81ac),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c589f2),
	.w1(32'h34ac76c0),
	.w2(32'h35079926),
	.w3(32'h3644e538),
	.w4(32'hb678c105),
	.w5(32'hb60cced4),
	.w6(32'h36125d65),
	.w7(32'h34c4d995),
	.w8(32'h3555d409),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35893920),
	.w1(32'hb6a1e7d5),
	.w2(32'hb6210f3d),
	.w3(32'h3563f908),
	.w4(32'hb6a5da9a),
	.w5(32'hb6a791c5),
	.w6(32'hb551c954),
	.w7(32'hb5d8bdf8),
	.w8(32'hb5082490),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3620ab6c),
	.w1(32'hb72cd747),
	.w2(32'hb69ca992),
	.w3(32'h35b5463c),
	.w4(32'hb67cc638),
	.w5(32'h36e3ed7d),
	.w6(32'hb706ece5),
	.w7(32'hb40926c4),
	.w8(32'h364ba7f0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74165d0),
	.w1(32'hb641c487),
	.w2(32'hb67df922),
	.w3(32'hb6a65931),
	.w4(32'hb5740d1d),
	.w5(32'hb5de0d94),
	.w6(32'h35cf8183),
	.w7(32'hb69bff5b),
	.w8(32'hb6974c56),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5200781),
	.w1(32'hb6934fc3),
	.w2(32'h360e7438),
	.w3(32'h33e3c589),
	.w4(32'hb6ca440c),
	.w5(32'h34aec248),
	.w6(32'hb64f8cfc),
	.w7(32'hb5ed1e7c),
	.w8(32'hb66c206c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb676caeb),
	.w1(32'h359c1999),
	.w2(32'hb6044c1e),
	.w3(32'hb641340b),
	.w4(32'h35ce5aa2),
	.w5(32'hb58e5765),
	.w6(32'h34f310ff),
	.w7(32'hb594771e),
	.w8(32'hb5b0e576),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34ff4de9),
	.w1(32'h36dad654),
	.w2(32'h361a45d0),
	.w3(32'hb655f857),
	.w4(32'h3453d8cc),
	.w5(32'hb48c025e),
	.w6(32'hb62b3ec0),
	.w7(32'hb6801a48),
	.w8(32'h35db2c04),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b53869),
	.w1(32'hb51df94a),
	.w2(32'h36fccc20),
	.w3(32'h359f0d51),
	.w4(32'h369739e1),
	.w5(32'h368afcb7),
	.w6(32'hb6d0ac22),
	.w7(32'hb68e9553),
	.w8(32'h36938a3a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f70af2),
	.w1(32'hb6abcc8c),
	.w2(32'h36b42e41),
	.w3(32'hb5f35679),
	.w4(32'hb75a441a),
	.w5(32'hb46e5064),
	.w6(32'hb4851535),
	.w7(32'h35028df6),
	.w8(32'h357cf38e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3666b274),
	.w1(32'h3380036b),
	.w2(32'h3592fb16),
	.w3(32'hb643e388),
	.w4(32'h35bcab3d),
	.w5(32'h359ce767),
	.w6(32'hb4db658b),
	.w7(32'h3356c4ec),
	.w8(32'h366f01e5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7602d93),
	.w1(32'hb757f14f),
	.w2(32'h36675ee8),
	.w3(32'h3614dcc1),
	.w4(32'hb58f55bb),
	.w5(32'hb7b5d125),
	.w6(32'h37a80a9e),
	.w7(32'h35ee170f),
	.w8(32'hb501de57),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ce44ad),
	.w1(32'h379479a8),
	.w2(32'h3775ab6e),
	.w3(32'h36cc61c0),
	.w4(32'h37ace35d),
	.w5(32'h3787ce37),
	.w6(32'h35925b18),
	.w7(32'h3735dd7d),
	.w8(32'h3729bf0f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb610281e),
	.w1(32'hb54ddf84),
	.w2(32'h35c51b48),
	.w3(32'h350b7056),
	.w4(32'hb64c4ed8),
	.w5(32'hb53b6df9),
	.w6(32'h3604c375),
	.w7(32'h35cf6897),
	.w8(32'h35ed63a5),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3635492a),
	.w1(32'hb69eadbd),
	.w2(32'hb619ba0b),
	.w3(32'hb51be0c5),
	.w4(32'hb6c70070),
	.w5(32'hb7251328),
	.w6(32'hb605a8b0),
	.w7(32'h357fdf08),
	.w8(32'h353e9004),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb651a773),
	.w1(32'hb60f98f0),
	.w2(32'hb551442e),
	.w3(32'hb7361b3b),
	.w4(32'hb5259868),
	.w5(32'h344a549c),
	.w6(32'hb6ca32cc),
	.w7(32'hb50c0d43),
	.w8(32'h35889a92),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4c51f63),
	.w1(32'h33a1d069),
	.w2(32'hb59c617e),
	.w3(32'hb42c5b92),
	.w4(32'h359cd11a),
	.w5(32'hb6263713),
	.w6(32'h35063fc5),
	.w7(32'h34464354),
	.w8(32'hb490c709),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e8259e),
	.w1(32'hb3bec9e1),
	.w2(32'h36ee8024),
	.w3(32'h3542fa4b),
	.w4(32'hb6d6ca61),
	.w5(32'h36c43f7d),
	.w6(32'hb69af04f),
	.w7(32'h35f38f7d),
	.w8(32'h362009e5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ec5353),
	.w1(32'hb71259f9),
	.w2(32'hb5f8b476),
	.w3(32'hb68d295c),
	.w4(32'hb70337d0),
	.w5(32'hb5bde54c),
	.w6(32'hb6f84296),
	.w7(32'hb7b0ac42),
	.w8(32'hb6eba801),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63f9d16),
	.w1(32'h36177582),
	.w2(32'hb6db2c8b),
	.w3(32'hb68d7775),
	.w4(32'hb6916ede),
	.w5(32'hb7375fe4),
	.w6(32'h37245c7e),
	.w7(32'hb6e8c84d),
	.w8(32'h34c771f5),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5922755),
	.w1(32'hb542ad10),
	.w2(32'hb4f3160a),
	.w3(32'hb6c3303d),
	.w4(32'hb4d01d22),
	.w5(32'h3405ac16),
	.w6(32'hb55e2dbe),
	.w7(32'hb591e563),
	.w8(32'hb569f362),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72dc7fb),
	.w1(32'hb70ee888),
	.w2(32'hb6955881),
	.w3(32'hb69ce978),
	.w4(32'hb729c993),
	.w5(32'hb74b5a12),
	.w6(32'hb57575e3),
	.w7(32'hb6b24387),
	.w8(32'hb702a0bd),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61b0e9f),
	.w1(32'hb60f9f2a),
	.w2(32'h3660f1c6),
	.w3(32'hb6741c82),
	.w4(32'h34c2bf28),
	.w5(32'h368e806a),
	.w6(32'h3642646e),
	.w7(32'h365677a1),
	.w8(32'hb5a2a22e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36045afa),
	.w1(32'hb5098606),
	.w2(32'h33d02df9),
	.w3(32'h361a0fdd),
	.w4(32'hb65fd4b6),
	.w5(32'hb5a294a1),
	.w6(32'h35c9fd05),
	.w7(32'h3496919c),
	.w8(32'h341009a9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33e68490),
	.w1(32'hb6aa2953),
	.w2(32'h36217b93),
	.w3(32'hb60d9bdf),
	.w4(32'hb658b3c1),
	.w5(32'h358db354),
	.w6(32'h35408432),
	.w7(32'hb5a1af0c),
	.w8(32'h35d2424b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36040442),
	.w1(32'h355065fe),
	.w2(32'h35aca578),
	.w3(32'h358fc7c7),
	.w4(32'hb48cf616),
	.w5(32'h342d984d),
	.w6(32'h36304062),
	.w7(32'h35f3dcc7),
	.w8(32'h358443c9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6131e44),
	.w1(32'h3721b82f),
	.w2(32'hb6a374d1),
	.w3(32'hb4e6ebf9),
	.w4(32'h373b3c21),
	.w5(32'h371e67eb),
	.w6(32'h36993623),
	.w7(32'h37460612),
	.w8(32'hb69d2f96),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37039635),
	.w1(32'hb631ba37),
	.w2(32'hb68791da),
	.w3(32'h36e01f9c),
	.w4(32'h373f5978),
	.w5(32'h376f7ba6),
	.w6(32'h36987eca),
	.w7(32'hb5ff51f6),
	.w8(32'hb6126d89),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f0187c),
	.w1(32'h35c9f6d7),
	.w2(32'h35d226e4),
	.w3(32'h36f2eb02),
	.w4(32'hb6121c81),
	.w5(32'h34613f22),
	.w6(32'h355d49b8),
	.w7(32'hb5c2cd2e),
	.w8(32'hb5aa89e2),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36479a67),
	.w1(32'h35294e30),
	.w2(32'h364c5a33),
	.w3(32'hb6a32db2),
	.w4(32'hb39cb96d),
	.w5(32'h35c47f1c),
	.w6(32'hb6a59b4e),
	.w7(32'hb64e8bd9),
	.w8(32'h34a833c3),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3662697d),
	.w1(32'h37317cfb),
	.w2(32'h36e2c5c8),
	.w3(32'h3659b029),
	.w4(32'h369fe816),
	.w5(32'hb539791a),
	.w6(32'h366207d4),
	.w7(32'h36d7f744),
	.w8(32'hb60eca05),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f2e42e),
	.w1(32'h36b86dab),
	.w2(32'hb5cc0ce8),
	.w3(32'h362c1cba),
	.w4(32'h362ae482),
	.w5(32'hb6d51a12),
	.w6(32'h36e6eda7),
	.w7(32'hb6785a6d),
	.w8(32'hb70d5f50),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7921eba),
	.w1(32'hb621373a),
	.w2(32'hb6bdeba5),
	.w3(32'h34fcabd7),
	.w4(32'h36f9cd17),
	.w5(32'hb7a2fc99),
	.w6(32'h37a548ac),
	.w7(32'hb6525bf3),
	.w8(32'hb6a29b4e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h352a922d),
	.w1(32'hb6722aeb),
	.w2(32'hb67e30f2),
	.w3(32'hb69fddde),
	.w4(32'hb6204d9a),
	.w5(32'hb6138f9d),
	.w6(32'hb6173983),
	.w7(32'hb66a95b4),
	.w8(32'h33d9a628),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5313bd0),
	.w1(32'h358d6085),
	.w2(32'h35a0f9e1),
	.w3(32'hb4e42e35),
	.w4(32'h3555cbed),
	.w5(32'hb33bdd77),
	.w6(32'h35f0e58e),
	.w7(32'h36150ea8),
	.w8(32'h361374a9),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66edf8a),
	.w1(32'hb664db4f),
	.w2(32'h36aec2d1),
	.w3(32'h353e86af),
	.w4(32'h36aa5b8a),
	.w5(32'h36fdf5f9),
	.w6(32'hb6c35003),
	.w7(32'hb6f77075),
	.w8(32'h35cfac1d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71445fc),
	.w1(32'hb68dd1f8),
	.w2(32'hb6e5d4dc),
	.w3(32'h35225585),
	.w4(32'h3731a7c7),
	.w5(32'h3661ff4f),
	.w6(32'hb67e2021),
	.w7(32'hb7529258),
	.w8(32'hb78bc824),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c68e03),
	.w1(32'h36bdf625),
	.w2(32'h34475a67),
	.w3(32'hb65a3a14),
	.w4(32'h35bc0245),
	.w5(32'hb66d4c07),
	.w6(32'hb69a956a),
	.w7(32'hb6b50bf0),
	.w8(32'hb67f75b8),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36940ec0),
	.w1(32'hb666c0ec),
	.w2(32'h36657692),
	.w3(32'h3654f635),
	.w4(32'h36ae6345),
	.w5(32'h3736dfd4),
	.w6(32'h369d8d4f),
	.w7(32'h3630fcde),
	.w8(32'h3391c7c4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59d085e),
	.w1(32'h35b488b7),
	.w2(32'h35af4d73),
	.w3(32'hb55cef98),
	.w4(32'h350b4fc4),
	.w5(32'h34ea7547),
	.w6(32'h35946d6f),
	.w7(32'h34c94b07),
	.w8(32'hb4dd8d00),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d49daf),
	.w1(32'hb5f6e943),
	.w2(32'hb631076f),
	.w3(32'hb599f2dd),
	.w4(32'h3480bfff),
	.w5(32'hb6902e87),
	.w6(32'hb54615ff),
	.w7(32'h34027167),
	.w8(32'hb5d7bcf9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb43d82d7),
	.w1(32'hb6a5ff26),
	.w2(32'h3568cf7d),
	.w3(32'hb656d9cd),
	.w4(32'hb67659e0),
	.w5(32'h359c0474),
	.w6(32'hb6629867),
	.w7(32'hb753f523),
	.w8(32'hb7196cb6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fd5fdd),
	.w1(32'hb7cb1a09),
	.w2(32'hb6ca0ee6),
	.w3(32'hb78a0063),
	.w4(32'hb763e087),
	.w5(32'hb71656d3),
	.w6(32'hb72be0d7),
	.w7(32'hb799c429),
	.w8(32'hb69b4be7),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4dcac37),
	.w1(32'hb6ad55c8),
	.w2(32'hb6833a98),
	.w3(32'h36248f4a),
	.w4(32'hb4c7c7e9),
	.w5(32'hb7150fb2),
	.w6(32'hb6cde9ce),
	.w7(32'hb747a488),
	.w8(32'hb7746655),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb463b3cd),
	.w1(32'h3479869a),
	.w2(32'h36e8faa5),
	.w3(32'h36698ecf),
	.w4(32'h36e081be),
	.w5(32'h3732a14b),
	.w6(32'hb62e5771),
	.w7(32'h3658809a),
	.w8(32'h36d3a3e5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb640db13),
	.w1(32'h36e3301a),
	.w2(32'hb6a60ffc),
	.w3(32'hb661e03a),
	.w4(32'h36a65902),
	.w5(32'hb725a0c0),
	.w6(32'hb485dc76),
	.w7(32'hb6da0060),
	.w8(32'hb5a392c4),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h357d4eb4),
	.w1(32'hb5acf0d1),
	.w2(32'hb5d81ecd),
	.w3(32'hb65668d1),
	.w4(32'hb4a8a79f),
	.w5(32'hb56b33a6),
	.w6(32'hb4a789f3),
	.w7(32'hb583385f),
	.w8(32'hb5e11d7f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6432b43),
	.w1(32'hb52bbdf6),
	.w2(32'hb5c5b447),
	.w3(32'hb6162002),
	.w4(32'hb4d550cf),
	.w5(32'hb50ddf90),
	.w6(32'hb5aa4513),
	.w7(32'hb66ca131),
	.w8(32'hb6355671),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360282df),
	.w1(32'h36eea527),
	.w2(32'hb68b6582),
	.w3(32'hb62727b2),
	.w4(32'h36a19fff),
	.w5(32'hb6c57fae),
	.w6(32'h36a78f24),
	.w7(32'hb6ef19cf),
	.w8(32'h365b1a90),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3635b689),
	.w1(32'hb6ba5ed6),
	.w2(32'hb54a480a),
	.w3(32'hb596b8dd),
	.w4(32'hb62abe27),
	.w5(32'hb5c4939d),
	.w6(32'hb6203834),
	.w7(32'h36ac34b5),
	.w8(32'hb61b3eae),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c379e1),
	.w1(32'hb4ffa803),
	.w2(32'hb5732366),
	.w3(32'hb65f1e68),
	.w4(32'h34fbd203),
	.w5(32'h357404ce),
	.w6(32'hb5f2c383),
	.w7(32'hb683bc48),
	.w8(32'hb6286807),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72e977b),
	.w1(32'h3715c963),
	.w2(32'hb73fc5b7),
	.w3(32'hb689f253),
	.w4(32'h370576fb),
	.w5(32'hb6e760f6),
	.w6(32'h35d9d5e6),
	.w7(32'hb72a8793),
	.w8(32'hb794567f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6517fda),
	.w1(32'hb42b2d90),
	.w2(32'h3728ca52),
	.w3(32'hb6925234),
	.w4(32'hb6ae4e9b),
	.w5(32'h36d114f5),
	.w6(32'hb70287cf),
	.w7(32'h3689ea54),
	.w8(32'hb67362bd),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb50a40df),
	.w1(32'hb6ded95b),
	.w2(32'hb6ad541d),
	.w3(32'h35c5d2d8),
	.w4(32'hb73593fc),
	.w5(32'hb698b4a4),
	.w6(32'hb67dea46),
	.w7(32'h3614e849),
	.w8(32'h36d0ee31),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72b403c),
	.w1(32'hb78dc350),
	.w2(32'hb6d80a44),
	.w3(32'hb76bc53b),
	.w4(32'hb75268fb),
	.w5(32'hb6ce36aa),
	.w6(32'hb735f635),
	.w7(32'hb78aa077),
	.w8(32'hb7945e98),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b738f3),
	.w1(32'hb55179dd),
	.w2(32'hb668f841),
	.w3(32'h35dfd6fe),
	.w4(32'hb5a583c7),
	.w5(32'hb6eee9b8),
	.w6(32'h3718f446),
	.w7(32'h360914bd),
	.w8(32'hb6d26ca2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35fd5a69),
	.w1(32'hb4faa6da),
	.w2(32'hb3908563),
	.w3(32'h35430980),
	.w4(32'hb64a4f84),
	.w5(32'hb5b1aa7b),
	.w6(32'h35107839),
	.w7(32'hb57bf2f6),
	.w8(32'hb4cd6751),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f174d8),
	.w1(32'hb6c5db42),
	.w2(32'h3643d85f),
	.w3(32'hb6ca98d0),
	.w4(32'hb6bf14e1),
	.w5(32'hb6201264),
	.w6(32'hb62ce749),
	.w7(32'hb6b3d38b),
	.w8(32'hb631d0a7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3662567c),
	.w1(32'h35c70073),
	.w2(32'hb56f70c6),
	.w3(32'h361ca6f2),
	.w4(32'h358437c9),
	.w5(32'hb581b501),
	.w6(32'hb3f46835),
	.w7(32'hb572686b),
	.w8(32'hb615e4c9),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5afba96),
	.w1(32'hb593a87b),
	.w2(32'hb547a200),
	.w3(32'hb4572a8f),
	.w4(32'hb4bedfcb),
	.w5(32'h349b066c),
	.w6(32'h36274bea),
	.w7(32'hb568705f),
	.w8(32'hb5c1ed6b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4a94641),
	.w1(32'hb46394bf),
	.w2(32'h34757c6a),
	.w3(32'h34f5f47c),
	.w4(32'hb64e3720),
	.w5(32'hb5a89225),
	.w6(32'h3559b1e4),
	.w7(32'hb531981b),
	.w8(32'hb4e1ddbc),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3587bd88),
	.w1(32'h361300ac),
	.w2(32'hb59d95b5),
	.w3(32'hb56e57bf),
	.w4(32'h369f5606),
	.w5(32'h34807e85),
	.w6(32'h3615aec4),
	.w7(32'hb502239f),
	.w8(32'hb500c313),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35fdb4f0),
	.w1(32'hb36d522b),
	.w2(32'h3650f3ea),
	.w3(32'hb6290011),
	.w4(32'hb5d7ba49),
	.w5(32'h35ec5259),
	.w6(32'hb58605c0),
	.w7(32'h367e4e96),
	.w8(32'h362c1a89),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5718606),
	.w1(32'hb443db7f),
	.w2(32'h3711ab94),
	.w3(32'hb5966150),
	.w4(32'h3695b733),
	.w5(32'h35ebf2c7),
	.w6(32'hb61f78f0),
	.w7(32'hb68e7de2),
	.w8(32'hb691d4da),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35304c84),
	.w1(32'hb68f1786),
	.w2(32'hb5d007a9),
	.w3(32'hb60233cf),
	.w4(32'hb6475dcd),
	.w5(32'hb68a636d),
	.w6(32'h3681e0dc),
	.w7(32'hb632df88),
	.w8(32'hb6d8d44c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364c22f6),
	.w1(32'h35ca7659),
	.w2(32'h36522847),
	.w3(32'h368dec65),
	.w4(32'h372632d1),
	.w5(32'h367d2119),
	.w6(32'h36b8b277),
	.w7(32'h35da2e21),
	.w8(32'h34d1891e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h338b9b94),
	.w1(32'h368c85c7),
	.w2(32'h35ff82b7),
	.w3(32'h354c7e82),
	.w4(32'h363945c4),
	.w5(32'hb5925d52),
	.w6(32'h36dbd910),
	.w7(32'h36a4eac0),
	.w8(32'h349ad77a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61fa1a2),
	.w1(32'hb4acc8c7),
	.w2(32'h34b703ec),
	.w3(32'hb66f6cfb),
	.w4(32'hb68b52bf),
	.w5(32'hb5cdb3f9),
	.w6(32'h35af5013),
	.w7(32'hb57c01d8),
	.w8(32'hb50dd3f6),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35992f66),
	.w1(32'hb5cc8485),
	.w2(32'hb584f84b),
	.w3(32'hb5aa7cdb),
	.w4(32'hb649a436),
	.w5(32'hb5ea73dd),
	.w6(32'hb330fdb1),
	.w7(32'hb5e9f93b),
	.w8(32'hb5ae94e3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3413d596),
	.w1(32'hb60a9cb8),
	.w2(32'hb5c83180),
	.w3(32'hb4cfb8cf),
	.w4(32'hb65d14eb),
	.w5(32'hb5a6dcfe),
	.w6(32'hb4d8a5d4),
	.w7(32'hb605d98e),
	.w8(32'hb5e6b3b3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7527507),
	.w1(32'hb71db21f),
	.w2(32'hb6e55908),
	.w3(32'hb73614fa),
	.w4(32'hb72f981a),
	.w5(32'hb69c6656),
	.w6(32'hb70a13b6),
	.w7(32'hb6f44216),
	.w8(32'hb6b8e828),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362d608c),
	.w1(32'hb6585d7f),
	.w2(32'h367e31f1),
	.w3(32'hb6542bb9),
	.w4(32'hb685a2aa),
	.w5(32'h35de6103),
	.w6(32'hb6367829),
	.w7(32'h3675bb7f),
	.w8(32'h336420b1),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bf1c53),
	.w1(32'hb68b1b0d),
	.w2(32'hb5e69440),
	.w3(32'hb68c4d58),
	.w4(32'hb6cd2456),
	.w5(32'hb618f1f1),
	.w6(32'hb7247c42),
	.w7(32'hb771385f),
	.w8(32'hb68b290d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb55326b9),
	.w1(32'hb5c498af),
	.w2(32'h35ae2e62),
	.w3(32'hb621e23d),
	.w4(32'h3583f996),
	.w5(32'h33513883),
	.w6(32'hb67c833f),
	.w7(32'hb521cd13),
	.w8(32'hb418c609),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4da1911),
	.w1(32'h34921a74),
	.w2(32'h352255f5),
	.w3(32'h349167ef),
	.w4(32'hb5d2c3d1),
	.w5(32'hb583504a),
	.w6(32'h361fc30c),
	.w7(32'h3569c711),
	.w8(32'h359468f4),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60653bf),
	.w1(32'h368c508a),
	.w2(32'h352c641c),
	.w3(32'hb57687a2),
	.w4(32'h363c64ba),
	.w5(32'hb47d3f5b),
	.w6(32'hb61911fe),
	.w7(32'hb59240ed),
	.w8(32'h367fd99f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e49da5),
	.w1(32'h36809d2b),
	.w2(32'h359e030f),
	.w3(32'hb680e634),
	.w4(32'h3643287b),
	.w5(32'h3572761c),
	.w6(32'h365dbc73),
	.w7(32'h356688fd),
	.w8(32'h3654d984),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7114f1e),
	.w1(32'hb6c5bd38),
	.w2(32'h35afe08c),
	.w3(32'hb72929ae),
	.w4(32'hb6abd1ed),
	.w5(32'h33888896),
	.w6(32'hb770fae6),
	.w7(32'hb78421e4),
	.w8(32'hb630aaa4),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h359c0e69),
	.w1(32'hb9d29179),
	.w2(32'hb94dcbec),
	.w3(32'h35cc7c9b),
	.w4(32'hba4106ef),
	.w5(32'hb9b1d372),
	.w6(32'hb96430a4),
	.w7(32'hb9e90d7b),
	.w8(32'h379e0016),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cfdcc1),
	.w1(32'hb8b62728),
	.w2(32'h3918631a),
	.w3(32'hba262734),
	.w4(32'hb8647b4d),
	.w5(32'h39135559),
	.w6(32'hb9caec8a),
	.w7(32'hb9893dc4),
	.w8(32'hb8648405),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule