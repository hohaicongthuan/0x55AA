module layer_10_featuremap_376(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c147a65),
	.w1(32'h3b86f70a),
	.w2(32'h3a7d56a1),
	.w3(32'hbbca106f),
	.w4(32'h3bb94210),
	.w5(32'hbc453cec),
	.w6(32'hbdb70374),
	.w7(32'hbb379f0c),
	.w8(32'hba9cdd1c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4ba190),
	.w1(32'hbc5b83a9),
	.w2(32'hbc91d2d4),
	.w3(32'hbccc014c),
	.w4(32'hbc156397),
	.w5(32'hbb709ee0),
	.w6(32'hbc759123),
	.w7(32'h3bb627b2),
	.w8(32'hbc1eb82d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66c65b),
	.w1(32'h3b6b49f7),
	.w2(32'hbc39dc61),
	.w3(32'h3b0e7ab8),
	.w4(32'h3ae4abbf),
	.w5(32'hbb8de85d),
	.w6(32'hbc590da7),
	.w7(32'hbb6f968e),
	.w8(32'h3ba2906a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fcc3b),
	.w1(32'hbd54c099),
	.w2(32'h3b473aaa),
	.w3(32'hb9f2b088),
	.w4(32'hbc7c97c0),
	.w5(32'h3bf75d52),
	.w6(32'hbb1fc499),
	.w7(32'h3b3dac3a),
	.w8(32'hbc5d545f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba69218),
	.w1(32'hb98dbf2d),
	.w2(32'hbb9e9d56),
	.w3(32'hbcc55b97),
	.w4(32'hbb7bd338),
	.w5(32'hb9b107a2),
	.w6(32'h3c679340),
	.w7(32'h3bc11277),
	.w8(32'h3bd9d5a7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991f013),
	.w1(32'hbcaf2b1a),
	.w2(32'h3b281048),
	.w3(32'h3a876204),
	.w4(32'hbb33f001),
	.w5(32'h3c6030e0),
	.w6(32'h3b83db2a),
	.w7(32'hbab6c1fe),
	.w8(32'hbab37d41),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbde91c),
	.w1(32'hbc86e2a8),
	.w2(32'hbc82b666),
	.w3(32'h3b1bdc77),
	.w4(32'hbd68dc8f),
	.w5(32'hbce080f9),
	.w6(32'h3c2ccfe3),
	.w7(32'hbbfcaf4c),
	.w8(32'hbc586f26),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd051827),
	.w1(32'hbc91e493),
	.w2(32'h3a40b74b),
	.w3(32'hbd0a7502),
	.w4(32'hbd094fa1),
	.w5(32'hbc47177b),
	.w6(32'hbca6bd1d),
	.w7(32'hbbc82c7d),
	.w8(32'hbc72c9cf),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2c25f5),
	.w1(32'h3cee58b3),
	.w2(32'hbc4aec6b),
	.w3(32'h3b2c34fa),
	.w4(32'hbbd73ed7),
	.w5(32'hbbdf2a10),
	.w6(32'h384442ff),
	.w7(32'h3abe9452),
	.w8(32'h3b368cca),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3d43ef),
	.w1(32'h3bba685a),
	.w2(32'hbcb5b9fc),
	.w3(32'hbc998bc4),
	.w4(32'h3cea4f7a),
	.w5(32'hba09a021),
	.w6(32'hbd9dca35),
	.w7(32'h3b30650a),
	.w8(32'hbcb5fd8c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4e993),
	.w1(32'hbc5eb062),
	.w2(32'hba45f939),
	.w3(32'h3ac668e0),
	.w4(32'hbc1ed8b4),
	.w5(32'h39bc65ba),
	.w6(32'hbc6f23c7),
	.w7(32'hba103310),
	.w8(32'hbba4df3d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06ad2c),
	.w1(32'h3c33d063),
	.w2(32'hbc7c8cde),
	.w3(32'hbc07ddb6),
	.w4(32'h3a25abbc),
	.w5(32'hbcc0a657),
	.w6(32'hbc6e3f00),
	.w7(32'h3ac48917),
	.w8(32'hbcc92482),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce097a),
	.w1(32'h3af23a94),
	.w2(32'hbcc0a64a),
	.w3(32'hbc7ad9d9),
	.w4(32'hbb73e4f5),
	.w5(32'hbc014e81),
	.w6(32'hbc68e704),
	.w7(32'hbc793e2b),
	.w8(32'hbc37a532),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc899110),
	.w1(32'hbb6ed4ce),
	.w2(32'hbc63beb3),
	.w3(32'h3c172ca1),
	.w4(32'h3cbf230d),
	.w5(32'hbd155122),
	.w6(32'hbc80df40),
	.w7(32'hba36b042),
	.w8(32'hba44d3d9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaba4f),
	.w1(32'hbbed51c4),
	.w2(32'hbc9c3302),
	.w3(32'hb984d59e),
	.w4(32'h3c9f86b1),
	.w5(32'hbbb8f328),
	.w6(32'hbc1b5d5f),
	.w7(32'h3c45b9fc),
	.w8(32'hbcb99b31),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd141d6a),
	.w1(32'hbc840717),
	.w2(32'hbd02ea3f),
	.w3(32'hbc9f0ab4),
	.w4(32'h3c7ac0ad),
	.w5(32'h3b14aea7),
	.w6(32'hbc6202c3),
	.w7(32'hbc08ae7d),
	.w8(32'hbdcea314),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9665a),
	.w1(32'hbc6bbc40),
	.w2(32'hbbc5911c),
	.w3(32'hbc342e6f),
	.w4(32'hb7ee1c94),
	.w5(32'h3b9988bd),
	.w6(32'h3c1b44c1),
	.w7(32'h3a977ada),
	.w8(32'hbac3a3e2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd34ba7c),
	.w1(32'hbc69dcaf),
	.w2(32'hbc567c11),
	.w3(32'hbcbc5c4c),
	.w4(32'hbce39aec),
	.w5(32'hbd079fb9),
	.w6(32'hbce9627c),
	.w7(32'hbb4e1f34),
	.w8(32'hbc6f211a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb4517f),
	.w1(32'hbbbe1602),
	.w2(32'hbc62d2c0),
	.w3(32'hbcc23254),
	.w4(32'h3b94628d),
	.w5(32'hbbaed469),
	.w6(32'hbcdbdc6c),
	.w7(32'hbca0a9d9),
	.w8(32'hbcd086b8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b5275),
	.w1(32'h3c339fc6),
	.w2(32'hbc01a267),
	.w3(32'h3c2dc320),
	.w4(32'hbd3dbf3d),
	.w5(32'h3b43df68),
	.w6(32'h3bfa609a),
	.w7(32'h3acd7c49),
	.w8(32'h3b0bfb17),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c3aa7),
	.w1(32'h38056218),
	.w2(32'hbc8726d5),
	.w3(32'hb9dce14a),
	.w4(32'h3b6aaa96),
	.w5(32'h3b8d9852),
	.w6(32'hba366fdc),
	.w7(32'h3b6b63ee),
	.w8(32'h3b82aac3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91f8a3),
	.w1(32'h3c5f093d),
	.w2(32'hbaba07ee),
	.w3(32'h3bd8bf2c),
	.w4(32'h3c228a41),
	.w5(32'h3b2d8f3e),
	.w6(32'hbd33b194),
	.w7(32'h3c0f09d8),
	.w8(32'hbb92751a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda2ce0e),
	.w1(32'hbc810b46),
	.w2(32'hbdc3408a),
	.w3(32'hbd3343da),
	.w4(32'h3cacb71e),
	.w5(32'hbcda15cf),
	.w6(32'hbdb19c50),
	.w7(32'hbca5104c),
	.w8(32'hbda15c03),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd94ad5d),
	.w1(32'h3a041172),
	.w2(32'hbcd476a8),
	.w3(32'hbc1d1dde),
	.w4(32'h3cee081c),
	.w5(32'hbc60b686),
	.w6(32'hbccbf980),
	.w7(32'h3c4b5aa5),
	.w8(32'hbcc4bf9b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd35be4b),
	.w1(32'h3cb43966),
	.w2(32'hbcabc8c7),
	.w3(32'hbcd3d5c9),
	.w4(32'h3d01c693),
	.w5(32'h3ab2f3b9),
	.w6(32'hbd813a00),
	.w7(32'hbb92edff),
	.w8(32'hbdf29ee8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baeec57),
	.w1(32'hbc1d946c),
	.w2(32'h3893bb71),
	.w3(32'h3a8187cf),
	.w4(32'h3c00c21d),
	.w5(32'hbba88725),
	.w6(32'h3b237cf4),
	.w7(32'hba87890d),
	.w8(32'hbb78c6d7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012adc),
	.w1(32'h3b6a8e4e),
	.w2(32'h3c2bae63),
	.w3(32'h3adba453),
	.w4(32'hba9bd6a2),
	.w5(32'h3b8f8957),
	.w6(32'h3bcdf697),
	.w7(32'h3b2d5d9c),
	.w8(32'h3b1753ad),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf45cb2),
	.w1(32'h3bcd74a3),
	.w2(32'hbd20faeb),
	.w3(32'hbc1a136f),
	.w4(32'h3c428447),
	.w5(32'hbdcc7b8e),
	.w6(32'h3bbf6c82),
	.w7(32'hbaaf9001),
	.w8(32'hbbe6069e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f1074),
	.w1(32'h3a8769ae),
	.w2(32'hbbd22821),
	.w3(32'hbac5c23e),
	.w4(32'h3c4b233a),
	.w5(32'hbc0eb178),
	.w6(32'hba2a4c9e),
	.w7(32'h3c0a58fc),
	.w8(32'hbbbf600e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d72dc),
	.w1(32'h3d0f3c5b),
	.w2(32'hbbd1be29),
	.w3(32'hba3e05bc),
	.w4(32'h3cbbcbbd),
	.w5(32'hbc2e5b71),
	.w6(32'hbc8d61f9),
	.w7(32'hb8c2ea6f),
	.w8(32'hbcc2a1dc),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35a77a),
	.w1(32'hbb421656),
	.w2(32'hbc8b9eec),
	.w3(32'hbbc865b7),
	.w4(32'hbb566f1d),
	.w5(32'h3c01b2fc),
	.w6(32'hbb8c5a2f),
	.w7(32'h3b4539df),
	.w8(32'h3b38de80),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7dd3b),
	.w1(32'h3b628b54),
	.w2(32'hbc400df6),
	.w3(32'hbb643485),
	.w4(32'hbc2aa9c7),
	.w5(32'hbd1f6084),
	.w6(32'h39851cf9),
	.w7(32'h3c5b585e),
	.w8(32'hbbfa7a70),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2865f4),
	.w1(32'hbbbd70c0),
	.w2(32'hbbfe55ad),
	.w3(32'h3b74add6),
	.w4(32'h3bbb4546),
	.w5(32'hbb6294fc),
	.w6(32'hbb073114),
	.w7(32'hbafd476d),
	.w8(32'hbca4f789),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc229270),
	.w1(32'hbd3f407e),
	.w2(32'hbc02cf80),
	.w3(32'hbb0eac66),
	.w4(32'hba528595),
	.w5(32'hbd1a7b98),
	.w6(32'hbc5d4482),
	.w7(32'hbadcfb0b),
	.w8(32'hbbe94230),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01be4f),
	.w1(32'hbb814782),
	.w2(32'h3befcc67),
	.w3(32'hbb670217),
	.w4(32'hbc10e4c2),
	.w5(32'hbc661ed3),
	.w6(32'h3b91dfed),
	.w7(32'hbc8fb891),
	.w8(32'hbd00b431),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f2eff),
	.w1(32'hbcad940f),
	.w2(32'hbb77c81b),
	.w3(32'hbb780608),
	.w4(32'hbbb7d82b),
	.w5(32'h3b6c54f1),
	.w6(32'h3a407e93),
	.w7(32'hbbfc223f),
	.w8(32'hbca1a29f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4f65fe),
	.w1(32'hb9bcc549),
	.w2(32'hbd05f7b9),
	.w3(32'h3aa43af1),
	.w4(32'hbda06c04),
	.w5(32'h3cab0e95),
	.w6(32'hbb724d7c),
	.w7(32'h3d29e3e2),
	.w8(32'hbc3b1d30),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0df247),
	.w1(32'h3cf6295d),
	.w2(32'hbdc67fc9),
	.w3(32'hbd1a4730),
	.w4(32'h3d5b23f3),
	.w5(32'hbc187f9f),
	.w6(32'hbd3c5c9c),
	.w7(32'h3d01492d),
	.w8(32'hbd3be866),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83aa17),
	.w1(32'h3d249e36),
	.w2(32'hbd534a8d),
	.w3(32'hbc3a54b1),
	.w4(32'h3d24acfd),
	.w5(32'hbd0fb716),
	.w6(32'hbcf09165),
	.w7(32'h3c6ee7b3),
	.w8(32'hbd34d905),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e4e57),
	.w1(32'h3b909480),
	.w2(32'hbadd57e8),
	.w3(32'hba0d8902),
	.w4(32'h3cc8fac4),
	.w5(32'h3ad0bf7b),
	.w6(32'hb98bb095),
	.w7(32'h3bdba938),
	.w8(32'h3c288708),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6643eb),
	.w1(32'hbc30b64e),
	.w2(32'h3bb8fe56),
	.w3(32'hbbec05d0),
	.w4(32'hbb862b7d),
	.w5(32'h3bb7c89a),
	.w6(32'h3addc352),
	.w7(32'h3b8f593e),
	.w8(32'h3ae1996f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47b7c5),
	.w1(32'h3c9ffd86),
	.w2(32'hbb913f0f),
	.w3(32'hbb5dea49),
	.w4(32'h3c7f7285),
	.w5(32'hbc063f6b),
	.w6(32'hbb9f2ca2),
	.w7(32'h3c292778),
	.w8(32'h3c1033a0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03561a),
	.w1(32'h3bdfba6b),
	.w2(32'hba046c35),
	.w3(32'hbc45f0b1),
	.w4(32'h3ca5f603),
	.w5(32'hbba3fb5a),
	.w6(32'hbcc46e03),
	.w7(32'h3c6882e7),
	.w8(32'hbc9f00e4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd03e966),
	.w1(32'hbb511eb4),
	.w2(32'hbd125483),
	.w3(32'hbd165223),
	.w4(32'h3b88c4e6),
	.w5(32'hbc98348d),
	.w6(32'hbd22be12),
	.w7(32'hbc8d864f),
	.w8(32'hbd1aff7e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce0070),
	.w1(32'h3d2b1b09),
	.w2(32'hbca73e02),
	.w3(32'h3b97011d),
	.w4(32'h3d2b4160),
	.w5(32'hbc54b90c),
	.w6(32'hbc916f31),
	.w7(32'hbaa1b800),
	.w8(32'hbcd88ed4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0dc60e),
	.w1(32'h3b5e68db),
	.w2(32'hbcbc166b),
	.w3(32'hbc7f364b),
	.w4(32'h3d0ccd8a),
	.w5(32'hbdb5570b),
	.w6(32'hbce8fe06),
	.w7(32'h3bc1168a),
	.w8(32'hbd8f195b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd30bf80),
	.w1(32'h3bfcd578),
	.w2(32'hbcc396fb),
	.w3(32'h3b6c0c64),
	.w4(32'h3caa548c),
	.w5(32'hbc9838d3),
	.w6(32'hbd064f38),
	.w7(32'hbbbc0dc2),
	.w8(32'hbc9e76d6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3bb1b3),
	.w1(32'hbd07562f),
	.w2(32'hbcde253a),
	.w3(32'hbd124203),
	.w4(32'hbd6fb037),
	.w5(32'hbcca22e0),
	.w6(32'hbcb28c5e),
	.w7(32'hbd13f7f2),
	.w8(32'hbd6ebadc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cbed6),
	.w1(32'hbc631353),
	.w2(32'hbb2681af),
	.w3(32'hbc2d1b14),
	.w4(32'h3b06d25e),
	.w5(32'hbbb0226f),
	.w6(32'hb9b70e28),
	.w7(32'hba3b4b9e),
	.w8(32'h3c4fc189),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb881896),
	.w1(32'hb9fd3bf7),
	.w2(32'hbd3dcb28),
	.w3(32'hbbefbc25),
	.w4(32'h3c148501),
	.w5(32'h3bfc89ca),
	.w6(32'h3c30c7b6),
	.w7(32'hbb5906c4),
	.w8(32'h3bd3e9cb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff02a2),
	.w1(32'h3b203ece),
	.w2(32'hb95a194f),
	.w3(32'h3ba5b3cf),
	.w4(32'hbad13ad2),
	.w5(32'h39575507),
	.w6(32'hb9e5a31b),
	.w7(32'hba8bed69),
	.w8(32'h3af2df13),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8017be),
	.w1(32'hbc8d1444),
	.w2(32'hbcbbd78a),
	.w3(32'h3cd5b8ce),
	.w4(32'hbc61b97e),
	.w5(32'hbc5d6d5b),
	.w6(32'hbc2f083d),
	.w7(32'h3c0e15f2),
	.w8(32'hbca6e806),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa39cec),
	.w1(32'h3c1cc19f),
	.w2(32'hbbef4bbf),
	.w3(32'h3b1f4a14),
	.w4(32'h3c183117),
	.w5(32'hbc18b2a2),
	.w6(32'hba88e7f1),
	.w7(32'hbbae0bb6),
	.w8(32'hbc6cf581),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0b5da7),
	.w1(32'hbdefd056),
	.w2(32'hbccd8251),
	.w3(32'hbc977876),
	.w4(32'hbc0c3bb4),
	.w5(32'hbd020394),
	.w6(32'hbca2e5af),
	.w7(32'hbc237be8),
	.w8(32'hbc37a28a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe910fc),
	.w1(32'h3b03f667),
	.w2(32'h3c318bcf),
	.w3(32'hbc32c665),
	.w4(32'hbbf3b2ec),
	.w5(32'hbc3feb00),
	.w6(32'hbc4b7034),
	.w7(32'h3b44b7b8),
	.w8(32'hbc37baed),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc587c),
	.w1(32'hbb7cf48c),
	.w2(32'h3b76a005),
	.w3(32'h3c1e42ef),
	.w4(32'h3c180a38),
	.w5(32'hbad7deec),
	.w6(32'h3b97dd71),
	.w7(32'h39444f3c),
	.w8(32'hbb46f2cf),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbc273),
	.w1(32'hbb82fe45),
	.w2(32'h3c8898de),
	.w3(32'hbb67f1d6),
	.w4(32'h3c1c5457),
	.w5(32'hbbd4cf50),
	.w6(32'hbbc86d48),
	.w7(32'h3bfb4ecc),
	.w8(32'h3ae9f020),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65ff7b),
	.w1(32'h3be636aa),
	.w2(32'h3c1e4a9e),
	.w3(32'hbb994397),
	.w4(32'h3c57a19d),
	.w5(32'hbb9d1c59),
	.w6(32'h3be5809c),
	.w7(32'h3c293302),
	.w8(32'hbb2d118f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4afd5),
	.w1(32'h3c224705),
	.w2(32'hbb8b6b78),
	.w3(32'h3c818cdc),
	.w4(32'hbb0eb967),
	.w5(32'hbaf91534),
	.w6(32'hbb5408cb),
	.w7(32'h3aebc32f),
	.w8(32'h39c936f3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b165b),
	.w1(32'h3ca7387e),
	.w2(32'h39c99c5a),
	.w3(32'hbab842ac),
	.w4(32'h3b63c7aa),
	.w5(32'h3b443263),
	.w6(32'hbab3d786),
	.w7(32'hbb835453),
	.w8(32'h3c11a844),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b644a),
	.w1(32'h3bce5a72),
	.w2(32'hbd27d05f),
	.w3(32'hbaee9247),
	.w4(32'h3bd06432),
	.w5(32'hbca250db),
	.w6(32'hbbcfa834),
	.w7(32'hbbf4665d),
	.w8(32'hbc36ff1c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2716d9),
	.w1(32'hbc0fec47),
	.w2(32'hbc253beb),
	.w3(32'hbca232cb),
	.w4(32'h3bc4d391),
	.w5(32'h3b29e30e),
	.w6(32'hbceb22d1),
	.w7(32'h3ca674e9),
	.w8(32'h3c67f08c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d9bbe),
	.w1(32'hbacdbfab),
	.w2(32'h3a15b750),
	.w3(32'hbb858de2),
	.w4(32'h3a6e358a),
	.w5(32'h37e88bc5),
	.w6(32'hbbcdaeba),
	.w7(32'h3b1bac8f),
	.w8(32'h3c05169b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9965a5e),
	.w1(32'hbbc87157),
	.w2(32'hbc30418a),
	.w3(32'h3c0c29c0),
	.w4(32'h3bf0c7a8),
	.w5(32'h3b6f915d),
	.w6(32'hbc46b2c0),
	.w7(32'hbc41daac),
	.w8(32'hbb9f3dd6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a6233),
	.w1(32'h3b9261fa),
	.w2(32'h3b1d6b6b),
	.w3(32'hbc95ba65),
	.w4(32'hbb9d3506),
	.w5(32'hbc35998c),
	.w6(32'h3c79ad96),
	.w7(32'hbbbb4972),
	.w8(32'hbbc057c5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c9103),
	.w1(32'h3cba522a),
	.w2(32'hbb3fe257),
	.w3(32'hbc12f46b),
	.w4(32'hba39b5eb),
	.w5(32'h3b3ddd29),
	.w6(32'h3c1c172e),
	.w7(32'h3c820f11),
	.w8(32'h3c0ab7ce),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4f1fc7),
	.w1(32'h3abb6c20),
	.w2(32'hbca9c2bf),
	.w3(32'hbcfad406),
	.w4(32'hbc9fbc86),
	.w5(32'hbcffc5d4),
	.w6(32'hbca4ef18),
	.w7(32'hba8ec032),
	.w8(32'h3b87425d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3d6c4a),
	.w1(32'hbc346242),
	.w2(32'hbd3dbaac),
	.w3(32'hbcb9e95d),
	.w4(32'h3c8ea2fe),
	.w5(32'hbcb192f3),
	.w6(32'hbd445db9),
	.w7(32'hbbf6a8e6),
	.w8(32'hbd238d70),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfbd24a),
	.w1(32'h3b934190),
	.w2(32'hbd269841),
	.w3(32'hbca3d392),
	.w4(32'h3c821123),
	.w5(32'hbca25939),
	.w6(32'hbd77c621),
	.w7(32'hbc843b27),
	.w8(32'hbd219218),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd32cabe),
	.w1(32'h3cfd8d5d),
	.w2(32'hbd445b5d),
	.w3(32'hbc5fb0c1),
	.w4(32'h3d818c67),
	.w5(32'hbb8539ea),
	.w6(32'hbd574a59),
	.w7(32'h3ca51571),
	.w8(32'hbd95ad5c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c788e73),
	.w1(32'hbc027c04),
	.w2(32'hbc8645e7),
	.w3(32'h3bb26873),
	.w4(32'h3ba45d42),
	.w5(32'h3b003754),
	.w6(32'hbbfddffc),
	.w7(32'hbaff94a5),
	.w8(32'hbc6cf47b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b2735),
	.w1(32'hbbeab629),
	.w2(32'hbb42efcc),
	.w3(32'hbb73c324),
	.w4(32'h3b84d455),
	.w5(32'h3ba48380),
	.w6(32'hbb4ce9ee),
	.w7(32'h3c014cee),
	.w8(32'hbae7367a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5edb59),
	.w1(32'hba14a9f7),
	.w2(32'h3b9210f4),
	.w3(32'hbb39129c),
	.w4(32'hba963ae9),
	.w5(32'hbc26eceb),
	.w6(32'h3b875910),
	.w7(32'h3b3ed5aa),
	.w8(32'h3c1cd8f0),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7367ab),
	.w1(32'h39395705),
	.w2(32'hbc02627a),
	.w3(32'hbb56178b),
	.w4(32'hbba30a6b),
	.w5(32'h3b98b35c),
	.w6(32'hbba7394b),
	.w7(32'h3b860a91),
	.w8(32'hbc2dfa68),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b752a47),
	.w1(32'h3be55016),
	.w2(32'h3b8d1fe3),
	.w3(32'h3d3b6f33),
	.w4(32'hbbf45142),
	.w5(32'h3a3cdacc),
	.w6(32'h3abf9e75),
	.w7(32'h3c0b1688),
	.w8(32'hbabe7f4c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca3dc1),
	.w1(32'hbc8c6fb6),
	.w2(32'h3beb901b),
	.w3(32'hbc2b2500),
	.w4(32'hbcef7557),
	.w5(32'hbc0d085b),
	.w6(32'hbbf91994),
	.w7(32'hbbaf559e),
	.w8(32'hbb264f7d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd392d29),
	.w1(32'hbd0494f7),
	.w2(32'hbccb2062),
	.w3(32'hbcd3f7f2),
	.w4(32'hbc76be9c),
	.w5(32'hbc948dc8),
	.w6(32'hbcd8e969),
	.w7(32'h3b2d941b),
	.w8(32'hbcd9a7ed),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd103306),
	.w1(32'hbb84c351),
	.w2(32'hbcf0e747),
	.w3(32'hbc85744b),
	.w4(32'h3c9dc53e),
	.w5(32'hbb93067b),
	.w6(32'hbce9e036),
	.w7(32'hbc927bbc),
	.w8(32'hbc8b9775),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0ec3d),
	.w1(32'hbb44c448),
	.w2(32'hbc93ff0c),
	.w3(32'hbbeb5e0a),
	.w4(32'h3bc0c327),
	.w5(32'hbc46972f),
	.w6(32'hbcc12e85),
	.w7(32'h3bc220eb),
	.w8(32'hbb9e5796),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac997b6),
	.w1(32'hbb7fcbc6),
	.w2(32'hbc60e967),
	.w3(32'hbb9e7a22),
	.w4(32'hbc3c66bb),
	.w5(32'hbb5d6adc),
	.w6(32'hbab8c146),
	.w7(32'hbb0e403b),
	.w8(32'hbc8c2691),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf51dc1),
	.w1(32'hbb111866),
	.w2(32'hbc564670),
	.w3(32'hbc31c1ea),
	.w4(32'h372fcd9e),
	.w5(32'hbae7f4ce),
	.w6(32'hbc8e8119),
	.w7(32'h3c8c04d9),
	.w8(32'hbc6af5af),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43ac70),
	.w1(32'h3a4f8953),
	.w2(32'hbc8b38a5),
	.w3(32'hbc9a2ce3),
	.w4(32'h3b886464),
	.w5(32'hbccc67f3),
	.w6(32'hbcecc99a),
	.w7(32'hbcb44660),
	.w8(32'hbcb4ed4b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57c9a3),
	.w1(32'h3c2313bb),
	.w2(32'h3a81de85),
	.w3(32'hb9f3fc36),
	.w4(32'h3c8d27c1),
	.w5(32'h3b2408a3),
	.w6(32'hbc1abeab),
	.w7(32'h3c28afae),
	.w8(32'hbc7e13f9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc61e3),
	.w1(32'hbb646da2),
	.w2(32'h3aa880c2),
	.w3(32'h3b61e902),
	.w4(32'hba11ea39),
	.w5(32'hbbdbdcdc),
	.w6(32'hbc143ab1),
	.w7(32'hbc013c69),
	.w8(32'hbbdde169),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c522a),
	.w1(32'hbc430e01),
	.w2(32'h3b6fb6b5),
	.w3(32'hbba45f64),
	.w4(32'hbc124a5c),
	.w5(32'h37ad4525),
	.w6(32'hbb20fb69),
	.w7(32'h3c83129b),
	.w8(32'h3a1ebe96),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b891646),
	.w1(32'hbbb2d466),
	.w2(32'hbb93d7de),
	.w3(32'hbb97ced2),
	.w4(32'h3b59130e),
	.w5(32'h3bd1ba35),
	.w6(32'hbb68bd74),
	.w7(32'h3a9a4557),
	.w8(32'hbb05e606),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5098e4),
	.w1(32'h3c62ce3a),
	.w2(32'hbc6baac4),
	.w3(32'hbcc04bbd),
	.w4(32'h3ce1b4a5),
	.w5(32'hbcdf9417),
	.w6(32'hbcd4519b),
	.w7(32'h3b4394d1),
	.w8(32'hbcb0fd60),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ac138),
	.w1(32'hb9ab91f7),
	.w2(32'h3a3ae3e2),
	.w3(32'h3b46cf9f),
	.w4(32'h3c85b9ed),
	.w5(32'h3c411502),
	.w6(32'h3c91c9f3),
	.w7(32'h3c516bbf),
	.w8(32'hbc2e798e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1b198f),
	.w1(32'hbc289bf2),
	.w2(32'h3c8d00eb),
	.w3(32'hbc204f29),
	.w4(32'h3c63c49b),
	.w5(32'h3bb84eca),
	.w6(32'hbad9d7e1),
	.w7(32'h3d21d4d7),
	.w8(32'hbc3c32b2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4b1f50),
	.w1(32'hbc32a32e),
	.w2(32'hbcf3c21d),
	.w3(32'hbd009da7),
	.w4(32'hbc719906),
	.w5(32'hbd151095),
	.w6(32'hbd7e9fd5),
	.w7(32'hbcb0760b),
	.w8(32'hbd02006c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba098577),
	.w1(32'h3c902155),
	.w2(32'hbb8db3fe),
	.w3(32'hbb29c39f),
	.w4(32'h3c6bf5e3),
	.w5(32'hbc1e1178),
	.w6(32'h3c82f242),
	.w7(32'h3b4d5efa),
	.w8(32'hbc7df754),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd26372b),
	.w1(32'hbcac7410),
	.w2(32'hbd01dd45),
	.w3(32'hbcc84d22),
	.w4(32'hbca83989),
	.w5(32'hbbb7a970),
	.w6(32'hbc663898),
	.w7(32'h3b476205),
	.w8(32'hbd1edc3b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade62fd),
	.w1(32'h3b60241f),
	.w2(32'hbc21e3fa),
	.w3(32'h3c073e54),
	.w4(32'h3cd02ef4),
	.w5(32'h3b8814c9),
	.w6(32'hbca5a8e5),
	.w7(32'hbc31f864),
	.w8(32'hbc70f766),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88d733),
	.w1(32'hbb70c21b),
	.w2(32'hbd540b1e),
	.w3(32'hbcaa0c82),
	.w4(32'h3bd39c10),
	.w5(32'hbc5be1c5),
	.w6(32'hbd0dba15),
	.w7(32'h3c460bfa),
	.w8(32'hbcc2ea33),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca19f6),
	.w1(32'h3b96e31e),
	.w2(32'hbbeb8e50),
	.w3(32'hbbb3bc04),
	.w4(32'h3ccfc503),
	.w5(32'hbb0f0c5a),
	.w6(32'hbc231e81),
	.w7(32'h3cc9ae82),
	.w8(32'hba19dbfd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc6449c),
	.w1(32'h3cb69a7b),
	.w2(32'hbc176dfc),
	.w3(32'hbc75fa90),
	.w4(32'h3c850142),
	.w5(32'hbbd5ef55),
	.w6(32'hbcae38e7),
	.w7(32'h3cce8010),
	.w8(32'hbc8b0311),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8da81d),
	.w1(32'h3b2d986d),
	.w2(32'h3ab75b43),
	.w3(32'hbb9a3085),
	.w4(32'hbc1eb374),
	.w5(32'hbbb26265),
	.w6(32'hbc90e96c),
	.w7(32'h3a2cc8d0),
	.w8(32'h3aad7de1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd213f),
	.w1(32'hbc3e6b2a),
	.w2(32'hbd15d864),
	.w3(32'hbc8d6884),
	.w4(32'hbb6e5b0c),
	.w5(32'hbc97adc8),
	.w6(32'hbd2d7bf9),
	.w7(32'hbbf78298),
	.w8(32'hbd24cc55),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc495bef),
	.w1(32'h3c0dcf83),
	.w2(32'hbca06e4c),
	.w3(32'h3bc61c2a),
	.w4(32'h3b3b9e8a),
	.w5(32'hbce91be8),
	.w6(32'hbc803ceb),
	.w7(32'h3c1784eb),
	.w8(32'hbcd8157e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9882a6),
	.w1(32'hbc86902d),
	.w2(32'hbcbc68dd),
	.w3(32'hbc24eb0d),
	.w4(32'h3c08cd24),
	.w5(32'hbbe0c870),
	.w6(32'hbd5f2e4d),
	.w7(32'hbbb37287),
	.w8(32'hbd1f29ab),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4bc72),
	.w1(32'h3cf56597),
	.w2(32'hbc5eac65),
	.w3(32'h3b66fba4),
	.w4(32'h3d7e5d23),
	.w5(32'h3c354c6b),
	.w6(32'hbc79f87b),
	.w7(32'h3ce93321),
	.w8(32'hbcf81b2f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a7891),
	.w1(32'h3c569072),
	.w2(32'hbc8a60ce),
	.w3(32'hbc075cac),
	.w4(32'h3cb30c85),
	.w5(32'h3addae70),
	.w6(32'hbd1ad76b),
	.w7(32'h3b05276f),
	.w8(32'hbd03c973),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd402b78),
	.w1(32'hbcb090fd),
	.w2(32'hbceb5762),
	.w3(32'hbc84fee2),
	.w4(32'h3aeea814),
	.w5(32'hbcab4d02),
	.w6(32'hbcb0bff0),
	.w7(32'h3ad94237),
	.w8(32'hbcb88cbe),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a609433),
	.w1(32'hba5f0735),
	.w2(32'h3becf8ad),
	.w3(32'h3959b3e8),
	.w4(32'h3ce42146),
	.w5(32'hbac4aeb3),
	.w6(32'h3baaf253),
	.w7(32'hbc2d71ce),
	.w8(32'h3d0374d4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6aecea),
	.w1(32'hbc9d226c),
	.w2(32'hbd128fe7),
	.w3(32'hbd11fe3a),
	.w4(32'h3c9ce3e9),
	.w5(32'hbcef189d),
	.w6(32'hbb612d10),
	.w7(32'h3d02d3a1),
	.w8(32'hbb81e49b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecf6d5),
	.w1(32'hbc075813),
	.w2(32'hbc74635b),
	.w3(32'hbc821ce3),
	.w4(32'h3981672a),
	.w5(32'hbc44f76d),
	.w6(32'hbc75a0b2),
	.w7(32'h3b946db7),
	.w8(32'hbcb4307e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a4291),
	.w1(32'h3ac85f9b),
	.w2(32'h3b91c8fc),
	.w3(32'h3bdaaff3),
	.w4(32'hba4baf00),
	.w5(32'h39dfa34d),
	.w6(32'h3c2f4eeb),
	.w7(32'hbb9ec0fd),
	.w8(32'h3aa40af8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90e385),
	.w1(32'hbc1bc38c),
	.w2(32'hbb933ec6),
	.w3(32'hbcbf8c8d),
	.w4(32'h3ba5613a),
	.w5(32'hbc14376f),
	.w6(32'hbc4642c1),
	.w7(32'h38ebf708),
	.w8(32'h3b53901e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9b847),
	.w1(32'h3b0cee2e),
	.w2(32'hbd05b184),
	.w3(32'hbc0f647e),
	.w4(32'h3a1de98a),
	.w5(32'hbcb99c89),
	.w6(32'hbce1bb46),
	.w7(32'hbc6696f4),
	.w8(32'hbc2b9d40),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14073f),
	.w1(32'h3c8b2951),
	.w2(32'hbaed863b),
	.w3(32'hbc0e86fd),
	.w4(32'h3cfcd48c),
	.w5(32'h3c0fb16f),
	.w6(32'hbc5a6bff),
	.w7(32'hba291081),
	.w8(32'hbcdc06d4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a2fbd),
	.w1(32'h3cb1876a),
	.w2(32'hbcc8e064),
	.w3(32'hbca602bf),
	.w4(32'h3cbc30f3),
	.w5(32'h3b2c3eaf),
	.w6(32'h3ba001e4),
	.w7(32'hbadc3a33),
	.w8(32'hbbc80714),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb35a21),
	.w1(32'hbc67ac8f),
	.w2(32'hbc999d22),
	.w3(32'hbc701409),
	.w4(32'h3c6e1546),
	.w5(32'hba8d9961),
	.w6(32'hbbb3875f),
	.w7(32'h3b865123),
	.w8(32'hbc9df678),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d7152),
	.w1(32'hbb1574a9),
	.w2(32'hbced8188),
	.w3(32'hbc14c60c),
	.w4(32'h3c0baeb2),
	.w5(32'h3bd5c447),
	.w6(32'hbc5704b4),
	.w7(32'hbb89ddc7),
	.w8(32'hbd038674),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc8bc4),
	.w1(32'hbc789f99),
	.w2(32'hbc9a91ac),
	.w3(32'hbc2e36fd),
	.w4(32'hbb143514),
	.w5(32'hbb8b672a),
	.w6(32'hbbe63370),
	.w7(32'h3bf520b9),
	.w8(32'hbc21e888),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87cbba),
	.w1(32'hbae6ed88),
	.w2(32'hbbe5c435),
	.w3(32'hbc2e4767),
	.w4(32'h3c6e5b07),
	.w5(32'hbcae060c),
	.w6(32'hbbef23bc),
	.w7(32'h3bf46a0b),
	.w8(32'hbc8f1937),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0aa9e),
	.w1(32'hbb5a609a),
	.w2(32'hbb34cbbf),
	.w3(32'h3ba12cb9),
	.w4(32'hbc89b35b),
	.w5(32'hb633a049),
	.w6(32'h3c3134e3),
	.w7(32'hbb920b61),
	.w8(32'hbbf693fb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2e3fa7),
	.w1(32'h3c2bf534),
	.w2(32'hbac644f0),
	.w3(32'h3b919af5),
	.w4(32'hbb1efc4e),
	.w5(32'hba265e7e),
	.w6(32'h3caa448b),
	.w7(32'h3c0fd640),
	.w8(32'hbc85c1b3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9c2af),
	.w1(32'hbb446778),
	.w2(32'h3c3ee82d),
	.w3(32'hbb3b9ebe),
	.w4(32'h3abed34c),
	.w5(32'hba4d097c),
	.w6(32'hb9fd99da),
	.w7(32'h3ac4fa1a),
	.w8(32'hba8276f9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58d199),
	.w1(32'h3abfcd0b),
	.w2(32'h3bb987d6),
	.w3(32'h3b8d5ed6),
	.w4(32'hbaaa71d2),
	.w5(32'h3be5ecf7),
	.w6(32'h38d686d0),
	.w7(32'h3a9189da),
	.w8(32'h3ba3f423),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc046b36),
	.w1(32'h3c120e14),
	.w2(32'hbc809665),
	.w3(32'hbd1414cb),
	.w4(32'h3c9754c4),
	.w5(32'hbc8f4679),
	.w6(32'hbc7433a8),
	.w7(32'h3bdf3529),
	.w8(32'hbc369ae3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21ca38),
	.w1(32'hbbc577c0),
	.w2(32'h3b1043ae),
	.w3(32'hba8b15cf),
	.w4(32'hbbc137f9),
	.w5(32'h3b8ddeff),
	.w6(32'hbc128faa),
	.w7(32'hbc1eaf3f),
	.w8(32'h3c491476),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb981230),
	.w1(32'hbba2ef0f),
	.w2(32'h3a075c73),
	.w3(32'hbc7ab01c),
	.w4(32'hbc4829b0),
	.w5(32'hbc5270af),
	.w6(32'hbc3af3e4),
	.w7(32'hbbca4ea6),
	.w8(32'hbb3c0467),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccff07f),
	.w1(32'hb96c1871),
	.w2(32'hbcb4bc12),
	.w3(32'hbb8406ad),
	.w4(32'h3c9277fd),
	.w5(32'h3c0b079b),
	.w6(32'hbcf4873a),
	.w7(32'h3bd80cd7),
	.w8(32'hbca61922),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30ad1e),
	.w1(32'hbc516f38),
	.w2(32'hbb25d259),
	.w3(32'hbaeea5c5),
	.w4(32'hbc187a8a),
	.w5(32'h3bee3426),
	.w6(32'h3aa5d047),
	.w7(32'hbbf7e943),
	.w8(32'h3a1c71ae),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99332a4),
	.w1(32'h3b5e6ba3),
	.w2(32'hbba91c1f),
	.w3(32'hbc5c3a95),
	.w4(32'h3c0a22aa),
	.w5(32'hb9b5e993),
	.w6(32'hbc4e4f5f),
	.w7(32'h3ccccc82),
	.w8(32'h3bf83d0f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cea31),
	.w1(32'hb8d3c748),
	.w2(32'hba8600e9),
	.w3(32'h3c2ca62f),
	.w4(32'h3cf30fff),
	.w5(32'h3840933a),
	.w6(32'h3c7583c1),
	.w7(32'hb9900e2d),
	.w8(32'h399147cf),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39799ed5),
	.w1(32'h3a23ae84),
	.w2(32'hbc7a003b),
	.w3(32'hbb2802eb),
	.w4(32'hbb8b958f),
	.w5(32'hbca96734),
	.w6(32'hbbb8b9d8),
	.w7(32'h395596b7),
	.w8(32'hbc8ea6b5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8f8aa),
	.w1(32'hbc365b60),
	.w2(32'hbcbdbe04),
	.w3(32'h392ee5b9),
	.w4(32'hbb8da397),
	.w5(32'hbd283ec0),
	.w6(32'hbd515f0e),
	.w7(32'hbd04866d),
	.w8(32'hbc392f4a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35a09e),
	.w1(32'hbbe83366),
	.w2(32'hbc8f2f5f),
	.w3(32'hbbc9006c),
	.w4(32'hbbd6fbcd),
	.w5(32'hbcc65094),
	.w6(32'hbc944d55),
	.w7(32'h3b192a3a),
	.w8(32'h3bba435e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2eff6d),
	.w1(32'hb937ff14),
	.w2(32'h39458779),
	.w3(32'hbbb9d718),
	.w4(32'h3acbc543),
	.w5(32'h3b2a446e),
	.w6(32'h3ae2eea1),
	.w7(32'h3bfa6f92),
	.w8(32'h3bfd78cf),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d59ee),
	.w1(32'hbb5e7c35),
	.w2(32'hbc020f48),
	.w3(32'h3bc0996e),
	.w4(32'hbb7909c6),
	.w5(32'h3b9f5978),
	.w6(32'hbc73845a),
	.w7(32'hbc5cb06a),
	.w8(32'hbc6355c8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d5ffa),
	.w1(32'h3bd125d1),
	.w2(32'hbbf974a3),
	.w3(32'hbc9f59a8),
	.w4(32'hbcf343f0),
	.w5(32'hbaa823ee),
	.w6(32'hbcd43cf3),
	.w7(32'hbbffd8fa),
	.w8(32'hbbd8b8e8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42db57),
	.w1(32'h3afbbd5b),
	.w2(32'hbbcac447),
	.w3(32'hbb8a0f57),
	.w4(32'h3bc8aaac),
	.w5(32'hbc528279),
	.w6(32'hbc482873),
	.w7(32'hbce414cf),
	.w8(32'hbb9a5226),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccd8934),
	.w1(32'h3a28a904),
	.w2(32'hbc851ef3),
	.w3(32'hbceeffca),
	.w4(32'h394a017d),
	.w5(32'h3c0f7b60),
	.w6(32'hbc9c4467),
	.w7(32'h3c75c79d),
	.w8(32'h396a9316),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bc872),
	.w1(32'hbcb6069d),
	.w2(32'hbd2247d9),
	.w3(32'hbcbdd6b1),
	.w4(32'hbd0eabc9),
	.w5(32'hbd190c7d),
	.w6(32'hbca75b12),
	.w7(32'h3b228d21),
	.w8(32'hbcdcdb73),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3d55e6),
	.w1(32'h3c321ab9),
	.w2(32'hbaf7c0c8),
	.w3(32'h3c985669),
	.w4(32'h3c8241e8),
	.w5(32'hbc023252),
	.w6(32'hbc14318a),
	.w7(32'h3c1f0a64),
	.w8(32'hbcaea5dc),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc522668),
	.w1(32'h3b512e5a),
	.w2(32'hbd1cddb7),
	.w3(32'hbc077072),
	.w4(32'hbc38d4ba),
	.w5(32'h3bde8c7c),
	.w6(32'hbbff3f36),
	.w7(32'h3bc7fa43),
	.w8(32'hbc865dd7),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce64245),
	.w1(32'hbd21bd63),
	.w2(32'hbc3682e8),
	.w3(32'hbbcdfe1b),
	.w4(32'hbbcc1bb0),
	.w5(32'hbc03bb02),
	.w6(32'hbc4952e7),
	.w7(32'h3b7204bf),
	.w8(32'hbc38caca),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdca4d8),
	.w1(32'h3b71867a),
	.w2(32'hbd36d007),
	.w3(32'hbbdf98e4),
	.w4(32'h3c7e0a05),
	.w5(32'hbaa342e9),
	.w6(32'hbd4b50c9),
	.w7(32'hb953279d),
	.w8(32'hbcd3c1c5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e089f),
	.w1(32'hbc672e31),
	.w2(32'hbca4a73a),
	.w3(32'hbc2a0c12),
	.w4(32'h3b2ce31d),
	.w5(32'hba4cf8f8),
	.w6(32'hbbf765a3),
	.w7(32'hba11a9c8),
	.w8(32'hbb85b2c1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ac2dc),
	.w1(32'h3aff6c4e),
	.w2(32'hbb9e8345),
	.w3(32'hbd132ee2),
	.w4(32'hbc82a7a0),
	.w5(32'h3c05ceb4),
	.w6(32'hbac7f775),
	.w7(32'hbb91b931),
	.w8(32'hbc3bb6d7),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc411eaf),
	.w1(32'h3c84df3c),
	.w2(32'hbbf036a4),
	.w3(32'hbbb21273),
	.w4(32'h3ca4b3c3),
	.w5(32'hbb9e9a85),
	.w6(32'hbcd24b2e),
	.w7(32'h3cfe4474),
	.w8(32'hbd0d4a67),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc455169),
	.w1(32'h3ba0638e),
	.w2(32'h3ae4cfc7),
	.w3(32'h3bc0bd20),
	.w4(32'h3cd5fefe),
	.w5(32'hbc039359),
	.w6(32'hbc821364),
	.w7(32'h3c36d611),
	.w8(32'hbc7b5d74),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8e5de),
	.w1(32'hba593c98),
	.w2(32'hbb01dcce),
	.w3(32'hbb5ccdb4),
	.w4(32'hbb204b3c),
	.w5(32'hbc25ddc9),
	.w6(32'hbc36cfec),
	.w7(32'hbcfb5f78),
	.w8(32'hbce9670a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58699e),
	.w1(32'h3b34fa51),
	.w2(32'h3b6500de),
	.w3(32'h3a12062d),
	.w4(32'hbcc3f63f),
	.w5(32'h3b2005f4),
	.w6(32'hba52d91b),
	.w7(32'hbb8950fd),
	.w8(32'hbc19990d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14b687),
	.w1(32'hbd18b2cf),
	.w2(32'hbd2b085c),
	.w3(32'hbc3e49a2),
	.w4(32'h3ba6bed1),
	.w5(32'h3a7c2a92),
	.w6(32'hbc241bb5),
	.w7(32'h3c4b9383),
	.w8(32'hbc0195c3),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc8e7c0),
	.w1(32'hbb37b8a1),
	.w2(32'hbcd28ef3),
	.w3(32'hbc2430e3),
	.w4(32'h3d12f0c4),
	.w5(32'hbbc568dd),
	.w6(32'hbcd2740c),
	.w7(32'h3afe36b2),
	.w8(32'hbcaead4b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3336a),
	.w1(32'h3c0098e9),
	.w2(32'hbc4e314d),
	.w3(32'hbd16e178),
	.w4(32'h3bb0ac83),
	.w5(32'hbb7a2bb4),
	.w6(32'hbcfe54a0),
	.w7(32'h3a9bd7d0),
	.w8(32'hbc9dcf30),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe44ec3),
	.w1(32'h3c86ea6e),
	.w2(32'h3cc832ec),
	.w3(32'h3bff0746),
	.w4(32'hbb2be882),
	.w5(32'h3c1db739),
	.w6(32'hbc4012df),
	.w7(32'hbbb943d3),
	.w8(32'hbb804b98),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd304c75),
	.w1(32'h3b38d718),
	.w2(32'hbc42574b),
	.w3(32'hbcb6885e),
	.w4(32'h3bda494c),
	.w5(32'hbc8efdfb),
	.w6(32'hbcc6f299),
	.w7(32'hbb096ec3),
	.w8(32'hbc684eea),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cced8),
	.w1(32'hbc67c551),
	.w2(32'hbc3d1cd6),
	.w3(32'hbc297fa1),
	.w4(32'h3c8ac2b6),
	.w5(32'hbbca425a),
	.w6(32'hbc3d44b8),
	.w7(32'hbc5401a6),
	.w8(32'hbc43953e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd045db8),
	.w1(32'hbcb0916f),
	.w2(32'hbcdc817a),
	.w3(32'hbcd1a1f5),
	.w4(32'hbca2ab1d),
	.w5(32'hbca2e0d8),
	.w6(32'h3c835edd),
	.w7(32'hbcabd826),
	.w8(32'hbc78273d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10655d),
	.w1(32'h3cee7672),
	.w2(32'hbc82b776),
	.w3(32'h3ab167a4),
	.w4(32'h3cd755e9),
	.w5(32'hbb64691e),
	.w6(32'hbc99c120),
	.w7(32'h3c2151ee),
	.w8(32'hbc815327),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdd96cd),
	.w1(32'hbb67ef07),
	.w2(32'h3c55fc60),
	.w3(32'hbc68e26c),
	.w4(32'h3bce442c),
	.w5(32'hbb10396e),
	.w6(32'hb69d93ae),
	.w7(32'h3bc74077),
	.w8(32'h3c8d27b6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba20c65),
	.w1(32'h3b2697a7),
	.w2(32'h3b93c558),
	.w3(32'h3b9baf7e),
	.w4(32'h3b9c020e),
	.w5(32'hbbe0127f),
	.w6(32'hbb5a9cdd),
	.w7(32'h3ba5bdd5),
	.w8(32'hb867ed53),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19152b),
	.w1(32'hb858ca9c),
	.w2(32'hbd715c0b),
	.w3(32'hbd6100cd),
	.w4(32'h3d0bd5be),
	.w5(32'h3c84d6bb),
	.w6(32'h3c814c6e),
	.w7(32'h3d1fe856),
	.w8(32'hbb88a541),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc408b23),
	.w1(32'h3caf85c7),
	.w2(32'hbc278345),
	.w3(32'hbc75cfe0),
	.w4(32'h3cead7d1),
	.w5(32'hbc74b058),
	.w6(32'hbd3fe056),
	.w7(32'h3cb782d8),
	.w8(32'hbc118ff7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h358189d2),
	.w1(32'h3cc335a8),
	.w2(32'hbbfa10e7),
	.w3(32'h3b5ec61f),
	.w4(32'h3c83d8c4),
	.w5(32'hbb76797c),
	.w6(32'hba878f8d),
	.w7(32'h3c6f4a85),
	.w8(32'hbc66c20a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc336205),
	.w1(32'hbba9cd4a),
	.w2(32'hbb82c9ab),
	.w3(32'hbc1e1479),
	.w4(32'hbbb354c6),
	.w5(32'hbb5cf880),
	.w6(32'hbc571995),
	.w7(32'hbc29ebfd),
	.w8(32'hbbc8acc4),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb641f75),
	.w1(32'h3b98722d),
	.w2(32'hbc5a5822),
	.w3(32'h3b63b2fa),
	.w4(32'hbb32c9c3),
	.w5(32'hbb8bdf9f),
	.w6(32'hbb4a5204),
	.w7(32'h387ef572),
	.w8(32'hbc1e0dd4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0f37e1),
	.w1(32'hbb8354dd),
	.w2(32'hbca2c189),
	.w3(32'hbc4f09a9),
	.w4(32'hba90435e),
	.w5(32'hbc8252a7),
	.w6(32'hbc8167ac),
	.w7(32'hba9b17bd),
	.w8(32'hbc8fabd3),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd27d5b0),
	.w1(32'h3b0f53f8),
	.w2(32'h3ca0ef40),
	.w3(32'hbbd5c70c),
	.w4(32'hbb9be96a),
	.w5(32'hbb5b8d0b),
	.w6(32'hbb2fdc4e),
	.w7(32'hbbc8a529),
	.w8(32'hbcfed2ce),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11cee7),
	.w1(32'h3c3b6564),
	.w2(32'hbbed0ab4),
	.w3(32'h3be9d6a8),
	.w4(32'h3cadb59b),
	.w5(32'hbc850489),
	.w6(32'hbbcdec24),
	.w7(32'h3c02e7d7),
	.w8(32'hbc4b0e5d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d7bdb),
	.w1(32'hbbbb31fd),
	.w2(32'h3a620234),
	.w3(32'h3b7b33b2),
	.w4(32'hbca8924c),
	.w5(32'h3b08b21c),
	.w6(32'hbcd7a694),
	.w7(32'hbc271d45),
	.w8(32'h3afddb73),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc071376),
	.w1(32'hbae9db4f),
	.w2(32'hbcda3be1),
	.w3(32'hbb44fae4),
	.w4(32'hbb9cc6c5),
	.w5(32'hbcd2aa67),
	.w6(32'hbc93eb7f),
	.w7(32'hbaaafcd5),
	.w8(32'hbdde963f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfced05),
	.w1(32'h3bbc3196),
	.w2(32'h3b510ae8),
	.w3(32'h3b35a89a),
	.w4(32'h3ba73083),
	.w5(32'hbd6e607d),
	.w6(32'hbd50b67a),
	.w7(32'hbb333b95),
	.w8(32'hbb99f7b9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f598e),
	.w1(32'h379d89df),
	.w2(32'h3cd056e9),
	.w3(32'hbb517c7b),
	.w4(32'hbbb052d8),
	.w5(32'hbaf6e805),
	.w6(32'hbb5e9db5),
	.w7(32'h3c263193),
	.w8(32'hbc198c22),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fbfd0),
	.w1(32'hbb2cfd24),
	.w2(32'h3b85f948),
	.w3(32'hbb149f2a),
	.w4(32'h3bb57376),
	.w5(32'hbc77d6e2),
	.w6(32'h3bd76cfa),
	.w7(32'h3becc137),
	.w8(32'hb9d97aa2),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf65c98),
	.w1(32'h3b6fdec9),
	.w2(32'hbce8a02d),
	.w3(32'hbcc00b52),
	.w4(32'h3baf1e7c),
	.w5(32'hbcd1f6be),
	.w6(32'hbd22e538),
	.w7(32'hbd7e1bb3),
	.w8(32'hbd156bbd),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98082c),
	.w1(32'hbb2684ee),
	.w2(32'hbc3e074a),
	.w3(32'hbb705bfb),
	.w4(32'h3bc00ef3),
	.w5(32'hbcd1affd),
	.w6(32'hbba90243),
	.w7(32'h3c81036a),
	.w8(32'hbcd0e310),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bc04a),
	.w1(32'h3b7f3139),
	.w2(32'hbb51b7b3),
	.w3(32'hbc0dcc02),
	.w4(32'h3c4e5f54),
	.w5(32'hbbeae85a),
	.w6(32'hbc7b75ca),
	.w7(32'hbbae856d),
	.w8(32'hbc6a0cda),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b0477),
	.w1(32'h3b456cdd),
	.w2(32'h3b48b79b),
	.w3(32'hbc20c3b7),
	.w4(32'hba5e3cab),
	.w5(32'hbc34136c),
	.w6(32'hbbda3d56),
	.w7(32'hb99c0890),
	.w8(32'hbba227df),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd03b970),
	.w1(32'h3c2137a0),
	.w2(32'hbd04ea33),
	.w3(32'hbc8b2471),
	.w4(32'h3cd829ae),
	.w5(32'hbc9bb606),
	.w6(32'hbd418cb4),
	.w7(32'hbc265c69),
	.w8(32'hbd453b1e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9381f),
	.w1(32'h3c1648f9),
	.w2(32'h3ca24fc3),
	.w3(32'hbc6691dd),
	.w4(32'h3b84cefd),
	.w5(32'hbc7f6426),
	.w6(32'hbca4991e),
	.w7(32'hbb75e05c),
	.w8(32'hbd4c78aa),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ae3a7),
	.w1(32'hbbbffc08),
	.w2(32'hbc7cff0b),
	.w3(32'hbce10d33),
	.w4(32'hb94b5e2b),
	.w5(32'hbc557228),
	.w6(32'hbd17f5be),
	.w7(32'hbc429c39),
	.w8(32'hbce4afae),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b970817),
	.w1(32'hbac92731),
	.w2(32'hbaf5cef0),
	.w3(32'h3c0eb5e2),
	.w4(32'h3a1c86d6),
	.w5(32'h3adf7eed),
	.w6(32'h3ba38216),
	.w7(32'hbd32632d),
	.w8(32'hbc0f7e17),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca45bb7),
	.w1(32'hbb68a756),
	.w2(32'hbb2a03b3),
	.w3(32'h3a7cfc3a),
	.w4(32'h3b186186),
	.w5(32'hbae0b529),
	.w6(32'h3a665671),
	.w7(32'hbc087540),
	.w8(32'hbb690b0f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c019125),
	.w1(32'h3bebe4b7),
	.w2(32'h3c228efa),
	.w3(32'h3c7cd2c5),
	.w4(32'h3b41715a),
	.w5(32'h3a842a09),
	.w6(32'h3b7dcaf1),
	.w7(32'h3c046826),
	.w8(32'h3b8ec66f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd91a42),
	.w1(32'hba1b9e1c),
	.w2(32'hbc026b8e),
	.w3(32'hbbfd5c6e),
	.w4(32'h3b09abcb),
	.w5(32'h3a99a680),
	.w6(32'hbc6e2301),
	.w7(32'h3a6fe5d7),
	.w8(32'hbc4e7ed1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ee69c),
	.w1(32'hbae46599),
	.w2(32'h3cb455f5),
	.w3(32'h3a770fab),
	.w4(32'h3b8a463a),
	.w5(32'hbba45b78),
	.w6(32'hbc08d5f4),
	.w7(32'hb94a0e25),
	.w8(32'hbb85cc6a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94d1ea),
	.w1(32'hbd1b9a9b),
	.w2(32'hbc8c750b),
	.w3(32'hbc905de0),
	.w4(32'h3b1de378),
	.w5(32'hbb9b34ca),
	.w6(32'hbcf04656),
	.w7(32'hbb998636),
	.w8(32'hbbc31b3f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9cdcf),
	.w1(32'h3c130196),
	.w2(32'h3bce5e2d),
	.w3(32'h3b76541f),
	.w4(32'hbaab7ad2),
	.w5(32'h3b4cde51),
	.w6(32'h3bc52660),
	.w7(32'h3d06a173),
	.w8(32'h3b06b474),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79fda6),
	.w1(32'h3c17060d),
	.w2(32'h3c19e4a2),
	.w3(32'h3c4e94f3),
	.w4(32'hbb1c3040),
	.w5(32'hbb795177),
	.w6(32'h3a605cad),
	.w7(32'hbcb61461),
	.w8(32'h3b249f91),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f2d5f),
	.w1(32'h3ad72f24),
	.w2(32'hbbf91fff),
	.w3(32'hbb88a4ca),
	.w4(32'hbcc48654),
	.w5(32'hbb074c03),
	.w6(32'hbb60cf14),
	.w7(32'h3a9ccd85),
	.w8(32'hbb4b02c8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc002bee),
	.w1(32'h3b952d6a),
	.w2(32'hbce2edcb),
	.w3(32'hbc8b2460),
	.w4(32'hba28ccc7),
	.w5(32'hbc4a2cd4),
	.w6(32'hbc840989),
	.w7(32'hbc3eb798),
	.w8(32'hbc93c4c4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92cf6b),
	.w1(32'h362de860),
	.w2(32'hbc868d1d),
	.w3(32'hbcc4555f),
	.w4(32'hbabffcb2),
	.w5(32'h3be7fae1),
	.w6(32'hbb71c6af),
	.w7(32'h3c447b9a),
	.w8(32'h3a400441),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa20e88),
	.w1(32'hbc00ce3a),
	.w2(32'h3b874efb),
	.w3(32'hbbc411e6),
	.w4(32'h3b1094a9),
	.w5(32'hbb496640),
	.w6(32'hbc270871),
	.w7(32'h3bedb44d),
	.w8(32'hbb78c376),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce6157d),
	.w1(32'h3b521ef9),
	.w2(32'hbcf5898c),
	.w3(32'hbc051526),
	.w4(32'h3bc8e8cd),
	.w5(32'hbce46511),
	.w6(32'hbc0a5058),
	.w7(32'h3c4f627a),
	.w8(32'hbd0b31b8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84e13e),
	.w1(32'h3c0a753a),
	.w2(32'hbcd5d586),
	.w3(32'h3c6caccf),
	.w4(32'h3d1732f4),
	.w5(32'hbc9f78d7),
	.w6(32'hbd36f411),
	.w7(32'h3cdb6fe4),
	.w8(32'hbcbb7a2a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8533bd),
	.w1(32'hbbdeaf9e),
	.w2(32'hbc6b7ce9),
	.w3(32'hbb15daf2),
	.w4(32'hbc0a9204),
	.w5(32'hbc75617f),
	.w6(32'h3b97abb7),
	.w7(32'hbbd4b9e9),
	.w8(32'hbaf75e7c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf1b65),
	.w1(32'hbbf3b033),
	.w2(32'h3bff5a85),
	.w3(32'h3d3ebcc2),
	.w4(32'h3b1747e9),
	.w5(32'hbbc04ce9),
	.w6(32'h3be453cd),
	.w7(32'h3bb62965),
	.w8(32'h3c077f2c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd01e08),
	.w1(32'h3d1a4c14),
	.w2(32'hbc855243),
	.w3(32'h3b278268),
	.w4(32'h3abc610e),
	.w5(32'h3ba0c8b4),
	.w6(32'hbb5f5418),
	.w7(32'h3bac9c9d),
	.w8(32'hbbd57d64),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47f551),
	.w1(32'h3b112abd),
	.w2(32'h3b279fab),
	.w3(32'hbc20659c),
	.w4(32'hbc18178e),
	.w5(32'hbbb0349e),
	.w6(32'h3ad07469),
	.w7(32'h3b661e71),
	.w8(32'hbb07226e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e742c),
	.w1(32'hbcdb85d8),
	.w2(32'hbbdd03f4),
	.w3(32'h3b7dedbf),
	.w4(32'hbbe10560),
	.w5(32'hbc55a95d),
	.w6(32'hbac15738),
	.w7(32'h3bcf5614),
	.w8(32'hba6d8571),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3efea),
	.w1(32'hbc1c83fc),
	.w2(32'hbba390ec),
	.w3(32'hbc07865e),
	.w4(32'h3c339dc8),
	.w5(32'h390906dd),
	.w6(32'hbca53e08),
	.w7(32'hbbd316b6),
	.w8(32'hbcb2c4c9),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbb00f1),
	.w1(32'h3a8acf95),
	.w2(32'hbd1bebbb),
	.w3(32'hbbfa27c5),
	.w4(32'h3c8569ff),
	.w5(32'hbc2ed094),
	.w6(32'hbc875432),
	.w7(32'hbc4cfa16),
	.w8(32'hbcae6143),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0fc20),
	.w1(32'h3cf50d72),
	.w2(32'hbc6a2f01),
	.w3(32'hba3fb85e),
	.w4(32'h3c214b86),
	.w5(32'hbbba6b31),
	.w6(32'h39fb1678),
	.w7(32'hbc589cfd),
	.w8(32'hbbf7c397),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbacd3f),
	.w1(32'hbca38f3e),
	.w2(32'hbd02b535),
	.w3(32'hbc9f759e),
	.w4(32'h3ba4b65c),
	.w5(32'hbc88a82f),
	.w6(32'hbcbfc08e),
	.w7(32'hbc83f90a),
	.w8(32'hbd0eca6c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4da2c8),
	.w1(32'hbcba624b),
	.w2(32'hbbb9b6ee),
	.w3(32'hbc946abe),
	.w4(32'h3ca7a0d3),
	.w5(32'h3c87de3c),
	.w6(32'h3b9755b0),
	.w7(32'hbc388a81),
	.w8(32'hbc901d43),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79fc7d),
	.w1(32'hbceed1f6),
	.w2(32'h3bc1a592),
	.w3(32'h3b39c825),
	.w4(32'hbb2e4441),
	.w5(32'h39011e22),
	.w6(32'h39b4a532),
	.w7(32'h3aa30e24),
	.w8(32'h3c67a89c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f0ee7),
	.w1(32'h3bccb5a0),
	.w2(32'hbbddfea3),
	.w3(32'hbcc6c796),
	.w4(32'hbcdd7f34),
	.w5(32'h3b633111),
	.w6(32'hbb9cc838),
	.w7(32'h3b11dee7),
	.w8(32'h3c382d20),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8db240),
	.w1(32'hbc18ca4e),
	.w2(32'hba1ab954),
	.w3(32'hb9f603fe),
	.w4(32'hbb01ee58),
	.w5(32'hbc18f200),
	.w6(32'h3b39bd2c),
	.w7(32'h3b939999),
	.w8(32'hbb4da8b3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9965cb),
	.w1(32'h3b1f07dd),
	.w2(32'hbcd02b38),
	.w3(32'hbcfc373b),
	.w4(32'hbbeed2ba),
	.w5(32'hbca1139d),
	.w6(32'hbc9c11d4),
	.w7(32'hbd05e481),
	.w8(32'hbc5d5eea),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfaa2a0),
	.w1(32'h3c984fe1),
	.w2(32'hbcb9c2f1),
	.w3(32'hbc9aced2),
	.w4(32'h3c888311),
	.w5(32'hbadb4d2b),
	.w6(32'hbdc2582f),
	.w7(32'h3cc0bd42),
	.w8(32'hbca26191),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3b8e70),
	.w1(32'h3ae48293),
	.w2(32'hbc95430f),
	.w3(32'hbc0434e0),
	.w4(32'h3c2637f5),
	.w5(32'hbc063ce9),
	.w6(32'hbc782922),
	.w7(32'hba857064),
	.w8(32'hbc5dbe6a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5fe101),
	.w1(32'hbb7a490b),
	.w2(32'hbc0c24ca),
	.w3(32'h3c4a8ed3),
	.w4(32'h3c552e9c),
	.w5(32'hbbcd5409),
	.w6(32'hba3dc945),
	.w7(32'h3d19ffe1),
	.w8(32'hbc90ff75),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd535fc2),
	.w1(32'hbbf15718),
	.w2(32'hbcfea11d),
	.w3(32'hbc4c58ac),
	.w4(32'h3cd2f80a),
	.w5(32'hbb08cf86),
	.w6(32'hbbdd968c),
	.w7(32'h3c3c94ea),
	.w8(32'hbce13c44),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a5419),
	.w1(32'hbb851c21),
	.w2(32'hbc406f28),
	.w3(32'h3ce726cc),
	.w4(32'hbc840132),
	.w5(32'hbc5355e6),
	.w6(32'hbc645c52),
	.w7(32'hbc587843),
	.w8(32'hbbd01a02),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd161d47),
	.w1(32'hbc073ee3),
	.w2(32'hbc5de07c),
	.w3(32'hbccf7943),
	.w4(32'h3953e2eb),
	.w5(32'hbacaff12),
	.w6(32'hbd178226),
	.w7(32'hbad686af),
	.w8(32'hbcc245e9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacb7a8),
	.w1(32'h37651efd),
	.w2(32'hbb056186),
	.w3(32'hbc2aaa31),
	.w4(32'hbbe08c13),
	.w5(32'hbb5e59a2),
	.w6(32'h3c0e21a9),
	.w7(32'hbc923ccf),
	.w8(32'h3c893dcd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba715c5),
	.w1(32'h3b2a7a5a),
	.w2(32'hbad17539),
	.w3(32'h3b5be494),
	.w4(32'h3adeba49),
	.w5(32'h3c87a65b),
	.w6(32'h3b7dbaf0),
	.w7(32'h3d127154),
	.w8(32'h3bf2e97d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce038cc),
	.w1(32'h3c43ad79),
	.w2(32'hbd0e42b5),
	.w3(32'hbca3e957),
	.w4(32'h3cfb4f8f),
	.w5(32'hbcbc87f3),
	.w6(32'hbd07fd41),
	.w7(32'hbc1a0a48),
	.w8(32'hbd2887cc),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1b26fc),
	.w1(32'h3c1cb3b3),
	.w2(32'hbd4b7c75),
	.w3(32'hbc3cadc5),
	.w4(32'h3ce49674),
	.w5(32'hbcae0937),
	.w6(32'hbcf4ecd6),
	.w7(32'hbcafdd94),
	.w8(32'hbd27dc35),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc6550),
	.w1(32'hbcaffae7),
	.w2(32'hbcbb7c8e),
	.w3(32'h3b4dddf0),
	.w4(32'h3ca385b2),
	.w5(32'hbaf9249d),
	.w6(32'hbcc1063a),
	.w7(32'h3c8514b7),
	.w8(32'hbcdbb572),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd43ec7),
	.w1(32'hbc85748d),
	.w2(32'hbc8003fa),
	.w3(32'hbc9b61a9),
	.w4(32'hbc9b229e),
	.w5(32'hbc789cc8),
	.w6(32'h3c57dc96),
	.w7(32'h39058a3c),
	.w8(32'h3b42f2cd),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda00020),
	.w1(32'hba7f513a),
	.w2(32'h3b6578a7),
	.w3(32'h3bcc6583),
	.w4(32'hbc319258),
	.w5(32'hbb67fc6f),
	.w6(32'hb8b4fc6b),
	.w7(32'h398f53e8),
	.w8(32'hbc67ecb6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb141ee0),
	.w1(32'hbc1e98ab),
	.w2(32'hbd317038),
	.w3(32'h3b565d81),
	.w4(32'hbae7666f),
	.w5(32'hbaaa57c6),
	.w6(32'hbb802121),
	.w7(32'hbafa4ff3),
	.w8(32'hbbb38aa0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c42f2),
	.w1(32'hbcd4ae2f),
	.w2(32'hbcf200b9),
	.w3(32'h3c06978c),
	.w4(32'hbbf963ca),
	.w5(32'hbcf04dcd),
	.w6(32'hbca6359b),
	.w7(32'h3a8a62cf),
	.w8(32'hbcbc4d17),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf98fca),
	.w1(32'hbc079605),
	.w2(32'hbcc80658),
	.w3(32'hbc37db3b),
	.w4(32'hbbb769c8),
	.w5(32'hbcfdbd92),
	.w6(32'hbcdbfdb1),
	.w7(32'h3d6c58d2),
	.w8(32'hbcb1e2ce),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0da969),
	.w1(32'hbceb8f82),
	.w2(32'hbcbfd13d),
	.w3(32'hbce698ec),
	.w4(32'hbc8abde6),
	.w5(32'hbb20d214),
	.w6(32'hbd158e92),
	.w7(32'hbc30d53d),
	.w8(32'hbc53984e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d62b9),
	.w1(32'h3c7a2ff5),
	.w2(32'hbb08df34),
	.w3(32'hbccc52d3),
	.w4(32'h3cedc588),
	.w5(32'hbbd498b1),
	.w6(32'hbcc568a5),
	.w7(32'h3c0752df),
	.w8(32'hbc0a11b9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a7df2),
	.w1(32'h3b9e6871),
	.w2(32'hbcdf756d),
	.w3(32'hbbe9bcb8),
	.w4(32'h3cd7218e),
	.w5(32'hbdf118d3),
	.w6(32'hbc8930ae),
	.w7(32'h3c754813),
	.w8(32'hbca35c0a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa0483),
	.w1(32'h3b8b3045),
	.w2(32'hb8903687),
	.w3(32'hbcdec6d9),
	.w4(32'hbbbc34b4),
	.w5(32'hbc72d9bc),
	.w6(32'hbbcefbec),
	.w7(32'hbc51a779),
	.w8(32'hbb3dd362),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af74c5c),
	.w1(32'hbb67d59c),
	.w2(32'h3c288154),
	.w3(32'hba843721),
	.w4(32'h3b12a88b),
	.w5(32'h3bb5fef1),
	.w6(32'hbbcb45ac),
	.w7(32'h3ca59d05),
	.w8(32'hbb0a836b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05ff6a),
	.w1(32'hbc49c870),
	.w2(32'h3a9771a2),
	.w3(32'h3b59588e),
	.w4(32'hbc08823b),
	.w5(32'h3b8eacf1),
	.w6(32'hbc0b31e0),
	.w7(32'hbc6c4117),
	.w8(32'h3b2b4853),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1521f0),
	.w1(32'hbbfb31fb),
	.w2(32'h3b149f7b),
	.w3(32'hbbdb8cbc),
	.w4(32'hbcb80037),
	.w5(32'hbbb7dd40),
	.w6(32'h3c02137c),
	.w7(32'h3bb737b4),
	.w8(32'hbb598eb5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8d5e5),
	.w1(32'hbc0fb78a),
	.w2(32'hb9a92427),
	.w3(32'hbbbbb0ee),
	.w4(32'h3ba7b854),
	.w5(32'h3ca1c3df),
	.w6(32'hbc118526),
	.w7(32'hbb75ab28),
	.w8(32'h3c1b162b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcda7975),
	.w1(32'hbb8e1ebe),
	.w2(32'hbcac285e),
	.w3(32'hbc1ece32),
	.w4(32'h3ca443b8),
	.w5(32'hbbf78dc2),
	.w6(32'hbc0981e7),
	.w7(32'hbb7f5d8f),
	.w8(32'hbc478960),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae5db2),
	.w1(32'h3cf92da4),
	.w2(32'hbc0ac0a9),
	.w3(32'hbbc1676f),
	.w4(32'h3c160800),
	.w5(32'hbacd9b8c),
	.w6(32'hbc641fa6),
	.w7(32'hbb7ef71d),
	.w8(32'hbcfb81a6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a832f9a),
	.w1(32'h3b37ea2a),
	.w2(32'h3c67fa17),
	.w3(32'hbc2caff0),
	.w4(32'hbc49e167),
	.w5(32'hba93a9d7),
	.w6(32'h3c2ec46c),
	.w7(32'hbc110485),
	.w8(32'hbaa907ee),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1f77c7),
	.w1(32'hbcfe8cca),
	.w2(32'hbcf55ecc),
	.w3(32'hbd087238),
	.w4(32'hbc13c428),
	.w5(32'hbc9e514c),
	.w6(32'hbcf8bc52),
	.w7(32'hbc99bcd5),
	.w8(32'hbccb1f78),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb133a31),
	.w1(32'hbcc28782),
	.w2(32'hbc8dc383),
	.w3(32'h3a07bba6),
	.w4(32'hbb6e06a3),
	.w5(32'hbc73d39c),
	.w6(32'hbc605306),
	.w7(32'h3b823c12),
	.w8(32'hbcf5eda2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f7c6a),
	.w1(32'h3b4a66f4),
	.w2(32'hbb832b6c),
	.w3(32'hbb117860),
	.w4(32'h3b9b2224),
	.w5(32'hbc21ae1c),
	.w6(32'h3b1e405b),
	.w7(32'h3986b266),
	.w8(32'h3be17058),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc230931),
	.w1(32'hbc43d387),
	.w2(32'h3b870754),
	.w3(32'hbc41dea5),
	.w4(32'hbb949817),
	.w5(32'hbcb0ca4f),
	.w6(32'h3a8f6e07),
	.w7(32'hb9fb06c2),
	.w8(32'h3ba2f131),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71a7b3),
	.w1(32'h39dab7e0),
	.w2(32'hbbb3a19a),
	.w3(32'h3bfe2c4e),
	.w4(32'h3a001ddb),
	.w5(32'hbc6b3302),
	.w6(32'hbc2ec585),
	.w7(32'hbbb1c6ff),
	.w8(32'h3b918277),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ddbf),
	.w1(32'h3bdc14d4),
	.w2(32'h3c7a85e7),
	.w3(32'hbb72b58b),
	.w4(32'h3b1163b9),
	.w5(32'hbb334132),
	.w6(32'hbbb848f8),
	.w7(32'hbb77a823),
	.w8(32'h3bc83f0e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4639ce),
	.w1(32'hbc2dd5f1),
	.w2(32'hbbef1585),
	.w3(32'hbb1ce3c4),
	.w4(32'h3adad9d9),
	.w5(32'hbbb20a9b),
	.w6(32'h3c09502f),
	.w7(32'h3b9c5aa9),
	.w8(32'hbadacf22),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2707),
	.w1(32'h3b96770c),
	.w2(32'h3c91fa4d),
	.w3(32'hb9bec54c),
	.w4(32'hbc3dc4e7),
	.w5(32'hbbda208b),
	.w6(32'h3c2a69a8),
	.w7(32'hbc4e10a0),
	.w8(32'h3ba4387a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc091763),
	.w1(32'h3a2bdacb),
	.w2(32'h3bb3183d),
	.w3(32'hbc6ddd56),
	.w4(32'hbc1d23d3),
	.w5(32'h3af69e8c),
	.w6(32'hbbcb4df9),
	.w7(32'hba70af91),
	.w8(32'hbb8a3b9c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf1593),
	.w1(32'hbbdf1bd1),
	.w2(32'hbc2e197d),
	.w3(32'hbc8e9524),
	.w4(32'h3c1cd3e4),
	.w5(32'h3bce1db4),
	.w6(32'hbc41b6a0),
	.w7(32'hbc9c4fe5),
	.w8(32'hbcbc026f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25ef08),
	.w1(32'hbbcaa1cd),
	.w2(32'hbc4ce078),
	.w3(32'hbc774986),
	.w4(32'h3b866c25),
	.w5(32'hbbd8d2be),
	.w6(32'hbc928449),
	.w7(32'h3ab5ee70),
	.w8(32'hbc76f7fe),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd13e48),
	.w1(32'hbc350828),
	.w2(32'hbc801eab),
	.w3(32'hbcb92b97),
	.w4(32'hbc6e064e),
	.w5(32'hbd0cfe64),
	.w6(32'hbc6fc045),
	.w7(32'hb98a500e),
	.w8(32'hbb6d9920),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f61af),
	.w1(32'h3bb9cc98),
	.w2(32'hbb14618b),
	.w3(32'h3c0e89a4),
	.w4(32'h3b659660),
	.w5(32'hbcc31801),
	.w6(32'hb790b148),
	.w7(32'hbaad1ef6),
	.w8(32'hbb2045b8),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d09ec),
	.w1(32'hbbf433d8),
	.w2(32'hba831990),
	.w3(32'h3b953261),
	.w4(32'hbbb839f3),
	.w5(32'h3b0903a4),
	.w6(32'hb9bd8e09),
	.w7(32'hbbf153cf),
	.w8(32'h3ab6a064),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6317b8),
	.w1(32'h3b4c43ca),
	.w2(32'h3b9bedf6),
	.w3(32'h39611588),
	.w4(32'h3c0dedbb),
	.w5(32'h3c3fcb17),
	.w6(32'h3b06ff94),
	.w7(32'hbc02cba2),
	.w8(32'h3b79662f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36ae95),
	.w1(32'h3b5cd50f),
	.w2(32'h3b906b3b),
	.w3(32'hbaa4c774),
	.w4(32'hbbc3279c),
	.w5(32'h3c837a30),
	.w6(32'h3baf4833),
	.w7(32'hbb2a89df),
	.w8(32'h3c85f7a8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd132b3b),
	.w1(32'hbc941f13),
	.w2(32'hbca499fc),
	.w3(32'hbcbbe8d3),
	.w4(32'h3bffe372),
	.w5(32'hbc8e4db8),
	.w6(32'hbcf9bb4a),
	.w7(32'hb9e98b0b),
	.w8(32'hbc432184),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe214ed),
	.w1(32'hbbaab917),
	.w2(32'hbc475973),
	.w3(32'hbbc13c21),
	.w4(32'hb9914df1),
	.w5(32'hbb4d2867),
	.w6(32'h3ce30418),
	.w7(32'hb9aa63a8),
	.w8(32'h3ba1b12c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c236e93),
	.w1(32'hbabe98ae),
	.w2(32'hbb676626),
	.w3(32'h3b925373),
	.w4(32'h3c4fc256),
	.w5(32'hbc07fdfe),
	.w6(32'h3ca13029),
	.w7(32'h3c130b2e),
	.w8(32'hbbc5fc01),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de253e),
	.w1(32'h3b6ad7db),
	.w2(32'hbc0a7005),
	.w3(32'hbaa8c8d5),
	.w4(32'h3b614b52),
	.w5(32'h3a76e33c),
	.w6(32'hb991abd2),
	.w7(32'h3c2ade5d),
	.w8(32'hba85b490),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d1562),
	.w1(32'hbc494cf7),
	.w2(32'hbb904422),
	.w3(32'h3b3dfb34),
	.w4(32'hbb1016a7),
	.w5(32'h3ac68b4c),
	.w6(32'hbb6ff052),
	.w7(32'h3b0502a6),
	.w8(32'hbb55d5d1),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89f7b0),
	.w1(32'hbb6d0712),
	.w2(32'hbb9ce523),
	.w3(32'hbc032dee),
	.w4(32'hbbefc177),
	.w5(32'hbc2e6d02),
	.w6(32'hbc10b7da),
	.w7(32'hbc5557c6),
	.w8(32'hbc9745ae),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61f9ae),
	.w1(32'h3b1930d1),
	.w2(32'hbb44e419),
	.w3(32'h3c1c5e6a),
	.w4(32'h3c187e00),
	.w5(32'hbaa1068d),
	.w6(32'hbbe9c104),
	.w7(32'hbb0bfef3),
	.w8(32'hbb54d300),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd02a0b6),
	.w1(32'h3b65e531),
	.w2(32'hbd03d3dc),
	.w3(32'hbc9cb76f),
	.w4(32'h3c467a3e),
	.w5(32'h3b3e0220),
	.w6(32'hbc83c42b),
	.w7(32'hbb900898),
	.w8(32'h3b6541f6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83e597),
	.w1(32'h3a8544e6),
	.w2(32'h3cb18796),
	.w3(32'h3b15b3de),
	.w4(32'hbb2ca904),
	.w5(32'hbadfa522),
	.w6(32'h3b4653d9),
	.w7(32'hbbd2e3c7),
	.w8(32'hbb194738),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25c8d9),
	.w1(32'h3cc2edf4),
	.w2(32'h3a0417ec),
	.w3(32'hbc08be45),
	.w4(32'h3c83f509),
	.w5(32'hbbd6497a),
	.w6(32'hbc8d0a6f),
	.w7(32'hbb45559e),
	.w8(32'hbcec3462),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule