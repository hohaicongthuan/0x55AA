module layer_8_featuremap_88(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b226846),
	.w1(32'hbcb0593a),
	.w2(32'hbc97cbb4),
	.w3(32'hbb3fb808),
	.w4(32'h3c46ef2c),
	.w5(32'hbcdff54d),
	.w6(32'h3a87e8c0),
	.w7(32'hbb2bab96),
	.w8(32'hbb1627d9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf4a0e4),
	.w1(32'h3bb908c9),
	.w2(32'hb9e28327),
	.w3(32'h3c37b3c8),
	.w4(32'hbc2a8719),
	.w5(32'h3c1f41f5),
	.w6(32'hbbf888c4),
	.w7(32'h3be6d5e2),
	.w8(32'h39405f0b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80dc9a),
	.w1(32'hbb76a48d),
	.w2(32'hbd146754),
	.w3(32'h3c42f233),
	.w4(32'h3ac84b4c),
	.w5(32'hbc0e235d),
	.w6(32'hbb8ad7b9),
	.w7(32'hbc2d073e),
	.w8(32'h3c7f733d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37ce40),
	.w1(32'h391d9212),
	.w2(32'hbc13ba4e),
	.w3(32'h3b7d84a1),
	.w4(32'hbca259dd),
	.w5(32'hbbe3355e),
	.w6(32'hbcd243f4),
	.w7(32'hbc8627ff),
	.w8(32'hbcccfe4d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc82aea),
	.w1(32'hbc48df79),
	.w2(32'hbbc82603),
	.w3(32'hbbefba98),
	.w4(32'hbb84fe0f),
	.w5(32'h3b7e5ff5),
	.w6(32'hbb052a5c),
	.w7(32'hbcce81e2),
	.w8(32'h3c931998),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd455c9),
	.w1(32'h3be9eac5),
	.w2(32'hbc25be09),
	.w3(32'hbca00c88),
	.w4(32'hbbc688d1),
	.w5(32'hbbfb43b7),
	.w6(32'hbbbf2cd3),
	.w7(32'h3becac36),
	.w8(32'hbb888db2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc900870),
	.w1(32'hbb8ded24),
	.w2(32'h3b9e27c7),
	.w3(32'hba9c4c0a),
	.w4(32'h3c5ad2b3),
	.w5(32'h3b196956),
	.w6(32'hbccc7ba9),
	.w7(32'hbc45edcf),
	.w8(32'hbaaf9e7a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb7f1b),
	.w1(32'hbc1cff21),
	.w2(32'hbc02a90a),
	.w3(32'hbbbaae52),
	.w4(32'hbc7a27fe),
	.w5(32'hbbb0ced8),
	.w6(32'hbc8f596b),
	.w7(32'h3c0d425d),
	.w8(32'hbc266ac4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0921da),
	.w1(32'hbc13556c),
	.w2(32'hbb779fa8),
	.w3(32'h39b6a341),
	.w4(32'h3c06dcf6),
	.w5(32'hbbbb90be),
	.w6(32'h3c18f134),
	.w7(32'h3be6ccc1),
	.w8(32'hbcdbc8f7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f9a9d),
	.w1(32'hbd3d0ae2),
	.w2(32'h3d0310ad),
	.w3(32'hbc05db3c),
	.w4(32'h3c1080c8),
	.w5(32'h3c36f156),
	.w6(32'hbcf8f0b2),
	.w7(32'hbbd6bef2),
	.w8(32'h3b250c99),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80fd67),
	.w1(32'hbbf0878d),
	.w2(32'hbbb6c971),
	.w3(32'hbc955c22),
	.w4(32'h3c68759d),
	.w5(32'hbccb0740),
	.w6(32'h3b722516),
	.w7(32'h3b59cf16),
	.w8(32'h3da41ac8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badae33),
	.w1(32'h3b6d887d),
	.w2(32'h3bfa4da9),
	.w3(32'h3c4476ff),
	.w4(32'h3d300c98),
	.w5(32'hbca6118d),
	.w6(32'h3c822133),
	.w7(32'hbaf9227d),
	.w8(32'hbbd43aa6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64ce70),
	.w1(32'hbb3df142),
	.w2(32'hbcb21bb5),
	.w3(32'h3d88fbcf),
	.w4(32'hbbc7a22c),
	.w5(32'h3bb36c39),
	.w6(32'h3be136ff),
	.w7(32'h3d248b5e),
	.w8(32'h3c7a58b7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49db37),
	.w1(32'hbb1aa6ac),
	.w2(32'hbcacd280),
	.w3(32'h3bbe11f9),
	.w4(32'hbcbfb05d),
	.w5(32'h3cce66d1),
	.w6(32'hbc358222),
	.w7(32'h3b3d661c),
	.w8(32'hbbb4560e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d07c1a5),
	.w1(32'hbccb8283),
	.w2(32'hbda0a7f8),
	.w3(32'h3c5f1644),
	.w4(32'hbcc368a8),
	.w5(32'hbbf5db08),
	.w6(32'hbb621451),
	.w7(32'hbd0c1784),
	.w8(32'h3bfd2a8c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17856c),
	.w1(32'hbd38e146),
	.w2(32'h3bb083ef),
	.w3(32'hbd800b4a),
	.w4(32'hbcceb002),
	.w5(32'h3d3a1832),
	.w6(32'h3c70361c),
	.w7(32'hbbf50701),
	.w8(32'h3c802b17),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e90af),
	.w1(32'h3c8917ab),
	.w2(32'h3c10ac25),
	.w3(32'h3a01d9cc),
	.w4(32'hb93228ca),
	.w5(32'hbb45b512),
	.w6(32'hbc8967e1),
	.w7(32'h3c78897e),
	.w8(32'hbced1585),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c410e86),
	.w1(32'h3c46f5a7),
	.w2(32'h3c22a2a8),
	.w3(32'h3c1b6f88),
	.w4(32'hbd07035d),
	.w5(32'hbbb9bee2),
	.w6(32'hbdd010f9),
	.w7(32'h3d04774e),
	.w8(32'h39b68c6d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cd666),
	.w1(32'hbdb9107e),
	.w2(32'hbcd0d2c4),
	.w3(32'hba88f0fd),
	.w4(32'hbc045caa),
	.w5(32'hbc849044),
	.w6(32'h3c2549d7),
	.w7(32'hbcf70597),
	.w8(32'hbd00bdae),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb0c44),
	.w1(32'hbc51feeb),
	.w2(32'h39df9ce7),
	.w3(32'h3c5ed31e),
	.w4(32'hbca7729d),
	.w5(32'hbb59b79f),
	.w6(32'hbc2b5cd8),
	.w7(32'h3cd3d659),
	.w8(32'h3c0464a4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9f25b),
	.w1(32'hbc573ab7),
	.w2(32'h3c7c320b),
	.w3(32'hbcbd6aee),
	.w4(32'hbd841171),
	.w5(32'hbb73152e),
	.w6(32'h3c8546d8),
	.w7(32'h3c8cda4f),
	.w8(32'hbda7b075),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3675f2),
	.w1(32'hbd3339de),
	.w2(32'h3bd63155),
	.w3(32'h3c519aaa),
	.w4(32'hbb3f34af),
	.w5(32'hbd7b486d),
	.w6(32'h3c1e9b3b),
	.w7(32'hbc957170),
	.w8(32'hbc4ef78a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bc92a),
	.w1(32'hbc4b3ce9),
	.w2(32'h3c466222),
	.w3(32'hbc39bf2f),
	.w4(32'hbc0e1d7a),
	.w5(32'h3cb07c5a),
	.w6(32'hbbf653cb),
	.w7(32'h3c2391a5),
	.w8(32'h3c573929),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7db49),
	.w1(32'hbda1a2ac),
	.w2(32'hbc973761),
	.w3(32'hbd072cc6),
	.w4(32'hbda18652),
	.w5(32'hbb77ff47),
	.w6(32'h3b920db1),
	.w7(32'hbd2b25f0),
	.w8(32'h3cf693ab),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0feb8c),
	.w1(32'h3c50ef38),
	.w2(32'h3c31caa9),
	.w3(32'hbc8ed054),
	.w4(32'hbc8dd71f),
	.w5(32'h3c0f3163),
	.w6(32'hbc8682be),
	.w7(32'h3bd1ba50),
	.w8(32'h3c4139b4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbac955),
	.w1(32'hbd0086db),
	.w2(32'hbc8a5866),
	.w3(32'hbc6f997c),
	.w4(32'h3c20c57b),
	.w5(32'hbcaeb100),
	.w6(32'hbb5f813c),
	.w7(32'hbba6f26b),
	.w8(32'hbd6e5e00),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfe15f1),
	.w1(32'hbbc72d66),
	.w2(32'hba4a4103),
	.w3(32'hbd15613b),
	.w4(32'h3bae3931),
	.w5(32'hbcd6ad48),
	.w6(32'h3afb28cf),
	.w7(32'hbc16aa09),
	.w8(32'h3c23ef2a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec511d),
	.w1(32'hbd0056ed),
	.w2(32'hbd15cf79),
	.w3(32'h3d027aeb),
	.w4(32'hbd7ef549),
	.w5(32'hbc288301),
	.w6(32'h3c4e4f21),
	.w7(32'h3d38caaa),
	.w8(32'h3aaef688),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceb350e),
	.w1(32'h3ca1ae00),
	.w2(32'hbc36a91d),
	.w3(32'hb8b2dcd3),
	.w4(32'h3a95cf39),
	.w5(32'hbbd5d01c),
	.w6(32'h3d10d4a5),
	.w7(32'h3c06e746),
	.w8(32'h3d258acb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc751078),
	.w1(32'hbd379beb),
	.w2(32'h3ca41774),
	.w3(32'hbd367fc0),
	.w4(32'hbb33c296),
	.w5(32'h3b0b0a23),
	.w6(32'hbba9c2cf),
	.w7(32'hbc693717),
	.w8(32'hbad64bd8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec3435),
	.w1(32'h3cde3e93),
	.w2(32'hbb1243e9),
	.w3(32'h3c547f9d),
	.w4(32'hbd055549),
	.w5(32'h3b148a05),
	.w6(32'h3c90fe8b),
	.w7(32'hbc5cd9c8),
	.w8(32'hbbd275fc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33bbab),
	.w1(32'hba9e5a1c),
	.w2(32'hbc69f99c),
	.w3(32'hbc2da0aa),
	.w4(32'hbc18f1d0),
	.w5(32'h3aa2dd8d),
	.w6(32'hbb88a66e),
	.w7(32'h3b5c1252),
	.w8(32'hbbb1462c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9317ff),
	.w1(32'h3c6279ac),
	.w2(32'hbba24596),
	.w3(32'hbcc1e74a),
	.w4(32'h3c1bbe86),
	.w5(32'hbb5cb087),
	.w6(32'hbc519c46),
	.w7(32'hbc4890b4),
	.w8(32'hbcd7643c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4eeff4),
	.w1(32'hbb50978f),
	.w2(32'hbd3dc76e),
	.w3(32'hbc8d923a),
	.w4(32'hbc49527d),
	.w5(32'h3c08d8bc),
	.w6(32'hbc1b4a0a),
	.w7(32'hbd4f12b2),
	.w8(32'h3b2ed3b5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3c671),
	.w1(32'h3b859cce),
	.w2(32'h3c06b771),
	.w3(32'hbc67b43b),
	.w4(32'hbbb50a31),
	.w5(32'h3c8d929e),
	.w6(32'hbca0ad47),
	.w7(32'h3c653caf),
	.w8(32'hbb8c2ea3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c78c6),
	.w1(32'hbbe462c1),
	.w2(32'hbc8420d4),
	.w3(32'hbd0ab4c4),
	.w4(32'hbc64c402),
	.w5(32'hbce28d40),
	.w6(32'h3bf9531c),
	.w7(32'h3cad1676),
	.w8(32'h3c7ac3f6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d2c45),
	.w1(32'hbb45ed6e),
	.w2(32'hbb622a2c),
	.w3(32'hbbb8901f),
	.w4(32'hbc2343bb),
	.w5(32'h3cb3b61d),
	.w6(32'h3d24bbf9),
	.w7(32'hbca9c8af),
	.w8(32'h3c52ba45),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc242965),
	.w1(32'hbc9dd619),
	.w2(32'hbbaa5e3c),
	.w3(32'hbc8af8e8),
	.w4(32'hb8b85c11),
	.w5(32'hbbcd8d64),
	.w6(32'h3b2a8440),
	.w7(32'hbc402ce5),
	.w8(32'hbc63ac98),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb0acfa),
	.w1(32'hbcc3ff9a),
	.w2(32'h3cad6d3b),
	.w3(32'hbc8fc694),
	.w4(32'hbce14042),
	.w5(32'hbcaafcec),
	.w6(32'hbae248a2),
	.w7(32'h3ad95c5c),
	.w8(32'h3bf316ec),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c7e82),
	.w1(32'hba40cc84),
	.w2(32'hbbb43a70),
	.w3(32'h3d12369e),
	.w4(32'hbc7b579e),
	.w5(32'hbc9021b2),
	.w6(32'h3ace65c3),
	.w7(32'h3c82c28b),
	.w8(32'h3ae685f3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34ea74),
	.w1(32'hba1ef795),
	.w2(32'hbcb2894c),
	.w3(32'hbd186221),
	.w4(32'hb9e2aa29),
	.w5(32'hbcbd8b02),
	.w6(32'hbcb6d475),
	.w7(32'h3a83ed32),
	.w8(32'h3b3f816f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c894993),
	.w1(32'h3c432985),
	.w2(32'hbce085a6),
	.w3(32'hbc8c8417),
	.w4(32'hbcb1b26c),
	.w5(32'hbc28f45a),
	.w6(32'h3b25112b),
	.w7(32'hbc937b44),
	.w8(32'h3c49a390),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41898f),
	.w1(32'h3bbdbc98),
	.w2(32'hba5819f0),
	.w3(32'hbc19c93a),
	.w4(32'h3c650f1d),
	.w5(32'h3ca6f85b),
	.w6(32'hbc930f36),
	.w7(32'hb9a1877b),
	.w8(32'hbcd7235f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfec5d7),
	.w1(32'h3cd11e41),
	.w2(32'hbc6c03d4),
	.w3(32'hbd00375e),
	.w4(32'h3c1c8aee),
	.w5(32'h3ba9165f),
	.w6(32'hbb1199a8),
	.w7(32'h3a3ce3ef),
	.w8(32'h3d1f553a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7bdd4),
	.w1(32'hbc000c79),
	.w2(32'h3c85a0bc),
	.w3(32'hbbfd54e9),
	.w4(32'h3c81d011),
	.w5(32'hbc8782b6),
	.w6(32'h3ce3c8e7),
	.w7(32'h3c3cc7dc),
	.w8(32'h3c09f649),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a8d76),
	.w1(32'h3c1f7ca3),
	.w2(32'hbccbb0c8),
	.w3(32'h3bd655c1),
	.w4(32'hbcdb0931),
	.w5(32'h3d0f27b4),
	.w6(32'hbbdb993e),
	.w7(32'h3c16dd56),
	.w8(32'h3c08ae9a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd466390),
	.w1(32'hbcca1217),
	.w2(32'h3cf8aa26),
	.w3(32'hbcb522c3),
	.w4(32'hbc9eb2f6),
	.w5(32'h3c3212ce),
	.w6(32'h3aac056a),
	.w7(32'hbc4ad291),
	.w8(32'hbc01b963),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc11ef),
	.w1(32'hbc202fa5),
	.w2(32'hbb99b2c2),
	.w3(32'hbb7cdaa1),
	.w4(32'hbbf3d687),
	.w5(32'hba0c8ef3),
	.w6(32'h3cbe34e5),
	.w7(32'hbb9a8e75),
	.w8(32'hbca7ad85),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be99e88),
	.w1(32'hbd0a15c6),
	.w2(32'hbc88e83c),
	.w3(32'h3c8ec6c1),
	.w4(32'hba7518d7),
	.w5(32'hbab1ea92),
	.w6(32'h3c13eb63),
	.w7(32'h3b68339d),
	.w8(32'hbd183e54),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd1f9b6),
	.w1(32'h38e65186),
	.w2(32'h3d159016),
	.w3(32'hbc55f33d),
	.w4(32'hbbc3736b),
	.w5(32'h3991dd16),
	.w6(32'h3c2c5132),
	.w7(32'h3d0d20e7),
	.w8(32'h3b5ab497),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc197831),
	.w1(32'h3cd5832c),
	.w2(32'hbc2849cf),
	.w3(32'hbc24be95),
	.w4(32'hbbd8679a),
	.w5(32'h3cdd94f0),
	.w6(32'hbca8867c),
	.w7(32'h3c5fe1da),
	.w8(32'hbbb4b523),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c043f01),
	.w1(32'hbc906569),
	.w2(32'h3bb7dc9c),
	.w3(32'hbcf00bb6),
	.w4(32'hbc23f836),
	.w5(32'h3c44ba5e),
	.w6(32'hbc3ef5de),
	.w7(32'h3d29209f),
	.w8(32'h3d2cc04e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82b9d7),
	.w1(32'hbd00e312),
	.w2(32'hbd2987fc),
	.w3(32'h3c6baf92),
	.w4(32'hbcbe3d6e),
	.w5(32'hbc71998b),
	.w6(32'h3cb04804),
	.w7(32'hbcdd498b),
	.w8(32'h3c098474),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6bf4b),
	.w1(32'hbcc8899e),
	.w2(32'hbbd13236),
	.w3(32'h3b75639c),
	.w4(32'h3c061042),
	.w5(32'hbb54d3a8),
	.w6(32'hbc3ccd95),
	.w7(32'hbb18896d),
	.w8(32'h3bcfa4e4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1af544),
	.w1(32'hbbedcff2),
	.w2(32'hbc0af1dc),
	.w3(32'h3977180d),
	.w4(32'hbc75e884),
	.w5(32'hbba287fa),
	.w6(32'hbab07e1a),
	.w7(32'hbcb89b2a),
	.w8(32'h3bef2545),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfb9dbf),
	.w1(32'hb99a1d64),
	.w2(32'hbd0d3153),
	.w3(32'h3afef0e1),
	.w4(32'hbc1a9ebb),
	.w5(32'h3bfc7f32),
	.w6(32'h3b334752),
	.w7(32'h3af89f81),
	.w8(32'hbb4f81d1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a33f8),
	.w1(32'h3d427185),
	.w2(32'h3ccc7067),
	.w3(32'hbc66346f),
	.w4(32'hbd5b9157),
	.w5(32'h3c67ed99),
	.w6(32'hbccc0ac1),
	.w7(32'h3c74b3f5),
	.w8(32'h3bddfaeb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca86e51),
	.w1(32'h3d2d65a6),
	.w2(32'h3c19dd71),
	.w3(32'h3c2ed762),
	.w4(32'hbc692c2f),
	.w5(32'h3bf2acad),
	.w6(32'hbc0faf1a),
	.w7(32'hbbc152b0),
	.w8(32'h3c07fbd9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f9764),
	.w1(32'hbd2a2ea8),
	.w2(32'h3c7cb598),
	.w3(32'h3c23ca31),
	.w4(32'h3c2cce78),
	.w5(32'hbbfbfa41),
	.w6(32'hbb4ee6af),
	.w7(32'h3c0c1a97),
	.w8(32'hb97a6bad),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc60718),
	.w1(32'h3b4323bd),
	.w2(32'h3c96086e),
	.w3(32'h3ce8f8ae),
	.w4(32'h3b1e00e3),
	.w5(32'hbc7633f4),
	.w6(32'hba027a34),
	.w7(32'hbbc1bb64),
	.w8(32'hbb50e0c9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd634d),
	.w1(32'hbcacfcb6),
	.w2(32'h3b5cab43),
	.w3(32'h3d436a2d),
	.w4(32'h3d05b2dd),
	.w5(32'hbcbce863),
	.w6(32'hbc5b8f8c),
	.w7(32'hbb7b10e4),
	.w8(32'h3c2aac3e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d32f28b),
	.w1(32'hb953a398),
	.w2(32'h3c0dde16),
	.w3(32'hbc812b4a),
	.w4(32'h3ba75ac6),
	.w5(32'hba8ad2b5),
	.w6(32'hbc9e914d),
	.w7(32'hbbd783a1),
	.w8(32'hb98f6d38),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2faa2f),
	.w1(32'h3bca407c),
	.w2(32'hbc4c6f7c),
	.w3(32'h3c4ec67c),
	.w4(32'hbbd6b178),
	.w5(32'hbaa095c5),
	.w6(32'h3c5c268f),
	.w7(32'h3c802120),
	.w8(32'h3cf0cb03),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc752a2),
	.w1(32'hbb9b1266),
	.w2(32'hbbdea5f3),
	.w3(32'hbc0a64af),
	.w4(32'hbd4fe86f),
	.w5(32'hb91b1f23),
	.w6(32'h3be1f8e9),
	.w7(32'h3a8d3437),
	.w8(32'h3a682f30),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba1d79),
	.w1(32'h3b845dbc),
	.w2(32'h3d54a514),
	.w3(32'h3b26624e),
	.w4(32'h3c52f93d),
	.w5(32'hbb6d6743),
	.w6(32'hbad68eca),
	.w7(32'hbc1c573d),
	.w8(32'hbc30b59c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbcf4e),
	.w1(32'h3b8e8bf6),
	.w2(32'h3c248040),
	.w3(32'h3b53ef0f),
	.w4(32'h3ccea2af),
	.w5(32'hbce43254),
	.w6(32'h3c842595),
	.w7(32'hbc373b66),
	.w8(32'hbb5fd7fa),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b7232),
	.w1(32'hbdb8aaf3),
	.w2(32'h3a233e86),
	.w3(32'hbb05b6b4),
	.w4(32'hbbb76fb8),
	.w5(32'hbb81ec1d),
	.w6(32'h3b6bcd91),
	.w7(32'h3abe9771),
	.w8(32'hb968cc57),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb23b5a),
	.w1(32'h3d0a0f73),
	.w2(32'h3b4e2dba),
	.w3(32'h3c6fe53d),
	.w4(32'h3c439c65),
	.w5(32'h3cb6de93),
	.w6(32'h3c24417f),
	.w7(32'hbbd54277),
	.w8(32'hbb99ca28),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3f25d),
	.w1(32'h3c46404d),
	.w2(32'h3d0c3ee8),
	.w3(32'hba6f74af),
	.w4(32'hbc8184ef),
	.w5(32'h3c0966cc),
	.w6(32'h3a1db0ce),
	.w7(32'hbca6c93e),
	.w8(32'h38be6830),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce10b36),
	.w1(32'h3bcc9c9e),
	.w2(32'hbc531000),
	.w3(32'h3b660677),
	.w4(32'hbbda61bb),
	.w5(32'h3bf8bbc0),
	.w6(32'h3c39b8e8),
	.w7(32'h3ccc0dbb),
	.w8(32'hbcb84dcb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce3fe4),
	.w1(32'h3aba3378),
	.w2(32'hbc7c1ab1),
	.w3(32'hbb0e02e0),
	.w4(32'hbc321b42),
	.w5(32'hbc5cf765),
	.w6(32'hba92a20d),
	.w7(32'hbb99797b),
	.w8(32'h3c90d1d9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c090f59),
	.w1(32'hb9ae806b),
	.w2(32'hbb66f8b1),
	.w3(32'h3b8f8fe3),
	.w4(32'hba1091a6),
	.w5(32'hbbd35175),
	.w6(32'hbc095dc5),
	.w7(32'hbccb86b5),
	.w8(32'hbc9b0136),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0e800),
	.w1(32'h3cf85dcc),
	.w2(32'hb9fa75f6),
	.w3(32'hbbff8e9f),
	.w4(32'hbbb0d8cb),
	.w5(32'hbc5fcc2d),
	.w6(32'h3cf7f68d),
	.w7(32'hbbedfee5),
	.w8(32'h3be70d88),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc497d9c),
	.w1(32'h3d8c6737),
	.w2(32'hbb59e4a1),
	.w3(32'h3c814d02),
	.w4(32'h3ced53db),
	.w5(32'hbb8d40b7),
	.w6(32'h3bf9427b),
	.w7(32'h3c8c7962),
	.w8(32'h3ba385ea),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b386978),
	.w1(32'hbc841501),
	.w2(32'hbb2ac4c4),
	.w3(32'hbc302a85),
	.w4(32'h3c4ff947),
	.w5(32'h3a2ffd11),
	.w6(32'h3c856989),
	.w7(32'hbc86339c),
	.w8(32'h3c489626),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba72b0a),
	.w1(32'h3a6cbe80),
	.w2(32'hbc35b521),
	.w3(32'h3c28d4d2),
	.w4(32'hbb51ea2f),
	.w5(32'hbb990eb6),
	.w6(32'hbbca7ce6),
	.w7(32'h3ba1dd84),
	.w8(32'h3c57e90e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedffa4),
	.w1(32'h3d0cbe03),
	.w2(32'hbb4037b1),
	.w3(32'hb99b7a5f),
	.w4(32'hbbe10f3c),
	.w5(32'hbc0fdf1f),
	.w6(32'hbb0da983),
	.w7(32'h3c70f2de),
	.w8(32'hbbf0122e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cd46c),
	.w1(32'hbca6ba7b),
	.w2(32'hbc09010a),
	.w3(32'h3b30a85c),
	.w4(32'h3bd54d01),
	.w5(32'h3b10fdfe),
	.w6(32'h3b7e09e0),
	.w7(32'h3c7f6245),
	.w8(32'hbca5e655),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc34119),
	.w1(32'hbbda5b0c),
	.w2(32'hbc9e3fd5),
	.w3(32'h3bddd679),
	.w4(32'h3cc3eb41),
	.w5(32'hbb112521),
	.w6(32'h3bd91fbb),
	.w7(32'h3c5cb8db),
	.w8(32'h3b14bc99),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc447dd7),
	.w1(32'h3c2831a9),
	.w2(32'h3c105b29),
	.w3(32'h3c02e70c),
	.w4(32'hbc0cb77f),
	.w5(32'hbb7fbd56),
	.w6(32'h3d063f96),
	.w7(32'h3cdf84a1),
	.w8(32'hbb857830),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c722c1e),
	.w1(32'hbc378db9),
	.w2(32'hbb747470),
	.w3(32'h3b11a272),
	.w4(32'hbc789c1f),
	.w5(32'h3ae53503),
	.w6(32'hbaecd2c4),
	.w7(32'hbb813550),
	.w8(32'h3c9b3c49),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c371665),
	.w1(32'h3bdbbf99),
	.w2(32'hbbab28c6),
	.w3(32'hbc48e38e),
	.w4(32'h3d343fd5),
	.w5(32'h3b9eada8),
	.w6(32'hbc23775a),
	.w7(32'hbbcfa01d),
	.w8(32'hbc26f5fe),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa46474),
	.w1(32'hbb304012),
	.w2(32'hbc389f21),
	.w3(32'h3ca21ce9),
	.w4(32'hbba1c44a),
	.w5(32'h3a652b7a),
	.w6(32'h3c974155),
	.w7(32'hbb57c84f),
	.w8(32'h3c559327),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba76aee),
	.w1(32'h3b57f87a),
	.w2(32'h3c3f122f),
	.w3(32'hba1d6869),
	.w4(32'h3c1d7dc8),
	.w5(32'h3cc880bb),
	.w6(32'h3b3fcd6f),
	.w7(32'hbba069a8),
	.w8(32'hba3c3123),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60263b),
	.w1(32'h3c6751a7),
	.w2(32'hbbdecaaf),
	.w3(32'h3b0e42f0),
	.w4(32'h3bb921f5),
	.w5(32'h3c8d50f1),
	.w6(32'h3c315493),
	.w7(32'h3dacd52f),
	.w8(32'h3cefa540),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb9243a),
	.w1(32'h3bd222cc),
	.w2(32'hbcb1e154),
	.w3(32'hbbadbe2d),
	.w4(32'hbd15ab8f),
	.w5(32'hbce9dba5),
	.w6(32'h3b3457c2),
	.w7(32'hbc037dc7),
	.w8(32'hbc59e70a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3469f1),
	.w1(32'hba1e7541),
	.w2(32'hbc84c043),
	.w3(32'h3cc1aabf),
	.w4(32'h3b068432),
	.w5(32'hbd0e258b),
	.w6(32'hbc8425e8),
	.w7(32'h3bea6dcf),
	.w8(32'hbd22f829),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b57e9),
	.w1(32'hbc4d372e),
	.w2(32'hbcb572c3),
	.w3(32'hbc65770b),
	.w4(32'hbb9b7add),
	.w5(32'h3c07feb2),
	.w6(32'h3bf66ba1),
	.w7(32'hbb831b63),
	.w8(32'hbbd172f9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb710aa7),
	.w1(32'h3bdad2b6),
	.w2(32'hbcc68aa4),
	.w3(32'h3c93c35b),
	.w4(32'h3b7e4e06),
	.w5(32'hbab586fc),
	.w6(32'hbc290284),
	.w7(32'hbc5d1ba5),
	.w8(32'hbb979261),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baec6a0),
	.w1(32'h3c4ff563),
	.w2(32'h3ce3a1a1),
	.w3(32'h3cf1c2b1),
	.w4(32'hbc8eafce),
	.w5(32'hbc5eb9d1),
	.w6(32'hbcc1b5ef),
	.w7(32'hbbdb5e85),
	.w8(32'hbc6d65b2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1e5e12),
	.w1(32'h3cbd2080),
	.w2(32'hbc7a20ea),
	.w3(32'h398b46fd),
	.w4(32'hbd77438a),
	.w5(32'h3c0f91e5),
	.w6(32'h3b54d1d5),
	.w7(32'hbcefe1c2),
	.w8(32'h39e3505b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9bce2),
	.w1(32'h3c202b78),
	.w2(32'hbbc699bb),
	.w3(32'hbcff3ef7),
	.w4(32'hbc890a85),
	.w5(32'h3aac0c66),
	.w6(32'hbaa4a243),
	.w7(32'hbbcdef7f),
	.w8(32'h3d5dbe65),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2404c2),
	.w1(32'hbb3b518f),
	.w2(32'hbbc285a6),
	.w3(32'h3bcbdf48),
	.w4(32'hbbcbc14a),
	.w5(32'h3c0fde8d),
	.w6(32'hba477c17),
	.w7(32'hbac44891),
	.w8(32'hbbe1561a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d8968),
	.w1(32'h3b8fb132),
	.w2(32'h3c4d4c08),
	.w3(32'hbc6553b4),
	.w4(32'h3c55464a),
	.w5(32'hbc84d45c),
	.w6(32'hbc1c486f),
	.w7(32'hbc355151),
	.w8(32'hbc24ee93),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cad0c),
	.w1(32'hbc7734a3),
	.w2(32'h3cbd6e35),
	.w3(32'h3b316454),
	.w4(32'hbd48f12a),
	.w5(32'h3c52b6a1),
	.w6(32'hbbc074d8),
	.w7(32'h3b94ceab),
	.w8(32'hbcb5a6a8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd18d460),
	.w1(32'hbc6e3990),
	.w2(32'hbafcbce3),
	.w3(32'hbb000e94),
	.w4(32'hbbbd3f16),
	.w5(32'h3ca57ea8),
	.w6(32'h3da9bb33),
	.w7(32'h3cbb6b8c),
	.w8(32'hb8d4321a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a984bd9),
	.w1(32'hbaf2e4bf),
	.w2(32'hbb21b279),
	.w3(32'h3b77ac59),
	.w4(32'h3c4e6e8d),
	.w5(32'h3c1d0872),
	.w6(32'h3ca78818),
	.w7(32'h3b394d74),
	.w8(32'h3bddd6ae),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc62dd6),
	.w1(32'h3bda0826),
	.w2(32'h3cb41b9f),
	.w3(32'h3ac07aeb),
	.w4(32'h3c42049f),
	.w5(32'h39d0c734),
	.w6(32'hbb6cc2b1),
	.w7(32'hbbd77e0a),
	.w8(32'hbc11f111),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cca1b3e),
	.w1(32'h3ca6ba3a),
	.w2(32'h3c056660),
	.w3(32'hbc316809),
	.w4(32'h3b96740a),
	.w5(32'h3c444053),
	.w6(32'h3d96c518),
	.w7(32'hbae68b79),
	.w8(32'h3b89b8bc),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd012e9f),
	.w1(32'hbd85483d),
	.w2(32'h3bf95f3f),
	.w3(32'hb9d5ebf4),
	.w4(32'hbd416081),
	.w5(32'hbc2622d1),
	.w6(32'hbc695e34),
	.w7(32'h3b6e5e2f),
	.w8(32'hbd40b5b4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd00fd67),
	.w1(32'h3aacf92b),
	.w2(32'h3d03a5cb),
	.w3(32'hbb02966c),
	.w4(32'h3ae6d368),
	.w5(32'h3c01bb0d),
	.w6(32'hba95da03),
	.w7(32'h3ad6e14e),
	.w8(32'hbc6023e5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd22bd4b),
	.w1(32'hbc27a76f),
	.w2(32'hbc4221d3),
	.w3(32'h3c0589fd),
	.w4(32'h3c947704),
	.w5(32'hbca46a75),
	.w6(32'h3c30d05e),
	.w7(32'h3bd5cf66),
	.w8(32'h3cc49775),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c183e44),
	.w1(32'h3c052c66),
	.w2(32'h3ca11b37),
	.w3(32'h3ad8b992),
	.w4(32'h3c8d2ffc),
	.w5(32'hbd366c2e),
	.w6(32'hbce985ec),
	.w7(32'hbc079cc3),
	.w8(32'h3cc34e26),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c9ea4),
	.w1(32'h3d3a4136),
	.w2(32'hbbd600ed),
	.w3(32'hbc79a2e6),
	.w4(32'hbcf27387),
	.w5(32'h3c0ecf3c),
	.w6(32'h3d0d82e4),
	.w7(32'h3cf35c84),
	.w8(32'hbcabc412),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b142384),
	.w1(32'h3c5ef647),
	.w2(32'h3d88c077),
	.w3(32'hbd162e38),
	.w4(32'hb9a41b89),
	.w5(32'hbb2292e0),
	.w6(32'hbd135913),
	.w7(32'hbb9da908),
	.w8(32'h3badd5ca),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a0b29),
	.w1(32'h3b8c4750),
	.w2(32'hbb1cd243),
	.w3(32'hbac622e5),
	.w4(32'hbd2942c0),
	.w5(32'hbb0d9a45),
	.w6(32'h3c48d221),
	.w7(32'hbd1dd0d1),
	.w8(32'h3c28ed15),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0db473),
	.w1(32'hbd086f90),
	.w2(32'hbc3afa74),
	.w3(32'hbb85f0f3),
	.w4(32'h395ff68e),
	.w5(32'hbd0e0b8c),
	.w6(32'h3cb81748),
	.w7(32'h3bd680f4),
	.w8(32'h3caef6e6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfa73f4),
	.w1(32'hbd367958),
	.w2(32'hbc8b3edb),
	.w3(32'hbcfe8adc),
	.w4(32'hbc4bd686),
	.w5(32'h3b1c96d0),
	.w6(32'hbc3aad5d),
	.w7(32'h3b9b292a),
	.w8(32'h3cda36f9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34b157),
	.w1(32'hbb56fe5b),
	.w2(32'hbb8e139a),
	.w3(32'hbc7f6dec),
	.w4(32'h3bc5dfc6),
	.w5(32'hbd5aea37),
	.w6(32'hbc1f6ba5),
	.w7(32'hbbb30c86),
	.w8(32'hbd30e3c7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cbafc4),
	.w1(32'hbca23145),
	.w2(32'hb90a4e12),
	.w3(32'hbcbea48b),
	.w4(32'hbadc58aa),
	.w5(32'h3c8b9ba4),
	.w6(32'hbcef83d9),
	.w7(32'hbd378239),
	.w8(32'h3d123003),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2c7c2a),
	.w1(32'hb7cf6953),
	.w2(32'h3b8adf08),
	.w3(32'h3b9b5058),
	.w4(32'h3c30a2bd),
	.w5(32'h3a96da3c),
	.w6(32'hbc744ea1),
	.w7(32'hbbefb17d),
	.w8(32'h3d0c0c1a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ceafe),
	.w1(32'hbceb3a58),
	.w2(32'h3c09117e),
	.w3(32'hbc3157f8),
	.w4(32'hbd3efc60),
	.w5(32'h3b715420),
	.w6(32'h3c2f29af),
	.w7(32'h3c31ef31),
	.w8(32'h3ce8167d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb611df),
	.w1(32'hbba9d0dc),
	.w2(32'h3ca5c2a2),
	.w3(32'hba404a5e),
	.w4(32'hbe01c4f4),
	.w5(32'hbce57b47),
	.w6(32'hbc28a9fd),
	.w7(32'h3c38aef8),
	.w8(32'h3cbc36b3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4461f3),
	.w1(32'h3cde2ddb),
	.w2(32'hbcb95988),
	.w3(32'hbc2f7fc1),
	.w4(32'h3bed9416),
	.w5(32'hbbfa39c8),
	.w6(32'h3da6b351),
	.w7(32'h3d90ca35),
	.w8(32'h3c0740a7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b3108),
	.w1(32'hbbd724f7),
	.w2(32'hbdd0231a),
	.w3(32'h3caa7417),
	.w4(32'hbd0712b0),
	.w5(32'hbd361bf7),
	.w6(32'h3c09248a),
	.w7(32'hbd36ab51),
	.w8(32'hbca47197),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a376455),
	.w1(32'hbce6f456),
	.w2(32'hbc976c66),
	.w3(32'h3c1d63b3),
	.w4(32'h3cde2846),
	.w5(32'h3bb6007f),
	.w6(32'h3c64e8b3),
	.w7(32'h3a8692e7),
	.w8(32'h3c24d7ad),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d075edd),
	.w1(32'hb797ab8e),
	.w2(32'h3b9f924b),
	.w3(32'hbc7d3df2),
	.w4(32'hbbeefe6f),
	.w5(32'h3b79f5ed),
	.w6(32'h3bd0a55d),
	.w7(32'hbce114bb),
	.w8(32'h3c6c8f95),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdecfd0),
	.w1(32'hbc02724c),
	.w2(32'h3c2dc0b5),
	.w3(32'hbc93ef51),
	.w4(32'hbd33282b),
	.w5(32'hbc1b41e7),
	.w6(32'h3b03f407),
	.w7(32'hbdb4ebc7),
	.w8(32'h3cf2c581),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b144d5e),
	.w1(32'h3c840df7),
	.w2(32'hbb65d980),
	.w3(32'h3bb415a5),
	.w4(32'hbbb971c6),
	.w5(32'hbcba8409),
	.w6(32'hbb75a23a),
	.w7(32'h3a506911),
	.w8(32'hbdd50a76),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdefb23),
	.w1(32'h3bad9afc),
	.w2(32'hbcd5f45a),
	.w3(32'h3d0e0721),
	.w4(32'hbd1391a5),
	.w5(32'h39ca5582),
	.w6(32'h3c3a51fa),
	.w7(32'hbcb55342),
	.w8(32'h3d186007),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c363a19),
	.w1(32'h3c9f3388),
	.w2(32'h3d2df25a),
	.w3(32'hbd870836),
	.w4(32'h3c447072),
	.w5(32'h3c97f736),
	.w6(32'hbd5b1cf2),
	.w7(32'h3bbd9f7f),
	.w8(32'h3c903c6f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce9f2f5),
	.w1(32'hbccc7d0c),
	.w2(32'h3c5a544b),
	.w3(32'hbd72afde),
	.w4(32'hbc0e7959),
	.w5(32'h3c70f48c),
	.w6(32'hbc118aab),
	.w7(32'h3cdc62cc),
	.w8(32'h3d129d12),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ad662),
	.w1(32'hbb0163df),
	.w2(32'h3d1d136e),
	.w3(32'hbc4b1089),
	.w4(32'h3bdaf3f9),
	.w5(32'h3c1ebe14),
	.w6(32'hbd16ecb0),
	.w7(32'hbc47bcc2),
	.w8(32'h3c11a5fd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb19900),
	.w1(32'hbbd81092),
	.w2(32'hbd361026),
	.w3(32'h3beb6fbc),
	.w4(32'h3c8b4cce),
	.w5(32'h3b26e256),
	.w6(32'hbc5ea95f),
	.w7(32'hbc32628f),
	.w8(32'h3b8958dc),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e9483),
	.w1(32'h3b1929b1),
	.w2(32'h3c850207),
	.w3(32'hbc1f9777),
	.w4(32'hbc95eae6),
	.w5(32'hbbe606d4),
	.w6(32'h3c4a81b3),
	.w7(32'h3b056898),
	.w8(32'h3be47e14),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1feb6d),
	.w1(32'hbd0bdc5c),
	.w2(32'hbb8cb102),
	.w3(32'hbc9f865c),
	.w4(32'hbd04824e),
	.w5(32'hbb489311),
	.w6(32'h3c7d216e),
	.w7(32'h3a786c42),
	.w8(32'h3bdb1c1e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10fc3f),
	.w1(32'hbc0802aa),
	.w2(32'hb99e445f),
	.w3(32'hbd0491ab),
	.w4(32'h3b711f56),
	.w5(32'hbbab435e),
	.w6(32'h3be60503),
	.w7(32'hbac466cb),
	.w8(32'h3b345738),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cdacb),
	.w1(32'hbb8a889e),
	.w2(32'h3b2a883b),
	.w3(32'hbbbb89cf),
	.w4(32'h3b8754d2),
	.w5(32'hbba2664a),
	.w6(32'hbb2b3afc),
	.w7(32'h3c1c5ad2),
	.w8(32'hb97c606d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule