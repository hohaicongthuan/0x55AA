module layer_8_featuremap_168(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbdf76),
	.w1(32'h3968046a),
	.w2(32'h3afe8188),
	.w3(32'hbc1c00a9),
	.w4(32'hbbefe8c2),
	.w5(32'hb9b49ad8),
	.w6(32'hbc1791c6),
	.w7(32'hbc0d242c),
	.w8(32'hbc2a9efc),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba659f),
	.w1(32'h3c537ea0),
	.w2(32'h3cbfaa65),
	.w3(32'h3b1433ca),
	.w4(32'h3c15182c),
	.w5(32'h3ca40d7c),
	.w6(32'h3a99799e),
	.w7(32'h3b11aa70),
	.w8(32'hbc0c31a6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c4e01),
	.w1(32'h3c1c638c),
	.w2(32'h3b999648),
	.w3(32'h3c76e106),
	.w4(32'h3c13dabf),
	.w5(32'h3c57e362),
	.w6(32'h3c7adb31),
	.w7(32'h3c0fac8e),
	.w8(32'h3b840671),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaea05),
	.w1(32'h3bd27a72),
	.w2(32'h39e78048),
	.w3(32'h38c792d0),
	.w4(32'h3b9fdcc6),
	.w5(32'h3b0026e8),
	.w6(32'hbae4e352),
	.w7(32'hbb699417),
	.w8(32'hbc146b5e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba685c90),
	.w1(32'hbbf310f5),
	.w2(32'hbc0f0a54),
	.w3(32'hba8241e1),
	.w4(32'hbc90ece6),
	.w5(32'hbc97d0a0),
	.w6(32'hbbd38937),
	.w7(32'hb70e409c),
	.w8(32'h3c473c9c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b7cf6),
	.w1(32'hbb831dbf),
	.w2(32'hbc2c7ef9),
	.w3(32'h3b0cdc97),
	.w4(32'h3b1e5070),
	.w5(32'h3b812de4),
	.w6(32'h3b9bdd72),
	.w7(32'hba37704b),
	.w8(32'hba7cb7cc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beac100),
	.w1(32'hbcc0025b),
	.w2(32'hbce4fee2),
	.w3(32'h3bfaaa0f),
	.w4(32'hbcb14ee6),
	.w5(32'hbccbf49e),
	.w6(32'hbc158381),
	.w7(32'hbc03ddd9),
	.w8(32'h3c19a940),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3bd77),
	.w1(32'h3b0acdf7),
	.w2(32'h3c3ad25e),
	.w3(32'h3b0aaa96),
	.w4(32'h3c24d274),
	.w5(32'h3ca52556),
	.w6(32'h3b98d306),
	.w7(32'h3b3a8958),
	.w8(32'h3b96bbd7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bef01),
	.w1(32'hbcb6505a),
	.w2(32'hbca1e80e),
	.w3(32'h3bbf841b),
	.w4(32'hbd056f50),
	.w5(32'hbd02bf0b),
	.w6(32'hbb063efa),
	.w7(32'hbbd404dd),
	.w8(32'h3c2c5a55),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc055e),
	.w1(32'hbb970710),
	.w2(32'h3c01dadd),
	.w3(32'hbb98dcc4),
	.w4(32'h3b44bfff),
	.w5(32'h3c035b9e),
	.w6(32'h3b9341f3),
	.w7(32'h3bbc5eb2),
	.w8(32'hbbcae8c3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc04c8),
	.w1(32'h3baf1a4f),
	.w2(32'h3c85754c),
	.w3(32'hbc308b99),
	.w4(32'hbbc77b1d),
	.w5(32'h3abe8259),
	.w6(32'hbc30e25e),
	.w7(32'hbc081904),
	.w8(32'h3ba2ea1e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab845ee),
	.w1(32'h3a0a615e),
	.w2(32'h3badb388),
	.w3(32'hbb8bea04),
	.w4(32'hbba8e1ca),
	.w5(32'h3b01d812),
	.w6(32'h3b6da9bc),
	.w7(32'h3b16237c),
	.w8(32'hbb9e844d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b931f4d),
	.w1(32'hbb14b431),
	.w2(32'hbb65c4ce),
	.w3(32'h3be77f92),
	.w4(32'h3b0d3bce),
	.w5(32'hbb341d8a),
	.w6(32'h3b582fdb),
	.w7(32'h3ba2c953),
	.w8(32'hbb41c2b2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5934f),
	.w1(32'h3bc0e848),
	.w2(32'h3b972ea0),
	.w3(32'hba8bd282),
	.w4(32'hbb27276f),
	.w5(32'h39ea98ef),
	.w6(32'h3bd1c101),
	.w7(32'h3a87b8a8),
	.w8(32'hbb0e7fd9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7831b),
	.w1(32'h3d0fee32),
	.w2(32'h3d0afbb2),
	.w3(32'h3a910896),
	.w4(32'h3d03a378),
	.w5(32'h3d0faa23),
	.w6(32'h3c6f9855),
	.w7(32'hb933ef3f),
	.w8(32'hbcc65efd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb448187),
	.w1(32'h3a92282d),
	.w2(32'h3bd55264),
	.w3(32'h392da380),
	.w4(32'h3be898a6),
	.w5(32'h3991f7b9),
	.w6(32'hb98f60cb),
	.w7(32'h3b9a1509),
	.w8(32'h3af752b3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa18300),
	.w1(32'hbb418b2d),
	.w2(32'hbbf0b9b6),
	.w3(32'hba894517),
	.w4(32'hbbc72a03),
	.w5(32'hbaf801a0),
	.w6(32'hb929e8b5),
	.w7(32'hbb72cb65),
	.w8(32'hb95b25fd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c24d6),
	.w1(32'h3c5d465b),
	.w2(32'h3c443bd6),
	.w3(32'h3bd941f2),
	.w4(32'h3c3ae068),
	.w5(32'h3c3257a0),
	.w6(32'h3c7331b3),
	.w7(32'h3c65b8c9),
	.w8(32'h3b3db317),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb732d38),
	.w1(32'h3cf29610),
	.w2(32'h3d17b246),
	.w3(32'hbd00585b),
	.w4(32'h3c048587),
	.w5(32'h3cb1f9f6),
	.w6(32'hbc838e80),
	.w7(32'hbbbb909f),
	.w8(32'h3b1de5c3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dafec),
	.w1(32'hbcbc4332),
	.w2(32'hbcd4a0bf),
	.w3(32'hbbda7b22),
	.w4(32'hbcb664c0),
	.w5(32'hbcf475b9),
	.w6(32'hbce0b287),
	.w7(32'hbced4bee),
	.w8(32'hbb01ba5a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79423f),
	.w1(32'h3b10a133),
	.w2(32'hbb39366e),
	.w3(32'hb962a9cc),
	.w4(32'h3b420b84),
	.w5(32'hbc2530e6),
	.w6(32'h3bd8c638),
	.w7(32'h3af12d05),
	.w8(32'hbc316cf7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2bbdf),
	.w1(32'h3b0637b7),
	.w2(32'hbb201dce),
	.w3(32'h3c0d6da2),
	.w4(32'h3c00637e),
	.w5(32'h3bde8374),
	.w6(32'h3bf7aaac),
	.w7(32'h3c3955d3),
	.w8(32'h3bc21a57),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a248ce1),
	.w1(32'h3cf59804),
	.w2(32'h3d158c45),
	.w3(32'hbc94dd98),
	.w4(32'h3bc8e166),
	.w5(32'h3cee8425),
	.w6(32'hbb7e77cd),
	.w7(32'hbc062ac3),
	.w8(32'h3bba4197),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fc75e),
	.w1(32'hbadefa31),
	.w2(32'h3aea846b),
	.w3(32'hba7b6dbc),
	.w4(32'h3c16d1b7),
	.w5(32'hb9e3e07c),
	.w6(32'h3b764a6b),
	.w7(32'h39264fd5),
	.w8(32'h3a4a35ff),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e5186),
	.w1(32'h394b3257),
	.w2(32'hba978a0a),
	.w3(32'hbc08346d),
	.w4(32'hbaa963e3),
	.w5(32'hbb2b87f6),
	.w6(32'hbb6b44d6),
	.w7(32'hba7c0303),
	.w8(32'hbb8b3715),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc548abf),
	.w1(32'hba2997c6),
	.w2(32'h3c18f76f),
	.w3(32'hbcce20d3),
	.w4(32'hbc6622e9),
	.w5(32'hbbce6e02),
	.w6(32'hbcea7ef4),
	.w7(32'hbca7b838),
	.w8(32'hbc9de33a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981ec49),
	.w1(32'hbb05871a),
	.w2(32'h3a8be331),
	.w3(32'hbb4980a0),
	.w4(32'hb966ef34),
	.w5(32'h3b5aee69),
	.w6(32'hbbd4f520),
	.w7(32'hbbefd702),
	.w8(32'hbc0e1ee0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf9e901),
	.w1(32'h3c03581c),
	.w2(32'h3db648b0),
	.w3(32'hbdb31bcf),
	.w4(32'hbd893cbb),
	.w5(32'h3a8bc0d2),
	.w6(32'hbdae21f7),
	.w7(32'hbd73f279),
	.w8(32'hbcdd66fa),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c0ca7),
	.w1(32'h3bcd91ac),
	.w2(32'h3bd73ff5),
	.w3(32'hbbd22a54),
	.w4(32'h3a9e287a),
	.w5(32'h3befaf16),
	.w6(32'h3b00149a),
	.w7(32'hbba8ffa2),
	.w8(32'hbb69dab3),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1bfe4),
	.w1(32'hbafa943f),
	.w2(32'h3bfb2183),
	.w3(32'h3b792971),
	.w4(32'h3b90cd0e),
	.w5(32'h3c3e2d7a),
	.w6(32'hb98fc64c),
	.w7(32'hbbd868ac),
	.w8(32'hbc224ef6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3a7c4),
	.w1(32'hbbc1d568),
	.w2(32'hbbc62576),
	.w3(32'h3bf3d237),
	.w4(32'hbc02d1f2),
	.w5(32'hb98b6584),
	.w6(32'h3aa3e07a),
	.w7(32'h3b099773),
	.w8(32'hbaf8c493),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5f48b),
	.w1(32'hbb29e0fc),
	.w2(32'h3bab8656),
	.w3(32'hbba5b5d5),
	.w4(32'hbc18f9ee),
	.w5(32'h3998a7bb),
	.w6(32'hbc46af61),
	.w7(32'hbb13b645),
	.w8(32'hbb92861f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffdb5f),
	.w1(32'h390e0b76),
	.w2(32'hba995418),
	.w3(32'h3b87823e),
	.w4(32'hbac00bf3),
	.w5(32'h3aa01e55),
	.w6(32'h3b672a4d),
	.w7(32'h3aa93e9e),
	.w8(32'hbb45d671),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52651e),
	.w1(32'hba45a5b4),
	.w2(32'h3b0b22f9),
	.w3(32'hbb20b5b3),
	.w4(32'hbabb79c2),
	.w5(32'h3a44cd14),
	.w6(32'hbbcdf76f),
	.w7(32'h3b7a3e39),
	.w8(32'h3b78fd40),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38189c),
	.w1(32'hbc5d52db),
	.w2(32'hbbfae0a3),
	.w3(32'hbb401647),
	.w4(32'hba4e15e7),
	.w5(32'hba1575b0),
	.w6(32'h3a4c3cbe),
	.w7(32'hbaaa47ee),
	.w8(32'hbb9b5cce),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc553543),
	.w1(32'hba61bb20),
	.w2(32'h3c4dfe15),
	.w3(32'hbc132da3),
	.w4(32'hbc17fbaf),
	.w5(32'h3acf912e),
	.w6(32'hbc5b0563),
	.w7(32'hbbd691bb),
	.w8(32'hb8c05ec7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb191e62),
	.w1(32'h3bb02fff),
	.w2(32'h3ad82188),
	.w3(32'hba89e293),
	.w4(32'h3bb11144),
	.w5(32'h3b83c509),
	.w6(32'h3b52228e),
	.w7(32'hbaddcc9a),
	.w8(32'hbb91c1ad),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59e8f9),
	.w1(32'h3d981e54),
	.w2(32'h3da0ccc2),
	.w3(32'hbb3eed5b),
	.w4(32'h3d7a8a2c),
	.w5(32'h3d8d1eb7),
	.w6(32'h3ce7b6d9),
	.w7(32'h3c1d5779),
	.w8(32'hbd1d96a6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6efede),
	.w1(32'h3b772dd7),
	.w2(32'hba600e2f),
	.w3(32'h3b9e36ac),
	.w4(32'h3b983b4e),
	.w5(32'h3a46ef47),
	.w6(32'h3ba506d2),
	.w7(32'hba777210),
	.w8(32'hbb3574f3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10968f),
	.w1(32'hbaf0dc1e),
	.w2(32'h3b40e4dd),
	.w3(32'hbae90ad6),
	.w4(32'hbab512b0),
	.w5(32'hbb16f316),
	.w6(32'hb9d78b75),
	.w7(32'h3b470601),
	.w8(32'h3be0f675),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c996c),
	.w1(32'h3c14e39a),
	.w2(32'h3c95296d),
	.w3(32'hbc1f9623),
	.w4(32'h3b1b11c6),
	.w5(32'h3c6c7e1e),
	.w6(32'hbb7868af),
	.w7(32'hb99b923c),
	.w8(32'hbc3f107e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c20c7),
	.w1(32'h3c192f02),
	.w2(32'h3c657378),
	.w3(32'h3c0c5009),
	.w4(32'h3c5a2e7b),
	.w5(32'h3c5f165b),
	.w6(32'h3c561ed8),
	.w7(32'h3be60b9e),
	.w8(32'h3c172e04),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c13e2),
	.w1(32'h3be218e7),
	.w2(32'h3acdc3eb),
	.w3(32'h3c692a5f),
	.w4(32'h3bfd9f92),
	.w5(32'h3b96db1d),
	.w6(32'h3bcaa99f),
	.w7(32'h3ac18cb4),
	.w8(32'h3ac02291),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb533064),
	.w1(32'h3b34152b),
	.w2(32'h3ba87f97),
	.w3(32'hbb231b32),
	.w4(32'h394987ff),
	.w5(32'h3b7b9bb2),
	.w6(32'hba718b9b),
	.w7(32'h3b1986d2),
	.w8(32'hbb3c69ca),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5456fc),
	.w1(32'hbbc6aa54),
	.w2(32'h3be46bfb),
	.w3(32'hbc34f975),
	.w4(32'hbbf4987d),
	.w5(32'h3c0a11e6),
	.w6(32'hbca16e29),
	.w7(32'hbc5f7f44),
	.w8(32'h3b0d77b2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cc847),
	.w1(32'hbc141349),
	.w2(32'hbc03350c),
	.w3(32'hba22ca8e),
	.w4(32'hbb8d6626),
	.w5(32'hba28934d),
	.w6(32'h3ab9b79b),
	.w7(32'hbb692426),
	.w8(32'h3b4edf9f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8505c),
	.w1(32'hba81988c),
	.w2(32'hbbbf3739),
	.w3(32'h39c79fc4),
	.w4(32'h3b15f56a),
	.w5(32'hbb2b2826),
	.w6(32'h3a8323be),
	.w7(32'hbb191a13),
	.w8(32'h3b61eb60),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6f063),
	.w1(32'h3b9ca7d6),
	.w2(32'h3c980545),
	.w3(32'hbc061488),
	.w4(32'hbb144bf6),
	.w5(32'hbab3c1e4),
	.w6(32'hbc710af4),
	.w7(32'hbc11c14d),
	.w8(32'hbc022e0d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e6a61),
	.w1(32'h3b4819a2),
	.w2(32'h3bafa9b0),
	.w3(32'hba9d2a52),
	.w4(32'h3b8ba190),
	.w5(32'h3ba6fc32),
	.w6(32'h3bdc1256),
	.w7(32'h3c3deea8),
	.w8(32'h3b3bb996),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9be4ec),
	.w1(32'h3ad82202),
	.w2(32'h3a46c442),
	.w3(32'hbc3258a9),
	.w4(32'hbaa2d332),
	.w5(32'h3b1a42a5),
	.w6(32'hbbc44ac9),
	.w7(32'hbb0bb5d6),
	.w8(32'hbbb6361f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41494a),
	.w1(32'h3c99b84b),
	.w2(32'h3d65465d),
	.w3(32'h3b5d1e10),
	.w4(32'h3c30064c),
	.w5(32'h3cc3bd19),
	.w6(32'h3b91fadd),
	.w7(32'h3c196833),
	.w8(32'hbcd8b1fb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c6ed1),
	.w1(32'h3c9a55fa),
	.w2(32'h3c7d312e),
	.w3(32'hbc86247b),
	.w4(32'h3c91d28e),
	.w5(32'h3cead65b),
	.w6(32'hbcbc9a8b),
	.w7(32'hbc65f735),
	.w8(32'hbbb87dc6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb429461),
	.w1(32'h3d87382d),
	.w2(32'h3db53ac6),
	.w3(32'hbba6d6ed),
	.w4(32'h3d7010a5),
	.w5(32'h3daef9b4),
	.w6(32'h3b7a4064),
	.w7(32'h3ab7671e),
	.w8(32'hbd314f05),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b930c9c),
	.w1(32'hbbaff132),
	.w2(32'h3c2187a9),
	.w3(32'h3bf1c5ac),
	.w4(32'h3b705990),
	.w5(32'h3c625023),
	.w6(32'h3c178275),
	.w7(32'h3c49a3a0),
	.w8(32'h3c1c252d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5406ee),
	.w1(32'h3c1a5ef2),
	.w2(32'hbacee4bb),
	.w3(32'h3b1c8f5c),
	.w4(32'h3b695d6c),
	.w5(32'hbb313174),
	.w6(32'h3bad27fd),
	.w7(32'h3b803cb4),
	.w8(32'h3b6857ad),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe88649),
	.w1(32'h3c00c314),
	.w2(32'h3cb2de1e),
	.w3(32'hbc91a2f9),
	.w4(32'hbbdcd45a),
	.w5(32'h3bf59171),
	.w6(32'hbbac0034),
	.w7(32'hbb044aff),
	.w8(32'h3b9807d3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37800b),
	.w1(32'hbb580ba8),
	.w2(32'hb8d426fa),
	.w3(32'h3b12e7a4),
	.w4(32'h3bb7f1c6),
	.w5(32'h3b4a4162),
	.w6(32'h3bcd22a0),
	.w7(32'h3aa5aa6d),
	.w8(32'h3b66c472),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c093923),
	.w1(32'h3c99938e),
	.w2(32'h3c0ab163),
	.w3(32'h3b91b152),
	.w4(32'h3ca430ea),
	.w5(32'h3c986f0e),
	.w6(32'h3c5f80b0),
	.w7(32'h3c104465),
	.w8(32'h3c557e9b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be91354),
	.w1(32'h3cb15866),
	.w2(32'h3ce5b577),
	.w3(32'h3c1829df),
	.w4(32'h3c8a2f91),
	.w5(32'h3cf0e1bb),
	.w6(32'h3b0962fc),
	.w7(32'h3bd1bea4),
	.w8(32'hb9a8092a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80bfdda),
	.w1(32'h3b3f864c),
	.w2(32'hbb233632),
	.w3(32'h3b103d21),
	.w4(32'h3b9ad2c8),
	.w5(32'hbb99b144),
	.w6(32'hbbd513f3),
	.w7(32'hbb5e9c90),
	.w8(32'hbc07424b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb63ea),
	.w1(32'hbb54419d),
	.w2(32'h3a3a4714),
	.w3(32'hbc15f188),
	.w4(32'h3b65bead),
	.w5(32'h3bda8a96),
	.w6(32'h3aa23cc8),
	.w7(32'hbb57ab0c),
	.w8(32'h398bd5d4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04d083),
	.w1(32'hbb79cb8c),
	.w2(32'hbb8ce000),
	.w3(32'h3b2f8253),
	.w4(32'hba24eeff),
	.w5(32'h3b36ed92),
	.w6(32'h3a064e09),
	.w7(32'hba9c6d14),
	.w8(32'h39a1364a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0484cc),
	.w1(32'hbc82ac6a),
	.w2(32'hbbc2bc73),
	.w3(32'hbb925398),
	.w4(32'hbc923606),
	.w5(32'hbba6008a),
	.w6(32'hbc736c01),
	.w7(32'hbc597f0a),
	.w8(32'hbabdf741),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f85c0),
	.w1(32'h3c27aa6d),
	.w2(32'h3c8532eb),
	.w3(32'h3bd86bfd),
	.w4(32'h3c6b82a1),
	.w5(32'h3c91a1cf),
	.w6(32'h3b9a6859),
	.w7(32'h3c65749b),
	.w8(32'h3c2ee30b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c398503),
	.w1(32'h3d60ce25),
	.w2(32'h3d870aa3),
	.w3(32'h3bfe1c81),
	.w4(32'h3d57d208),
	.w5(32'h3d8a5cc8),
	.w6(32'h3ca0fdf7),
	.w7(32'h3c5283b5),
	.w8(32'hbcccd714),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ad3b4),
	.w1(32'h3af36652),
	.w2(32'h3c3df0fa),
	.w3(32'h3c4ff8e0),
	.w4(32'hbab304ea),
	.w5(32'h3b8a900c),
	.w6(32'h3a38ab56),
	.w7(32'h3bd16300),
	.w8(32'h3c0c7450),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8f895),
	.w1(32'h3b29564f),
	.w2(32'hbaaf4c68),
	.w3(32'h3b40ad7f),
	.w4(32'hba66918a),
	.w5(32'hba8896b8),
	.w6(32'h3b4612dd),
	.w7(32'h3ab47fc7),
	.w8(32'h3b09459d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27ab8e),
	.w1(32'hbbb0b83b),
	.w2(32'hbc039309),
	.w3(32'hbbcba628),
	.w4(32'hbbc173a4),
	.w5(32'hbc5d54a6),
	.w6(32'hbae83c8b),
	.w7(32'hbb3d8ea2),
	.w8(32'hbb6518e3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37596f),
	.w1(32'h3888f9b2),
	.w2(32'hba30bec6),
	.w3(32'hbb34c512),
	.w4(32'hbb8812eb),
	.w5(32'hbb981e9c),
	.w6(32'h3b34fd27),
	.w7(32'h38ef6001),
	.w8(32'hb9c06ea2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4496c8),
	.w1(32'h3c3a40eb),
	.w2(32'h3cf42103),
	.w3(32'hbca92c03),
	.w4(32'hbba90686),
	.w5(32'h3c550254),
	.w6(32'hbcb889ca),
	.w7(32'hbc932141),
	.w8(32'hbc365a7d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb956f9e),
	.w1(32'h3a5372e0),
	.w2(32'hbab2fae5),
	.w3(32'h3a16bff6),
	.w4(32'hbb681e33),
	.w5(32'hba9eddc8),
	.w6(32'hb9a2e81e),
	.w7(32'hbbc699cd),
	.w8(32'h3c1dd87c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95cd50),
	.w1(32'h3a97c55e),
	.w2(32'h3bac6812),
	.w3(32'h3c539359),
	.w4(32'hbb1b8cf8),
	.w5(32'h39bd530d),
	.w6(32'hbb893637),
	.w7(32'hbc2141ee),
	.w8(32'hbbb1f1a8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdda718),
	.w1(32'hbbf8c39b),
	.w2(32'h3aa6ccbe),
	.w3(32'hba4e3c2f),
	.w4(32'h3b030f69),
	.w5(32'h3bbaef25),
	.w6(32'hba9e3137),
	.w7(32'hbb044489),
	.w8(32'hba985a87),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe087a2),
	.w1(32'hbab8d965),
	.w2(32'h3b50ef06),
	.w3(32'hbc0f35ed),
	.w4(32'hbb417771),
	.w5(32'hbba38cc3),
	.w6(32'hba87ddc9),
	.w7(32'hbbda439a),
	.w8(32'hbb3b13ae),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec1125),
	.w1(32'h3be0e00a),
	.w2(32'hbb371433),
	.w3(32'h3a041f7b),
	.w4(32'h3bb9eda2),
	.w5(32'h39f04a82),
	.w6(32'h3b7f47c2),
	.w7(32'h3aa89d40),
	.w8(32'h3b8e707b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9072103),
	.w1(32'h3bbdef88),
	.w2(32'h3b29fd5c),
	.w3(32'hbacb0284),
	.w4(32'h3b5b55d4),
	.w5(32'h3bbed27a),
	.w6(32'hbb4ccf93),
	.w7(32'hbbb7d6f2),
	.w8(32'hbb10e204),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4640cc),
	.w1(32'h3b8dc04c),
	.w2(32'hba842f02),
	.w3(32'h3ae2b583),
	.w4(32'h3b0d5f22),
	.w5(32'hb8bf8143),
	.w6(32'h3bb427e1),
	.w7(32'h39ec1f9c),
	.w8(32'hba320ceb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb903048),
	.w1(32'h3c9325e5),
	.w2(32'h3cd6d60e),
	.w3(32'hbc6abd67),
	.w4(32'h3b3e8ba9),
	.w5(32'h3c56a9de),
	.w6(32'hbbed39ae),
	.w7(32'hbabadc57),
	.w8(32'hbc00e42c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc322270),
	.w1(32'hba860452),
	.w2(32'h3bc6afa5),
	.w3(32'hbbeffb1d),
	.w4(32'h39edd55b),
	.w5(32'h3c133f53),
	.w6(32'h3b8d8eb2),
	.w7(32'h3a878f22),
	.w8(32'h3c23d18b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e3117),
	.w1(32'hb7c2743e),
	.w2(32'hba2c0bfa),
	.w3(32'h3b6ca28a),
	.w4(32'h3b5f51e1),
	.w5(32'h3ad63f78),
	.w6(32'h3bbc2da5),
	.w7(32'h3b59bb43),
	.w8(32'h3b026ff5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00e202),
	.w1(32'h3b1d12ea),
	.w2(32'h3b8c04ba),
	.w3(32'h3a34c32e),
	.w4(32'hba409607),
	.w5(32'h3b801911),
	.w6(32'h3a2f37c9),
	.w7(32'hbae5223a),
	.w8(32'h39912f8a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20c899),
	.w1(32'h3bc1c1bc),
	.w2(32'hba8841dd),
	.w3(32'h390cc79c),
	.w4(32'hba4034c0),
	.w5(32'hbb05cba6),
	.w6(32'hbb603d0b),
	.w7(32'hbbb2605a),
	.w8(32'hba083c8f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25f3fb),
	.w1(32'h39c69117),
	.w2(32'h3c0c0f64),
	.w3(32'hbc2bf2e9),
	.w4(32'hbc125a48),
	.w5(32'h3b64e331),
	.w6(32'hbc89bede),
	.w7(32'hbc8ad371),
	.w8(32'hbc3191a3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b74ff),
	.w1(32'hbbc77e0c),
	.w2(32'hbc9677dd),
	.w3(32'hbc1c7d73),
	.w4(32'hbb185b28),
	.w5(32'hbbfbc314),
	.w6(32'hbb91f9a0),
	.w7(32'hbc01d863),
	.w8(32'hbcc01f97),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e0f56),
	.w1(32'h3c1a658e),
	.w2(32'h3c5b1398),
	.w3(32'hbcaae191),
	.w4(32'hbc43100e),
	.w5(32'h3b889110),
	.w6(32'hbcd63261),
	.w7(32'hbcbf7f53),
	.w8(32'hbc8ca01c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54f0e1),
	.w1(32'h3ac6cdba),
	.w2(32'h3c6635e9),
	.w3(32'hbc480218),
	.w4(32'hbb2f3bc5),
	.w5(32'h3c38bb17),
	.w6(32'hbc9c34b7),
	.w7(32'hbc875986),
	.w8(32'hbc4bf7c9),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53d9df),
	.w1(32'h3ad1e5fa),
	.w2(32'h3ab6b597),
	.w3(32'h3b6cbbd4),
	.w4(32'h3aa762a4),
	.w5(32'h3b0b4ae3),
	.w6(32'h3b30c4e6),
	.w7(32'h3b3391d2),
	.w8(32'h3b4f5b2a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16bf6c),
	.w1(32'h3a0236c1),
	.w2(32'h3a6cbdef),
	.w3(32'h3b3cdabf),
	.w4(32'h3bcbb342),
	.w5(32'h3bd295c2),
	.w6(32'hbb380577),
	.w7(32'hbb8759da),
	.w8(32'hb9e2007d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ad892),
	.w1(32'h3a6b2c07),
	.w2(32'h3b687092),
	.w3(32'hba259090),
	.w4(32'hb8d525e4),
	.w5(32'h3abf4d4f),
	.w6(32'h3b56957d),
	.w7(32'h3b0f4b93),
	.w8(32'h3aa152b6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9fbb7),
	.w1(32'h3b7ef827),
	.w2(32'h3c1fab58),
	.w3(32'hbbb58002),
	.w4(32'h3b175d86),
	.w5(32'h3bb9b57b),
	.w6(32'hbc019a2e),
	.w7(32'hbc1db9e2),
	.w8(32'hbc0cf6a8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e8510),
	.w1(32'h3b273e12),
	.w2(32'hbb6b7e7d),
	.w3(32'hbb1d4e5b),
	.w4(32'hbaaf9092),
	.w5(32'h3b15b21c),
	.w6(32'hb9a46231),
	.w7(32'hbb8736ec),
	.w8(32'hbbb99637),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8900eb),
	.w1(32'hbbc33e0f),
	.w2(32'hbbd3107b),
	.w3(32'hbbdacb3c),
	.w4(32'hbb988b62),
	.w5(32'h39e4db66),
	.w6(32'hba64e50a),
	.w7(32'h3ab498e1),
	.w8(32'h3aae12bb),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a915155),
	.w1(32'hbc8cf258),
	.w2(32'hbc8e4c1d),
	.w3(32'h3bd7efcb),
	.w4(32'hbc68892a),
	.w5(32'hbcb3819b),
	.w6(32'hbc053663),
	.w7(32'hbb794f75),
	.w8(32'h3bdd06e4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9abe5),
	.w1(32'h3b88ed58),
	.w2(32'h3b8f9da2),
	.w3(32'h3a8f1f99),
	.w4(32'h3ab87aab),
	.w5(32'h3b751d61),
	.w6(32'h3a0a5e71),
	.w7(32'h3a54a83f),
	.w8(32'h3b82a621),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab14d7c),
	.w1(32'h3b8dea61),
	.w2(32'h3b4460e7),
	.w3(32'h3ad8e734),
	.w4(32'h3a9f53c9),
	.w5(32'h3bbed43d),
	.w6(32'h3b77b72e),
	.w7(32'h3b316962),
	.w8(32'hbbad1ad4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a265b),
	.w1(32'h3b5e6fbd),
	.w2(32'h3b96decc),
	.w3(32'hbc18a6a3),
	.w4(32'h3b03e63f),
	.w5(32'h3b1133c7),
	.w6(32'h3a5f1d0e),
	.w7(32'hba0a8569),
	.w8(32'h3b383ad2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33fb78),
	.w1(32'h3c9ba0c8),
	.w2(32'h3c22cdc7),
	.w3(32'hbc82b33b),
	.w4(32'h3bb0d560),
	.w5(32'h3b9724f4),
	.w6(32'hbc4263e1),
	.w7(32'hbc6a57b0),
	.w8(32'hbca41b5d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb547970),
	.w1(32'h3ba08e22),
	.w2(32'h3c1fbdc6),
	.w3(32'h3b381588),
	.w4(32'h3c2151b4),
	.w5(32'h3c0d5aa5),
	.w6(32'h3b966946),
	.w7(32'h3bfdef7a),
	.w8(32'h3a09c2d4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15e2a6),
	.w1(32'hba7ecaac),
	.w2(32'h3be757d5),
	.w3(32'h3b3fab23),
	.w4(32'h3b162f88),
	.w5(32'h3c119ce1),
	.w6(32'h3abb04e2),
	.w7(32'h3ba72d17),
	.w8(32'hbafb614e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6425f),
	.w1(32'h3b60c98e),
	.w2(32'h3ba2b383),
	.w3(32'h3b8dd468),
	.w4(32'hbbfa751a),
	.w5(32'h3b5b2357),
	.w6(32'h3ac799bc),
	.w7(32'h3b7c8bc7),
	.w8(32'hbb784968),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39415b9b),
	.w1(32'h3b0368b2),
	.w2(32'h3b994a21),
	.w3(32'h3b5d074e),
	.w4(32'h3a081522),
	.w5(32'h3b96f67d),
	.w6(32'h3bbf77ce),
	.w7(32'h3b212208),
	.w8(32'h39995446),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983ce82),
	.w1(32'hbb20aaa4),
	.w2(32'h3bf35691),
	.w3(32'hb9c642fc),
	.w4(32'hbaa98726),
	.w5(32'h3c284f24),
	.w6(32'hbb9907f5),
	.w7(32'hbb7889a7),
	.w8(32'hbb6bd777),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08385f),
	.w1(32'hbb6340e9),
	.w2(32'hbb9d1d1c),
	.w3(32'hbaa5d230),
	.w4(32'hbb91f9bf),
	.w5(32'hbc12f46d),
	.w6(32'hbbdf17e1),
	.w7(32'hbb761bf8),
	.w8(32'hbb5619fe),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2777f9),
	.w1(32'h3a5561dd),
	.w2(32'hb9b87a69),
	.w3(32'h3b508e2d),
	.w4(32'h3b80e7f5),
	.w5(32'h3ab8c30b),
	.w6(32'hbae69984),
	.w7(32'hbb5c0fe3),
	.w8(32'hba3b573b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7444d5),
	.w1(32'hbb359b2f),
	.w2(32'hbace8a63),
	.w3(32'hbbe14c5b),
	.w4(32'h3933bd0c),
	.w5(32'h3bb6ebf2),
	.w6(32'h3b0f327a),
	.w7(32'h3b0ae5d9),
	.w8(32'h3b761970),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcca72f),
	.w1(32'h3d158ea7),
	.w2(32'h3d560865),
	.w3(32'hbc20879e),
	.w4(32'h3cf1bee3),
	.w5(32'h3d5aed22),
	.w6(32'hbbe3a932),
	.w7(32'hbc829247),
	.w8(32'hbd1d11a6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41a902),
	.w1(32'h3ba80819),
	.w2(32'h3c15931f),
	.w3(32'hbbebeb68),
	.w4(32'h3a3b3252),
	.w5(32'h3b06dda0),
	.w6(32'hbbe443ad),
	.w7(32'hbba9978a),
	.w8(32'hbbcda796),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8700f),
	.w1(32'h3b91ebbd),
	.w2(32'h3b88e111),
	.w3(32'h3b0c42ba),
	.w4(32'h3baf4d09),
	.w5(32'h3c05e36f),
	.w6(32'h3bb656b2),
	.w7(32'h3b5f674b),
	.w8(32'h39004c8e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb645a6a),
	.w1(32'h3a97c08f),
	.w2(32'h3b9b7849),
	.w3(32'h3c26e5c9),
	.w4(32'h3b93d796),
	.w5(32'h3b09cc64),
	.w6(32'h3c1d65e0),
	.w7(32'h3be9fbe4),
	.w8(32'h3b8a3533),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96206f),
	.w1(32'h3ce8822a),
	.w2(32'h3d1a1709),
	.w3(32'hbbb7d5e2),
	.w4(32'h3c7808ac),
	.w5(32'h3cc922db),
	.w6(32'h3b50a49a),
	.w7(32'h3ab73302),
	.w8(32'hbc6fc93c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945cd5d),
	.w1(32'hbbc5ed8b),
	.w2(32'hbc1251fb),
	.w3(32'h3a45975c),
	.w4(32'hbc41b4b7),
	.w5(32'hbc5ca6cd),
	.w6(32'h3b33289e),
	.w7(32'h39ccce4d),
	.w8(32'hbb7aa0d0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5cd97a),
	.w1(32'hbbbad8d3),
	.w2(32'hbc057dda),
	.w3(32'h3bd75574),
	.w4(32'hbbbe656a),
	.w5(32'hbc2f5e04),
	.w6(32'h3c085865),
	.w7(32'h3b87473d),
	.w8(32'h3c45d797),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7dcdf7),
	.w1(32'hbbaf3b5c),
	.w2(32'h3b3a5f3b),
	.w3(32'h3bf97572),
	.w4(32'h3b6afb74),
	.w5(32'h38a8e9f3),
	.w6(32'h3c87f186),
	.w7(32'h3c0490bd),
	.w8(32'h3c5a3df4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7185f9),
	.w1(32'h3a6aa5af),
	.w2(32'hbb875e7e),
	.w3(32'hb9c7622c),
	.w4(32'hba9eb0ac),
	.w5(32'h3a1dac3d),
	.w6(32'hb741711d),
	.w7(32'hbb41fc7f),
	.w8(32'hbbe6ae58),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf63db),
	.w1(32'h3a8adddf),
	.w2(32'hb9101b94),
	.w3(32'hbb927829),
	.w4(32'hbb01f61d),
	.w5(32'h3b8a77e9),
	.w6(32'h3ad672de),
	.w7(32'h3a8f5a91),
	.w8(32'h3b065a5c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61e6cc),
	.w1(32'h3d38fed6),
	.w2(32'h3d5b1daa),
	.w3(32'hbafce67e),
	.w4(32'h3d18ad1d),
	.w5(32'h3d48def5),
	.w6(32'h3c793014),
	.w7(32'h3c31be8e),
	.w8(32'hbc83c001),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e6a87),
	.w1(32'h3b6d29f0),
	.w2(32'h3c10190b),
	.w3(32'h3c6bec60),
	.w4(32'h3aa0ece3),
	.w5(32'h3b8e3607),
	.w6(32'h3bc479e1),
	.w7(32'h3c08b159),
	.w8(32'h3b8bae82),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8107c9),
	.w1(32'hbb8323c0),
	.w2(32'h3b0938f4),
	.w3(32'hba3db8e3),
	.w4(32'hbb86d11e),
	.w5(32'h3a299f72),
	.w6(32'hbb89ab92),
	.w7(32'h3b08d4a8),
	.w8(32'h3b7637c4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f7b74),
	.w1(32'hbb103a5b),
	.w2(32'h3a982d4c),
	.w3(32'hb90ecf57),
	.w4(32'hbb1e14e5),
	.w5(32'hba6e5327),
	.w6(32'h3a1de43c),
	.w7(32'h3aca127c),
	.w8(32'hbab87b93),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba72dd9),
	.w1(32'h3b1a5d1c),
	.w2(32'h3a17257f),
	.w3(32'h3b427038),
	.w4(32'h3bbfb9f5),
	.w5(32'h3b03e83f),
	.w6(32'h3b52630a),
	.w7(32'h3b400645),
	.w8(32'h3ba81971),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bdc71),
	.w1(32'hbb294378),
	.w2(32'hbaf34bda),
	.w3(32'h3c0bc277),
	.w4(32'h3b52a9d0),
	.w5(32'h3af38619),
	.w6(32'hbb71adc1),
	.w7(32'h3b12c690),
	.w8(32'h3916d5dc),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a6e2a),
	.w1(32'hbbc82496),
	.w2(32'h3bbad864),
	.w3(32'hbc5abf32),
	.w4(32'hbc1e3ee7),
	.w5(32'hbb3bfbf0),
	.w6(32'hbc765955),
	.w7(32'hbc523c57),
	.w8(32'hbbbe56ae),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c14c8),
	.w1(32'hbca112b0),
	.w2(32'hbc71707a),
	.w3(32'hbb22761e),
	.w4(32'hbc8fa563),
	.w5(32'hbc63c08b),
	.w6(32'hbc24f9d8),
	.w7(32'hba9f70c2),
	.w8(32'h3c68859a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef69ff),
	.w1(32'hbbdc42f4),
	.w2(32'hb980249f),
	.w3(32'h3be27c3b),
	.w4(32'hbb03bae3),
	.w5(32'hba77bdd8),
	.w6(32'h3bb49919),
	.w7(32'h3bf8c8df),
	.w8(32'h3bb3862c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb207eb6),
	.w1(32'hbb8a7a63),
	.w2(32'hbb5ec05b),
	.w3(32'hbc14297d),
	.w4(32'hb85415c7),
	.w5(32'h3ac8bfa7),
	.w6(32'hbb2b4890),
	.w7(32'hbab63197),
	.w8(32'hbbc03f25),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc6cf9),
	.w1(32'h3a08f25b),
	.w2(32'h392b5ffe),
	.w3(32'hba43ae4b),
	.w4(32'h3b16639f),
	.w5(32'hbb996a2b),
	.w6(32'h3aed6e3d),
	.w7(32'h3ae57819),
	.w8(32'h3b1a0d13),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94e19c),
	.w1(32'h3a99e9b2),
	.w2(32'h3b205980),
	.w3(32'hbc458238),
	.w4(32'hbb2c81aa),
	.w5(32'hb9cb3cef),
	.w6(32'hbac3e282),
	.w7(32'hb9f386bc),
	.w8(32'hbade8957),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e7590),
	.w1(32'hbb460c7d),
	.w2(32'hbaa4eebf),
	.w3(32'hba4cbc0a),
	.w4(32'hbbaba88f),
	.w5(32'h3a8687fa),
	.w6(32'h3b44a48d),
	.w7(32'h3b5bbb0d),
	.w8(32'h3bf60148),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule