module layer_8_featuremap_148(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d23d3),
	.w1(32'hbb5c1e24),
	.w2(32'h3b0fa9a7),
	.w3(32'hbafdfd35),
	.w4(32'h3c2f2856),
	.w5(32'h3c5c5798),
	.w6(32'hbb33cbe7),
	.w7(32'h3c6ca7a8),
	.w8(32'h3c6bd55e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf38e06),
	.w1(32'hbb14b4f4),
	.w2(32'hbb421271),
	.w3(32'h3c5a3c09),
	.w4(32'hbbb64214),
	.w5(32'h3bde7086),
	.w6(32'h3ca25ad1),
	.w7(32'hbbb2c9fb),
	.w8(32'h3ba2ce7b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d80ba),
	.w1(32'h39495ba5),
	.w2(32'h3aa42884),
	.w3(32'hbafc5ab7),
	.w4(32'hbb99e603),
	.w5(32'hbc147247),
	.w6(32'hbb508a1d),
	.w7(32'hbb579279),
	.w8(32'hbb5083d0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b47a6),
	.w1(32'h3b5c1f7c),
	.w2(32'h3a465915),
	.w3(32'h3bed1ad9),
	.w4(32'h3c6f3fcf),
	.w5(32'h3bd0749e),
	.w6(32'h3ac0aeed),
	.w7(32'h3c6a9336),
	.w8(32'h3ba8541c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad282b6),
	.w1(32'h3c3104c9),
	.w2(32'hbb9aeccc),
	.w3(32'h3bd57a52),
	.w4(32'hbb2e7c21),
	.w5(32'h3bf05de5),
	.w6(32'h3c59b8df),
	.w7(32'hbb03449a),
	.w8(32'h39a10c53),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c177f),
	.w1(32'hbb1e456e),
	.w2(32'hbc1e6e3d),
	.w3(32'h3c190ccf),
	.w4(32'h3ae8270a),
	.w5(32'h3a1a9f4a),
	.w6(32'h3b7f05f4),
	.w7(32'hbb9052b8),
	.w8(32'hbad8f4e7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb01757),
	.w1(32'h3b5e806e),
	.w2(32'h3bd03efc),
	.w3(32'hbba11bd7),
	.w4(32'h3b18b1da),
	.w5(32'h3bb59e36),
	.w6(32'h3b7842ff),
	.w7(32'h3b9d9c17),
	.w8(32'hbb320602),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb89586),
	.w1(32'hbb4b676b),
	.w2(32'h3b0bdcb2),
	.w3(32'h3bac7a64),
	.w4(32'h3ab23672),
	.w5(32'hba735e31),
	.w6(32'hbb6ba71f),
	.w7(32'h3aab11b7),
	.w8(32'hbb98d34d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2f82c),
	.w1(32'hba25f6c2),
	.w2(32'hbaab9b81),
	.w3(32'h3902ce8c),
	.w4(32'h3a400af4),
	.w5(32'hbb0e6055),
	.w6(32'h3b4d5282),
	.w7(32'h3cbc95f2),
	.w8(32'h3c6e7989),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1c32f),
	.w1(32'h3a84ad2f),
	.w2(32'h3c8af871),
	.w3(32'hbaf0d311),
	.w4(32'hbb27b319),
	.w5(32'hbb81cfac),
	.w6(32'h3c9065c9),
	.w7(32'h3b7f0acc),
	.w8(32'hbc1622e5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42dd4b),
	.w1(32'hba9f05ff),
	.w2(32'hbc0d7342),
	.w3(32'hbc265e03),
	.w4(32'hbb4a04dd),
	.w5(32'hbc125640),
	.w6(32'hbcaa41a0),
	.w7(32'hbbf842a1),
	.w8(32'h398171e3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae759bc),
	.w1(32'h3bb270b2),
	.w2(32'hbad60cd7),
	.w3(32'h3bb8b8bf),
	.w4(32'h3beb9828),
	.w5(32'h3baece99),
	.w6(32'h3bca8ef4),
	.w7(32'h3b1539a8),
	.w8(32'hba6dd601),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07982e),
	.w1(32'hb9a48ba0),
	.w2(32'h38008eeb),
	.w3(32'h3b933575),
	.w4(32'hb89bd7fc),
	.w5(32'hb91dd5af),
	.w6(32'h3b20fbf4),
	.w7(32'hb9220202),
	.w8(32'hb98d8bbc),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb800c1a2),
	.w1(32'hb98e9dd6),
	.w2(32'h3a4cdb82),
	.w3(32'hb9526b90),
	.w4(32'h3a86b62f),
	.w5(32'h39ca62ce),
	.w6(32'hb9b62ae6),
	.w7(32'h3a395154),
	.w8(32'hb901b4dc),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3601556c),
	.w1(32'hb9ecb58f),
	.w2(32'h3acb0e72),
	.w3(32'hb8ef54f7),
	.w4(32'h3adb830e),
	.w5(32'h3ab5ec42),
	.w6(32'hb9f5a077),
	.w7(32'h3ac9c8a3),
	.w8(32'h3a8c1170),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92c8a7),
	.w1(32'h3a0a5866),
	.w2(32'hba96c905),
	.w3(32'h3a41804d),
	.w4(32'hba69481b),
	.w5(32'hba7ddfa1),
	.w6(32'h39ee168c),
	.w7(32'hbaa81423),
	.w8(32'hbad7942b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5772c),
	.w1(32'hbaf94089),
	.w2(32'h39c49a47),
	.w3(32'hba9589fd),
	.w4(32'h39f7146d),
	.w5(32'h39d0eb5a),
	.w6(32'hbaf7a78e),
	.w7(32'hb9073125),
	.w8(32'hb8a6c4f6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3874d),
	.w1(32'h3a6aba7b),
	.w2(32'hbaaaa0b5),
	.w3(32'h3ab639db),
	.w4(32'hbaec7a17),
	.w5(32'hbaab17ec),
	.w6(32'h3a6e9f2b),
	.w7(32'hbab122db),
	.w8(32'hbaa1b391),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6dac6),
	.w1(32'hb9f7f7a0),
	.w2(32'hba93177d),
	.w3(32'hbad86fb3),
	.w4(32'hbaf202ad),
	.w5(32'hbaac5791),
	.w6(32'hbb00e0da),
	.w7(32'hbb0ee9e0),
	.w8(32'hbacb6a85),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79d032),
	.w1(32'hba9168a1),
	.w2(32'hbac036d4),
	.w3(32'hb9c0b4df),
	.w4(32'hba7b0c19),
	.w5(32'hb9ca40de),
	.w6(32'hba16be8d),
	.w7(32'hbacb05a7),
	.w8(32'hba8fff16),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacf6cc),
	.w1(32'hbae01ce9),
	.w2(32'hba43cb56),
	.w3(32'hba597f32),
	.w4(32'hbb0bebd8),
	.w5(32'hba8385a4),
	.w6(32'hbab8f4e7),
	.w7(32'hba909902),
	.w8(32'hb8984662),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba952c0e),
	.w1(32'hba9e8446),
	.w2(32'hb9ef7e0f),
	.w3(32'hba8e10f9),
	.w4(32'hba32cc11),
	.w5(32'hba49d4f5),
	.w6(32'hba8d1d34),
	.w7(32'hba77d06d),
	.w8(32'hba7792e4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60c858),
	.w1(32'hba7baae7),
	.w2(32'h3b0070ce),
	.w3(32'hbaa6120d),
	.w4(32'h3ab16df1),
	.w5(32'h3a93e306),
	.w6(32'hbaf19e80),
	.w7(32'h3868ec6d),
	.w8(32'hb9dcc714),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fd7a9),
	.w1(32'h3b11cb09),
	.w2(32'hba7eb3e1),
	.w3(32'h3b1e5e2c),
	.w4(32'hba7b2c9a),
	.w5(32'hba24454f),
	.w6(32'h3ab918a3),
	.w7(32'hba99a822),
	.w8(32'hba56e667),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c3463),
	.w1(32'hba1ea8bd),
	.w2(32'h3a194115),
	.w3(32'hb9f88a9b),
	.w4(32'h3890ee52),
	.w5(32'h38837928),
	.w6(32'hba497a68),
	.w7(32'h399fa724),
	.w8(32'hb81de023),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391a393b),
	.w1(32'hb956d2ca),
	.w2(32'h39a93a36),
	.w3(32'hb9e1bf9b),
	.w4(32'h3a93e916),
	.w5(32'h3a58b4af),
	.w6(32'hba05da7e),
	.w7(32'h3a645f4c),
	.w8(32'h3a6d75d1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c23713),
	.w1(32'h37962df5),
	.w2(32'hbacbc2a6),
	.w3(32'h3aa6dafb),
	.w4(32'hb9e2fca9),
	.w5(32'hba84ddea),
	.w6(32'h3a9095d7),
	.w7(32'hbaa31d73),
	.w8(32'hbae3933f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e0f31),
	.w1(32'hbb77242c),
	.w2(32'h3b1bea49),
	.w3(32'hbb8693ed),
	.w4(32'hbb517bae),
	.w5(32'h3a8ee1a2),
	.w6(32'hbba1b56d),
	.w7(32'hbb48c540),
	.w8(32'h39f57f60),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add763f),
	.w1(32'h3ada198d),
	.w2(32'h3a027e2a),
	.w3(32'h3aa8610e),
	.w4(32'h3a45f02c),
	.w5(32'h399cee4f),
	.w6(32'h3a979ee4),
	.w7(32'h395bef51),
	.w8(32'hb97e2f11),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991dd9c),
	.w1(32'h3a594d32),
	.w2(32'hbadde3a0),
	.w3(32'h3a6d3344),
	.w4(32'hba6d82da),
	.w5(32'hb8dc3ef3),
	.w6(32'h39dfb56f),
	.w7(32'hba850654),
	.w8(32'hb8cd15be),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41ee70),
	.w1(32'hba9077e2),
	.w2(32'h39cb1eb7),
	.w3(32'hba202314),
	.w4(32'h3a0d7ee5),
	.w5(32'h3968f1c5),
	.w6(32'hb80f1841),
	.w7(32'h399b00a6),
	.w8(32'hb88d2f2d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940f7f5),
	.w1(32'h3906ea09),
	.w2(32'hba1ff22a),
	.w3(32'h397d1e42),
	.w4(32'hbaabeccc),
	.w5(32'hbaa73191),
	.w6(32'h382c10b0),
	.w7(32'hba727447),
	.w8(32'hba64396d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b259b),
	.w1(32'hb9d83688),
	.w2(32'h3a4c4a9b),
	.w3(32'hbaa57dc8),
	.w4(32'h3aa526ff),
	.w5(32'h3aa1c438),
	.w6(32'hba545a1f),
	.w7(32'h3a9bc322),
	.w8(32'h3ab49a30),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab41eb0),
	.w1(32'h3a6618e1),
	.w2(32'h3a676caa),
	.w3(32'h3aadd0e5),
	.w4(32'hb6ae3fd4),
	.w5(32'h398f53b5),
	.w6(32'h3ab50f8c),
	.w7(32'h38bf4e47),
	.w8(32'h391a3000),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a565fd8),
	.w1(32'h3a75a36a),
	.w2(32'hbab79882),
	.w3(32'h3a0f2c52),
	.w4(32'hba41f094),
	.w5(32'hba450c98),
	.w6(32'h39f2387b),
	.w7(32'hba7264bb),
	.w8(32'hba7c9082),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca6629),
	.w1(32'hbae2a0d6),
	.w2(32'h3a26ffd9),
	.w3(32'hba7c3e84),
	.w4(32'hb95f296a),
	.w5(32'hb9589fd8),
	.w6(32'hbac9bbb4),
	.w7(32'hba0eaad3),
	.w8(32'hb9d8698c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26a6f3),
	.w1(32'h3a8e3ee8),
	.w2(32'h3a96a58e),
	.w3(32'h38f604b6),
	.w4(32'h3ade6088),
	.w5(32'h3ab85fc8),
	.w6(32'h39d69f0d),
	.w7(32'h3ab7c844),
	.w8(32'h3a736314),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a684fe3),
	.w1(32'h3ab78661),
	.w2(32'h39cf087c),
	.w3(32'h3ac2eae7),
	.w4(32'h39d125f2),
	.w5(32'hb981d07f),
	.w6(32'h3ab2a8b9),
	.w7(32'h388fbf44),
	.w8(32'hba2a8c30),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d34737),
	.w1(32'h37b537b5),
	.w2(32'hbae30b20),
	.w3(32'hb96ecdef),
	.w4(32'hbad9c675),
	.w5(32'hba857f7f),
	.w6(32'hba02071a),
	.w7(32'hbae17629),
	.w8(32'hbacc18b4),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6a0bb),
	.w1(32'hba88e43d),
	.w2(32'h392c4398),
	.w3(32'hba45a7af),
	.w4(32'h39c3544d),
	.w5(32'h39ab572d),
	.w6(32'hba9775dd),
	.w7(32'hb779a452),
	.w8(32'hb91431b5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02ed3b),
	.w1(32'hb98214c4),
	.w2(32'hb9676c62),
	.w3(32'hb8847116),
	.w4(32'h399d4fa5),
	.w5(32'h3a5490c1),
	.w6(32'hba3f3401),
	.w7(32'hba31f753),
	.w8(32'hb81737ec),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d885f),
	.w1(32'hbabff352),
	.w2(32'hba356cbd),
	.w3(32'h394d2178),
	.w4(32'hba54b767),
	.w5(32'hba1cc8a6),
	.w6(32'hba50e32b),
	.w7(32'hba858b7d),
	.w8(32'hba87d1d0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06e52b),
	.w1(32'hb8dee65a),
	.w2(32'hba5d4d98),
	.w3(32'h39decbef),
	.w4(32'hba8844c6),
	.w5(32'hbae3674e),
	.w6(32'hb8ef78e0),
	.w7(32'hbab26c1c),
	.w8(32'hbaff185f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72cd4c),
	.w1(32'hba89e525),
	.w2(32'h38e34b42),
	.w3(32'hbabe2f7a),
	.w4(32'h390ec713),
	.w5(32'h390d7f61),
	.w6(32'hbaf79e03),
	.w7(32'hb76e50b1),
	.w8(32'hb92347a7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1eb82),
	.w1(32'hba0ee0ba),
	.w2(32'h39d8328e),
	.w3(32'hb9ba92d0),
	.w4(32'h38d3c699),
	.w5(32'hb99d780b),
	.w6(32'hba4410d6),
	.w7(32'hb9c53dc7),
	.w8(32'hba90f093),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd3cae),
	.w1(32'hb9f96545),
	.w2(32'hb9eafeab),
	.w3(32'h39bd285d),
	.w4(32'hba64c6e9),
	.w5(32'hb98611dd),
	.w6(32'hba360044),
	.w7(32'hba865da1),
	.w8(32'h39e7d772),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba36fc),
	.w1(32'h3aa8defd),
	.w2(32'h3956f44b),
	.w3(32'h3a19bc69),
	.w4(32'h38eca769),
	.w5(32'hb9b27231),
	.w6(32'h3ac442a1),
	.w7(32'hb9026c8e),
	.w8(32'hb9686873),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951749a),
	.w1(32'hb99ba440),
	.w2(32'h3a52d3d6),
	.w3(32'hba645efc),
	.w4(32'h38963e84),
	.w5(32'h38d06c2f),
	.w6(32'hba95b3b1),
	.w7(32'hb94f4f61),
	.w8(32'hba6b7261),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a88a83),
	.w1(32'hb97827ff),
	.w2(32'hbaeb4fbe),
	.w3(32'h3a650094),
	.w4(32'hbb2f63bd),
	.w5(32'hbafa965c),
	.w6(32'hb9bc69ee),
	.w7(32'hbaf67c11),
	.w8(32'hbac84a82),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab32ace),
	.w1(32'hba9555cd),
	.w2(32'h39e40c45),
	.w3(32'hbad42b4b),
	.w4(32'hb9485a85),
	.w5(32'hba4e1895),
	.w6(32'hba9d96fc),
	.w7(32'hba1cc114),
	.w8(32'hbabdcb50),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99965e4),
	.w1(32'h3a803396),
	.w2(32'h3a3e63a3),
	.w3(32'h392327b3),
	.w4(32'h39fbc444),
	.w5(32'h3a89353f),
	.w6(32'hb9564696),
	.w7(32'h3a1bed61),
	.w8(32'h3aae5527),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fb3c4),
	.w1(32'h3a5ba03d),
	.w2(32'h3aa2fd5c),
	.w3(32'h3a29176c),
	.w4(32'h380ea5e2),
	.w5(32'hb9bfe304),
	.w6(32'h3a25c13d),
	.w7(32'h384f3bf4),
	.w8(32'hb9977a1b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5156ca),
	.w1(32'h3a080aa1),
	.w2(32'hbab9e9ef),
	.w3(32'h3a1926f9),
	.w4(32'hbb05857c),
	.w5(32'hbb119558),
	.w6(32'h3930498d),
	.w7(32'hbaf02630),
	.w8(32'hbb15584e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec1250),
	.w1(32'hba8d1cb9),
	.w2(32'h362d9423),
	.w3(32'hbae90805),
	.w4(32'h39cfd0ad),
	.w5(32'hb9419872),
	.w6(32'hbaea957e),
	.w7(32'h38cb3a53),
	.w8(32'hba16e037),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9040a),
	.w1(32'hba1f184a),
	.w2(32'hbaa46672),
	.w3(32'hb985d738),
	.w4(32'hbacc2670),
	.w5(32'hbaefbcb4),
	.w6(32'hba1534d6),
	.w7(32'hbacc1523),
	.w8(32'hbac28254),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82204b),
	.w1(32'hba90a251),
	.w2(32'hbab2a1dc),
	.w3(32'hbb0b75b4),
	.w4(32'hbb0adfec),
	.w5(32'hbaa3f131),
	.w6(32'hbae6c770),
	.w7(32'hbaeb7116),
	.w8(32'hba5de8b4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1762ed),
	.w1(32'hba9c91df),
	.w2(32'h39918ab7),
	.w3(32'hbad3cdf8),
	.w4(32'h3a19cbed),
	.w5(32'hb58d0e90),
	.w6(32'hbaa9facc),
	.w7(32'h39821a0e),
	.w8(32'hba0690ab),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f726f),
	.w1(32'hba476663),
	.w2(32'h39d5d37d),
	.w3(32'hb9c17d4c),
	.w4(32'h39f0777f),
	.w5(32'h3a38beef),
	.w6(32'hbaa7bcf2),
	.w7(32'hba4386a9),
	.w8(32'hba596a0c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ebf15),
	.w1(32'h39b8c977),
	.w2(32'h37023102),
	.w3(32'h39bc4fdc),
	.w4(32'h3829aded),
	.w5(32'hb93792f9),
	.w6(32'hba577b5f),
	.w7(32'hb9b6215d),
	.w8(32'hba221f3b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab9a72),
	.w1(32'hba0c469a),
	.w2(32'hba81f272),
	.w3(32'hb917028b),
	.w4(32'hbae16830),
	.w5(32'hba589fa3),
	.w6(32'hb9fc1627),
	.w7(32'hb938cf17),
	.w8(32'h3a53e179),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3955a3ce),
	.w1(32'hba9cbc81),
	.w2(32'h39d8254a),
	.w3(32'hbb011b6c),
	.w4(32'hb92897d6),
	.w5(32'hb9c91764),
	.w6(32'hb9aa4c30),
	.w7(32'hb9885874),
	.w8(32'hb9f12dc5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7580a),
	.w1(32'h38cdca34),
	.w2(32'hb813a02f),
	.w3(32'h399f8491),
	.w4(32'hb99b1cf1),
	.w5(32'hba354ee0),
	.w6(32'hb7bc3539),
	.w7(32'hb9007fb0),
	.w8(32'hb9d0d88d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9a666),
	.w1(32'hba0e0694),
	.w2(32'hb99f9206),
	.w3(32'hba56b9f8),
	.w4(32'hba140b71),
	.w5(32'hba7fe5c3),
	.w6(32'hba555cbe),
	.w7(32'hba16ab6d),
	.w8(32'hba544e91),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e63e4),
	.w1(32'hbaaa7b5e),
	.w2(32'hba5b555c),
	.w3(32'hbad134cf),
	.w4(32'hba8e88ae),
	.w5(32'hba46d2e9),
	.w6(32'hbaace4f4),
	.w7(32'hbab364da),
	.w8(32'hbaa926e7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54d14e),
	.w1(32'hba695e7d),
	.w2(32'h3a85b593),
	.w3(32'hba40e9c8),
	.w4(32'h36c9a5ce),
	.w5(32'hba64c9d0),
	.w6(32'hba892b0d),
	.w7(32'hb8bb3d5f),
	.w8(32'hba80ea74),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9386c13),
	.w1(32'hb9933e31),
	.w2(32'hba9518f9),
	.w3(32'hba5c6372),
	.w4(32'hba9fa588),
	.w5(32'hbabfa9ce),
	.w6(32'hba5c5644),
	.w7(32'hbae036e8),
	.w8(32'hbaface60),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcc367),
	.w1(32'hba8a5776),
	.w2(32'hbb0a5bc7),
	.w3(32'hba4e73b3),
	.w4(32'hba882ce1),
	.w5(32'hb9e1686a),
	.w6(32'hba9f2f78),
	.w7(32'hba8d2ef5),
	.w8(32'hba155e8a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6a147),
	.w1(32'hba4997d6),
	.w2(32'hb8334ee4),
	.w3(32'hb99573dd),
	.w4(32'h39cfa308),
	.w5(32'hb86bcfd0),
	.w6(32'hb9637632),
	.w7(32'h3901e618),
	.w8(32'hba7824d4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba779649),
	.w1(32'h37538319),
	.w2(32'hba7d524f),
	.w3(32'h3a26898b),
	.w4(32'hba606a3d),
	.w5(32'hbaa32e1a),
	.w6(32'hb9b11fc4),
	.w7(32'hbaab7708),
	.w8(32'hbaf2ee8b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ccb04),
	.w1(32'hba185daa),
	.w2(32'h3a8deaac),
	.w3(32'hbac796ec),
	.w4(32'hb76f54be),
	.w5(32'h386e2727),
	.w6(32'hbb0f862b),
	.w7(32'hb9f8a34a),
	.w8(32'hba96782f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8a0fa),
	.w1(32'h3a5b01bd),
	.w2(32'h3abe0c29),
	.w3(32'hb7bbf86e),
	.w4(32'h3b122ad9),
	.w5(32'h3a454c7f),
	.w6(32'hb9be3846),
	.w7(32'h3a6711a6),
	.w8(32'hba071bf8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a424f5c),
	.w1(32'h3b1d5aa3),
	.w2(32'hba760fca),
	.w3(32'h3ad4c5d3),
	.w4(32'hbab0772b),
	.w5(32'hba09f3a2),
	.w6(32'h3a507cef),
	.w7(32'hbaaf2a5a),
	.w8(32'hba713f6c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7696c5),
	.w1(32'hbb0b566a),
	.w2(32'h394cb249),
	.w3(32'hbabb3d91),
	.w4(32'hb8c3a6f6),
	.w5(32'hba05c1db),
	.w6(32'hbacabdf4),
	.w7(32'hb97f52d1),
	.w8(32'hba2ef374),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b63bff),
	.w1(32'h39c493c5),
	.w2(32'h38739361),
	.w3(32'hb8ac2a55),
	.w4(32'h394392bf),
	.w5(32'h399cfc88),
	.w6(32'hb93d6e26),
	.w7(32'hb7fc3be3),
	.w8(32'hb92f86bb),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972c6ce),
	.w1(32'hb9a1de76),
	.w2(32'hba9cac84),
	.w3(32'hb9239446),
	.w4(32'hbb004c26),
	.w5(32'hba8153db),
	.w6(32'hb99216e7),
	.w7(32'hbacca9ea),
	.w8(32'hba250003),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940f068),
	.w1(32'hb91c26a9),
	.w2(32'hba6a55c1),
	.w3(32'hba9307fe),
	.w4(32'hba91c468),
	.w5(32'hba857a65),
	.w6(32'hba042be7),
	.w7(32'hba8656f4),
	.w8(32'hba88e644),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dc6a9),
	.w1(32'hb9ec178c),
	.w2(32'hb63fc7fe),
	.w3(32'hba3b36e2),
	.w4(32'h36cbe5de),
	.w5(32'h3701312f),
	.w6(32'hba1f3991),
	.w7(32'h3742484b),
	.w8(32'h374c2da1),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f79689),
	.w1(32'hb8df3ec1),
	.w2(32'hb8b580fc),
	.w3(32'hb95c0880),
	.w4(32'hb95ba777),
	.w5(32'hb8ce9aae),
	.w6(32'hb967f2bf),
	.w7(32'hb9330c16),
	.w8(32'hb8a61669),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cd45fc),
	.w1(32'hb7aa7bdc),
	.w2(32'hb89335c7),
	.w3(32'hb802df65),
	.w4(32'hb66c8c7c),
	.w5(32'hb744a4f9),
	.w6(32'hb8aae272),
	.w7(32'hb8849222),
	.w8(32'hb88840c3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bbfa80),
	.w1(32'h36f2e853),
	.w2(32'h37e8cb0c),
	.w3(32'h376e497e),
	.w4(32'hb7442dd5),
	.w5(32'hb5d5e1f6),
	.w6(32'hb6cc7773),
	.w7(32'hb7ce964d),
	.w8(32'hb5350470),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cc87df),
	.w1(32'hb700a27b),
	.w2(32'hb37f8901),
	.w3(32'hb7b30c04),
	.w4(32'hb7843f38),
	.w5(32'hb68430da),
	.w6(32'hb6669a99),
	.w7(32'hb6ec06c3),
	.w8(32'h3458a96b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ac2bc4),
	.w1(32'h374f0cc3),
	.w2(32'h3845e441),
	.w3(32'h383ed546),
	.w4(32'h3851424d),
	.w5(32'h37ec40e8),
	.w6(32'hb81d4135),
	.w7(32'hb89117ec),
	.w8(32'hb8e40715),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9302c87),
	.w1(32'hb945e07d),
	.w2(32'hb90b8c63),
	.w3(32'hb8e51c55),
	.w4(32'hb92f390a),
	.w5(32'hb7d322a1),
	.w6(32'hb957f2b8),
	.w7(32'hb94f03b0),
	.w8(32'hb854de92),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba380abe),
	.w1(32'hba171ccd),
	.w2(32'hb9de50f9),
	.w3(32'hba4b49d5),
	.w4(32'hba150661),
	.w5(32'hb840b8cb),
	.w6(32'hba560afb),
	.w7(32'hba323e7c),
	.w8(32'hb8ff6767),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba831a),
	.w1(32'hb98ff84f),
	.w2(32'hb90aef07),
	.w3(32'hb9e7bc37),
	.w4(32'hb9f1038d),
	.w5(32'hb7a93529),
	.w6(32'hba229454),
	.w7(32'hba14913b),
	.w8(32'hb93e9b06),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b800d),
	.w1(32'hb990d49c),
	.w2(32'hb911baff),
	.w3(32'hb9599d67),
	.w4(32'hb9aa5027),
	.w5(32'hb8464569),
	.w6(32'hb94c29c0),
	.w7(32'hb9950c48),
	.w8(32'h38430d99),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb720fe8d),
	.w1(32'hb690bb47),
	.w2(32'h35d04c19),
	.w3(32'h37435a94),
	.w4(32'hb6992160),
	.w5(32'hb6c785c5),
	.w6(32'hb3f3d672),
	.w7(32'h35631dbd),
	.w8(32'hb54b58d5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3f682e1),
	.w1(32'h36c9c4cf),
	.w2(32'hb6f4f76f),
	.w3(32'h35eada19),
	.w4(32'h35369472),
	.w5(32'h36298952),
	.w6(32'h35405355),
	.w7(32'hb63782b0),
	.w8(32'h3615d023),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3712c261),
	.w1(32'h362d1506),
	.w2(32'hb5189f0f),
	.w3(32'h36eecaaa),
	.w4(32'h36b34e3e),
	.w5(32'h366044b1),
	.w6(32'h379d34f8),
	.w7(32'h3807bcd7),
	.w8(32'h37da3483),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3604bbbe),
	.w1(32'hb72665fc),
	.w2(32'hb7cc7192),
	.w3(32'hb76b4e23),
	.w4(32'hb7d2bf61),
	.w5(32'hb7b1f1dc),
	.w6(32'h370bccda),
	.w7(32'h36fb5b71),
	.w8(32'hb7c56278),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35625e60),
	.w1(32'hb763208a),
	.w2(32'hb83e2004),
	.w3(32'h382b93cf),
	.w4(32'h3759394d),
	.w5(32'hb789551c),
	.w6(32'h373d9c20),
	.w7(32'h37fd5525),
	.w8(32'h3805d514),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38021da1),
	.w1(32'h36f24dda),
	.w2(32'h37d3e59f),
	.w3(32'h37a501d9),
	.w4(32'hb39ef6a6),
	.w5(32'h37877fa0),
	.w6(32'h36a93813),
	.w7(32'h360c7d37),
	.w8(32'h37294be9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379f94e5),
	.w1(32'h37c69408),
	.w2(32'h38164a78),
	.w3(32'h38826a78),
	.w4(32'h3842fb55),
	.w5(32'h38c7bc44),
	.w6(32'hb565353c),
	.w7(32'hb76e04a8),
	.w8(32'hb662e607),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb831cd9d),
	.w1(32'hb8c52546),
	.w2(32'hb8ade64e),
	.w3(32'hb8238402),
	.w4(32'hb75110df),
	.w5(32'h35dec83d),
	.w6(32'hb7b8a613),
	.w7(32'hb7f6cb5c),
	.w8(32'h383364e4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8479048),
	.w1(32'hb8131bfd),
	.w2(32'hb807ad4b),
	.w3(32'h37b9a511),
	.w4(32'h3822b0c2),
	.w5(32'hb7b5696f),
	.w6(32'hb3f32b24),
	.w7(32'h37c74da6),
	.w8(32'h36fe150c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb836065b),
	.w1(32'hb8950f72),
	.w2(32'hb89e2f08),
	.w3(32'hb873e1df),
	.w4(32'hb88e2ed9),
	.w5(32'hb8c20188),
	.w6(32'h36ce82cc),
	.w7(32'h3646906b),
	.w8(32'hb889ba50),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb51afa93),
	.w1(32'h36ecbcff),
	.w2(32'hb85bf9b3),
	.w3(32'h377a9eaa),
	.w4(32'h38c383a9),
	.w5(32'h375a6db3),
	.w6(32'h37ead46f),
	.w7(32'h38d04902),
	.w8(32'h38a6b0de),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h359e8fd6),
	.w1(32'h36144880),
	.w2(32'h36cf4443),
	.w3(32'h3756af46),
	.w4(32'hb745fe92),
	.w5(32'hb72e90a8),
	.w6(32'h37569dea),
	.w7(32'hb650e4b6),
	.w8(32'hb5ec9711),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d6db2a),
	.w1(32'h372b280d),
	.w2(32'hb6458d45),
	.w3(32'hb4acd88d),
	.w4(32'h36a972c8),
	.w5(32'h369a1a10),
	.w6(32'h36de4691),
	.w7(32'h3636fe33),
	.w8(32'h371259b7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c96f62),
	.w1(32'h3616857f),
	.w2(32'h3512da0a),
	.w3(32'hb605ac2b),
	.w4(32'hb6d1841a),
	.w5(32'hb592f62f),
	.w6(32'h36243022),
	.w7(32'hb5c58898),
	.w8(32'h358f21d2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3501e124),
	.w1(32'h374e9712),
	.w2(32'h36c292cf),
	.w3(32'hb6142168),
	.w4(32'hb61d1d1e),
	.w5(32'h37122be7),
	.w6(32'hb62a2c27),
	.w7(32'hb70802d2),
	.w8(32'h36897803),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81414a4),
	.w1(32'hb6a63f14),
	.w2(32'h372bf0f1),
	.w3(32'hb84795ba),
	.w4(32'hb7b3b845),
	.w5(32'hb7d0acf2),
	.w6(32'hb800a2d7),
	.w7(32'hb6eb20eb),
	.w8(32'hb825be4f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3835627b),
	.w1(32'h36d25d92),
	.w2(32'h369a1143),
	.w3(32'hb6cd79e2),
	.w4(32'hb7dcd9d4),
	.w5(32'hb6456420),
	.w6(32'h382b85c9),
	.w7(32'h38705e6c),
	.w8(32'h38e03320),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bcf2c2),
	.w1(32'hb885c9fd),
	.w2(32'h36d44844),
	.w3(32'hb829af60),
	.w4(32'h385d83ec),
	.w5(32'h389fb23a),
	.w6(32'hb8ec480c),
	.w7(32'hb8313bd0),
	.w8(32'hb8462486),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74091aa),
	.w1(32'hb79de586),
	.w2(32'hb526a98d),
	.w3(32'h377e4bdd),
	.w4(32'h37e22f23),
	.w5(32'h36c7deee),
	.w6(32'h36a8319b),
	.w7(32'h371ea472),
	.w8(32'hb7510d0a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8479c25),
	.w1(32'hb8a1f6c7),
	.w2(32'h38aa1d86),
	.w3(32'hb8effb88),
	.w4(32'hb9797932),
	.w5(32'h392c2a62),
	.w6(32'hb9ae70a6),
	.w7(32'hb980694a),
	.w8(32'h37970277),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3827a452),
	.w1(32'h3838111a),
	.w2(32'h37ecb2a1),
	.w3(32'h386c0420),
	.w4(32'h377f704e),
	.w5(32'hb7b953e2),
	.w6(32'h37c28e55),
	.w7(32'hb86e9a9d),
	.w8(32'hb804d28f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38006dc9),
	.w1(32'hb76a7d92),
	.w2(32'hb7ecbc3d),
	.w3(32'hb734602b),
	.w4(32'h38ac41a9),
	.w5(32'h36f09489),
	.w6(32'hb7609a28),
	.w7(32'h372e7bd0),
	.w8(32'hb8120ce9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a20c27),
	.w1(32'hb83fe853),
	.w2(32'hb839dccb),
	.w3(32'h377f5c60),
	.w4(32'h37a24737),
	.w5(32'hb7c036ba),
	.w6(32'h364b69e7),
	.w7(32'hb8008764),
	.w8(32'hb8853e02),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380c64f6),
	.w1(32'h38b99e31),
	.w2(32'hb8790364),
	.w3(32'hb85b4e3e),
	.w4(32'h38805529),
	.w5(32'hb8d3ddf9),
	.w6(32'hb8c05297),
	.w7(32'h389470dc),
	.w8(32'h381d5961),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f30975),
	.w1(32'hb91bed09),
	.w2(32'hb8ab08e5),
	.w3(32'hb92fc510),
	.w4(32'hb92b4448),
	.w5(32'hb93ae523),
	.w6(32'hb98c5d3f),
	.w7(32'hb93d926c),
	.w8(32'hb950eb6b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f2cbd8),
	.w1(32'hb8d1f0f6),
	.w2(32'hb7fe7acb),
	.w3(32'hb8b7ef1c),
	.w4(32'hb8a1b7a4),
	.w5(32'hb78f7d7d),
	.w6(32'hb90d4049),
	.w7(32'hb8faffbb),
	.w8(32'hb85d83af),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79572dc),
	.w1(32'h3731674f),
	.w2(32'hb7dcb3e0),
	.w3(32'h377d0b16),
	.w4(32'h37d020b6),
	.w5(32'hb7785fef),
	.w6(32'h3787288e),
	.w7(32'h3810c447),
	.w8(32'hb805e30c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72a798c),
	.w1(32'h36c70832),
	.w2(32'hb4d02b32),
	.w3(32'hb4e8524d),
	.w4(32'h3650d94e),
	.w5(32'hb619a322),
	.w6(32'hb7c33851),
	.w7(32'h370291e1),
	.w8(32'h36cef4dc),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3701e928),
	.w1(32'h371ba2f4),
	.w2(32'hb7a1aaaf),
	.w3(32'hb5e3b88b),
	.w4(32'hb697ee04),
	.w5(32'hb77c4f52),
	.w6(32'h375bb384),
	.w7(32'h371bb826),
	.w8(32'hb7cd5386),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378b0d5b),
	.w1(32'h3725be09),
	.w2(32'hb6458511),
	.w3(32'h37fe6671),
	.w4(32'hb53dc7ab),
	.w5(32'h377c1a77),
	.w6(32'hb6fe2eac),
	.w7(32'hb755b99c),
	.w8(32'hb67078e2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb802fda3),
	.w1(32'hb82439af),
	.w2(32'hb82da6ac),
	.w3(32'hb738dbe4),
	.w4(32'h37e31b8b),
	.w5(32'hb895af35),
	.w6(32'hb8a44db3),
	.w7(32'hb7d7cbfe),
	.w8(32'hb8a441bf),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8407efd),
	.w1(32'hb8f27431),
	.w2(32'hb890111b),
	.w3(32'hb7841d58),
	.w4(32'hb86210b1),
	.w5(32'hb7107680),
	.w6(32'hb85bd8d1),
	.w7(32'hb87353b3),
	.w8(32'hb5d7cf02),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h357ca192),
	.w1(32'hb4913ca1),
	.w2(32'hb6d48054),
	.w3(32'hb5d62910),
	.w4(32'h3699b9c8),
	.w5(32'hb5f05e2d),
	.w6(32'h3568506d),
	.w7(32'h3587865d),
	.w8(32'h36ec7fd3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ffdb56),
	.w1(32'hb69fba80),
	.w2(32'hb781c3e8),
	.w3(32'hb73707d5),
	.w4(32'h364bc037),
	.w5(32'hb7c2e588),
	.w6(32'hb789363c),
	.w7(32'h36ba9936),
	.w8(32'hb77eac51),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59856f0),
	.w1(32'hb7bdd0d6),
	.w2(32'hb8178502),
	.w3(32'h37d4a99e),
	.w4(32'hb6bcd22e),
	.w5(32'hb79c6e09),
	.w6(32'hb69dd605),
	.w7(32'hb84ba7ec),
	.w8(32'hb82f1a5c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e3d2c),
	.w1(32'hb9801b97),
	.w2(32'hb9002599),
	.w3(32'hb9b9aa0c),
	.w4(32'hb98a0534),
	.w5(32'hb90ac8e8),
	.w6(32'hb9ed075a),
	.w7(32'hb968fe74),
	.w8(32'hb68da408),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371cfb21),
	.w1(32'h3750c057),
	.w2(32'hb602042d),
	.w3(32'hb711bdd6),
	.w4(32'hb68bc2bb),
	.w5(32'hb71e398d),
	.w6(32'hb4aa425e),
	.w7(32'hb6c39358),
	.w8(32'h3702c94a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363d0557),
	.w1(32'h368c873c),
	.w2(32'h36824203),
	.w3(32'hb7b68159),
	.w4(32'hb8005a81),
	.w5(32'hb183b42e),
	.w6(32'hb7c378e8),
	.w7(32'hb79e9d65),
	.w8(32'hb8247e39),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38174b1f),
	.w1(32'h37c6ccfd),
	.w2(32'hb5fa9be2),
	.w3(32'h3668514e),
	.w4(32'h378ff948),
	.w5(32'h36cc51c4),
	.w6(32'h377a3aea),
	.w7(32'h37959f6c),
	.w8(32'hb72ca832),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d86df0),
	.w1(32'hb795ba1c),
	.w2(32'h385c9b98),
	.w3(32'h3699038c),
	.w4(32'hb7e63895),
	.w5(32'hb70c270f),
	.w6(32'h378e4147),
	.w7(32'hb7ccfa9b),
	.w8(32'h36afe0ec),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7621f6c),
	.w1(32'h36f1ddf9),
	.w2(32'hb729352e),
	.w3(32'hb8481d86),
	.w4(32'hb7d6384a),
	.w5(32'hb8a9b22f),
	.w6(32'hb8cc2289),
	.w7(32'hb855a75f),
	.w8(32'hb89e2801),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9667abf),
	.w1(32'hb907ddc3),
	.w2(32'hb8b96ec6),
	.w3(32'hb97137ec),
	.w4(32'hb9808f08),
	.w5(32'hb9297bd9),
	.w6(32'hb9a46459),
	.w7(32'hb9a59a9e),
	.w8(32'hb996f726),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule