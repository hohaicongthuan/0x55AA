module layer_6_featuremap_103(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21a258),
	.w1(32'hbadbcde9),
	.w2(32'h3b7e3392),
	.w3(32'hbb0ecb43),
	.w4(32'h3a25e249),
	.w5(32'hbb16f7c2),
	.w6(32'hbbf8c857),
	.w7(32'hbc28cd73),
	.w8(32'hbba6c50c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a324ef2),
	.w1(32'h3bd191fe),
	.w2(32'h3c3b5084),
	.w3(32'hbbd1ae44),
	.w4(32'hbbea3096),
	.w5(32'hbbe6a892),
	.w6(32'hbc90825c),
	.w7(32'hbbe21e17),
	.w8(32'hbc247028),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c816296),
	.w1(32'hbb0e182f),
	.w2(32'h3ab129d9),
	.w3(32'h3ba7708d),
	.w4(32'hbc274953),
	.w5(32'hba414c06),
	.w6(32'hbb4c4112),
	.w7(32'hbb910dba),
	.w8(32'hbbe03bd0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c812fc6),
	.w1(32'h386c5558),
	.w2(32'hbbd374a9),
	.w3(32'h3bcc107b),
	.w4(32'h3b307ab4),
	.w5(32'h3b4f5991),
	.w6(32'h3af40e19),
	.w7(32'h3a465b5b),
	.w8(32'hbb4332ac),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24e1ca),
	.w1(32'h3d4c91c6),
	.w2(32'h3da9b934),
	.w3(32'h3d04eafe),
	.w4(32'h3d6a8fd8),
	.w5(32'h3d349451),
	.w6(32'hbdb59db1),
	.w7(32'hbe1339be),
	.w8(32'hbdd0f8c8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4fccb7),
	.w1(32'h3a457348),
	.w2(32'h3b49ae72),
	.w3(32'h392fe36f),
	.w4(32'hb9e1cfe6),
	.w5(32'hbaf1bbdf),
	.w6(32'hbb8075fa),
	.w7(32'hbc01ac52),
	.w8(32'hbb970718),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ea396),
	.w1(32'hbbb83100),
	.w2(32'hbc3b595e),
	.w3(32'h3b9b4956),
	.w4(32'h3a87a146),
	.w5(32'hba3d5c84),
	.w6(32'h3c4fbdb9),
	.w7(32'h3c31eba3),
	.w8(32'h3bcead7e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde923f),
	.w1(32'hbc3c7fc0),
	.w2(32'hbb73eb67),
	.w3(32'hbc201262),
	.w4(32'hbc291bc4),
	.w5(32'hbcd4b501),
	.w6(32'h3c7cbf56),
	.w7(32'h3c88ba93),
	.w8(32'h3cfb0136),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3ea7b),
	.w1(32'h3a6072fe),
	.w2(32'hbcb96d52),
	.w3(32'h3c8d55f9),
	.w4(32'hba075123),
	.w5(32'hbb9d8d4e),
	.w6(32'h3bae2d00),
	.w7(32'h3c5ca747),
	.w8(32'h3ca2f434),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78af11),
	.w1(32'h3b28f319),
	.w2(32'h3bb3b678),
	.w3(32'h3b874d0b),
	.w4(32'h3aeeaa11),
	.w5(32'h3b4b369b),
	.w6(32'h39d41876),
	.w7(32'hba95378a),
	.w8(32'h3b01ecdd),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f5726),
	.w1(32'h3c96e626),
	.w2(32'h3be51a65),
	.w3(32'h3c86644d),
	.w4(32'h3c110b08),
	.w5(32'h3c253f11),
	.w6(32'h3c75ba6a),
	.w7(32'h3b783084),
	.w8(32'h3c654a58),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc76704),
	.w1(32'h3b2bdc89),
	.w2(32'h3ba19316),
	.w3(32'h3b0a9f35),
	.w4(32'h3bdc14be),
	.w5(32'hbb476a0b),
	.w6(32'h3b9f01d2),
	.w7(32'h3c3f5036),
	.w8(32'h3c637e2f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3664d6),
	.w1(32'hba0bb2f1),
	.w2(32'h3b5bf7c8),
	.w3(32'hba4bf73d),
	.w4(32'h39221b00),
	.w5(32'hba26e292),
	.w6(32'hbbfe1e14),
	.w7(32'hbb6d6937),
	.w8(32'hbbb350a8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c422e1c),
	.w1(32'h3c83c42b),
	.w2(32'h3d223e7a),
	.w3(32'h3c3654b1),
	.w4(32'h3c6ae97f),
	.w5(32'hbb37a96e),
	.w6(32'hbc94ef6d),
	.w7(32'hbce629ac),
	.w8(32'hbd2af6d3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccbf21b),
	.w1(32'h3ac7d5e6),
	.w2(32'hba9b4f7e),
	.w3(32'h3befe8f6),
	.w4(32'hb926b0f5),
	.w5(32'hbac6d84e),
	.w6(32'h3b2d688e),
	.w7(32'hbb3e384c),
	.w8(32'hbb384427),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36f6fb),
	.w1(32'h3a7844fc),
	.w2(32'hbb23aac1),
	.w3(32'h3b199c46),
	.w4(32'hba896fc4),
	.w5(32'hbb3dfe31),
	.w6(32'h3bdb5a30),
	.w7(32'h3bb58086),
	.w8(32'h3aa75916),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7ad9e),
	.w1(32'h3bfa991e),
	.w2(32'h3c0e37ac),
	.w3(32'h3b2c430b),
	.w4(32'hbaeec4dc),
	.w5(32'h3c29c866),
	.w6(32'h3b97d327),
	.w7(32'hbc38acc2),
	.w8(32'hbc27aa32),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb503d80),
	.w1(32'hbb8e8cce),
	.w2(32'hbb6b69a0),
	.w3(32'hbb96532b),
	.w4(32'hbb274ee0),
	.w5(32'hbb00c85d),
	.w6(32'hbb2697fd),
	.w7(32'hba0425a5),
	.w8(32'hba55acdc),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a51b5e),
	.w1(32'h3bc59c01),
	.w2(32'h3bd08f9c),
	.w3(32'h3b910a13),
	.w4(32'h3b62bc2d),
	.w5(32'h3b16c60f),
	.w6(32'h3c0ce95a),
	.w7(32'h3b7e4dc9),
	.w8(32'h3b80e051),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b900c50),
	.w1(32'hbc1db099),
	.w2(32'hbbc7c5c4),
	.w3(32'hbb7d9eee),
	.w4(32'h3b277347),
	.w5(32'h3b240e74),
	.w6(32'h3af2c3f6),
	.w7(32'hbc1cdf7b),
	.w8(32'hbbb924cc),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5288b8),
	.w1(32'h3aa34441),
	.w2(32'hba9a32fa),
	.w3(32'h3b06013f),
	.w4(32'h39c5c130),
	.w5(32'hbacf1705),
	.w6(32'h3ab5b889),
	.w7(32'hba733014),
	.w8(32'hbb2439ba),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba01df4),
	.w1(32'h3b3304d7),
	.w2(32'h3c539073),
	.w3(32'h3c353cd2),
	.w4(32'h3c34ae23),
	.w5(32'h3c95008f),
	.w6(32'hbbe7c4ba),
	.w7(32'hbb973e63),
	.w8(32'hbc7e9d9d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dc2c7),
	.w1(32'hbc09aa3b),
	.w2(32'h3c6767ce),
	.w3(32'h3bbe11dd),
	.w4(32'h391767aa),
	.w5(32'h3b6799ec),
	.w6(32'h3b8258bc),
	.w7(32'hbc13ff46),
	.w8(32'hbc91ac16),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc562d7),
	.w1(32'hbcbaf7f3),
	.w2(32'hbcac5424),
	.w3(32'hbcc9cea7),
	.w4(32'hbd1247f2),
	.w5(32'hbc8b5266),
	.w6(32'h3d8412b8),
	.w7(32'h3d87e59e),
	.w8(32'h3d24f835),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcafdc9a),
	.w1(32'h3c61ac64),
	.w2(32'h3d192761),
	.w3(32'hbb1b7a02),
	.w4(32'h3cdb1a93),
	.w5(32'h3cf23722),
	.w6(32'h3cceb090),
	.w7(32'h3d282efa),
	.w8(32'h3ce1c625),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0870f3),
	.w1(32'hbbcf29dd),
	.w2(32'hbc1ad744),
	.w3(32'h3b1231c0),
	.w4(32'hbc1897cf),
	.w5(32'hbbdc1cc7),
	.w6(32'hbad4152d),
	.w7(32'hbc0d9935),
	.w8(32'h3bb6153a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad94b73),
	.w1(32'h3c6ef552),
	.w2(32'h3c82088d),
	.w3(32'h3bdc6349),
	.w4(32'h3c27193c),
	.w5(32'h3b8e8131),
	.w6(32'h3cf25534),
	.w7(32'h3ce06afa),
	.w8(32'h3cac11b0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0418d2),
	.w1(32'h39adacdd),
	.w2(32'hbb009381),
	.w3(32'hba5cc6ff),
	.w4(32'h3ac3802a),
	.w5(32'hbae750f9),
	.w6(32'h3b23b3d9),
	.w7(32'hb99d15c6),
	.w8(32'hbb2aafa0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f0308),
	.w1(32'h3b9edcab),
	.w2(32'h3a5e879e),
	.w3(32'h38378c76),
	.w4(32'h3918d3fd),
	.w5(32'hbab8adcc),
	.w6(32'h3af7eae4),
	.w7(32'hba0367db),
	.w8(32'hba4acd20),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c020b19),
	.w1(32'hbc824bfc),
	.w2(32'hbce6d6b6),
	.w3(32'hbc931425),
	.w4(32'hbd0ea4a2),
	.w5(32'hbd0c94cf),
	.w6(32'h3bf0f5eb),
	.w7(32'h3b6fab7a),
	.w8(32'hbb6f45fc),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d3166),
	.w1(32'hbce9b1f8),
	.w2(32'hbd20e488),
	.w3(32'hbc0c0e42),
	.w4(32'hbc7de9ef),
	.w5(32'hbc9fe035),
	.w6(32'h3d29c60c),
	.w7(32'h3d495469),
	.w8(32'h3cdf6456),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fe457),
	.w1(32'hbc881a28),
	.w2(32'hbc95f3fc),
	.w3(32'h3b059405),
	.w4(32'hbbec80d5),
	.w5(32'h3b0322eb),
	.w6(32'h3ca35299),
	.w7(32'h3cc30be9),
	.w8(32'h3d2540e6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a903b),
	.w1(32'hbbe21896),
	.w2(32'hbc6ba8c9),
	.w3(32'h3b51a84a),
	.w4(32'hbc2c757e),
	.w5(32'hbaf233e8),
	.w6(32'hbb9dfcec),
	.w7(32'h3c068ca7),
	.w8(32'h3c404203),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0931f5),
	.w1(32'h3c0262a3),
	.w2(32'h3adc6008),
	.w3(32'h3ae2c452),
	.w4(32'hbb72803e),
	.w5(32'h3bfd9c6c),
	.w6(32'hbc18cb03),
	.w7(32'hbc508714),
	.w8(32'h3b059480),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe661e),
	.w1(32'h3b5bb015),
	.w2(32'h3b80c21b),
	.w3(32'h3bce7d5e),
	.w4(32'h3b19aff9),
	.w5(32'h3b3e994c),
	.w6(32'hbbcf5e64),
	.w7(32'hbbe77bed),
	.w8(32'hbaaa3446),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b235917),
	.w1(32'h3b6a1bfd),
	.w2(32'hb98b87fd),
	.w3(32'h3bf60039),
	.w4(32'h3c80b168),
	.w5(32'h3bd7c643),
	.w6(32'hbba062f9),
	.w7(32'hbc7e3571),
	.w8(32'hbc098503),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39c7af),
	.w1(32'h38984cff),
	.w2(32'h3b2637e4),
	.w3(32'h3bb760d2),
	.w4(32'h3bb3acfc),
	.w5(32'hbb083751),
	.w6(32'hba382212),
	.w7(32'hbbcc1381),
	.w8(32'hbabcfbd3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae14b40),
	.w1(32'h3b55447b),
	.w2(32'h3bb0f554),
	.w3(32'h3b08dd92),
	.w4(32'h3b50411e),
	.w5(32'h3ab3c219),
	.w6(32'h3a31b3f7),
	.w7(32'hbacf3ef4),
	.w8(32'hbab60ccf),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6522fc),
	.w1(32'hbc971944),
	.w2(32'h3b9fcbf7),
	.w3(32'hbc3bddf4),
	.w4(32'hbc618da9),
	.w5(32'hbc518ee1),
	.w6(32'h3cb86ab1),
	.w7(32'h3d417d17),
	.w8(32'h3cdea2fb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80a2c1),
	.w1(32'h3d3b2f67),
	.w2(32'h3d46cd88),
	.w3(32'h3bb11ca4),
	.w4(32'h3cc3aef4),
	.w5(32'h3c7b5555),
	.w6(32'hbd05d0c8),
	.w7(32'hbd7ca03f),
	.w8(32'hbd943e37),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d7861),
	.w1(32'h3ab28bab),
	.w2(32'h3b244924),
	.w3(32'h3c82c5ae),
	.w4(32'hbbc8c663),
	.w5(32'hbca9cbef),
	.w6(32'h3b6b9aa4),
	.w7(32'h3b9fe723),
	.w8(32'h3cca0a63),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb165996),
	.w1(32'h3bc8e590),
	.w2(32'h3aefec91),
	.w3(32'h3c1353a1),
	.w4(32'h3b5c7067),
	.w5(32'h3b49950f),
	.w6(32'h3c024b7b),
	.w7(32'h3bab8ca9),
	.w8(32'h3b909b60),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54dba3),
	.w1(32'h3b959a3f),
	.w2(32'h3ae2f311),
	.w3(32'h3be3403e),
	.w4(32'h3bff3052),
	.w5(32'h3b9809b9),
	.w6(32'h3bae920f),
	.w7(32'h3b48512f),
	.w8(32'h3b950923),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c673098),
	.w1(32'h3a37a4e8),
	.w2(32'hbb9fe489),
	.w3(32'h3c8809c1),
	.w4(32'hbaccc0d4),
	.w5(32'hbc92154d),
	.w6(32'h3cb6217b),
	.w7(32'h3ca44e0d),
	.w8(32'h3c5a1cd9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad54cee),
	.w1(32'h3c0b2d6a),
	.w2(32'h3c0ef6ae),
	.w3(32'h3bd3bdea),
	.w4(32'h3b88ce2e),
	.w5(32'hba07186c),
	.w6(32'h3c04fbe8),
	.w7(32'h3b6461a2),
	.w8(32'hbc08c45d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2da36),
	.w1(32'hba138aa5),
	.w2(32'hbc24e26e),
	.w3(32'hbad7c308),
	.w4(32'h3ca9b679),
	.w5(32'hba40e112),
	.w6(32'hbd20e437),
	.w7(32'hbd661106),
	.w8(32'hbcea12aa),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca71f34),
	.w1(32'h3be7293a),
	.w2(32'h3c902235),
	.w3(32'hbc0ecb0f),
	.w4(32'hbc165abe),
	.w5(32'hbc57a751),
	.w6(32'hbbb717d9),
	.w7(32'h3b033d50),
	.w8(32'h3c439906),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0616b8),
	.w1(32'h3caccc33),
	.w2(32'h3c39327d),
	.w3(32'h3c142552),
	.w4(32'hba8bd520),
	.w5(32'hbb031fec),
	.w6(32'h3b72239e),
	.w7(32'h3ba72c83),
	.w8(32'h3aa08d4c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c199b7c),
	.w1(32'h3c31ea1e),
	.w2(32'h3bc9b85c),
	.w3(32'h3ba670eb),
	.w4(32'h3bc2b709),
	.w5(32'h3a2dfab0),
	.w6(32'hba890878),
	.w7(32'hbad60ad1),
	.w8(32'hbb6f7f2d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39988ed7),
	.w1(32'h3c964f1c),
	.w2(32'h3d0a7365),
	.w3(32'hbc60f783),
	.w4(32'h3bd7f7d5),
	.w5(32'h3cca5fc6),
	.w6(32'hbcab861b),
	.w7(32'hbd7d90b0),
	.w8(32'hbd2e2dde),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1784ab),
	.w1(32'h3c6b690e),
	.w2(32'h3c173624),
	.w3(32'h3c5c6ee4),
	.w4(32'h3c234b84),
	.w5(32'h3bb876de),
	.w6(32'h3c61507e),
	.w7(32'h3c54c3da),
	.w8(32'h3c0d1966),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c256672),
	.w1(32'h3c0670e0),
	.w2(32'h3c6b6b25),
	.w3(32'h3c0ae702),
	.w4(32'h3bd1f890),
	.w5(32'h3c594aa2),
	.w6(32'h3bf3515a),
	.w7(32'h3b96c1d5),
	.w8(32'h3c1b6b27),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbbcf81),
	.w1(32'h3c685377),
	.w2(32'h3c0fbba8),
	.w3(32'h3c83a267),
	.w4(32'h3c15033b),
	.w5(32'h3bf39cab),
	.w6(32'h3c7d118c),
	.w7(32'h3bb4ac61),
	.w8(32'hbb2604c6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fa8b9),
	.w1(32'h3c121ba9),
	.w2(32'h3bfb4236),
	.w3(32'hbba7410c),
	.w4(32'hbbbd3207),
	.w5(32'hba8c4e84),
	.w6(32'hbb853232),
	.w7(32'h3bcc6c57),
	.w8(32'h3bcc2105),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7546f),
	.w1(32'hbbc5d4d0),
	.w2(32'hbc1bbbb9),
	.w3(32'hbbbd0015),
	.w4(32'hbbd1203f),
	.w5(32'hbbe21b64),
	.w6(32'hbb48f1ad),
	.w7(32'h3a93dc28),
	.w8(32'h3a8c5923),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fda19),
	.w1(32'hbc5501ed),
	.w2(32'hbc0936d2),
	.w3(32'hbb408ddf),
	.w4(32'hbb9bca2a),
	.w5(32'hbb73937c),
	.w6(32'hbbc567b2),
	.w7(32'h3a872ed8),
	.w8(32'h3b080797),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14a8c1),
	.w1(32'h3c035c08),
	.w2(32'h3c0e232e),
	.w3(32'h3be9a9b2),
	.w4(32'h3bc399b7),
	.w5(32'h3be851db),
	.w6(32'h3bb83f36),
	.w7(32'h3b9a2637),
	.w8(32'h3bc61aff),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9010106),
	.w1(32'h3becf976),
	.w2(32'h3ca1852d),
	.w3(32'h3bc94544),
	.w4(32'h3c486a1b),
	.w5(32'h3a282319),
	.w6(32'h3b5c875b),
	.w7(32'h3c9c1934),
	.w8(32'h3acc02f7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ddf0b),
	.w1(32'hba8ac01f),
	.w2(32'hbb8739bf),
	.w3(32'h3a7e2a60),
	.w4(32'h3a23afb4),
	.w5(32'h3aed2e2d),
	.w6(32'h3b21a02c),
	.w7(32'h3aa84f01),
	.w8(32'h3a63e91c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe99625),
	.w1(32'hbb951136),
	.w2(32'hbc7c5b88),
	.w3(32'hbc9b585c),
	.w4(32'hbbb6b734),
	.w5(32'h3c2b8175),
	.w6(32'hbc2d3e2b),
	.w7(32'hbbc99f93),
	.w8(32'hbbf532e1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f66c8),
	.w1(32'hbbb74765),
	.w2(32'h3a8e991a),
	.w3(32'hbacf602f),
	.w4(32'hbaaadd10),
	.w5(32'hbb89cffd),
	.w6(32'hbad1fa03),
	.w7(32'h3a8d7955),
	.w8(32'hbba8beff),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2c6fc),
	.w1(32'h3ba5b8a5),
	.w2(32'h3c4cfc4c),
	.w3(32'h3ba196ba),
	.w4(32'h3c3d10c8),
	.w5(32'h3d036d5f),
	.w6(32'h3bc0d354),
	.w7(32'h3c981e8c),
	.w8(32'h3ca7948f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c744602),
	.w1(32'h3c60b820),
	.w2(32'h3c3d1254),
	.w3(32'hbb2904d9),
	.w4(32'hbc1013ca),
	.w5(32'hbcd79dde),
	.w6(32'h3bbaef29),
	.w7(32'h3bfbf813),
	.w8(32'hbc552dd7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd65788),
	.w1(32'hbc066076),
	.w2(32'h3acd2fef),
	.w3(32'hbbf7b057),
	.w4(32'h3bb31344),
	.w5(32'h3c234977),
	.w6(32'hbc1e4cf1),
	.w7(32'h3b143e72),
	.w8(32'h3bf5ae98),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule