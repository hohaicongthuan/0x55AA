module layer_6_featuremap_105(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d0a04),
	.w1(32'h3b30374f),
	.w2(32'hbaef4e66),
	.w3(32'h3b38ed2c),
	.w4(32'h3b7933e6),
	.w5(32'hba568cd7),
	.w6(32'h3a92b7fd),
	.w7(32'h3b8939c3),
	.w8(32'h3a7735d9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcad9a),
	.w1(32'h3b212596),
	.w2(32'h3ba4ea6e),
	.w3(32'hb9ec05c5),
	.w4(32'hbabd582e),
	.w5(32'hbad027fd),
	.w6(32'hbb51ddcb),
	.w7(32'hbb33532f),
	.w8(32'hbb09255a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988d367),
	.w1(32'hbc23dabb),
	.w2(32'hbb87af06),
	.w3(32'h3c5c9b76),
	.w4(32'h3c514ace),
	.w5(32'h3c6c6138),
	.w6(32'h3bed5aef),
	.w7(32'h3bb54bd5),
	.w8(32'h3beff931),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0ea1b),
	.w1(32'hbb8f3b0e),
	.w2(32'h3ab3fc7c),
	.w3(32'hbc0c96a3),
	.w4(32'hbc4223ad),
	.w5(32'hbba0d659),
	.w6(32'h3a844c8f),
	.w7(32'hba892754),
	.w8(32'h3b09f4d2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15e9f7),
	.w1(32'hbb509da7),
	.w2(32'h3b1b0d7e),
	.w3(32'h3b1650eb),
	.w4(32'h3b8c5e10),
	.w5(32'h3b9b935c),
	.w6(32'h3b4f1be5),
	.w7(32'h3ba19bba),
	.w8(32'h3b605600),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9abf16),
	.w1(32'hb9417124),
	.w2(32'hbb59c7a7),
	.w3(32'h3b372918),
	.w4(32'h3a9a1dd0),
	.w5(32'hbb0678c3),
	.w6(32'h3abe4b0b),
	.w7(32'hba615a0f),
	.w8(32'hbb75fe26),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab284a),
	.w1(32'h3c8579e9),
	.w2(32'h3c5b3e6a),
	.w3(32'h3c19ca09),
	.w4(32'h3c719a94),
	.w5(32'h3c0587a8),
	.w6(32'h3c00e6b4),
	.w7(32'h3c757eb7),
	.w8(32'h3c0f431e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08725c),
	.w1(32'hbb134feb),
	.w2(32'hbaef5c9a),
	.w3(32'hbb1d26b7),
	.w4(32'h3a9f36c8),
	.w5(32'h3a19e8d8),
	.w6(32'hbbe8d941),
	.w7(32'hbbaa12fd),
	.w8(32'hbaeb1a9f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a3a1f),
	.w1(32'hbc1b819f),
	.w2(32'hbb43c8e4),
	.w3(32'h3abff885),
	.w4(32'hbbc1a291),
	.w5(32'hbb369365),
	.w6(32'h3ae25b75),
	.w7(32'hbb629db7),
	.w8(32'hbb5a5cf8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81df0e),
	.w1(32'hbad96f8e),
	.w2(32'hbc054cd3),
	.w3(32'h3b82b9d0),
	.w4(32'hb9f4fef5),
	.w5(32'hbbadabf0),
	.w6(32'h3badd9b7),
	.w7(32'hba82c46d),
	.w8(32'hbbfe1f40),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd24bc9),
	.w1(32'hbc9c8b14),
	.w2(32'hbc56135f),
	.w3(32'hbc098343),
	.w4(32'hbbe346f5),
	.w5(32'hbbc9dcd2),
	.w6(32'hbc2b31b0),
	.w7(32'hbbbf300a),
	.w8(32'hbbdb2d4f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d16ab),
	.w1(32'h3bd1b245),
	.w2(32'h3b81f1fa),
	.w3(32'hba8f4062),
	.w4(32'hbb0ac57a),
	.w5(32'hb9a2ddb2),
	.w6(32'h39be546b),
	.w7(32'hbac87737),
	.w8(32'hbb3cbf65),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40d447),
	.w1(32'hbaff5407),
	.w2(32'h3865267a),
	.w3(32'hbaefdc51),
	.w4(32'hbacbd56d),
	.w5(32'hba7e62c0),
	.w6(32'hbaf962a2),
	.w7(32'hba0081dc),
	.w8(32'h3a048856),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c1acd),
	.w1(32'hbcc09d8d),
	.w2(32'hbc3daa66),
	.w3(32'hb8fd0c8d),
	.w4(32'h3771ccea),
	.w5(32'hbba26736),
	.w6(32'hbb8dbf57),
	.w7(32'hbbb8af31),
	.w8(32'hbc2268d5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba673479),
	.w1(32'hbac35a12),
	.w2(32'hb96f2f6a),
	.w3(32'hba887566),
	.w4(32'hbb0e39cf),
	.w5(32'hbb17cd3e),
	.w6(32'h3b80b7a8),
	.w7(32'h3b45003f),
	.w8(32'h3b319f81),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03eda4),
	.w1(32'hbbafd34e),
	.w2(32'hbb05d41d),
	.w3(32'hbb227493),
	.w4(32'hbaa19988),
	.w5(32'hba7eaad9),
	.w6(32'h3b1a4dac),
	.w7(32'h3b6b89ea),
	.w8(32'h3b571371),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01d3df),
	.w1(32'hbceccfb7),
	.w2(32'h3b842d1b),
	.w3(32'hbbac57cd),
	.w4(32'h3c862076),
	.w5(32'h3ca6f4c2),
	.w6(32'h3cc43287),
	.w7(32'h3c90e2fb),
	.w8(32'h3c68c057),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3872be89),
	.w1(32'hba80fc71),
	.w2(32'hbaf157f3),
	.w3(32'h39ea1678),
	.w4(32'h39118cf0),
	.w5(32'hbaa8d5cb),
	.w6(32'h397c3699),
	.w7(32'hb9b32245),
	.w8(32'hbb049e6a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c4358),
	.w1(32'hbb48c500),
	.w2(32'h3b17b4a1),
	.w3(32'hbb0eb6b4),
	.w4(32'hbb1a6c0f),
	.w5(32'h3b439c1f),
	.w6(32'hbb1b1409),
	.w7(32'hbab8c796),
	.w8(32'h3b24261d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb39b26),
	.w1(32'hbc19b7ee),
	.w2(32'hbc085a54),
	.w3(32'hba363223),
	.w4(32'hbb54dbd5),
	.w5(32'hbb4d6b78),
	.w6(32'h3b617e4f),
	.w7(32'hb9aa0973),
	.w8(32'hbabebddb),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0779),
	.w1(32'h3a398123),
	.w2(32'h3aa11d7e),
	.w3(32'hba6b3123),
	.w4(32'h3a1e2895),
	.w5(32'h3b806be1),
	.w6(32'hbac49f9f),
	.w7(32'hba6d35f3),
	.w8(32'hb8e6c380),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f23ec),
	.w1(32'hbcb323ec),
	.w2(32'hbbdd67e8),
	.w3(32'hbb8a87b6),
	.w4(32'hbaf22b20),
	.w5(32'h3b83a468),
	.w6(32'h3b2e9901),
	.w7(32'h3b96a6db),
	.w8(32'h3be53feb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4cd252),
	.w1(32'hb8f1c80d),
	.w2(32'hba8ffc17),
	.w3(32'hba9d00a1),
	.w4(32'hba8f8e79),
	.w5(32'h3a1a9cc0),
	.w6(32'hbbda6ac8),
	.w7(32'hbc0076c2),
	.w8(32'hbba6fb0a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51b4fc),
	.w1(32'hbcddc26c),
	.w2(32'hbc864000),
	.w3(32'hbb979925),
	.w4(32'h3bdf7873),
	.w5(32'h3aec2795),
	.w6(32'hbc0a542b),
	.w7(32'h3c5ab822),
	.w8(32'h3b5a6331),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc771518),
	.w1(32'hbc7efc8c),
	.w2(32'hba0c750e),
	.w3(32'hbc90aa22),
	.w4(32'hbc9cfc36),
	.w5(32'hb925becc),
	.w6(32'h3cca5673),
	.w7(32'h3cb04f7e),
	.w8(32'h3c9f8bfb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc828e36),
	.w1(32'hbcca19e9),
	.w2(32'hbc7f4283),
	.w3(32'hbccac17a),
	.w4(32'hbcfaa900),
	.w5(32'hbc82a6e1),
	.w6(32'hbb8e09ee),
	.w7(32'hbc318beb),
	.w8(32'hbbb7a85e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb1a27),
	.w1(32'hbb83bcbd),
	.w2(32'hbbe8225d),
	.w3(32'h3be8f70e),
	.w4(32'h3bf73693),
	.w5(32'h3b0f7a69),
	.w6(32'hbb7cb5bb),
	.w7(32'h3b18d045),
	.w8(32'hbaa3e427),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb082f76),
	.w1(32'hbb221398),
	.w2(32'h3acf4e0e),
	.w3(32'h3921d567),
	.w4(32'hb98a1a8b),
	.w5(32'h3b056ede),
	.w6(32'h3a652a93),
	.w7(32'h3a83862e),
	.w8(32'h3baf681a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae15e6),
	.w1(32'hbaae3844),
	.w2(32'hb8f59963),
	.w3(32'hba03296c),
	.w4(32'hb92db30d),
	.w5(32'h3a1264fe),
	.w6(32'h39c6c049),
	.w7(32'h39766d49),
	.w8(32'h3ae2e6f7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1bf18),
	.w1(32'h3c526d39),
	.w2(32'hbc9e304d),
	.w3(32'hbd8021d4),
	.w4(32'hbd566172),
	.w5(32'hbd09c0f0),
	.w6(32'hbd304491),
	.w7(32'hbd46f1f4),
	.w8(32'hbc15fb0a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba37b5b),
	.w1(32'h3985eb0d),
	.w2(32'h3b68386b),
	.w3(32'h3b82358b),
	.w4(32'h3b913603),
	.w5(32'h3b9ccc79),
	.w6(32'h3b53b567),
	.w7(32'h3b9f14d1),
	.w8(32'h3c04a710),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b79b87),
	.w1(32'hbb460543),
	.w2(32'h3b66091d),
	.w3(32'hbb1e7260),
	.w4(32'hbb5eee1b),
	.w5(32'hba849531),
	.w6(32'h3acf9765),
	.w7(32'h3b9aad30),
	.w8(32'h3b0536cf),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f9d3c),
	.w1(32'hba7a7c9f),
	.w2(32'hbac86963),
	.w3(32'h3aac0406),
	.w4(32'h3b06cc62),
	.w5(32'hbacaba0d),
	.w6(32'h390e316b),
	.w7(32'h3a75b8cb),
	.w8(32'h3a5e9b9f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a2050),
	.w1(32'hba781527),
	.w2(32'hbae35f4a),
	.w3(32'hbb4b2243),
	.w4(32'hbab6ad4e),
	.w5(32'hba32847a),
	.w6(32'hbafbcdd7),
	.w7(32'hbb290473),
	.w8(32'hbb3c0a6c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3aef2),
	.w1(32'hb9df5104),
	.w2(32'hbb236480),
	.w3(32'h3acc5abd),
	.w4(32'hb9ddd33d),
	.w5(32'hba52ebd3),
	.w6(32'h399bbd7d),
	.w7(32'hbadd03a7),
	.w8(32'hbb293d4d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac518e0),
	.w1(32'hba425fcf),
	.w2(32'h3a87c6e7),
	.w3(32'hbb45bbc8),
	.w4(32'hbb65699f),
	.w5(32'h3be8d6c4),
	.w6(32'h3b8df189),
	.w7(32'hbb2b85e1),
	.w8(32'h3bb75fa4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafda9db),
	.w1(32'h3821a68e),
	.w2(32'hba8ba3c6),
	.w3(32'h3b35d4df),
	.w4(32'h3b11fa74),
	.w5(32'hbaea4ca0),
	.w6(32'h3b167ba0),
	.w7(32'h3ac11009),
	.w8(32'hbb3d218e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fdce2),
	.w1(32'h3c1a331a),
	.w2(32'h3c08d89c),
	.w3(32'h3a42a81f),
	.w4(32'h3b0e0918),
	.w5(32'h3be2ec7e),
	.w6(32'h3c5d0750),
	.w7(32'h3c1c4906),
	.w8(32'h3c0d823d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b324cd4),
	.w1(32'h3a562f1d),
	.w2(32'hb934e110),
	.w3(32'hbacd6a3b),
	.w4(32'hbaa8fb9c),
	.w5(32'h39d7e1ea),
	.w6(32'h38403843),
	.w7(32'h3b133263),
	.w8(32'h3bbae16f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd220260),
	.w1(32'hbd1db3a0),
	.w2(32'hbc5b46d6),
	.w3(32'h3d0ebb03),
	.w4(32'h3cef8a0f),
	.w5(32'h3c8d9510),
	.w6(32'h3ccd31ef),
	.w7(32'h3ca77503),
	.w8(32'h3c448248),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba08f4c),
	.w1(32'hbba299bd),
	.w2(32'hbbe96e2f),
	.w3(32'h3b1c6f1f),
	.w4(32'hbba3a842),
	.w5(32'hbc0f3ee9),
	.w6(32'h3bf5c578),
	.w7(32'h3aff53a7),
	.w8(32'hbb9060b0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c059215),
	.w1(32'h3b59e5d0),
	.w2(32'h3b6fc3cf),
	.w3(32'hba8bdeb1),
	.w4(32'h3a785172),
	.w5(32'h3bd738eb),
	.w6(32'hb982cb21),
	.w7(32'hbaecc69e),
	.w8(32'h3accb2d2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e4a56),
	.w1(32'h3affe4fc),
	.w2(32'h39ae4757),
	.w3(32'h3a869302),
	.w4(32'h399486f9),
	.w5(32'h3a6aa7fe),
	.w6(32'h3aabb7d9),
	.w7(32'hba34c18b),
	.w8(32'hb9c56f9e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba85837),
	.w1(32'h3ca4642b),
	.w2(32'h3ba05fa4),
	.w3(32'hbd7bc710),
	.w4(32'hbd530529),
	.w5(32'hbc001db6),
	.w6(32'hbca8afd5),
	.w7(32'hbcb6fcd8),
	.w8(32'h3c6e25e1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc926cbd),
	.w1(32'hbcb9e9c1),
	.w2(32'hbb4ff39c),
	.w3(32'h3c025b5a),
	.w4(32'h3c59cad1),
	.w5(32'h3c886aec),
	.w6(32'h3b958ab5),
	.w7(32'h3c2fef0b),
	.w8(32'h3c53fe05),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f713f9),
	.w1(32'h3aa70a36),
	.w2(32'h3b4dd2ff),
	.w3(32'h3b1fdb62),
	.w4(32'h3b405496),
	.w5(32'h3a87acea),
	.w6(32'h3b4274bb),
	.w7(32'h3b5bcd17),
	.w8(32'h3b3bde1a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22b86c),
	.w1(32'h3b84defb),
	.w2(32'h3c24fc59),
	.w3(32'h39590439),
	.w4(32'hba94bf27),
	.w5(32'hbb9cdc25),
	.w6(32'hbac1523a),
	.w7(32'hba905b90),
	.w8(32'h3b970a24),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f95e8),
	.w1(32'hbbd5338e),
	.w2(32'hbad51f3c),
	.w3(32'hbcbdd718),
	.w4(32'hbc8c972a),
	.w5(32'hbbdde5f1),
	.w6(32'hbc8ab733),
	.w7(32'hbc801ebe),
	.w8(32'hbb60aeff),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad50f6e),
	.w1(32'h3b5bd5de),
	.w2(32'h3bc0cedd),
	.w3(32'h3c490f37),
	.w4(32'h3c2ce165),
	.w5(32'h3c072ff2),
	.w6(32'h3c50a6f4),
	.w7(32'h3c2a5a5a),
	.w8(32'h3bd50bce),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ddcdc),
	.w1(32'hbc3f2a8c),
	.w2(32'hbc867cba),
	.w3(32'h3c1f1753),
	.w4(32'hbbd0625f),
	.w5(32'hbc8c312c),
	.w6(32'h3be879eb),
	.w7(32'h3baf1f59),
	.w8(32'hba32e0c7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab484e9),
	.w1(32'hbc22cc1a),
	.w2(32'hbbc12c2f),
	.w3(32'hbc17bc39),
	.w4(32'hbc46b3d7),
	.w5(32'hbbc476dd),
	.w6(32'hb960d7ca),
	.w7(32'hbb987c65),
	.w8(32'h39cde692),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e41aa),
	.w1(32'hbc3d7c56),
	.w2(32'hbc195df6),
	.w3(32'hbafa054e),
	.w4(32'hbc13847c),
	.w5(32'hbbcdd09d),
	.w6(32'h3b33dadd),
	.w7(32'hbbc20e8a),
	.w8(32'hbb8cc950),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1935f8),
	.w1(32'hbcaf1340),
	.w2(32'h3c253da5),
	.w3(32'hba76b235),
	.w4(32'h3c42bad6),
	.w5(32'h3c960bcb),
	.w6(32'hba85b67e),
	.w7(32'h3c687a67),
	.w8(32'h3cb151b2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a6cf0),
	.w1(32'h3c3291db),
	.w2(32'h3c404fbe),
	.w3(32'h3c8d5e2b),
	.w4(32'h3c8e22a5),
	.w5(32'h3c652e98),
	.w6(32'h3c5960a0),
	.w7(32'h3cab3bc5),
	.w8(32'h3c915e1e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f0392),
	.w1(32'h3897c9e3),
	.w2(32'hbab99cf2),
	.w3(32'hba79e678),
	.w4(32'hbb8f941d),
	.w5(32'hbb8356e8),
	.w6(32'hbb887364),
	.w7(32'hbb9a2e97),
	.w8(32'hbbaa57a2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14fc67),
	.w1(32'hbceba8bf),
	.w2(32'hbcbff647),
	.w3(32'hbd0f748e),
	.w4(32'hbd201f79),
	.w5(32'hbbffffd0),
	.w6(32'hbd01b424),
	.w7(32'hbd1b369a),
	.w8(32'hba0cc7a8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87058b),
	.w1(32'h3b1a1b4e),
	.w2(32'hbb76d498),
	.w3(32'h3bfb3d0c),
	.w4(32'h3b820ef4),
	.w5(32'hbbc032ae),
	.w6(32'h3c58e3ea),
	.w7(32'h3c06e45b),
	.w8(32'h39334343),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4b76d),
	.w1(32'hbc30f665),
	.w2(32'hbbf36543),
	.w3(32'h3a3a4e65),
	.w4(32'hbc87deed),
	.w5(32'hbc579d04),
	.w6(32'hbc2d83f3),
	.w7(32'hbcdd0e41),
	.w8(32'hbc758f9d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdb1b7),
	.w1(32'h3b24f634),
	.w2(32'hbb324c34),
	.w3(32'h3b4abeee),
	.w4(32'h3a03bb7f),
	.w5(32'hbb00f58f),
	.w6(32'h3a87b597),
	.w7(32'hbb848a10),
	.w8(32'hbc1328ac),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2ad8a9),
	.w1(32'hbd25b6f8),
	.w2(32'h3b676423),
	.w3(32'hbbf34f70),
	.w4(32'hbd080420),
	.w5(32'h3c05eaa7),
	.w6(32'h3ca5fba4),
	.w7(32'h3c5f8b92),
	.w8(32'h3ca3e3b7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badeffb),
	.w1(32'hbc80e78d),
	.w2(32'hbc4f99fa),
	.w3(32'hbbd36fcc),
	.w4(32'hbca865ab),
	.w5(32'hbc5eb8d0),
	.w6(32'hbc9b79f9),
	.w7(32'hbcd755ab),
	.w8(32'hbcaae6df),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccac66f),
	.w1(32'hbd26057a),
	.w2(32'hbd0ca504),
	.w3(32'hbbaad462),
	.w4(32'hbcf10e02),
	.w5(32'h3c06c351),
	.w6(32'h3a342bb8),
	.w7(32'hbc7b6641),
	.w8(32'h3cfe8050),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d835dbf),
	.w1(32'h3d552003),
	.w2(32'hbbd0357c),
	.w3(32'hbd0afcb6),
	.w4(32'hbd196447),
	.w5(32'hbc8a6cb8),
	.w6(32'hbd1c2cd9),
	.w7(32'hbd74bbfa),
	.w8(32'hbb574cef),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83c065),
	.w1(32'hbad89220),
	.w2(32'hbb92792b),
	.w3(32'hbbcd4ae1),
	.w4(32'hbbe2babe),
	.w5(32'hbbafb363),
	.w6(32'hbc2e4bba),
	.w7(32'hbc375e24),
	.w8(32'hbc4b5b74),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule