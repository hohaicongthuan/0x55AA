module layer_10_featuremap_136(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5517bae),
	.w1(32'hb5c438a9),
	.w2(32'hb48565fb),
	.w3(32'hb5ba7784),
	.w4(32'hb5968a6e),
	.w5(32'h32e01a28),
	.w6(32'hb57321b2),
	.w7(32'h363eda1e),
	.w8(32'h345b20c1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dc7ec8),
	.w1(32'hb8ae027d),
	.w2(32'hb8a72f11),
	.w3(32'h38a54b2a),
	.w4(32'hb63c5e83),
	.w5(32'h3902b19f),
	.w6(32'h38d47982),
	.w7(32'h37c93f8b),
	.w8(32'h38957640),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3410630b),
	.w1(32'hb5e71e91),
	.w2(32'hb6088586),
	.w3(32'h35931bb3),
	.w4(32'h353a9a53),
	.w5(32'hb64ae0ff),
	.w6(32'hb667b041),
	.w7(32'hb5a61963),
	.w8(32'hb61990f3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cc76d8),
	.w1(32'h356327b8),
	.w2(32'h37688d40),
	.w3(32'h37f28718),
	.w4(32'h36eea007),
	.w5(32'h38051058),
	.w6(32'h37fdb670),
	.w7(32'hb842daec),
	.w8(32'hb80b7d98),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h354e2510),
	.w1(32'hb6b3d77b),
	.w2(32'hb67ea6bd),
	.w3(32'hb65d4141),
	.w4(32'hb5ceb75c),
	.w5(32'hb5701129),
	.w6(32'hb614fa16),
	.w7(32'h320cde3e),
	.w8(32'h35a2f632),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb663b4fa),
	.w1(32'hb5859cd9),
	.w2(32'h34f58c49),
	.w3(32'hb68d12b1),
	.w4(32'hb674c1f8),
	.w5(32'hb525fe75),
	.w6(32'hb6d06bf1),
	.w7(32'hb65c59a2),
	.w8(32'hb61dc40a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e23537),
	.w1(32'hb80c7dc9),
	.w2(32'hb855a9ce),
	.w3(32'hb9ce81c0),
	.w4(32'hb994ad35),
	.w5(32'hba1c107f),
	.w6(32'hb994f949),
	.w7(32'hba01c5fd),
	.w8(32'hba4ec38b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39edc5f2),
	.w1(32'hba687545),
	.w2(32'hba679a05),
	.w3(32'hb7ad8d04),
	.w4(32'hba0e9b8c),
	.w5(32'hba6bcacf),
	.w6(32'hb9e7d951),
	.w7(32'h3961a820),
	.w8(32'hba7e312d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae6c6f),
	.w1(32'h39909e18),
	.w2(32'h398f059f),
	.w3(32'h39cf5fe4),
	.w4(32'h39b40e67),
	.w5(32'h3986f5b0),
	.w6(32'h399991c1),
	.w7(32'h39988c92),
	.w8(32'h39778113),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39809c8b),
	.w1(32'h391eb192),
	.w2(32'h39d319e2),
	.w3(32'hb890b922),
	.w4(32'hb9188c7a),
	.w5(32'h382876b6),
	.w6(32'hb9dc2077),
	.w7(32'hba88b18f),
	.w8(32'hba91a234),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3796f7d3),
	.w1(32'h396debe9),
	.w2(32'hb904764c),
	.w3(32'h37c36f45),
	.w4(32'h3926e939),
	.w5(32'hb8d1d51e),
	.w6(32'h3804f6c0),
	.w7(32'hb8685dae),
	.w8(32'hb932761c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fcca39),
	.w1(32'hb8c222da),
	.w2(32'h39d855f5),
	.w3(32'hba4650ed),
	.w4(32'hb9bee7a6),
	.w5(32'hba214c03),
	.w6(32'hba07c60a),
	.w7(32'hba4802d2),
	.w8(32'hbaa83611),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944336f),
	.w1(32'h3933fbbf),
	.w2(32'hb87e2ee9),
	.w3(32'hb9ff59b0),
	.w4(32'hb99b0a8e),
	.w5(32'hba3f4ff9),
	.w6(32'hb99f610b),
	.w7(32'hb9dcada5),
	.w8(32'hba61fb3a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa3a53),
	.w1(32'hb993e2ee),
	.w2(32'hb9fbe3df),
	.w3(32'hb9d5258e),
	.w4(32'hb9cb8484),
	.w5(32'hb9e86866),
	.w6(32'hb9d63ab4),
	.w7(32'hb9ad6d37),
	.w8(32'hb9c37a82),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fbdfc6),
	.w1(32'hb886fde0),
	.w2(32'hb89eccbd),
	.w3(32'h38ea7f1b),
	.w4(32'hb892153e),
	.w5(32'hb887b176),
	.w6(32'h39acea2a),
	.w7(32'hb8d5faa3),
	.w8(32'hb9689c33),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0d361),
	.w1(32'h3a751fe9),
	.w2(32'hb9b3cb51),
	.w3(32'h392c5c9c),
	.w4(32'h39ce11c4),
	.w5(32'hb9e1e254),
	.w6(32'hb99eabdd),
	.w7(32'hb93b9054),
	.w8(32'hba1ae456),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399612b9),
	.w1(32'hb8e3578e),
	.w2(32'hb90edef0),
	.w3(32'h3a10ef67),
	.w4(32'hb847f5d4),
	.w5(32'hb908a16a),
	.w6(32'h3923effa),
	.w7(32'hb95d087c),
	.w8(32'hb9b96f1c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96cf062),
	.w1(32'h38dcf20b),
	.w2(32'hba1e04b8),
	.w3(32'hb90253b2),
	.w4(32'hba2326f2),
	.w5(32'hba7ce701),
	.w6(32'hba1b800c),
	.w7(32'hba3db7c9),
	.w8(32'hba76e719),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8abf168),
	.w1(32'h3904367d),
	.w2(32'h37dcf9df),
	.w3(32'hb91c1048),
	.w4(32'hb961fa1c),
	.w5(32'hb95997bf),
	.w6(32'hb9121152),
	.w7(32'hb96376db),
	.w8(32'hb98ad395),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3503a960),
	.w1(32'hb61b6298),
	.w2(32'hb6582cc8),
	.w3(32'hb60afe3b),
	.w4(32'h36316894),
	.w5(32'hb69576e6),
	.w6(32'hb618a540),
	.w7(32'hb4d74f91),
	.w8(32'hb69c9f2c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6369a6c),
	.w1(32'h3688d6af),
	.w2(32'h35848945),
	.w3(32'hb606d26d),
	.w4(32'h36f1afec),
	.w5(32'h367d7fd3),
	.w6(32'h3656838a),
	.w7(32'h371b0896),
	.w8(32'h36d85418),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372fe4b1),
	.w1(32'hb896dfa9),
	.w2(32'h3796d724),
	.w3(32'h37b20322),
	.w4(32'hb7710a6b),
	.w5(32'h390d2250),
	.w6(32'h385ef3fb),
	.w7(32'hb7981db7),
	.w8(32'h38c49fa3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f1fcd),
	.w1(32'h3a840dd5),
	.w2(32'h38db2948),
	.w3(32'hb99bcd04),
	.w4(32'h3a060918),
	.w5(32'hba0dd4a2),
	.w6(32'hba27fbe0),
	.w7(32'hba7b9642),
	.w8(32'hba1e76b5),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c6cf5),
	.w1(32'hb728818b),
	.w2(32'hb786ca4f),
	.w3(32'h38b1f5ea),
	.w4(32'hb918d81d),
	.w5(32'hb8ca04dc),
	.w6(32'hb97530b6),
	.w7(32'hb9ed1eba),
	.w8(32'hb9b35a1a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9974465),
	.w1(32'hb9878c99),
	.w2(32'hb98d35e7),
	.w3(32'hb91d8314),
	.w4(32'hb8449571),
	.w5(32'h39fcada1),
	.w6(32'h39850692),
	.w7(32'h38354b95),
	.w8(32'h39d30a9f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38985581),
	.w1(32'h381d9239),
	.w2(32'hb80630ba),
	.w3(32'h3741b0ff),
	.w4(32'h371a78d7),
	.w5(32'hb6ea648f),
	.w6(32'hb86db558),
	.w7(32'hb8add231),
	.w8(32'hb8681807),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fe28f9),
	.w1(32'hb74040a4),
	.w2(32'hb76bb785),
	.w3(32'hb77a4a44),
	.w4(32'hb711e523),
	.w5(32'hb6abfc52),
	.w6(32'hb737792a),
	.w7(32'hb63678de),
	.w8(32'hb755ddc2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43b6b9),
	.w1(32'h3a6ec815),
	.w2(32'h39b6c471),
	.w3(32'h3a5e6492),
	.w4(32'h3989272f),
	.w5(32'hb9b2c7e2),
	.w6(32'hb7f8e719),
	.w7(32'h38b68a74),
	.w8(32'hba2422fa),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d97f0d),
	.w1(32'hb95930c0),
	.w2(32'hb91b374e),
	.w3(32'hb9f22945),
	.w4(32'hb9f9e9ca),
	.w5(32'hb99662ed),
	.w6(32'hba039441),
	.w7(32'hba2bed4b),
	.w8(32'hba2094a2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a522ed8),
	.w1(32'h39b45476),
	.w2(32'hb8da017d),
	.w3(32'h3a92e29b),
	.w4(32'h3a0f548d),
	.w5(32'h3999b763),
	.w6(32'h3a2c74a9),
	.w7(32'h39221a3a),
	.w8(32'hb9407b86),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7954072),
	.w1(32'hb78d5d36),
	.w2(32'hb7cc3ce5),
	.w3(32'hb7723d34),
	.w4(32'hb793b1e2),
	.w5(32'hb7c87ced),
	.w6(32'hb7552305),
	.w7(32'hb7ed9a7f),
	.w8(32'hb83b3839),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e368aa),
	.w1(32'hb8339adc),
	.w2(32'hb88ff471),
	.w3(32'h387e0d3b),
	.w4(32'hb87eb0a2),
	.w5(32'hb8b0ceac),
	.w6(32'h3849386c),
	.w7(32'hb8d769a7),
	.w8(32'hb90cd630),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926c80b),
	.w1(32'hb9c2735c),
	.w2(32'hba098dc8),
	.w3(32'hb8ad25ed),
	.w4(32'hb9f4a911),
	.w5(32'hba30b151),
	.w6(32'hb98e8dcd),
	.w7(32'hba451b2a),
	.w8(32'hba876601),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3965356f),
	.w1(32'h38c7b3cd),
	.w2(32'hb8f95541),
	.w3(32'h39842432),
	.w4(32'h399da1fb),
	.w5(32'h39827a71),
	.w6(32'h398b9a97),
	.w7(32'h39afae87),
	.w8(32'h398f7cd7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6846ff9),
	.w1(32'h38971ff4),
	.w2(32'h3908fc55),
	.w3(32'hb7caeed7),
	.w4(32'h3669cb3b),
	.w5(32'hb824c6a4),
	.w6(32'hb88895bd),
	.w7(32'hb8a68f82),
	.w8(32'hb9091929),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93fbdbb),
	.w1(32'hb96a6f4a),
	.w2(32'hb959c6a6),
	.w3(32'hb8944030),
	.w4(32'hb9039447),
	.w5(32'hb9ab6801),
	.w6(32'hb808e41b),
	.w7(32'hb9876c16),
	.w8(32'hb99bfec4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cbadf),
	.w1(32'hb96a2525),
	.w2(32'h399ad554),
	.w3(32'h38aee092),
	.w4(32'hb91ee819),
	.w5(32'h3627483b),
	.w6(32'h39bc1ba8),
	.w7(32'hba290f14),
	.w8(32'hba53e303),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3910b397),
	.w1(32'hb925c873),
	.w2(32'h39ebab6a),
	.w3(32'h3a39bc1c),
	.w4(32'h3868b58a),
	.w5(32'h3a841361),
	.w6(32'h3a63b7d5),
	.w7(32'hb6c1624e),
	.w8(32'h3a01323d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c58ab),
	.w1(32'hb9844164),
	.w2(32'h39a6add0),
	.w3(32'h39cb98eb),
	.w4(32'h39f45981),
	.w5(32'h3aa4cd9a),
	.w6(32'h3a0cfbb1),
	.w7(32'h3a106301),
	.w8(32'h3aae2419),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ed56fd),
	.w1(32'hb8df2e5a),
	.w2(32'h3856efd5),
	.w3(32'h37d2ac33),
	.w4(32'hb8236a22),
	.w5(32'h3917116e),
	.w6(32'h38ad8244),
	.w7(32'hb82ea412),
	.w8(32'h38cbd93f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d56a2),
	.w1(32'h3968865e),
	.w2(32'h3970d183),
	.w3(32'h38f0f0b9),
	.w4(32'h388ac578),
	.w5(32'h38f37159),
	.w6(32'hb7808e9b),
	.w7(32'hb8710a7b),
	.w8(32'h38f4d983),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cc2c5c),
	.w1(32'h3886500b),
	.w2(32'h36f282fd),
	.w3(32'h37684906),
	.w4(32'h38b010bb),
	.w5(32'h3813e38b),
	.w6(32'h389f71c0),
	.w7(32'h39029164),
	.w8(32'h38944919),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb930083e),
	.w1(32'hb8e5c17b),
	.w2(32'hb9780ccf),
	.w3(32'hb8e4dc70),
	.w4(32'hb9257afd),
	.w5(32'hb9378da7),
	.w6(32'hb8696715),
	.w7(32'hb9050da9),
	.w8(32'hb9335330),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383f5707),
	.w1(32'h3a3c8a41),
	.w2(32'hb8a07cb6),
	.w3(32'hba399c4c),
	.w4(32'hb9b9ec68),
	.w5(32'hba9d17c1),
	.w6(32'hbade05fe),
	.w7(32'hbab2b544),
	.w8(32'hbad0ab0b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e7247),
	.w1(32'h3905099d),
	.w2(32'h38e6aaf0),
	.w3(32'h39d4f165),
	.w4(32'h3878ef14),
	.w5(32'h39b7d162),
	.w6(32'h397d7294),
	.w7(32'hb8b5d56a),
	.w8(32'h391877fc),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab4c1c),
	.w1(32'h38a7a8f2),
	.w2(32'h389072d5),
	.w3(32'h397e0091),
	.w4(32'h398df618),
	.w5(32'h38d0fc38),
	.w6(32'hb6e27f0f),
	.w7(32'hb8a4ebd2),
	.w8(32'h394efc9d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa1370),
	.w1(32'h3aaac362),
	.w2(32'h3aa36f18),
	.w3(32'h3a8b6a9e),
	.w4(32'h3a9857ee),
	.w5(32'h3a9f8cea),
	.w6(32'h3a72b91a),
	.w7(32'h3a2cf601),
	.w8(32'h3a895566),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ffcf23),
	.w1(32'h3a0b0d27),
	.w2(32'h3a45a7a5),
	.w3(32'hb9ab0af4),
	.w4(32'hb8abb988),
	.w5(32'hb96f5e24),
	.w6(32'hb9eca8c0),
	.w7(32'hba0de910),
	.w8(32'hba2796b9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e22244),
	.w1(32'h3727cbe3),
	.w2(32'h39048b17),
	.w3(32'hb98f35d5),
	.w4(32'hb80c6466),
	.w5(32'h38b92328),
	.w6(32'hb924c547),
	.w7(32'hb964683b),
	.w8(32'h3904fff3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961d761),
	.w1(32'h39e2b3f3),
	.w2(32'h3a22562b),
	.w3(32'h3838f3c5),
	.w4(32'h3a23973b),
	.w5(32'h3a24e7d3),
	.w6(32'h39c4eb25),
	.w7(32'h3a2c1a57),
	.w8(32'h3a39cca5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6c4d1),
	.w1(32'hb9b00638),
	.w2(32'hb9a68dd3),
	.w3(32'hba252181),
	.w4(32'hb9c60222),
	.w5(32'hb98aa714),
	.w6(32'hba1ab982),
	.w7(32'hb95659c0),
	.w8(32'h384457f1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38824223),
	.w1(32'h39a455d6),
	.w2(32'hb9561be3),
	.w3(32'hb856ee8c),
	.w4(32'h37ac3176),
	.w5(32'hb99cc87f),
	.w6(32'hb9ce1e26),
	.w7(32'hb9a65f4b),
	.w8(32'hb98050bb),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b38cc4),
	.w1(32'hb8144f23),
	.w2(32'hb979b42e),
	.w3(32'hb6cdb303),
	.w4(32'h37006bc1),
	.w5(32'hb946c380),
	.w6(32'hb84ae164),
	.w7(32'h37fe15c0),
	.w8(32'hb8da1a7c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b16eb1),
	.w1(32'h39d70a00),
	.w2(32'hb8fa3781),
	.w3(32'hba01dad7),
	.w4(32'hb98e9ccc),
	.w5(32'hba2ce14a),
	.w6(32'hb9a2a896),
	.w7(32'hba1eaa02),
	.w8(32'hba904efa),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9785c83),
	.w1(32'hb81b7a5f),
	.w2(32'hb963228e),
	.w3(32'hb99e8f9c),
	.w4(32'hb98ae909),
	.w5(32'hb98e104f),
	.w6(32'hb9bda9ae),
	.w7(32'hb8134797),
	.w8(32'hb986e684),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f0b3a1),
	.w1(32'hb6fbc7ae),
	.w2(32'h37039cb7),
	.w3(32'h37be4c63),
	.w4(32'h37a02338),
	.w5(32'h38310d9f),
	.w6(32'h3825292d),
	.w7(32'h37aea166),
	.w8(32'h38211c0b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5654a3e),
	.w1(32'hb55729aa),
	.w2(32'h3561fb37),
	.w3(32'hb4ba5ef1),
	.w4(32'h368e5c53),
	.w5(32'h36f23570),
	.w6(32'h36026793),
	.w7(32'h35375e08),
	.w8(32'h36db6b04),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37854ff5),
	.w1(32'hb7f02dcb),
	.w2(32'hb6b95677),
	.w3(32'h3893c574),
	.w4(32'h37764b03),
	.w5(32'h387769bd),
	.w6(32'h37d15293),
	.w7(32'hb7027765),
	.w8(32'h37d229c0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb935be0f),
	.w1(32'hb920fa38),
	.w2(32'hb8c80be4),
	.w3(32'hb7690d19),
	.w4(32'hb88dee13),
	.w5(32'h38807b77),
	.w6(32'h37d0fec9),
	.w7(32'hb822a059),
	.w8(32'h385a576c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8478cc2),
	.w1(32'hb7dd3bb7),
	.w2(32'hb84e6ff3),
	.w3(32'hb818f745),
	.w4(32'h379767e2),
	.w5(32'h37fdb614),
	.w6(32'hb8f6e6ed),
	.w7(32'hb8ce8079),
	.w8(32'hb89397ba),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38695908),
	.w1(32'h3980a422),
	.w2(32'hb929c73a),
	.w3(32'hb61ad7aa),
	.w4(32'h36fa93f5),
	.w5(32'hb9bb0162),
	.w6(32'hb978ebe0),
	.w7(32'hb957c032),
	.w8(32'hb9d84bd9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9783a1c),
	.w1(32'h3a188995),
	.w2(32'hb8aaae72),
	.w3(32'hb9c26639),
	.w4(32'hb8f6637b),
	.w5(32'hba04345d),
	.w6(32'hba675b87),
	.w7(32'hb977e8cb),
	.w8(32'hba24adea),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376fcd3c),
	.w1(32'h37467efc),
	.w2(32'hb688ab15),
	.w3(32'hb7c773e5),
	.w4(32'hb7972bd0),
	.w5(32'hb78e2fb0),
	.w6(32'hb846d5e9),
	.w7(32'hb81b89c8),
	.w8(32'hb7e994fd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65a8f97),
	.w1(32'hb608240c),
	.w2(32'hb4afbaf4),
	.w3(32'h34f0a18a),
	.w4(32'hb62bf0dc),
	.w5(32'hb491aff5),
	.w6(32'hb6ac8b22),
	.w7(32'hb32d0a4a),
	.w8(32'h35ed5287),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71b30f1),
	.w1(32'hb72570b2),
	.w2(32'hb886ce91),
	.w3(32'hb6e90b2d),
	.w4(32'hb81a62f2),
	.w5(32'hb83dc6d9),
	.w6(32'hb8160b1f),
	.w7(32'hb82bdf62),
	.w8(32'hb8882edb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a97b3c),
	.w1(32'h36016dfc),
	.w2(32'hb6e45a5d),
	.w3(32'hb6cb0e8c),
	.w4(32'hb680925e),
	.w5(32'hb70282af),
	.w6(32'hb6c7a7e1),
	.w7(32'hb68bf42c),
	.w8(32'hb6cfecb3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982dc56),
	.w1(32'h3aa604db),
	.w2(32'h3a62c118),
	.w3(32'hba2e7cf1),
	.w4(32'hb7a33651),
	.w5(32'hba5bdce6),
	.w6(32'hba52c0c2),
	.w7(32'hba8563dc),
	.w8(32'hbaeefa32),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88a963c),
	.w1(32'hb88303ed),
	.w2(32'hba429bfb),
	.w3(32'hb8d0b598),
	.w4(32'hb9362bbb),
	.w5(32'hba464793),
	.w6(32'hba093b0e),
	.w7(32'hb92c23d7),
	.w8(32'hb9b4eaa3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2180da),
	.w1(32'hb959fe0f),
	.w2(32'hba36a68d),
	.w3(32'hb9eaa03e),
	.w4(32'hba0719ed),
	.w5(32'hba442a26),
	.w6(32'hba312c22),
	.w7(32'hba12c2cd),
	.w8(32'hb9e52519),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ecd47c),
	.w1(32'h36cafa7c),
	.w2(32'h39548329),
	.w3(32'h39c44674),
	.w4(32'h392b3eb5),
	.w5(32'h3a35946a),
	.w6(32'h3a461c74),
	.w7(32'hb5fd70d2),
	.w8(32'h39b82d0f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5166afc),
	.w1(32'h341e664e),
	.w2(32'hb5daea56),
	.w3(32'hb4ac975b),
	.w4(32'h368a8c0a),
	.w5(32'hb658bda4),
	.w6(32'hb59899c1),
	.w7(32'h369c0d9e),
	.w8(32'h3475fac0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36181a55),
	.w1(32'h362b0747),
	.w2(32'hb721e694),
	.w3(32'h362f18cc),
	.w4(32'h365ab1ca),
	.w5(32'hb6a31d49),
	.w6(32'hb59c1b55),
	.w7(32'h362d8056),
	.w8(32'hb6d6afe8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3681c9f4),
	.w1(32'h372b10c7),
	.w2(32'hb7131f71),
	.w3(32'hb50ceb0f),
	.w4(32'hb4d7e3d6),
	.w5(32'hb78edbb9),
	.w6(32'h365d6bff),
	.w7(32'h37087d02),
	.w8(32'h36e26c9c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59d934d),
	.w1(32'h38f7becb),
	.w2(32'hb8a63a8f),
	.w3(32'hb780ff36),
	.w4(32'hb8279485),
	.w5(32'hb98c0463),
	.w6(32'hb7ca167e),
	.w7(32'hb695425b),
	.w8(32'hb91bf6d5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb797f012),
	.w1(32'hb82c8251),
	.w2(32'hb7d05b32),
	.w3(32'hb8880042),
	.w4(32'hb816149c),
	.w5(32'h37098b7c),
	.w6(32'hb79c0211),
	.w7(32'h37754a18),
	.w8(32'h365632c5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8764a3a),
	.w1(32'h3750435f),
	.w2(32'h39944557),
	.w3(32'hb9d0fa02),
	.w4(32'hb856596e),
	.w5(32'hb933a1d8),
	.w6(32'hb94881bf),
	.w7(32'hb95276ec),
	.w8(32'hba1d18a6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9407521),
	.w1(32'hb9ae165b),
	.w2(32'h3808d76b),
	.w3(32'hb9850537),
	.w4(32'hb94c9677),
	.w5(32'hb9f457d7),
	.w6(32'hb8d5e0ea),
	.w7(32'hb988e438),
	.w8(32'hba018e0e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ddc8f4),
	.w1(32'h39106392),
	.w2(32'h38cf3375),
	.w3(32'h37e89224),
	.w4(32'h3908ee66),
	.w5(32'h3997e643),
	.w6(32'hb8d4d841),
	.w7(32'hb866216f),
	.w8(32'h384df5e4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f6083b),
	.w1(32'h38e1b353),
	.w2(32'hb71908cd),
	.w3(32'hb8a8e304),
	.w4(32'hb5b77604),
	.w5(32'hb91c4fa6),
	.w6(32'hb97b1af9),
	.w7(32'h340efd86),
	.w8(32'hb91de173),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8804ca3),
	.w1(32'h399b39b9),
	.w2(32'h3a0c8e13),
	.w3(32'hb959557e),
	.w4(32'h3849f8d4),
	.w5(32'hb902b6e9),
	.w6(32'h37640999),
	.w7(32'hb9a077bc),
	.w8(32'hba534fc6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39960fc8),
	.w1(32'h399469eb),
	.w2(32'hb7af7873),
	.w3(32'h395b1bc4),
	.w4(32'h38ac25b3),
	.w5(32'hb818de6e),
	.w6(32'hb844cf91),
	.w7(32'hb901ff71),
	.w8(32'hb9b07048),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92981aa),
	.w1(32'h37b3c89f),
	.w2(32'h37db857e),
	.w3(32'hb92a281f),
	.w4(32'hb8e62624),
	.w5(32'hb96b9bac),
	.w6(32'hb8b1c130),
	.w7(32'hb9695fc2),
	.w8(32'hb9db832c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3698519c),
	.w1(32'h3644f02d),
	.w2(32'hb67ead63),
	.w3(32'h35ff87ea),
	.w4(32'hb5e52bc6),
	.w5(32'hb6ff5eef),
	.w6(32'h35e6dbc3),
	.w7(32'hb6b49b0b),
	.w8(32'hb7127af6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36568215),
	.w1(32'hb698f914),
	.w2(32'hb6d2c438),
	.w3(32'h35a8997b),
	.w4(32'hb6a1662c),
	.w5(32'hb5e1116f),
	.w6(32'hb69bcdba),
	.w7(32'hb6000b3e),
	.w8(32'h35ee12f3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b53390),
	.w1(32'h370c3412),
	.w2(32'hb557cb13),
	.w3(32'hb6865a2e),
	.w4(32'h36e54553),
	.w5(32'hb48684c0),
	.w6(32'h371e1294),
	.w7(32'h35d1bb4a),
	.w8(32'hb5b14adc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38785515),
	.w1(32'hb7e26b5c),
	.w2(32'h3811ad1b),
	.w3(32'h38bf4169),
	.w4(32'h385367a1),
	.w5(32'h38c306ab),
	.w6(32'h38bc5077),
	.w7(32'h380c09b7),
	.w8(32'h38c0ad0c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39736d6c),
	.w1(32'h383d9dc8),
	.w2(32'h3897a8fc),
	.w3(32'h39539d95),
	.w4(32'h39450644),
	.w5(32'h399d9789),
	.w6(32'h390da347),
	.w7(32'h38950125),
	.w8(32'h39a4e1c4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eabb59),
	.w1(32'h374fa024),
	.w2(32'h3841d53a),
	.w3(32'h3818a67c),
	.w4(32'h37c67e1f),
	.w5(32'h382b7c93),
	.w6(32'hb786e0ac),
	.w7(32'hb7590acc),
	.w8(32'h36b56820),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f44811),
	.w1(32'hb8afc606),
	.w2(32'hb992de4f),
	.w3(32'h3890763d),
	.w4(32'h38b579f0),
	.w5(32'hb801ffb8),
	.w6(32'h389ae2f4),
	.w7(32'hb8390f84),
	.w8(32'hb93a6571),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c81152),
	.w1(32'hb9b02fb8),
	.w2(32'hb930d91f),
	.w3(32'hb98f1d50),
	.w4(32'hb9b00a9c),
	.w5(32'hb9d0dcea),
	.w6(32'hb95bcf3f),
	.w7(32'hb966842a),
	.w8(32'hb9aec62a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998242b),
	.w1(32'h3892d932),
	.w2(32'h39c0afeb),
	.w3(32'h3a21bcc7),
	.w4(32'h39d9bdbf),
	.w5(32'h3a01a51f),
	.w6(32'h3a1b44b7),
	.w7(32'h39a0b5e3),
	.w8(32'h3984d610),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371823ca),
	.w1(32'h3a3564a0),
	.w2(32'h3a743d0d),
	.w3(32'hb8032120),
	.w4(32'h39dd14d1),
	.w5(32'hb90e9f23),
	.w6(32'hb7452789),
	.w7(32'hba681b3a),
	.w8(32'hba956730),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d2f2f),
	.w1(32'hb90f3a76),
	.w2(32'h398d1461),
	.w3(32'h394cd4dc),
	.w4(32'hb89db3f2),
	.w5(32'h39e56053),
	.w6(32'h39a9befb),
	.w7(32'hb7c5ed9f),
	.w8(32'h3928bcbc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995c7fe),
	.w1(32'h392f356f),
	.w2(32'hba3808fb),
	.w3(32'hb96f825e),
	.w4(32'h3569b8ae),
	.w5(32'hba26a90b),
	.w6(32'hba163016),
	.w7(32'hb9b073ae),
	.w8(32'hba134b96),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aadba8),
	.w1(32'h3a3f493f),
	.w2(32'h3991b7e5),
	.w3(32'h3937dc2f),
	.w4(32'h39b12907),
	.w5(32'hb8d9ab51),
	.w6(32'h3831743d),
	.w7(32'hb854bc74),
	.w8(32'hb9914880),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3970428d),
	.w1(32'hb962ee55),
	.w2(32'h38d148a4),
	.w3(32'h39c04a9e),
	.w4(32'h38f011a6),
	.w5(32'h39319cb7),
	.w6(32'h39dcc621),
	.w7(32'hb5b1fd6c),
	.w8(32'h39108aa3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba072eb9),
	.w1(32'hb9e2b963),
	.w2(32'hb9ebd7b6),
	.w3(32'hba146d28),
	.w4(32'hb9b2cd7e),
	.w5(32'hba3c9848),
	.w6(32'hb9965696),
	.w7(32'hb9f5aa37),
	.w8(32'hb9defc12),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba455228),
	.w1(32'hb8558f81),
	.w2(32'h38e19f8a),
	.w3(32'hba1b870e),
	.w4(32'h392b8a69),
	.w5(32'hb93659d9),
	.w6(32'hba1d8a28),
	.w7(32'h39b38fd5),
	.w8(32'h39105e2a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943df43),
	.w1(32'h39fee762),
	.w2(32'h3aab89fc),
	.w3(32'hba2b3839),
	.w4(32'h38ca5805),
	.w5(32'h3a0dace8),
	.w6(32'h382548be),
	.w7(32'h39c6bf1d),
	.w8(32'h3980d099),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3892c358),
	.w1(32'hb96831c2),
	.w2(32'hba2efab4),
	.w3(32'hb82e42e0),
	.w4(32'hb69f4c0d),
	.w5(32'hba84fbc4),
	.w6(32'h38cc515d),
	.w7(32'hba99f90e),
	.w8(32'hb9f51481),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a809b21),
	.w1(32'hbaad03c3),
	.w2(32'hb95e2c76),
	.w3(32'h39fb6014),
	.w4(32'hba4e2c38),
	.w5(32'h3a263e7e),
	.w6(32'h39a9be6f),
	.w7(32'hba2a8149),
	.w8(32'h3a6a169b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ff7b2),
	.w1(32'h3990e1ab),
	.w2(32'h385469b6),
	.w3(32'hb8a1f50c),
	.w4(32'h39d74a1e),
	.w5(32'h39df15ea),
	.w6(32'h390f8ef3),
	.w7(32'h37803127),
	.w8(32'h38c5a446),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3869840f),
	.w1(32'h39433bd7),
	.w2(32'h3a601043),
	.w3(32'hba266395),
	.w4(32'h3964b05e),
	.w5(32'hb902eef1),
	.w6(32'hb9959493),
	.w7(32'hba8851bc),
	.w8(32'hba451817),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4953f),
	.w1(32'hba92af79),
	.w2(32'hb981d74e),
	.w3(32'hbae3b26f),
	.w4(32'hba866a55),
	.w5(32'hba89e3bd),
	.w6(32'hbaa38bc3),
	.w7(32'hbab3029b),
	.w8(32'hb99bfe23),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd928e),
	.w1(32'hba4aaf76),
	.w2(32'hb9e224d0),
	.w3(32'hb9160e05),
	.w4(32'hb961b083),
	.w5(32'hba536df1),
	.w6(32'h3a32b3f8),
	.w7(32'hba22a13a),
	.w8(32'hba72c06c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c63d2f),
	.w1(32'hb994f0b4),
	.w2(32'h382c44a5),
	.w3(32'hb90d9d3e),
	.w4(32'hba0762f9),
	.w5(32'hb9f0b04a),
	.w6(32'h38fdd022),
	.w7(32'hba04141f),
	.w8(32'hba2418a1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb892625e),
	.w1(32'hb745a76f),
	.w2(32'h37d35ad1),
	.w3(32'hb6603517),
	.w4(32'hb5f89537),
	.w5(32'h37c10541),
	.w6(32'h3687096f),
	.w7(32'h3716e811),
	.w8(32'h380fb9b9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a1930),
	.w1(32'h39a89a07),
	.w2(32'hb8813dd1),
	.w3(32'h39a4cf60),
	.w4(32'h39b5cdc7),
	.w5(32'h38d34b92),
	.w6(32'h369fe722),
	.w7(32'h37ea2afa),
	.w8(32'h380f5c1c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a2606),
	.w1(32'hba05908a),
	.w2(32'hb8ce0287),
	.w3(32'hba4bac4c),
	.w4(32'hba2f23d3),
	.w5(32'hb9de2f52),
	.w6(32'hb9ee4cda),
	.w7(32'hba0fe8c0),
	.w8(32'hb9ecc9ba),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac0216),
	.w1(32'h3a2e57d5),
	.w2(32'h3a62cf6c),
	.w3(32'h3950ae23),
	.w4(32'h3a32ab60),
	.w5(32'h3a7a2eb7),
	.w6(32'h39a40a9c),
	.w7(32'h3a235081),
	.w8(32'h3a8a3dfb),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b07029),
	.w1(32'h3979edf9),
	.w2(32'h399c1d5c),
	.w3(32'h39f271a6),
	.w4(32'h3963a569),
	.w5(32'h39f6aae5),
	.w6(32'h398be9d2),
	.w7(32'h38483c3c),
	.w8(32'h3975a578),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e605e7),
	.w1(32'hb9bf1b03),
	.w2(32'hb966d8ec),
	.w3(32'h38a4b483),
	.w4(32'h37d311bf),
	.w5(32'h39b2e781),
	.w6(32'hb90695d3),
	.w7(32'hb9313f9f),
	.w8(32'h390453f7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a0b988),
	.w1(32'hb9a9bfc1),
	.w2(32'hb98a44b9),
	.w3(32'h3a0a4349),
	.w4(32'h38c814c6),
	.w5(32'h38a79782),
	.w6(32'hb83dc3f0),
	.w7(32'hb9a8502a),
	.w8(32'hb8dcc0a2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca4f53),
	.w1(32'h3a862cfc),
	.w2(32'hb69f748b),
	.w3(32'h39bd9095),
	.w4(32'h3a1a0912),
	.w5(32'hb780324a),
	.w6(32'hb9677d69),
	.w7(32'h388e8761),
	.w8(32'hb911aeab),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395c2276),
	.w1(32'h38eae18c),
	.w2(32'h393bbea4),
	.w3(32'h39610ea6),
	.w4(32'h396a5a5a),
	.w5(32'h399fc805),
	.w6(32'h390bd96f),
	.w7(32'h39229a0b),
	.w8(32'h3986bd1c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bf18af),
	.w1(32'h3741622a),
	.w2(32'hb741c468),
	.w3(32'h385f88db),
	.w4(32'hb5d58c13),
	.w5(32'hb5b6d5a8),
	.w6(32'h3624ee0f),
	.w7(32'hb837adf5),
	.w8(32'hb727caeb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78aa7b4),
	.w1(32'hb8a5088c),
	.w2(32'hb90d70a8),
	.w3(32'h3516d98f),
	.w4(32'hb88e3617),
	.w5(32'hb8f50f87),
	.w6(32'hb5c648bf),
	.w7(32'hb7ed6f37),
	.w8(32'hb8946f6b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b392d8),
	.w1(32'hb55d17ef),
	.w2(32'h35942f58),
	.w3(32'h350fc5d6),
	.w4(32'h34215617),
	.w5(32'hb6c48f41),
	.w6(32'hb47f3fb4),
	.w7(32'hb53a9e99),
	.w8(32'hb6bb9da9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379cc0b1),
	.w1(32'hb7948b8d),
	.w2(32'hb6793b25),
	.w3(32'h37c2ec9c),
	.w4(32'hb6d62499),
	.w5(32'hb67cd9ae),
	.w6(32'h3774cc23),
	.w7(32'hb80ee096),
	.w8(32'h379922de),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9347726),
	.w1(32'hb9c77c86),
	.w2(32'hb9e72911),
	.w3(32'hb94ada9d),
	.w4(32'hb9d4a053),
	.w5(32'hb993a986),
	.w6(32'hb996ce11),
	.w7(32'hb9ba8ee8),
	.w8(32'hb9cefaf4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3897c716),
	.w1(32'hb733f563),
	.w2(32'h380eb237),
	.w3(32'h37f86c74),
	.w4(32'hb8a99c0a),
	.w5(32'h37989db5),
	.w6(32'hb88673e2),
	.w7(32'hb93f5922),
	.w8(32'hb81c828f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3811fe0b),
	.w1(32'h386cb6c1),
	.w2(32'h393f05d6),
	.w3(32'hb91fd06f),
	.w4(32'hb82a9d52),
	.w5(32'hb8f126b3),
	.w6(32'hb8c6ff37),
	.w7(32'hb98f0daa),
	.w8(32'hb9e79817),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39717518),
	.w1(32'hb8ac2691),
	.w2(32'h38bfcd8f),
	.w3(32'h3961642d),
	.w4(32'h38e5e6ed),
	.w5(32'h3998aebe),
	.w6(32'h3982979d),
	.w7(32'h36386941),
	.w8(32'h39576a30),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6aed919),
	.w1(32'hb63928ad),
	.w2(32'hb6ecc513),
	.w3(32'hb6cb19ae),
	.w4(32'hb64ac717),
	.w5(32'hb6772120),
	.w6(32'hb70cf322),
	.w7(32'hb6bad234),
	.w8(32'hb7156cae),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380da0a6),
	.w1(32'h378099a3),
	.w2(32'h382df760),
	.w3(32'h376f3305),
	.w4(32'h3734e002),
	.w5(32'h3807c973),
	.w6(32'h378bed34),
	.w7(32'h374044a0),
	.w8(32'h37d11932),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3747dac3),
	.w1(32'h37033ed5),
	.w2(32'hb6559d0c),
	.w3(32'hb5ee7b62),
	.w4(32'h357df9ae),
	.w5(32'hb720f2f4),
	.w6(32'h36b9604c),
	.w7(32'h365cfbc3),
	.w8(32'hb7acd32c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74cd20e),
	.w1(32'hb9e552b9),
	.w2(32'hb9ca3027),
	.w3(32'hb66c9dd9),
	.w4(32'hb9aed2c9),
	.w5(32'hb9e2fb8f),
	.w6(32'hb9848cfe),
	.w7(32'h39697e07),
	.w8(32'h385add08),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38af2acf),
	.w1(32'h39aee445),
	.w2(32'hb9472e17),
	.w3(32'h3a4d8de2),
	.w4(32'h39d8c3d1),
	.w5(32'hb9a45438),
	.w6(32'h395850b9),
	.w7(32'hb96093cd),
	.w8(32'hb93661bb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e7e19f),
	.w1(32'h38661749),
	.w2(32'h3925c2bd),
	.w3(32'hba009444),
	.w4(32'hb9dbf87b),
	.w5(32'hba871446),
	.w6(32'hba0552d8),
	.w7(32'hba375049),
	.w8(32'hba3b2a5d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39453761),
	.w1(32'h396cb1ca),
	.w2(32'h3962e0ec),
	.w3(32'hb93350ca),
	.w4(32'h383df385),
	.w5(32'hb9059b7b),
	.w6(32'h3981d3fb),
	.w7(32'hb9283c6b),
	.w8(32'hb8fcc91d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b68903),
	.w1(32'hb98b01f5),
	.w2(32'hb858bdfc),
	.w3(32'hba0abbec),
	.w4(32'hb94037cd),
	.w5(32'hb9fc38b9),
	.w6(32'hb98e2cea),
	.w7(32'hba0f9d16),
	.w8(32'hba1287c6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b0e37),
	.w1(32'h3aec896b),
	.w2(32'h3a3794e2),
	.w3(32'hba18074f),
	.w4(32'h380aa22e),
	.w5(32'hb84ffb1d),
	.w6(32'hb8cd10c9),
	.w7(32'hba13c730),
	.w8(32'hb9f6c7b4),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80f98c),
	.w1(32'hb9f527a2),
	.w2(32'hba8ed917),
	.w3(32'hb9a9f2c6),
	.w4(32'hb999f3f5),
	.w5(32'hba704ebb),
	.w6(32'hba2ff650),
	.w7(32'hba69dda0),
	.w8(32'hbac40757),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ebb6c),
	.w1(32'h397aa887),
	.w2(32'hb9e297cb),
	.w3(32'hb949befc),
	.w4(32'hba160975),
	.w5(32'hba94e579),
	.w6(32'hb85d954c),
	.w7(32'hb9b684a2),
	.w8(32'hb9a9661c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b78199),
	.w1(32'h3a37649f),
	.w2(32'h3a088529),
	.w3(32'hbab42510),
	.w4(32'hb9155b93),
	.w5(32'hba0e074c),
	.w6(32'hb985940b),
	.w7(32'hba1ed885),
	.w8(32'hbab0b8cb),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b059b8),
	.w1(32'hb98ed895),
	.w2(32'hb9681d21),
	.w3(32'hba42c3fa),
	.w4(32'hba0e5045),
	.w5(32'hb9a083ed),
	.w6(32'h387aacac),
	.w7(32'hb989a00d),
	.w8(32'hb8d4f203),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0808fd),
	.w1(32'h39d110ba),
	.w2(32'h3a08e1e3),
	.w3(32'hba3815ae),
	.w4(32'h391e6e98),
	.w5(32'hb86a903e),
	.w6(32'hb97478e4),
	.w7(32'hb7ebd3dc),
	.w8(32'h39136988),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4f84e),
	.w1(32'h3a5ab6eb),
	.w2(32'h399ec6a9),
	.w3(32'hba006ef5),
	.w4(32'h3a3e1ad6),
	.w5(32'hb9353d71),
	.w6(32'h3a74ae89),
	.w7(32'h38a41847),
	.w8(32'h397eef45),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bebd0),
	.w1(32'h3a09dca0),
	.w2(32'h3a3cd6b4),
	.w3(32'h3a3acc68),
	.w4(32'h396c13a5),
	.w5(32'h394fcda2),
	.w6(32'hb92780fd),
	.w7(32'hb91bf445),
	.w8(32'h39507f57),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a3d9b),
	.w1(32'h37d28bf0),
	.w2(32'hb94bbcc0),
	.w3(32'hba025b58),
	.w4(32'hba3f2696),
	.w5(32'hb9b78aec),
	.w6(32'h3a2b6030),
	.w7(32'h39a6449d),
	.w8(32'hb8c7cfb1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee79d4),
	.w1(32'hb9aea040),
	.w2(32'h3605442b),
	.w3(32'hb919588b),
	.w4(32'hb9fda293),
	.w5(32'hb9d7625d),
	.w6(32'hb90e56ee),
	.w7(32'hb906ca4c),
	.w8(32'hb866d08f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c07196),
	.w1(32'hb9fc29bd),
	.w2(32'hba2d1b55),
	.w3(32'h3a04902b),
	.w4(32'hb9be38cf),
	.w5(32'hb97c4325),
	.w6(32'h39d1f83c),
	.w7(32'hb93fcaee),
	.w8(32'hb8a07d7b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10f56f),
	.w1(32'h39958d7b),
	.w2(32'hba043c18),
	.w3(32'hb9fb0879),
	.w4(32'hba0788ed),
	.w5(32'h38e7b2f7),
	.w6(32'h38c7dd04),
	.w7(32'hb9d76433),
	.w8(32'hb9c75933),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86fd2fa),
	.w1(32'h394cd409),
	.w2(32'h39cea8f2),
	.w3(32'h39f1353b),
	.w4(32'hb8a58e4e),
	.w5(32'hb9894bef),
	.w6(32'h390517b7),
	.w7(32'h39bf3bf4),
	.w8(32'h393259a4),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905de01),
	.w1(32'hba2273d0),
	.w2(32'hba00f9f6),
	.w3(32'hb9fac5e3),
	.w4(32'hb7798425),
	.w5(32'h38e3a9ea),
	.w6(32'hb7d59238),
	.w7(32'hb9393f9e),
	.w8(32'h398d4d2f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba362390),
	.w1(32'h39efe27b),
	.w2(32'h3a1216f0),
	.w3(32'h39c32335),
	.w4(32'h3a325cf0),
	.w5(32'h39b6a7d1),
	.w6(32'h3a15a3e1),
	.w7(32'h3988920c),
	.w8(32'h3954ea0a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d619a),
	.w1(32'h392364b4),
	.w2(32'h39967410),
	.w3(32'h3a0cef7e),
	.w4(32'h39acf7d2),
	.w5(32'h38e33935),
	.w6(32'h39ac996d),
	.w7(32'hb893312d),
	.w8(32'h39169c3c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9571c),
	.w1(32'h39dbb3bf),
	.w2(32'h3a20b475),
	.w3(32'hba19afe3),
	.w4(32'h38de4ccb),
	.w5(32'h383a50dd),
	.w6(32'hb55f8bed),
	.w7(32'h39ca0a61),
	.w8(32'h39295323),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c02d5e),
	.w1(32'hba18c923),
	.w2(32'hba207995),
	.w3(32'h38696dca),
	.w4(32'hba24e7c9),
	.w5(32'hb9fc879b),
	.w6(32'hb9133329),
	.w7(32'hb9dc76d7),
	.w8(32'hb9a1692e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05881b),
	.w1(32'h3a9151e9),
	.w2(32'h3b170cf8),
	.w3(32'hba3fe33e),
	.w4(32'hbab8c699),
	.w5(32'hbabba59c),
	.w6(32'hb985c6ca),
	.w7(32'hba7adfc8),
	.w8(32'h38a8c043),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abf608),
	.w1(32'h39d88443),
	.w2(32'h3a28c7ec),
	.w3(32'hba5642bf),
	.w4(32'h39d47fd8),
	.w5(32'h39add66c),
	.w6(32'hb9b6f35e),
	.w7(32'hb790f772),
	.w8(32'hb98710ca),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84a89d),
	.w1(32'h39ffd082),
	.w2(32'h3a4260b6),
	.w3(32'h3a164fe1),
	.w4(32'hb80c7982),
	.w5(32'hb8bd4ded),
	.w6(32'h3919dbf3),
	.w7(32'hb9970d06),
	.w8(32'hb9c45dc6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e52cff),
	.w1(32'h3a1114dc),
	.w2(32'h39d369c9),
	.w3(32'hb6242897),
	.w4(32'h3767b307),
	.w5(32'h383d2306),
	.w6(32'hb8fbad4b),
	.w7(32'h39cc077d),
	.w8(32'hb95448fe),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ada76b),
	.w1(32'h3a589314),
	.w2(32'h3a5c49d7),
	.w3(32'h394cee79),
	.w4(32'hba34e29a),
	.w5(32'hba77f18f),
	.w6(32'h3ac61174),
	.w7(32'h3b16691e),
	.w8(32'h3ae6e4c4),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83bfac),
	.w1(32'hba482968),
	.w2(32'h3882b3ed),
	.w3(32'hbaf1768a),
	.w4(32'hba9847db),
	.w5(32'hba28a0ee),
	.w6(32'hbaa70f8c),
	.w7(32'hba37efaa),
	.w8(32'hb950e065),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7a29d),
	.w1(32'h3a6ccc6b),
	.w2(32'h3b0030e0),
	.w3(32'h3a97fd19),
	.w4(32'h3a331922),
	.w5(32'h3a640068),
	.w6(32'h388d26f2),
	.w7(32'h3963390a),
	.w8(32'h3a966c22),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a602b8c),
	.w1(32'hba3c2e77),
	.w2(32'hba60e0b2),
	.w3(32'h39754a18),
	.w4(32'hb968c57b),
	.w5(32'hb8a8e3bc),
	.w6(32'hba7cb985),
	.w7(32'hbaa81fd7),
	.w8(32'hb9a26a59),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b104c8),
	.w1(32'hba05be3f),
	.w2(32'hba455403),
	.w3(32'h39b7de2e),
	.w4(32'h39971143),
	.w5(32'hb917cd91),
	.w6(32'hb9cca2d3),
	.w7(32'hba721e9b),
	.w8(32'hb939bc6d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d46ce),
	.w1(32'hb9e71d9f),
	.w2(32'hb96856cb),
	.w3(32'hb8fc0f65),
	.w4(32'hb94f3d04),
	.w5(32'hb906cfed),
	.w6(32'hb96165ff),
	.w7(32'hba09cb7e),
	.w8(32'hba0e57b3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9802073),
	.w1(32'h38d0cdc0),
	.w2(32'h39a7744e),
	.w3(32'hb9362fa4),
	.w4(32'hb8db4f47),
	.w5(32'hb90c975f),
	.w6(32'h39650c36),
	.w7(32'h3995e7e1),
	.w8(32'h39458a91),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91938b9),
	.w1(32'h3a9cd7e0),
	.w2(32'h39f782fc),
	.w3(32'hb9e5cfba),
	.w4(32'h3a12bf43),
	.w5(32'hba26d0e6),
	.w6(32'h3a96b048),
	.w7(32'h3a479f11),
	.w8(32'h3a3ef3e1),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfdc9a),
	.w1(32'hb98ebb5f),
	.w2(32'h3aa2547e),
	.w3(32'h3a08c271),
	.w4(32'hb9fdc497),
	.w5(32'h394d717c),
	.w6(32'hb9186c81),
	.w7(32'h3ad0a393),
	.w8(32'h3ab150d5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd03f4),
	.w1(32'hb998f12a),
	.w2(32'hb96faa82),
	.w3(32'h3a7295fe),
	.w4(32'hb8451535),
	.w5(32'hb94ea838),
	.w6(32'hb66ecf3f),
	.w7(32'hb9439aac),
	.w8(32'h390c9019),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39230a17),
	.w1(32'h3a034fcc),
	.w2(32'h39f646d4),
	.w3(32'hb8d93352),
	.w4(32'h3752ede4),
	.w5(32'h3826bafd),
	.w6(32'h3a10e0a9),
	.w7(32'h3a0cb3b6),
	.w8(32'h39f82ed1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb807886b),
	.w1(32'hb95ad7b8),
	.w2(32'hb9e66ab2),
	.w3(32'hb9120a37),
	.w4(32'hb8a96e56),
	.w5(32'hb9ed64bf),
	.w6(32'hb9b74455),
	.w7(32'hba55f1c8),
	.w8(32'hba39c745),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8095ed),
	.w1(32'h38a438fb),
	.w2(32'h386170e2),
	.w3(32'hba466e77),
	.w4(32'h389259ae),
	.w5(32'hb8b6ab10),
	.w6(32'h39798fb2),
	.w7(32'hb9359cdc),
	.w8(32'hb9015502),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eba7aa),
	.w1(32'hb9a60e16),
	.w2(32'hb94b4ce4),
	.w3(32'hba134de7),
	.w4(32'hba21aeb9),
	.w5(32'hba17db7d),
	.w6(32'hb92fc706),
	.w7(32'hb98edd80),
	.w8(32'hb994299c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370a1fa2),
	.w1(32'hb9edbac5),
	.w2(32'hb94439e0),
	.w3(32'hba20d1d6),
	.w4(32'hb95833d6),
	.w5(32'hb920ce14),
	.w6(32'hb904f995),
	.w7(32'hba50e428),
	.w8(32'hb9cefbac),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9494c5e),
	.w1(32'hba175d32),
	.w2(32'hba3ce335),
	.w3(32'hba135af6),
	.w4(32'hb8204c89),
	.w5(32'h372bdd8f),
	.w6(32'hb9c10e53),
	.w7(32'hba5bd846),
	.w8(32'hba03e7af),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ac031),
	.w1(32'h37d600b6),
	.w2(32'hb8176cd8),
	.w3(32'hb9b905db),
	.w4(32'hba084624),
	.w5(32'hb994cfe4),
	.w6(32'hb99c3f71),
	.w7(32'hba02c98b),
	.w8(32'hba11c331),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1949f9),
	.w1(32'hba17223c),
	.w2(32'hba104462),
	.w3(32'hba134770),
	.w4(32'hba09dd8b),
	.w5(32'hb97e8641),
	.w6(32'h38fedf19),
	.w7(32'h37cb4638),
	.w8(32'h38fbb266),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9541754),
	.w1(32'h3ab44edb),
	.w2(32'h3a1df1f3),
	.w3(32'hba0ab714),
	.w4(32'h3aac9f3a),
	.w5(32'h3a25585f),
	.w6(32'h3a8918c8),
	.w7(32'h3a01bb16),
	.w8(32'h3a847975),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a956f60),
	.w1(32'h3a940914),
	.w2(32'hb8e8bae7),
	.w3(32'h3a8ec62c),
	.w4(32'h3880147c),
	.w5(32'hbab9062c),
	.w6(32'hba2085e1),
	.w7(32'hba723c73),
	.w8(32'hb9cdd3be),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b88be6),
	.w1(32'h3971f78f),
	.w2(32'h3a6bff4a),
	.w3(32'hb9c566ed),
	.w4(32'hb951fa11),
	.w5(32'hb9fb4753),
	.w6(32'hb9904a15),
	.w7(32'hb9069ff2),
	.w8(32'h39a940d0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3920aea6),
	.w1(32'h398ee9b7),
	.w2(32'hb9f5dc09),
	.w3(32'hba514853),
	.w4(32'hba200a61),
	.w5(32'h39d3bba6),
	.w6(32'hb9aad62c),
	.w7(32'hb9e0c6de),
	.w8(32'hba7a4cdd),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff3a5f),
	.w1(32'hba3b1ce6),
	.w2(32'hb9d2ef60),
	.w3(32'hb967e81b),
	.w4(32'hb90a791a),
	.w5(32'hb9cc954f),
	.w6(32'hbabb1e03),
	.w7(32'hbaa307cc),
	.w8(32'hb9ea0991),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d003d),
	.w1(32'h3a74e0cc),
	.w2(32'h3a08b7f9),
	.w3(32'h3a90c452),
	.w4(32'h396ba189),
	.w5(32'hb88cd2a5),
	.w6(32'h39c7a0d7),
	.w7(32'h399ebf20),
	.w8(32'h3962c9d6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997492b),
	.w1(32'hb9a8a65f),
	.w2(32'hb9d29bd1),
	.w3(32'hb9ae2a37),
	.w4(32'hba1b9636),
	.w5(32'hb9f7db57),
	.w6(32'hb98abdd3),
	.w7(32'hb9f17102),
	.w8(32'hb9d92e75),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef0ea7),
	.w1(32'h392cba98),
	.w2(32'h3a0523ee),
	.w3(32'hb9e8e4ca),
	.w4(32'h395a24a1),
	.w5(32'h38ed0bfd),
	.w6(32'h39c512b0),
	.w7(32'h3a11a83c),
	.w8(32'h3a05c08f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f1a7eb),
	.w1(32'h3a8e58ae),
	.w2(32'h3af3a549),
	.w3(32'hb9369e3e),
	.w4(32'h389eb2a0),
	.w5(32'hbaa71d83),
	.w6(32'h399508e7),
	.w7(32'h3aab3c84),
	.w8(32'h38e7cc53),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9134473),
	.w1(32'h3a3cdf8b),
	.w2(32'h3a4afcca),
	.w3(32'hba62851c),
	.w4(32'hb91466d9),
	.w5(32'hba0f9ffc),
	.w6(32'h393eb551),
	.w7(32'h3928b83e),
	.w8(32'h38a15866),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e82f5),
	.w1(32'h394be518),
	.w2(32'hba38f624),
	.w3(32'hba6bfea9),
	.w4(32'h38f81e97),
	.w5(32'hba1df928),
	.w6(32'h3a05e984),
	.w7(32'hb963e5ac),
	.w8(32'hb9b988ce),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d16b28),
	.w1(32'h39b77198),
	.w2(32'h394f4501),
	.w3(32'hb8be3ede),
	.w4(32'h38c680e0),
	.w5(32'hb77b6134),
	.w6(32'h3a201c29),
	.w7(32'h3a031c89),
	.w8(32'h39ef45da),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a15bdc),
	.w1(32'h397312ad),
	.w2(32'h39156d3d),
	.w3(32'hb8972e0a),
	.w4(32'h3a5487c0),
	.w5(32'h3a7a474f),
	.w6(32'hb9aec7e5),
	.w7(32'hb991e75f),
	.w8(32'hb98ced33),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d167ce),
	.w1(32'h396a1f1e),
	.w2(32'h3a01bd30),
	.w3(32'h3a87f56d),
	.w4(32'h39de69b6),
	.w5(32'h39c81258),
	.w6(32'h38afd413),
	.w7(32'hb7557738),
	.w8(32'h37ea6807),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81a44c6),
	.w1(32'hb94bb92c),
	.w2(32'h39e833c1),
	.w3(32'hb89c0375),
	.w4(32'hba08f624),
	.w5(32'hb9cf06c3),
	.w6(32'h3a968f8a),
	.w7(32'h3a9f3a90),
	.w8(32'hba0a0b0b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39244aaa),
	.w1(32'h38f76f29),
	.w2(32'hb8faa9b9),
	.w3(32'hb9368d86),
	.w4(32'h37d30a4a),
	.w5(32'hb9e580d4),
	.w6(32'h398efedf),
	.w7(32'hb994b363),
	.w8(32'hb9988c72),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdaaf4),
	.w1(32'h39ff07d3),
	.w2(32'h39d06486),
	.w3(32'hba20ed74),
	.w4(32'hb9ee965b),
	.w5(32'hba84e804),
	.w6(32'hba088d7d),
	.w7(32'hba0604e7),
	.w8(32'hba28d7a5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24c131),
	.w1(32'h3aa5014c),
	.w2(32'h3a910de6),
	.w3(32'hb900abfc),
	.w4(32'h3a0a100a),
	.w5(32'h39abd2ab),
	.w6(32'h37868f57),
	.w7(32'hb9c8c42d),
	.w8(32'hb9555332),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40a858),
	.w1(32'hba39c6ed),
	.w2(32'hb9b8a435),
	.w3(32'hba98898d),
	.w4(32'hba4f08ed),
	.w5(32'hba6c481d),
	.w6(32'hba85c70a),
	.w7(32'hbac29a85),
	.w8(32'hbabc84be),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b4ee1),
	.w1(32'h3a91cdb2),
	.w2(32'h377123e9),
	.w3(32'hba221ef2),
	.w4(32'hb807f1aa),
	.w5(32'hba422793),
	.w6(32'h3aa4fb66),
	.w7(32'h3abb86dd),
	.w8(32'h3a8ac5d3),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8ec46),
	.w1(32'h3a67a5a5),
	.w2(32'h39d6a6d4),
	.w3(32'h38699053),
	.w4(32'h3a5f301f),
	.w5(32'h39df295a),
	.w6(32'h3a5a85e0),
	.w7(32'h39f49fd6),
	.w8(32'h3a8fcc81),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33e730),
	.w1(32'h396515d8),
	.w2(32'h39902ecb),
	.w3(32'h3a35e78b),
	.w4(32'hb777cc3f),
	.w5(32'hb8c49cb7),
	.w6(32'h390d5677),
	.w7(32'h3983cbe8),
	.w8(32'h39cfe85f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3972b1ab),
	.w1(32'h39b495fa),
	.w2(32'h3a3730c5),
	.w3(32'hb9705707),
	.w4(32'hb9a594af),
	.w5(32'hba5af212),
	.w6(32'h3a0cb60f),
	.w7(32'h3a61ca6b),
	.w8(32'hb910d535),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb909aec2),
	.w1(32'h3901354e),
	.w2(32'hb8a9d13b),
	.w3(32'hb9fec4b2),
	.w4(32'h39f75ebd),
	.w5(32'h398b2aea),
	.w6(32'hb8a0707d),
	.w7(32'hb9c8ef34),
	.w8(32'hba135d80),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e8903),
	.w1(32'h393c3cba),
	.w2(32'h38a98a17),
	.w3(32'h39d51b54),
	.w4(32'h38df6c32),
	.w5(32'hb8147c67),
	.w6(32'hb7d5d15b),
	.w7(32'h38d35bf9),
	.w8(32'hba0b9929),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a80d64),
	.w1(32'h38cafb36),
	.w2(32'h39933fed),
	.w3(32'hb93ca1e8),
	.w4(32'hb9951874),
	.w5(32'hb9cddda3),
	.w6(32'h3986173e),
	.w7(32'h39412352),
	.w8(32'h38eb8fa7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba172d90),
	.w1(32'h39dd377d),
	.w2(32'h3a6883b6),
	.w3(32'hba5def77),
	.w4(32'hb7bc1ee3),
	.w5(32'h3995e8d6),
	.w6(32'h39aa6f01),
	.w7(32'h39fb937b),
	.w8(32'h3948b764),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a300c43),
	.w1(32'h389f9cbc),
	.w2(32'h382b4399),
	.w3(32'h39a64121),
	.w4(32'h39bef732),
	.w5(32'hb71b8788),
	.w6(32'h3a1b4be1),
	.w7(32'h395762fd),
	.w8(32'hb7e6b3f1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9407653),
	.w1(32'hb97bd1cc),
	.w2(32'hb89c6e8b),
	.w3(32'hb930172c),
	.w4(32'hba0386e8),
	.w5(32'hb9667c46),
	.w6(32'hb88be698),
	.w7(32'hb8969c33),
	.w8(32'hb8b78d1f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb683afd7),
	.w1(32'hb733dc10),
	.w2(32'hba21fa98),
	.w3(32'hb9e92514),
	.w4(32'hb9c61a46),
	.w5(32'hba657578),
	.w6(32'hb8c177d9),
	.w7(32'hb9083931),
	.w8(32'hba082210),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd3d50),
	.w1(32'hb81ff4be),
	.w2(32'h397a6963),
	.w3(32'hba0fe1dd),
	.w4(32'hb9313982),
	.w5(32'hb97cdcae),
	.w6(32'h3974c8f9),
	.w7(32'h395a39a4),
	.w8(32'h3917adc3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80ed847),
	.w1(32'hb81aef96),
	.w2(32'h38c04a87),
	.w3(32'hba088412),
	.w4(32'hb98b8d7a),
	.w5(32'hba52c464),
	.w6(32'hb9ec3672),
	.w7(32'hba0a03d8),
	.w8(32'hba1dd170),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9362170),
	.w1(32'h3ad13ffe),
	.w2(32'hb97bbb24),
	.w3(32'hb885a586),
	.w4(32'hba5a08d7),
	.w5(32'hba335cc4),
	.w6(32'h3b35f635),
	.w7(32'h3b079333),
	.w8(32'h3a55f4f8),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e9c64),
	.w1(32'hb79a5e24),
	.w2(32'hb978299c),
	.w3(32'hb9c5f286),
	.w4(32'hb9ce665f),
	.w5(32'hb9b12f92),
	.w6(32'hb79e302b),
	.w7(32'hb98740d3),
	.w8(32'hb7bf569e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9412bb1),
	.w1(32'h39933bd7),
	.w2(32'hb9b7ff75),
	.w3(32'hb9868f01),
	.w4(32'h38d1aa11),
	.w5(32'hba1c21fc),
	.w6(32'h3a02a099),
	.w7(32'hb987f3cc),
	.w8(32'hb9c5c444),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6e833),
	.w1(32'h39eabe14),
	.w2(32'hba238330),
	.w3(32'hba14b521),
	.w4(32'hba1aea22),
	.w5(32'hbaa7ff31),
	.w6(32'h3a882ad5),
	.w7(32'h3a954fb2),
	.w8(32'h3a00b5d1),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9acb49d),
	.w1(32'hb94356eb),
	.w2(32'hb98b6924),
	.w3(32'hba863bdf),
	.w4(32'hb9336a96),
	.w5(32'hb97dd932),
	.w6(32'hb9b98480),
	.w7(32'hb9fa6a96),
	.w8(32'hba2982dd),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c9e2e),
	.w1(32'hb90e8f09),
	.w2(32'hb881f8bc),
	.w3(32'hb8bf0876),
	.w4(32'h39d7176e),
	.w5(32'h3a51abff),
	.w6(32'hb972ab76),
	.w7(32'hb98bbe79),
	.w8(32'hba44c99f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09002e),
	.w1(32'hb8d1260d),
	.w2(32'h3a00a4dd),
	.w3(32'h38f8a512),
	.w4(32'hb9959bc8),
	.w5(32'hb9012f95),
	.w6(32'h38c959c3),
	.w7(32'hb9aced9f),
	.w8(32'hb99c06c8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e93642),
	.w1(32'hb99e16bb),
	.w2(32'hb957ceaa),
	.w3(32'hba1fd364),
	.w4(32'h3766530e),
	.w5(32'h383d980d),
	.w6(32'hb9c9639c),
	.w7(32'hb9e3275c),
	.w8(32'hb9463915),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f00479),
	.w1(32'hb92e0b48),
	.w2(32'h3985fe7f),
	.w3(32'h39f4bb1b),
	.w4(32'h38d30ef3),
	.w5(32'hb9cda562),
	.w6(32'h39eda978),
	.w7(32'hb9b4d819),
	.w8(32'hb9a87324),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebe45a),
	.w1(32'hb9fa24c5),
	.w2(32'hb9c4eba1),
	.w3(32'hba507ec6),
	.w4(32'hb9d78882),
	.w5(32'hb97f62b7),
	.w6(32'hba4c97d7),
	.w7(32'hba937194),
	.w8(32'hbacec0d7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75e783),
	.w1(32'h39c795b8),
	.w2(32'h3a3a0064),
	.w3(32'h39a3f837),
	.w4(32'h3a6f20a1),
	.w5(32'h3a8e622a),
	.w6(32'hb949ce07),
	.w7(32'hb9bc11b7),
	.w8(32'h394fb483),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9074375),
	.w1(32'h3a900a5b),
	.w2(32'h39b041c8),
	.w3(32'hb808e0c0),
	.w4(32'h39d4cf01),
	.w5(32'hb9cf7d95),
	.w6(32'h39eaa22c),
	.w7(32'h386fa4ed),
	.w8(32'hba333ee4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa5eab),
	.w1(32'hb99d3596),
	.w2(32'hb97d513b),
	.w3(32'h39fe21b3),
	.w4(32'hb960cda4),
	.w5(32'hb910232a),
	.w6(32'hb90c463d),
	.w7(32'hb9ef5d21),
	.w8(32'hb9bd081e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987fe05),
	.w1(32'h39642ab1),
	.w2(32'h388bad70),
	.w3(32'hb8bf1a0e),
	.w4(32'h390fa1f0),
	.w5(32'h387f319e),
	.w6(32'h3a0d6c99),
	.w7(32'h39828c5f),
	.w8(32'h39a3c1db),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2a65e),
	.w1(32'hb9fb3da1),
	.w2(32'hb9a91e15),
	.w3(32'hb9ebe35a),
	.w4(32'hb9e4455f),
	.w5(32'hba8b7a30),
	.w6(32'hb9148a90),
	.w7(32'hba33d927),
	.w8(32'hba8bd56f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4e3fa),
	.w1(32'hb88451c9),
	.w2(32'hba103e40),
	.w3(32'hb999a4e3),
	.w4(32'hba157e74),
	.w5(32'hba992c1c),
	.w6(32'hb9cd03ff),
	.w7(32'hba4cbfba),
	.w8(32'hba8f56ce),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba495f1a),
	.w1(32'h39529886),
	.w2(32'h3a330253),
	.w3(32'hba76c16a),
	.w4(32'h399a587b),
	.w5(32'hb8854d88),
	.w6(32'h39b3c509),
	.w7(32'hb9e969ca),
	.w8(32'hb9b3f2ef),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993549a),
	.w1(32'hba104d2b),
	.w2(32'hb8fa5584),
	.w3(32'h3998fed1),
	.w4(32'hb9e699c2),
	.w5(32'hb9118f97),
	.w6(32'h39cd7d7e),
	.w7(32'h3844fd0e),
	.w8(32'h39b5bf99),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d401b2),
	.w1(32'hb950015b),
	.w2(32'hb6eda5d3),
	.w3(32'hb9120c60),
	.w4(32'h39eabd45),
	.w5(32'h3a9119da),
	.w6(32'hb5ee9796),
	.w7(32'hb979255b),
	.w8(32'h39273d34),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cefc89),
	.w1(32'hb92f7101),
	.w2(32'h3945602a),
	.w3(32'h38d9ab84),
	.w4(32'hb9217250),
	.w5(32'hb95bf05b),
	.w6(32'hb8bb4f38),
	.w7(32'hb9dc629a),
	.w8(32'hb9b4d176),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d68a6a),
	.w1(32'hb9b9b86d),
	.w2(32'hb99941d0),
	.w3(32'hba17111f),
	.w4(32'hba33a55d),
	.w5(32'hba006ecb),
	.w6(32'h39460454),
	.w7(32'hba26fedb),
	.w8(32'h3805277e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33110b),
	.w1(32'hb96167d3),
	.w2(32'h3a205950),
	.w3(32'h398118d9),
	.w4(32'hb978399f),
	.w5(32'h3a221226),
	.w6(32'hb993b19e),
	.w7(32'h3919ec92),
	.w8(32'hb98d6aa7),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03a2d7),
	.w1(32'h3a494a30),
	.w2(32'h39a4fbb5),
	.w3(32'h3a2af524),
	.w4(32'h3906722b),
	.w5(32'hba4120ca),
	.w6(32'h3a282ad4),
	.w7(32'h3a65c97a),
	.w8(32'h3a60c1a0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50ba41),
	.w1(32'hb99cf292),
	.w2(32'hb82c3689),
	.w3(32'h39be0b1d),
	.w4(32'hb97e5825),
	.w5(32'hb9f3873d),
	.w6(32'h399bc87b),
	.w7(32'hba050363),
	.w8(32'hb9e23fa9),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1253a6),
	.w1(32'h39212c99),
	.w2(32'hb89f9d05),
	.w3(32'hba501850),
	.w4(32'h362e66c3),
	.w5(32'hba33a01b),
	.w6(32'hb99088da),
	.w7(32'hba2b3850),
	.w8(32'hb97aad43),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f2fe7),
	.w1(32'h3a841df5),
	.w2(32'h3a84cd1e),
	.w3(32'hb940b1ff),
	.w4(32'h398b08d7),
	.w5(32'hb73fa6b5),
	.w6(32'h3aba4087),
	.w7(32'h3af792ba),
	.w8(32'h3a4fec16),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6facd6),
	.w1(32'h389474bd),
	.w2(32'h3a2b7c11),
	.w3(32'h39d67a44),
	.w4(32'hb9f12528),
	.w5(32'hba454a58),
	.w6(32'hb9edac2d),
	.w7(32'hb8bb1c46),
	.w8(32'hb9982493),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8928e1f),
	.w1(32'hb93935f5),
	.w2(32'hb941a535),
	.w3(32'hb88ec17d),
	.w4(32'hba30926c),
	.w5(32'hba917cff),
	.w6(32'h38008201),
	.w7(32'hba608811),
	.w8(32'hba8985be),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a06060),
	.w1(32'hb8c471c3),
	.w2(32'hb948b306),
	.w3(32'hb9c45121),
	.w4(32'hb9f78d92),
	.w5(32'hb9ff3ae7),
	.w6(32'hb88a0a14),
	.w7(32'hb97e475a),
	.w8(32'hb9eecd8e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937a8bb),
	.w1(32'h37d5e15e),
	.w2(32'hb95e5043),
	.w3(32'hb95d0f5c),
	.w4(32'hb995936b),
	.w5(32'hb9caacc7),
	.w6(32'h3829d698),
	.w7(32'hb933f429),
	.w8(32'hb8ad5efc),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97fa154),
	.w1(32'h39c5a076),
	.w2(32'h3a1bce48),
	.w3(32'hb98e6d4c),
	.w4(32'hb7072b3b),
	.w5(32'hb92e9433),
	.w6(32'h39295847),
	.w7(32'h38174aca),
	.w8(32'hb916dc76),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38318ff9),
	.w1(32'hb9a793d7),
	.w2(32'hb8b8c0f0),
	.w3(32'hb9786952),
	.w4(32'hb9c6116c),
	.w5(32'hb9b94e06),
	.w6(32'hba008ca0),
	.w7(32'hba41de54),
	.w8(32'hba1ff3fd),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f15cf0),
	.w1(32'hba1f6f11),
	.w2(32'hba1ba94a),
	.w3(32'hba61d82a),
	.w4(32'hba0c9dd8),
	.w5(32'hb9984f45),
	.w6(32'hb9f48a07),
	.w7(32'hba658063),
	.w8(32'hba25de09),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17a77f),
	.w1(32'h37a632b4),
	.w2(32'hb92db8b9),
	.w3(32'hb9f54ff6),
	.w4(32'hb998dcb4),
	.w5(32'hb9aea98e),
	.w6(32'h37106633),
	.w7(32'hb93c91cd),
	.w8(32'hb90451a0),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb932064d),
	.w1(32'hb958623a),
	.w2(32'hba17051d),
	.w3(32'hb94b561f),
	.w4(32'hb97a6f1a),
	.w5(32'hba47693d),
	.w6(32'h3992b326),
	.w7(32'h37cb93e2),
	.w8(32'h39f13dc7),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f836d),
	.w1(32'h39ad9a0c),
	.w2(32'h3a3f9733),
	.w3(32'hb93dabd0),
	.w4(32'hb80fd1de),
	.w5(32'hb9198d13),
	.w6(32'h39743ee7),
	.w7(32'h39ff40d2),
	.w8(32'h3a1d7d6c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a383e),
	.w1(32'h3adb7ee2),
	.w2(32'hba1e8ee0),
	.w3(32'hb9eb8f6f),
	.w4(32'hb9239722),
	.w5(32'hbb256ea1),
	.w6(32'h3a0b047b),
	.w7(32'h3962b93c),
	.w8(32'hba92fc40),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8930be9),
	.w1(32'h39b5f93c),
	.w2(32'h39b763ef),
	.w3(32'hba62e0f6),
	.w4(32'hb9a0c0f1),
	.w5(32'hba5fdfdf),
	.w6(32'hb8a7ef49),
	.w7(32'hb9751ec8),
	.w8(32'hb9e1c281),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f38dc),
	.w1(32'hb91d0b4f),
	.w2(32'hba14a7bf),
	.w3(32'hba24ded2),
	.w4(32'hb9e849e5),
	.w5(32'hba5f20b6),
	.w6(32'hb9f25a97),
	.w7(32'hba94df8c),
	.w8(32'hbaafd92d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ff24b),
	.w1(32'hb897a1b1),
	.w2(32'hba55123d),
	.w3(32'hba486fa5),
	.w4(32'hb9a5c6bd),
	.w5(32'hba90856c),
	.w6(32'hb95bb156),
	.w7(32'hb9bcd328),
	.w8(32'hb908a7b0),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52c939),
	.w1(32'h37c57915),
	.w2(32'hb9bac10a),
	.w3(32'hba9d4966),
	.w4(32'hb9d97f9e),
	.w5(32'hba19da7b),
	.w6(32'hb77242ef),
	.w7(32'hb9802acb),
	.w8(32'hb94d5494),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c9e2c9),
	.w1(32'hb8e6352a),
	.w2(32'hb9630bc1),
	.w3(32'hb959b074),
	.w4(32'hb9d214d5),
	.w5(32'hb9de2cca),
	.w6(32'h383fb60b),
	.w7(32'hb92d9c74),
	.w8(32'hb98507af),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971fc51),
	.w1(32'hb8bf0e47),
	.w2(32'hb9734191),
	.w3(32'hb9fcdd5b),
	.w4(32'hb9f65df6),
	.w5(32'hb9f4ebd5),
	.w6(32'h38e20fd3),
	.w7(32'hb957c0cd),
	.w8(32'hb9395465),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997b433),
	.w1(32'h3a7f8de7),
	.w2(32'h3a8bfa14),
	.w3(32'hba48aa0c),
	.w4(32'hb9f59ede),
	.w5(32'hbabcbff7),
	.w6(32'hba02ca1b),
	.w7(32'hba826283),
	.w8(32'hb9d283c2),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c0db8),
	.w1(32'h3a758b90),
	.w2(32'h3a4978d8),
	.w3(32'hb8bcb633),
	.w4(32'h3a82aac4),
	.w5(32'h38ab50c7),
	.w6(32'h3a7c0f63),
	.w7(32'h3a5e30bc),
	.w8(32'h3a28921b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5c23d),
	.w1(32'h39e4f6f5),
	.w2(32'h3a5ed270),
	.w3(32'hba3093bc),
	.w4(32'hb9589843),
	.w5(32'hb932750f),
	.w6(32'h39fc1875),
	.w7(32'h39c9aad7),
	.w8(32'h3a0f9049),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a5da6),
	.w1(32'hb7303925),
	.w2(32'h39fac9e0),
	.w3(32'h367f2065),
	.w4(32'hb99dae00),
	.w5(32'hb9294e36),
	.w6(32'h395d5d64),
	.w7(32'h3941b459),
	.w8(32'h39c2cc2b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce10fc),
	.w1(32'hb942f214),
	.w2(32'hb94af7f5),
	.w3(32'hb929ed6d),
	.w4(32'hba1a7161),
	.w5(32'hba1823d7),
	.w6(32'hb98d4b43),
	.w7(32'hb9a2b752),
	.w8(32'hb9a63a57),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba011e13),
	.w1(32'h39b0427c),
	.w2(32'h3acd3918),
	.w3(32'hba49dec1),
	.w4(32'hb9de5722),
	.w5(32'hba683aba),
	.w6(32'hb94dc73b),
	.w7(32'hba45f1a3),
	.w8(32'h37bc56c6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39230be0),
	.w1(32'h38bf189e),
	.w2(32'h391298d7),
	.w3(32'hb98db97e),
	.w4(32'hb8dde77d),
	.w5(32'hb99a3d60),
	.w6(32'h39cf47e1),
	.w7(32'hb8ec75ac),
	.w8(32'h398100bc),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a860f6),
	.w1(32'h3a28a810),
	.w2(32'hb97e54a8),
	.w3(32'hba6f3565),
	.w4(32'hb721148f),
	.w5(32'hba3cf49b),
	.w6(32'hba9472de),
	.w7(32'hbab056db),
	.w8(32'hbac3e131),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a3734),
	.w1(32'h3c95e5fd),
	.w2(32'hbc2d3843),
	.w3(32'hb9b007b6),
	.w4(32'h3b850909),
	.w5(32'hbc4e7fc2),
	.w6(32'h3c57044c),
	.w7(32'hbb7de553),
	.w8(32'hbc1054c6),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c0504),
	.w1(32'h3cb31e02),
	.w2(32'hb9649722),
	.w3(32'hbc265544),
	.w4(32'h3be2bbd5),
	.w5(32'hbb404dc2),
	.w6(32'h3c46d9a0),
	.w7(32'h3b43f6a5),
	.w8(32'hbbc8247e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule