module layer_10_featuremap_301(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c060e37),
	.w1(32'h3c95e006),
	.w2(32'h3bfd5f61),
	.w3(32'h3c01d17f),
	.w4(32'h3c092527),
	.w5(32'h3bf15cc9),
	.w6(32'hbbcdb5b3),
	.w7(32'h3c96c3dc),
	.w8(32'h3b87a20c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b9d2c),
	.w1(32'hba52700f),
	.w2(32'hbc92689c),
	.w3(32'hbbc60f3f),
	.w4(32'hbc3a59fb),
	.w5(32'hbbce6b60),
	.w6(32'hbc8079a0),
	.w7(32'hbcaa3f63),
	.w8(32'hbc243aaf),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23855d),
	.w1(32'hbbd23d84),
	.w2(32'hba4923b1),
	.w3(32'hbb806619),
	.w4(32'hbb282add),
	.w5(32'hba3cd576),
	.w6(32'hbba07283),
	.w7(32'hbc0157a0),
	.w8(32'h3ba89716),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fdc32),
	.w1(32'h3bdc830a),
	.w2(32'hbb0664b2),
	.w3(32'hbb89c525),
	.w4(32'hbb58a87a),
	.w5(32'h3bcb9d42),
	.w6(32'h3ba030d6),
	.w7(32'hbac8c446),
	.w8(32'h3b6f3b4f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ea480),
	.w1(32'h3afd10bc),
	.w2(32'hbc750d95),
	.w3(32'h3b8fb50f),
	.w4(32'h3a4fed57),
	.w5(32'hba6ccb29),
	.w6(32'hbb5332bf),
	.w7(32'hbc243ed0),
	.w8(32'h3b25f1db),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39834b05),
	.w1(32'h3b1e0cc3),
	.w2(32'hbb984a8a),
	.w3(32'hb9c6aab4),
	.w4(32'h3bcff766),
	.w5(32'hbbe6d948),
	.w6(32'h3c026e5f),
	.w7(32'h3ada71c8),
	.w8(32'hbb557bec),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc216b67),
	.w1(32'h381d9dad),
	.w2(32'hbb958028),
	.w3(32'hbc5adb06),
	.w4(32'hbc558c1b),
	.w5(32'hbc23044f),
	.w6(32'hbbeb6234),
	.w7(32'hbc3486b4),
	.w8(32'hbc86104b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37f6ce),
	.w1(32'h3d0cc493),
	.w2(32'h3cd701b1),
	.w3(32'hbc31df4b),
	.w4(32'h3af0dba1),
	.w5(32'h3b9d54db),
	.w6(32'hbc43c6ce),
	.w7(32'h3d53f9d6),
	.w8(32'h3c82766d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1e3dd),
	.w1(32'h3b879982),
	.w2(32'h3ba3a5ac),
	.w3(32'h3be2642e),
	.w4(32'h3b2db948),
	.w5(32'hbb2c9e23),
	.w6(32'h3c040e4d),
	.w7(32'h3b56dd9c),
	.w8(32'h3a87ae34),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ca8e0),
	.w1(32'h3b7f255f),
	.w2(32'hbb2f8d56),
	.w3(32'hbb119d6d),
	.w4(32'h3bc79763),
	.w5(32'h3bb50afe),
	.w6(32'h3c12211c),
	.w7(32'h3bc8e83c),
	.w8(32'h3c4af599),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37e81c),
	.w1(32'h3bcbf1cf),
	.w2(32'hbb414c60),
	.w3(32'hbb739852),
	.w4(32'hbaf58373),
	.w5(32'h3a5ca77a),
	.w6(32'h3b338faf),
	.w7(32'h39fcaa55),
	.w8(32'h3b0d5b3a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61dff8),
	.w1(32'hba86d00f),
	.w2(32'hbb1384b4),
	.w3(32'hbc232ac7),
	.w4(32'hbbcc52bf),
	.w5(32'h3b88d4bd),
	.w6(32'hbb65545b),
	.w7(32'hbb82489d),
	.w8(32'hbc018515),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95c05d),
	.w1(32'h3c6c3cae),
	.w2(32'h3c0cec73),
	.w3(32'h3aef57df),
	.w4(32'h3c9e9015),
	.w5(32'h3bffce14),
	.w6(32'hbc698c5b),
	.w7(32'h3c730cd4),
	.w8(32'h3bcc20ca),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921cbed),
	.w1(32'hbbe90f62),
	.w2(32'hba88b5c8),
	.w3(32'hbb720a52),
	.w4(32'hbbe38c56),
	.w5(32'hbc238e2b),
	.w6(32'hbb8a0667),
	.w7(32'hbbbed9d1),
	.w8(32'hb98dce48),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf8bfd),
	.w1(32'h3b59d8b6),
	.w2(32'h3ab87b71),
	.w3(32'hbb7dc43e),
	.w4(32'hbc050e18),
	.w5(32'h3c08b0a6),
	.w6(32'h3b83503d),
	.w7(32'hbc43c36d),
	.w8(32'h3bd21efd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcee551),
	.w1(32'hbc1abf58),
	.w2(32'hbc4c044e),
	.w3(32'h3b61075a),
	.w4(32'hbae589e4),
	.w5(32'hb84ffcc8),
	.w6(32'hbab92b6b),
	.w7(32'hba22b293),
	.w8(32'h3c0df3f2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66afa4),
	.w1(32'hbbca99e4),
	.w2(32'hbc0baad7),
	.w3(32'h3c39cdb8),
	.w4(32'h3c37271f),
	.w5(32'h3b4b832f),
	.w6(32'h3a966bd8),
	.w7(32'h3aa2d929),
	.w8(32'h3b978db4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01722c),
	.w1(32'hbc276edc),
	.w2(32'h3a312bc1),
	.w3(32'hbad1dd4b),
	.w4(32'h3b30b947),
	.w5(32'h3bbd7bab),
	.w6(32'h3bf6ce60),
	.w7(32'h3bd92d1c),
	.w8(32'h3c8c7a7b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeab6cd),
	.w1(32'hb92fe19a),
	.w2(32'hba59298d),
	.w3(32'hbbd0d2b6),
	.w4(32'hbbdba6d3),
	.w5(32'h3c19d45b),
	.w6(32'hbb33ae39),
	.w7(32'h3971dc46),
	.w8(32'h3c7a71a8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81830a),
	.w1(32'hbbc35012),
	.w2(32'hbb8289cb),
	.w3(32'h3bb6594c),
	.w4(32'hbada056b),
	.w5(32'h3c3f5e37),
	.w6(32'h3b89d8d2),
	.w7(32'hbb8546e7),
	.w8(32'h3c5f1cb4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b4611),
	.w1(32'hbc083926),
	.w2(32'hbc2b9d3c),
	.w3(32'h3c75c241),
	.w4(32'h3c1d35b2),
	.w5(32'hbb352de4),
	.w6(32'h3bdf6af4),
	.w7(32'hbbb48d1a),
	.w8(32'hb9daa7df),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2344f6),
	.w1(32'h3bc41c7a),
	.w2(32'h3b689f61),
	.w3(32'h39d53eeb),
	.w4(32'hb9c5f4a0),
	.w5(32'h3b19101a),
	.w6(32'h3b58c92e),
	.w7(32'h3b51d9d3),
	.w8(32'h3b930609),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f84ce),
	.w1(32'hbcf05cb6),
	.w2(32'hba4a9620),
	.w3(32'hbc918024),
	.w4(32'hbac59d90),
	.w5(32'h3bd6085f),
	.w6(32'h3b89d8b0),
	.w7(32'h3ae2d0d6),
	.w8(32'h3c33ca6a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cf89b),
	.w1(32'h3b57e461),
	.w2(32'hbba5b781),
	.w3(32'h3afec935),
	.w4(32'h3c2a79ff),
	.w5(32'hbb7c21c6),
	.w6(32'hbbc5f5cd),
	.w7(32'hbb2c81bf),
	.w8(32'hba4a022e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4fab3),
	.w1(32'h3add284e),
	.w2(32'h3c118312),
	.w3(32'h3c499692),
	.w4(32'h3b0cc859),
	.w5(32'hbc67c5ef),
	.w6(32'h3aadb513),
	.w7(32'h39780f65),
	.w8(32'hbb951faf),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52afcf),
	.w1(32'hbbf479df),
	.w2(32'hbb18c4e1),
	.w3(32'h3b7c7a68),
	.w4(32'h3b2a3b2f),
	.w5(32'h3a0bd40a),
	.w6(32'h3be9729f),
	.w7(32'hbbda7ecc),
	.w8(32'h3abe2573),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9844a),
	.w1(32'h3b43d63d),
	.w2(32'h3b0b9684),
	.w3(32'h3b5f9cad),
	.w4(32'h3ae5860f),
	.w5(32'h3c82bf09),
	.w6(32'h3bc2800e),
	.w7(32'h3a337002),
	.w8(32'h3c72237c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c366fd3),
	.w1(32'h3c8f38e1),
	.w2(32'h3bfb0448),
	.w3(32'h3c1b650e),
	.w4(32'h3cd48dfe),
	.w5(32'h3b41a422),
	.w6(32'h3c4b8ff8),
	.w7(32'h3c92215b),
	.w8(32'h3b6dff44),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc566b6),
	.w1(32'hbb7f0ab8),
	.w2(32'hbbe34a04),
	.w3(32'h3b513d9a),
	.w4(32'hbab00981),
	.w5(32'h3b35b6de),
	.w6(32'h3b4faa27),
	.w7(32'hbbcf94f8),
	.w8(32'h3ba1e1e6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1706eb),
	.w1(32'h3bf59193),
	.w2(32'h3bcc91ad),
	.w3(32'h3ba8c36b),
	.w4(32'h3c385969),
	.w5(32'hbb02ebef),
	.w6(32'hbbd443c2),
	.w7(32'hbb76cd43),
	.w8(32'hbc5dd28a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2738e),
	.w1(32'h3bfcd414),
	.w2(32'h3b60d68a),
	.w3(32'hbc1da595),
	.w4(32'h3b1cfabd),
	.w5(32'h3b4cfc4d),
	.w6(32'h3c3ef5c9),
	.w7(32'hb9bb64dd),
	.w8(32'h3b355b16),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb602066),
	.w1(32'hb9b0f43a),
	.w2(32'h3c09614f),
	.w3(32'h39b4ba70),
	.w4(32'h3b358c4f),
	.w5(32'hbbdc51ed),
	.w6(32'h3af37d39),
	.w7(32'h3c524e45),
	.w8(32'hba296bc2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc020165),
	.w1(32'hbbe8d783),
	.w2(32'h3c2897d3),
	.w3(32'h387df312),
	.w4(32'hbc023ba0),
	.w5(32'h3c18d56f),
	.w6(32'hbc59453b),
	.w7(32'h3adeeaf6),
	.w8(32'h3c28a409),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92cfa9),
	.w1(32'hbb169d17),
	.w2(32'hbc28206f),
	.w3(32'h3c4e9d61),
	.w4(32'h3a8d16ef),
	.w5(32'hbb82dbbc),
	.w6(32'h3b82dca0),
	.w7(32'hbc2286b6),
	.w8(32'hbb9d70d4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ba29d),
	.w1(32'h39e8548a),
	.w2(32'h3ab703bb),
	.w3(32'h39a65430),
	.w4(32'h3ae9c1db),
	.w5(32'h3c3acaf3),
	.w6(32'hbb25745d),
	.w7(32'h3b496c05),
	.w8(32'h3ba477b3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1b5c4),
	.w1(32'hbc04b2e0),
	.w2(32'hbbb2ed6c),
	.w3(32'h3b436c14),
	.w4(32'hbaa5b9d6),
	.w5(32'h3b8704c8),
	.w6(32'hbbffe3b4),
	.w7(32'hbc138066),
	.w8(32'h3b9a6e79),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a513ba),
	.w1(32'h3c01bd09),
	.w2(32'hbc8c82f6),
	.w3(32'h3b36f2e3),
	.w4(32'hbc8ca977),
	.w5(32'hbc92bd57),
	.w6(32'hbc2beb6e),
	.w7(32'hbca77480),
	.w8(32'hbc11934b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15974e),
	.w1(32'h3c480bca),
	.w2(32'hbc0c6e44),
	.w3(32'h3c4fa0bc),
	.w4(32'hbb4df299),
	.w5(32'hbc323ed2),
	.w6(32'h3bc931ba),
	.w7(32'hbc9f634f),
	.w8(32'hbc4b2b52),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c7075),
	.w1(32'h3c6fe73d),
	.w2(32'hbb6161d5),
	.w3(32'h3bcef136),
	.w4(32'h3bc5eb4b),
	.w5(32'h3c196ded),
	.w6(32'h3afc6d41),
	.w7(32'hbbc50516),
	.w8(32'hbc0356b3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67b4c9),
	.w1(32'h3bab6a17),
	.w2(32'hbc6f797f),
	.w3(32'h3a0f2878),
	.w4(32'hbb4b523c),
	.w5(32'hbb23a031),
	.w6(32'h38ad7e0c),
	.w7(32'hbbe081cf),
	.w8(32'hbb84952c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bc8e5),
	.w1(32'hbb11dd87),
	.w2(32'hb9e98995),
	.w3(32'hbb8d1052),
	.w4(32'hbb434d9d),
	.w5(32'hbc02e3f7),
	.w6(32'hbb6c8452),
	.w7(32'hba23053b),
	.w8(32'hbb70da92),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2ef7d),
	.w1(32'hbbde5e4f),
	.w2(32'hbc117551),
	.w3(32'hbbbc39a0),
	.w4(32'hbabde5f2),
	.w5(32'hbbcb737b),
	.w6(32'h3a633ba5),
	.w7(32'hbb97df36),
	.w8(32'h3b2d9375),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71b3d9),
	.w1(32'h3bd162f1),
	.w2(32'h39edfe70),
	.w3(32'hbbed1d0e),
	.w4(32'hbc6ce906),
	.w5(32'h3a85bfaa),
	.w6(32'h3a92b5a4),
	.w7(32'hbc1bc1df),
	.w8(32'hba90640d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64a22c),
	.w1(32'hbc0f6645),
	.w2(32'h3a2b7d0d),
	.w3(32'hbc0f90cf),
	.w4(32'hba6653a3),
	.w5(32'h3c05bce6),
	.w6(32'h3c052a78),
	.w7(32'h3bbeced7),
	.w8(32'h3ca53fd4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c149c6b),
	.w1(32'h3c61b72a),
	.w2(32'h3c6ec6c2),
	.w3(32'h3b3d20df),
	.w4(32'h3b538fb1),
	.w5(32'hbb3c1e32),
	.w6(32'h3b8e9541),
	.w7(32'h3ba099a9),
	.w8(32'h3b7a7cf4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93efa1),
	.w1(32'hbb9da388),
	.w2(32'h3c0295e0),
	.w3(32'h39dda323),
	.w4(32'h3c3d590f),
	.w5(32'h3ad3fd6a),
	.w6(32'h3be0803b),
	.w7(32'h3b677340),
	.w8(32'h3bdb05eb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa574b9),
	.w1(32'hbbb81a14),
	.w2(32'hbb3395f7),
	.w3(32'hbba1e0c3),
	.w4(32'hbbdb19b9),
	.w5(32'hbbded5f1),
	.w6(32'hbba52ba6),
	.w7(32'hbbd567ae),
	.w8(32'hbb2ce73e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89fd8f),
	.w1(32'hbb7efab9),
	.w2(32'h3b11dbda),
	.w3(32'hbb86e744),
	.w4(32'h3b872041),
	.w5(32'h3bd5d007),
	.w6(32'h3c468b5c),
	.w7(32'h3cad8c0a),
	.w8(32'h3c030c3f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4367ae),
	.w1(32'h3b8442c6),
	.w2(32'hbaba4bae),
	.w3(32'hbc870b98),
	.w4(32'hbb14de87),
	.w5(32'hbb7f3789),
	.w6(32'hbc2f8b9c),
	.w7(32'h3a35ce26),
	.w8(32'h3995cb51),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d527df),
	.w1(32'h3c1f6a26),
	.w2(32'hba0aae08),
	.w3(32'h3b7fb91f),
	.w4(32'hbb5330d7),
	.w5(32'hba87783b),
	.w6(32'h3becde6f),
	.w7(32'h3b10dfc7),
	.w8(32'hb900c7e2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8870d9),
	.w1(32'hbb663e29),
	.w2(32'h3a1bf60e),
	.w3(32'h3ba7d05b),
	.w4(32'hbad8088c),
	.w5(32'h38bf28c8),
	.w6(32'h3bb41f25),
	.w7(32'hbbb10f7f),
	.w8(32'hba1c9d88),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5b20e),
	.w1(32'hbbf5a46d),
	.w2(32'h3b0d82ae),
	.w3(32'h3b13f5e7),
	.w4(32'h3b9ef8a0),
	.w5(32'h3be05672),
	.w6(32'hbb6f8251),
	.w7(32'hbbcae35e),
	.w8(32'h3ad3d03f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18ffa9),
	.w1(32'h3acd5235),
	.w2(32'h3b981e6b),
	.w3(32'hbb2b7394),
	.w4(32'h3a027236),
	.w5(32'hbb83111b),
	.w6(32'hbc04ec81),
	.w7(32'h3a5830cd),
	.w8(32'h3b2ff6a6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6c3b1),
	.w1(32'hbc1e9d32),
	.w2(32'hbbbfe3ed),
	.w3(32'hbc2725fd),
	.w4(32'hbb0ca0a7),
	.w5(32'h3bf131d3),
	.w6(32'hbb58da35),
	.w7(32'h3bc15fad),
	.w8(32'h3c932867),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca9a1),
	.w1(32'hbbcdfb38),
	.w2(32'hba8eabd2),
	.w3(32'h3b0bb9de),
	.w4(32'hb92869a1),
	.w5(32'h3bc050fe),
	.w6(32'hba10c00a),
	.w7(32'hbb9bcd54),
	.w8(32'h3c08de91),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7621b),
	.w1(32'hbc0ad1a8),
	.w2(32'hbb93d192),
	.w3(32'h3b841f29),
	.w4(32'h3b26d951),
	.w5(32'hbb60ef20),
	.w6(32'hba99b0d1),
	.w7(32'hbbeae5fb),
	.w8(32'hbb592b48),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac94890),
	.w1(32'hbb5f0b37),
	.w2(32'h3bd2180b),
	.w3(32'hbadb5e1c),
	.w4(32'hbac7560e),
	.w5(32'hbb3bef54),
	.w6(32'h3ad05490),
	.w7(32'h3b17b0db),
	.w8(32'hba78d2d7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94b495),
	.w1(32'h3be0f23a),
	.w2(32'hbade54d7),
	.w3(32'hbb6bcb6d),
	.w4(32'hbb938c2d),
	.w5(32'hbc088986),
	.w6(32'hbc030efb),
	.w7(32'hbb8c7a4b),
	.w8(32'hbbaf6d7d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb616428),
	.w1(32'h3bb64035),
	.w2(32'h39d6b8e6),
	.w3(32'h3b99e8fa),
	.w4(32'hbb7d1b76),
	.w5(32'hbc769ef7),
	.w6(32'h3c1f1351),
	.w7(32'hbab7c3c0),
	.w8(32'h3c1b3d0d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad10f61),
	.w1(32'h3c51d4ac),
	.w2(32'h3c2d5a65),
	.w3(32'hbc6f020b),
	.w4(32'hbc3fcf9e),
	.w5(32'h3c22f69a),
	.w6(32'h3badac1b),
	.w7(32'hbbc5532c),
	.w8(32'h3c1a903e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeaecc3),
	.w1(32'h3b9df965),
	.w2(32'hba6966fb),
	.w3(32'h3b83540d),
	.w4(32'hb9025687),
	.w5(32'h3beb8885),
	.w6(32'h3c6d9e33),
	.w7(32'h3b6841ae),
	.w8(32'h3c4eea44),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba71717),
	.w1(32'h3b51460f),
	.w2(32'hb9da3618),
	.w3(32'hbafb27e4),
	.w4(32'h3c4854c2),
	.w5(32'hbb4e9489),
	.w6(32'hb73e7d77),
	.w7(32'h3bd500ef),
	.w8(32'h3a6c93f4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7420e),
	.w1(32'hbb895b17),
	.w2(32'hbb03995c),
	.w3(32'hbb378662),
	.w4(32'h3a67039f),
	.w5(32'h390e113d),
	.w6(32'hbb913616),
	.w7(32'h3934babb),
	.w8(32'h3b0dec9f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eff048),
	.w1(32'hbb8b5f3c),
	.w2(32'hbb7443cf),
	.w3(32'hbb5790b5),
	.w4(32'hbb6e0e70),
	.w5(32'hbb52ec23),
	.w6(32'hbb839848),
	.w7(32'hbb46fc6a),
	.w8(32'h3bcafa8a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ee31f),
	.w1(32'hbb078ad6),
	.w2(32'h3ae986ed),
	.w3(32'hba956fe1),
	.w4(32'hbafed19f),
	.w5(32'h3b834ff4),
	.w6(32'h3b180b2b),
	.w7(32'h3af8fc60),
	.w8(32'hbb203246),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d73e8),
	.w1(32'hbb7199c1),
	.w2(32'hba33d856),
	.w3(32'h3adb1712),
	.w4(32'h3bb862e4),
	.w5(32'h3b752295),
	.w6(32'hbb0fbbdd),
	.w7(32'h3a1e989f),
	.w8(32'hba0e9c17),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae249c0),
	.w1(32'h3c900339),
	.w2(32'h3afb6162),
	.w3(32'hbcb4df3d),
	.w4(32'hbc203ac8),
	.w5(32'hbb4cac66),
	.w6(32'hbc56b599),
	.w7(32'h3c914a1a),
	.w8(32'h3bb55985),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37de63),
	.w1(32'hbc4ac9ab),
	.w2(32'hbb5ed5e9),
	.w3(32'hbb3aeac9),
	.w4(32'h3b5656e8),
	.w5(32'h3c30f462),
	.w6(32'hbb5ff4e9),
	.w7(32'hbc5a580c),
	.w8(32'h3c1331c0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc106098),
	.w1(32'hbc9a9075),
	.w2(32'h39167fab),
	.w3(32'hbaa21e33),
	.w4(32'hbc25e4e9),
	.w5(32'h3bf1feef),
	.w6(32'hb983f61a),
	.w7(32'hbbf88373),
	.w8(32'h3a9a9cb3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c409410),
	.w1(32'h3bdd26a2),
	.w2(32'h3ba7fe7d),
	.w3(32'h3bfb9e5b),
	.w4(32'h3a35fc1c),
	.w5(32'hbbf9ff7e),
	.w6(32'hbb91b03c),
	.w7(32'hbbadf5ea),
	.w8(32'hbc4925a9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc372ad),
	.w1(32'h3c30c051),
	.w2(32'h3b30860f),
	.w3(32'h3a6c5620),
	.w4(32'hbbd8ee3d),
	.w5(32'hbbc151f2),
	.w6(32'h3b678d10),
	.w7(32'hba49e14b),
	.w8(32'hbc2d6e55),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf791fe),
	.w1(32'hbaa9ecc4),
	.w2(32'hb98e8808),
	.w3(32'hbc138833),
	.w4(32'h3b627c80),
	.w5(32'hbbe8d985),
	.w6(32'hbc6bc7f5),
	.w7(32'h3c248e48),
	.w8(32'hbb9bb203),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ef3fa),
	.w1(32'h3baf893f),
	.w2(32'h3bb3f648),
	.w3(32'hbc13818b),
	.w4(32'hbbcdb6d7),
	.w5(32'h3b8fecf5),
	.w6(32'hbc442f80),
	.w7(32'hbacb37cf),
	.w8(32'h3bdb4ffb),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d3387),
	.w1(32'h3a1be069),
	.w2(32'hbbcfb5b7),
	.w3(32'h3b6c6918),
	.w4(32'hba0e2501),
	.w5(32'h3c4f97c8),
	.w6(32'h3c20a579),
	.w7(32'hbb6e810e),
	.w8(32'h3c8d1a9a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ee71b6),
	.w1(32'h3ba5efae),
	.w2(32'hbbe98b6b),
	.w3(32'h3bf40631),
	.w4(32'hbbde9082),
	.w5(32'h3baf4ae0),
	.w6(32'hbbd75e74),
	.w7(32'hbba7399b),
	.w8(32'h3b666a29),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e3f1d6),
	.w1(32'hbb45eb05),
	.w2(32'h3a8cb8d1),
	.w3(32'hbbe40388),
	.w4(32'hbace4a9f),
	.w5(32'h3bfe1323),
	.w6(32'h3a362978),
	.w7(32'h3bc770bf),
	.w8(32'h3aebd7f2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6aafc),
	.w1(32'h3aa490b4),
	.w2(32'h3ad731a1),
	.w3(32'hbbbb7b08),
	.w4(32'hbb0f8191),
	.w5(32'h3b61bf5d),
	.w6(32'hbc095bd4),
	.w7(32'h3c0258ce),
	.w8(32'h3c37218d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c0c63),
	.w1(32'h3b948f5a),
	.w2(32'h3b38a5cc),
	.w3(32'h3c35b261),
	.w4(32'h3bae0160),
	.w5(32'h3c4276f7),
	.w6(32'h3b043b28),
	.w7(32'h3b4f6e09),
	.w8(32'hbb95076c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb840e3f),
	.w1(32'h3bfaf497),
	.w2(32'hbb246e10),
	.w3(32'hbc0de61b),
	.w4(32'h3ba3dde5),
	.w5(32'h3bbc25de),
	.w6(32'hba62adb9),
	.w7(32'h3c48fa39),
	.w8(32'h3bc3d752),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba194f33),
	.w1(32'h3c22bc9e),
	.w2(32'hbb331653),
	.w3(32'hbb74c964),
	.w4(32'h3c561438),
	.w5(32'h3b037c9c),
	.w6(32'hba32aed9),
	.w7(32'h3bc7f96f),
	.w8(32'hbc838004),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b359473),
	.w1(32'h3bb4b305),
	.w2(32'h3b6bd593),
	.w3(32'hbc06e7a3),
	.w4(32'hbb8373e1),
	.w5(32'h3b2998f5),
	.w6(32'hbb54632b),
	.w7(32'h3ba0d121),
	.w8(32'h3a3cbb2c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6699fd),
	.w1(32'h3b8c1c8e),
	.w2(32'hbafba87e),
	.w3(32'hbbd1dd7a),
	.w4(32'hbbaaa1f4),
	.w5(32'h3a015d7f),
	.w6(32'h3bc57084),
	.w7(32'h3b9c9d6e),
	.w8(32'h3bdcf5f7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbc012),
	.w1(32'h3b364b35),
	.w2(32'hbb0c1b36),
	.w3(32'hbc11527d),
	.w4(32'hb9d2bdcb),
	.w5(32'hbbe90244),
	.w6(32'hbb7376eb),
	.w7(32'h3bac3910),
	.w8(32'h398abc3d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96eb7f),
	.w1(32'hbc66ee6c),
	.w2(32'hbc93ec92),
	.w3(32'hbbb0bd8b),
	.w4(32'hbc0bf12b),
	.w5(32'h3b208aab),
	.w6(32'hbbfb7d6d),
	.w7(32'hbc84a8d0),
	.w8(32'h3b889785),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae96ae4),
	.w1(32'hbb451e5f),
	.w2(32'hba942f93),
	.w3(32'h3b0229e3),
	.w4(32'h3b53e00e),
	.w5(32'h3b365da9),
	.w6(32'hbb11cdda),
	.w7(32'h3b0d1a88),
	.w8(32'h3b6cefb0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84aa91),
	.w1(32'h3b5c9441),
	.w2(32'h3b86b437),
	.w3(32'hbbb1de1f),
	.w4(32'h3c0b58e7),
	.w5(32'hbbc1d013),
	.w6(32'h3c24ca5a),
	.w7(32'h3c443f23),
	.w8(32'hbab700ac),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afe755),
	.w1(32'hbb010412),
	.w2(32'hbc2c9f7b),
	.w3(32'h39100696),
	.w4(32'hbc28e835),
	.w5(32'hbbac5d3a),
	.w6(32'hb8d2768d),
	.w7(32'hbc883614),
	.w8(32'hbc4bd00f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a7f6c),
	.w1(32'h3a958561),
	.w2(32'h3b3e8f71),
	.w3(32'h3bc76e0c),
	.w4(32'h3c024e4d),
	.w5(32'h3ad7a2ea),
	.w6(32'hba5f910a),
	.w7(32'hba5dee2c),
	.w8(32'h3a9422cb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77c1d9),
	.w1(32'h3ba97725),
	.w2(32'h3b5fe0b4),
	.w3(32'h3c489181),
	.w4(32'h3be68bd0),
	.w5(32'h3bee4662),
	.w6(32'h3892d765),
	.w7(32'hbbaef9c1),
	.w8(32'hbc604e1f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc710345),
	.w1(32'hbc41f5f4),
	.w2(32'h3a9b24b6),
	.w3(32'hbbfb0151),
	.w4(32'h3c407f8f),
	.w5(32'h3c5eb312),
	.w6(32'h3b19da5a),
	.w7(32'h3c46ac53),
	.w8(32'h3ca17eca),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19770c),
	.w1(32'hbbb499c8),
	.w2(32'hbbeaf4ea),
	.w3(32'h3c4dc0d6),
	.w4(32'h3c752f83),
	.w5(32'h3b01a6ac),
	.w6(32'hbc2bff2b),
	.w7(32'hbc14191f),
	.w8(32'hbb16d8e2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68723c),
	.w1(32'hbc46172c),
	.w2(32'hbb6ffcad),
	.w3(32'hbc922a5d),
	.w4(32'hbc7b2945),
	.w5(32'h3afc4158),
	.w6(32'hbba1854c),
	.w7(32'h3886cf14),
	.w8(32'h3b58016f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c747c),
	.w1(32'hbbdb77ba),
	.w2(32'hbc20d61a),
	.w3(32'h3b1ad9a6),
	.w4(32'h3ae4e5c8),
	.w5(32'hb90cb801),
	.w6(32'hbc13ef7b),
	.w7(32'hbb57dc91),
	.w8(32'hbbe64067),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b48bdd),
	.w1(32'hbbccc252),
	.w2(32'h3a9edeb3),
	.w3(32'hbbb9dc6b),
	.w4(32'hbc48436c),
	.w5(32'hb98d4b5f),
	.w6(32'hbb4cee29),
	.w7(32'hbadef184),
	.w8(32'h3b9bd9ef),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e8874),
	.w1(32'hbb1d567d),
	.w2(32'hb8ff3f60),
	.w3(32'hbc157c0b),
	.w4(32'hbbf6a1bf),
	.w5(32'hbbd2f2c2),
	.w6(32'hbbe2e3eb),
	.w7(32'hbb4d2714),
	.w8(32'hbc498330),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc809a5),
	.w1(32'h3c487387),
	.w2(32'h3b4ac23a),
	.w3(32'h3a8368ae),
	.w4(32'hbc4652bf),
	.w5(32'h3c51e50e),
	.w6(32'hbc39c5a2),
	.w7(32'hbcbe5f93),
	.w8(32'h3af79b34),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b4f72),
	.w1(32'hbb8bcc7c),
	.w2(32'hbc343b35),
	.w3(32'hbb826e53),
	.w4(32'hbb9960dd),
	.w5(32'hbc8e8eb4),
	.w6(32'h3995b196),
	.w7(32'hbc10e287),
	.w8(32'hbc4072e4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b0792),
	.w1(32'hbc5274fd),
	.w2(32'h3c29dd71),
	.w3(32'hbc000a8a),
	.w4(32'hba90d5db),
	.w5(32'h3c34cffc),
	.w6(32'hbb709a59),
	.w7(32'h3bd6e8f1),
	.w8(32'h3ccc51f7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d6c60),
	.w1(32'h3c5a0cd2),
	.w2(32'h3adfbdc5),
	.w3(32'hbbeea061),
	.w4(32'hbc50da1c),
	.w5(32'h3a351804),
	.w6(32'h3bc8c853),
	.w7(32'h3b1989e4),
	.w8(32'hba1164ef),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78b619),
	.w1(32'hbd08364f),
	.w2(32'hbcb8a28b),
	.w3(32'hbbaa9fc9),
	.w4(32'hbccc3aa7),
	.w5(32'hbb2b436f),
	.w6(32'hbc14ae36),
	.w7(32'hbc96b308),
	.w8(32'hbabde48e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d927b),
	.w1(32'h3a4500a0),
	.w2(32'hbc9a4af7),
	.w3(32'hbc1ec345),
	.w4(32'hbd0f5edc),
	.w5(32'hbcb61585),
	.w6(32'hbc4136f9),
	.w7(32'hbd3766ec),
	.w8(32'hbcbbaa74),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52bb4d),
	.w1(32'h3bd8d464),
	.w2(32'h3b007596),
	.w3(32'h3bb1d1fe),
	.w4(32'h3b6ba495),
	.w5(32'hbadd8b6e),
	.w6(32'h3b88aeb2),
	.w7(32'hbae60b9a),
	.w8(32'hbb9a343f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc088466),
	.w1(32'hbba2b6e4),
	.w2(32'hbbd5614b),
	.w3(32'hbcd0ea53),
	.w4(32'hbca37f17),
	.w5(32'hba37737a),
	.w6(32'hbc6fd1fb),
	.w7(32'hbc608348),
	.w8(32'hbb1f437a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61a069),
	.w1(32'hbbf572a2),
	.w2(32'hbc451095),
	.w3(32'hbb81284f),
	.w4(32'hbc3627e1),
	.w5(32'hbc4b4244),
	.w6(32'hbc1f99ca),
	.w7(32'hbc3c7801),
	.w8(32'h3a4ad215),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba77349),
	.w1(32'hbbf687f4),
	.w2(32'hbc545b93),
	.w3(32'hbca1b936),
	.w4(32'hbcc77531),
	.w5(32'h3b65b8d2),
	.w6(32'hbc187693),
	.w7(32'hbc478509),
	.w8(32'hbc512829),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf61730),
	.w1(32'hbb12d4a5),
	.w2(32'h3ac07aee),
	.w3(32'h3c780d1a),
	.w4(32'h3c21d9fa),
	.w5(32'hbbc8f1d8),
	.w6(32'h3b4d1cf6),
	.w7(32'h3c065ad2),
	.w8(32'hbbaac047),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3cb47),
	.w1(32'hbc0c690d),
	.w2(32'hbb991314),
	.w3(32'hbc90ddf3),
	.w4(32'hbb9a8a2a),
	.w5(32'h3b41c932),
	.w6(32'hbc64dfd5),
	.w7(32'h3b24110f),
	.w8(32'h3a10afa3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbd533),
	.w1(32'hbb17878a),
	.w2(32'h3b80edb6),
	.w3(32'h3b825ada),
	.w4(32'hbbc8b418),
	.w5(32'h3b72a43d),
	.w6(32'h3b2b3e52),
	.w7(32'hbba1c822),
	.w8(32'h3caf0b46),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a6346),
	.w1(32'h3ca6175f),
	.w2(32'h3bad306e),
	.w3(32'h3b631cb9),
	.w4(32'hbb9f42f7),
	.w5(32'h3be932e3),
	.w6(32'h3cac6ad2),
	.w7(32'h3c394b90),
	.w8(32'h3c8b3d0e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8357ab),
	.w1(32'h3b88e112),
	.w2(32'h3c65c414),
	.w3(32'h3c1bb4f8),
	.w4(32'h3bb48614),
	.w5(32'hbb53cb43),
	.w6(32'h3c0a19a4),
	.w7(32'h3c164ac3),
	.w8(32'hbc0bd0b7),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eeaa4),
	.w1(32'h3bd4d1b5),
	.w2(32'h3bb2d192),
	.w3(32'h3b6f0727),
	.w4(32'h3c7a19c8),
	.w5(32'h3b928c2f),
	.w6(32'hbb97ab4c),
	.w7(32'h3b70a520),
	.w8(32'h3b7a9164),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be37e71),
	.w1(32'h3c0b68aa),
	.w2(32'h3b4e27c8),
	.w3(32'h3b3a0118),
	.w4(32'hba3aec88),
	.w5(32'hbbdc811e),
	.w6(32'h3b9cebd2),
	.w7(32'hbad4abe1),
	.w8(32'hbbcb097a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28eb1c),
	.w1(32'hbb29f660),
	.w2(32'h3af147a9),
	.w3(32'h3c36d6a9),
	.w4(32'h3be3b6ce),
	.w5(32'h3be4c5a6),
	.w6(32'h3c42aa37),
	.w7(32'h3bd3d166),
	.w8(32'h3b140caf),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7a432),
	.w1(32'hbba2f01a),
	.w2(32'h3ab201cf),
	.w3(32'hbb6edf69),
	.w4(32'hbb8f635d),
	.w5(32'h3bae1b18),
	.w6(32'h3b7b844a),
	.w7(32'h3ab9b666),
	.w8(32'hbbcb1b31),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe89331),
	.w1(32'hbc725fbe),
	.w2(32'hbb1bcda0),
	.w3(32'h3adf4b0b),
	.w4(32'hbb02d403),
	.w5(32'hbaea5127),
	.w6(32'hbb4087d3),
	.w7(32'hbc44affe),
	.w8(32'hbb3e2607),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b176408),
	.w1(32'h3ba97094),
	.w2(32'hbae25efb),
	.w3(32'hbba0d173),
	.w4(32'hbb7ea4f8),
	.w5(32'h3b9bcfed),
	.w6(32'h3b74efcb),
	.w7(32'h3ae2e285),
	.w8(32'h3c720973),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e50e5),
	.w1(32'h3bc62640),
	.w2(32'h3bbd89cb),
	.w3(32'hbb087359),
	.w4(32'h3ac21a8a),
	.w5(32'hbc44e85d),
	.w6(32'h3bee6293),
	.w7(32'h3baeefbe),
	.w8(32'hbbfb8835),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd13b2),
	.w1(32'hbbc783de),
	.w2(32'hbc23b6df),
	.w3(32'hbc845424),
	.w4(32'hbc4d5907),
	.w5(32'h3b415d08),
	.w6(32'hbc2abedc),
	.w7(32'hbc4a151b),
	.w8(32'h3c16c8d6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be54505),
	.w1(32'hbb2fab8b),
	.w2(32'hbb54d4db),
	.w3(32'hbb81fe63),
	.w4(32'hbb8a6add),
	.w5(32'h3c060f15),
	.w6(32'h3aa0979e),
	.w7(32'hbb33c9eb),
	.w8(32'h3c815edd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c653ab8),
	.w1(32'h3be15c7f),
	.w2(32'h38dec0a2),
	.w3(32'h3c1cc1ae),
	.w4(32'hbbab1b1f),
	.w5(32'h3bcfe43b),
	.w6(32'h3c526704),
	.w7(32'hbaea3001),
	.w8(32'hbb55f5b2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeeed22),
	.w1(32'hb98d1c3e),
	.w2(32'hbaa7be58),
	.w3(32'hbc38b27c),
	.w4(32'h3a660953),
	.w5(32'hbbefef5a),
	.w6(32'hbbb1aefc),
	.w7(32'hb8cc1cd5),
	.w8(32'hbc535477),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d5fa4),
	.w1(32'hbbcf78f5),
	.w2(32'hbb613124),
	.w3(32'hbbb6f874),
	.w4(32'hbabb2d37),
	.w5(32'hbc4e4be9),
	.w6(32'hbc39aed5),
	.w7(32'h3c6c93de),
	.w8(32'hbc51b450),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ab330),
	.w1(32'h3c027c4b),
	.w2(32'h399dbe3b),
	.w3(32'h3c095fba),
	.w4(32'h3c9208f3),
	.w5(32'h3baa3706),
	.w6(32'hbc5e386c),
	.w7(32'h3c0a37e9),
	.w8(32'hbc71430b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69d2af),
	.w1(32'hbc265583),
	.w2(32'h3bc79a17),
	.w3(32'h3c6a0036),
	.w4(32'h3bf937f4),
	.w5(32'hbb0d95b1),
	.w6(32'h3b8e4ece),
	.w7(32'h3c41030e),
	.w8(32'hbc63fbf4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc198bed),
	.w1(32'hbb1a4088),
	.w2(32'h3a0e1355),
	.w3(32'h3b5c9cca),
	.w4(32'h3c4be2ae),
	.w5(32'hbbd2b047),
	.w6(32'hb964b22b),
	.w7(32'h3c8b13ae),
	.w8(32'hbb3e1d6a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e335e),
	.w1(32'hbc189073),
	.w2(32'hbb72be2d),
	.w3(32'hbad4fae8),
	.w4(32'hbb849750),
	.w5(32'h3b63d3e4),
	.w6(32'hbb91655c),
	.w7(32'h3af6ff72),
	.w8(32'h3bcad556),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb844ac6d),
	.w1(32'h3a61b549),
	.w2(32'hb9ef6146),
	.w3(32'h3b90f890),
	.w4(32'hbb2c76d1),
	.w5(32'hbad39888),
	.w6(32'h3bcd6d19),
	.w7(32'h3a16853b),
	.w8(32'hbc339695),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8a1a2),
	.w1(32'hbc6dfea7),
	.w2(32'h3b184c12),
	.w3(32'h3b6d0a2c),
	.w4(32'h38861058),
	.w5(32'h3bfb6fba),
	.w6(32'h38720afc),
	.w7(32'hbbab8ca6),
	.w8(32'h3c2c115d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10764c),
	.w1(32'hb92b1fb1),
	.w2(32'h3c8de041),
	.w3(32'h3b50f9bb),
	.w4(32'h3c487497),
	.w5(32'h3b3ec7ec),
	.w6(32'h3c02bae9),
	.w7(32'h3cba8014),
	.w8(32'h3bfb5d4d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba97cc9),
	.w1(32'hbbfa12e6),
	.w2(32'hba2fd992),
	.w3(32'h3bb14c8d),
	.w4(32'hbad98fbe),
	.w5(32'h3ba11b31),
	.w6(32'hb96ee85d),
	.w7(32'h3b739f51),
	.w8(32'hba8d7058),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22e2da),
	.w1(32'hbb575084),
	.w2(32'hbbe45c25),
	.w3(32'hbc0f4195),
	.w4(32'hbc0ea493),
	.w5(32'h3c308e3c),
	.w6(32'hbbe956d9),
	.w7(32'hb854107f),
	.w8(32'h3cb509d5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ad55b),
	.w1(32'h3c710bfa),
	.w2(32'h3b3549e6),
	.w3(32'h3b15a309),
	.w4(32'hba610544),
	.w5(32'hba05d803),
	.w6(32'h3c87cdb9),
	.w7(32'hba67fc9d),
	.w8(32'h3bfdbada),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecfe55),
	.w1(32'hbc01cde9),
	.w2(32'hbbb445b3),
	.w3(32'h3b8fc7cf),
	.w4(32'hbc2dceaa),
	.w5(32'h3ba565d7),
	.w6(32'h3b5812ef),
	.w7(32'h3c294d80),
	.w8(32'h3c5508b1),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc9583),
	.w1(32'h3b335a55),
	.w2(32'h3ba69b5d),
	.w3(32'hb9178ca2),
	.w4(32'hbbc5383f),
	.w5(32'hbbc42354),
	.w6(32'h3aa86e64),
	.w7(32'hbade44bd),
	.w8(32'hbb86360e),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdde9a2),
	.w1(32'hbc04fa9e),
	.w2(32'h3a632c58),
	.w3(32'hbc92280b),
	.w4(32'hbbb131cf),
	.w5(32'h3b1da97c),
	.w6(32'h3ba14d4f),
	.w7(32'h3bbb0832),
	.w8(32'h3ce1207c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2e216),
	.w1(32'h3c458a70),
	.w2(32'h3bb910b9),
	.w3(32'hbac43c59),
	.w4(32'hbc071260),
	.w5(32'hb9fa3264),
	.w6(32'hba9f8905),
	.w7(32'hbb6a0194),
	.w8(32'h3992ccb2),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a720ef5),
	.w1(32'h3ac36445),
	.w2(32'h3be6149c),
	.w3(32'hbb33bedb),
	.w4(32'h3b210b2f),
	.w5(32'h3b5858fe),
	.w6(32'h3c3f199c),
	.w7(32'h3ba8ad31),
	.w8(32'h3c1f3da2),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd12bf6),
	.w1(32'hbb8b8b9e),
	.w2(32'h3be7ce83),
	.w3(32'hbc4fdd40),
	.w4(32'hbc4ca87e),
	.w5(32'h3b0a38f3),
	.w6(32'h3bcfdbfc),
	.w7(32'h3ba83d0a),
	.w8(32'h3c89c5de),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99dd1b),
	.w1(32'h3baff9b4),
	.w2(32'h3b08a675),
	.w3(32'h3b7f1b7a),
	.w4(32'hbb0f2390),
	.w5(32'h3ac36fcc),
	.w6(32'h3c075f1b),
	.w7(32'h3b97a017),
	.w8(32'hbc4b7932),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb86893),
	.w1(32'hba8290b2),
	.w2(32'hb91ab357),
	.w3(32'hbc50282a),
	.w4(32'hbc659ecc),
	.w5(32'h3b8b656a),
	.w6(32'hbc4bc6dd),
	.w7(32'h3bca9631),
	.w8(32'h3a7c941c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb798e22),
	.w1(32'h3b0b2a86),
	.w2(32'h3c18f76e),
	.w3(32'h3ca3ece5),
	.w4(32'h3c8eac3f),
	.w5(32'hba460c63),
	.w6(32'h3ac84611),
	.w7(32'h3c584f55),
	.w8(32'hbb0d3f4f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b847b8a),
	.w1(32'hbace1394),
	.w2(32'h3a3f0cd5),
	.w3(32'hbb68a6a6),
	.w4(32'h3adb6ca9),
	.w5(32'hbb42cf4f),
	.w6(32'hbcb97f7b),
	.w7(32'hbbef781c),
	.w8(32'hbbc84a9a),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c3e04),
	.w1(32'hbb8d00cc),
	.w2(32'hbbbd885d),
	.w3(32'hbbfd635e),
	.w4(32'hbbda273d),
	.w5(32'hbbc48b5f),
	.w6(32'hbb77ec9f),
	.w7(32'hbb9ad973),
	.w8(32'h3ad19658),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd95570),
	.w1(32'hbbbdbe0c),
	.w2(32'h3a57debd),
	.w3(32'h3ba0f487),
	.w4(32'h39b44636),
	.w5(32'h3b631c05),
	.w6(32'hbb1f8a4e),
	.w7(32'h3aa6664d),
	.w8(32'hb92da8bd),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82a366),
	.w1(32'h3c150643),
	.w2(32'h3c32821d),
	.w3(32'h3c3997a6),
	.w4(32'h3b166618),
	.w5(32'hb8acdc3e),
	.w6(32'h3c11d27d),
	.w7(32'h3baa5373),
	.w8(32'hbb8e906b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42c604),
	.w1(32'hbb9ea24a),
	.w2(32'hbb825734),
	.w3(32'h3bbad165),
	.w4(32'h3b74bbe9),
	.w5(32'hba8637ac),
	.w6(32'hba0384ed),
	.w7(32'h3bea74e9),
	.w8(32'hbb8980dd),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb099d25),
	.w1(32'hba7e0030),
	.w2(32'hbba16b03),
	.w3(32'h3bf1ade1),
	.w4(32'hbc01bff2),
	.w5(32'hbb4faed1),
	.w6(32'hbb198cd0),
	.w7(32'hbc580ac4),
	.w8(32'hbbbef037),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac117c),
	.w1(32'h3b4762fa),
	.w2(32'hbaa4c1e4),
	.w3(32'h3c842137),
	.w4(32'h3b1a35ae),
	.w5(32'hb9dab27a),
	.w6(32'h3ba56edc),
	.w7(32'h3bd9be3e),
	.w8(32'h3bd489d5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16f694),
	.w1(32'hbc401bbe),
	.w2(32'hbaccb8f1),
	.w3(32'h3bfb183f),
	.w4(32'h3c083acf),
	.w5(32'h3c08ecbf),
	.w6(32'hbc2b1e30),
	.w7(32'h3b68b1ed),
	.w8(32'h3c8790d5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d029a),
	.w1(32'h3c5f4c25),
	.w2(32'h3b8d953f),
	.w3(32'hbc0db5ab),
	.w4(32'hbc48373c),
	.w5(32'h3c08f91b),
	.w6(32'h3be59edb),
	.w7(32'hb9daaeee),
	.w8(32'h3c57bdcb),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d5cae),
	.w1(32'h3b2d0b50),
	.w2(32'h3b0955e5),
	.w3(32'h3b333efa),
	.w4(32'h3b932e06),
	.w5(32'hbb266c76),
	.w6(32'h3b79f822),
	.w7(32'h3b879afb),
	.w8(32'h3afb49a0),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c4db6),
	.w1(32'hbc49d04f),
	.w2(32'h3a18f2e8),
	.w3(32'h3b33e92e),
	.w4(32'hbbe059a3),
	.w5(32'hbaa9cdd4),
	.w6(32'hbc44c89c),
	.w7(32'hbb9bc40f),
	.w8(32'h3b1676ed),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba043cf),
	.w1(32'h3bcf6523),
	.w2(32'h3c3ed4c1),
	.w3(32'hbba3e9d2),
	.w4(32'h3c24b36a),
	.w5(32'h3bac6523),
	.w6(32'hbbcaa87e),
	.w7(32'h3b241839),
	.w8(32'hbada5b74),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8009e1),
	.w1(32'hbba2de11),
	.w2(32'hbbaa4b25),
	.w3(32'hbb65047a),
	.w4(32'hbbeb2a7a),
	.w5(32'hbbf4e061),
	.w6(32'h3920c97b),
	.w7(32'hbc3ba5d9),
	.w8(32'h3b3f06b8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde6f4f),
	.w1(32'h3c33925c),
	.w2(32'h3a86e1fe),
	.w3(32'hbb82907e),
	.w4(32'hbc17a220),
	.w5(32'h3beb58f7),
	.w6(32'h3c3a0f96),
	.w7(32'hbb9481d8),
	.w8(32'h3c14364e),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb9d82),
	.w1(32'h3bb149ba),
	.w2(32'h3c8a7bf3),
	.w3(32'h3c868736),
	.w4(32'h3c07e064),
	.w5(32'hbbd6e77a),
	.w6(32'h3c640cd4),
	.w7(32'h3c45c22d),
	.w8(32'hbbf35b3c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38489d),
	.w1(32'hbc3009e4),
	.w2(32'hbb9f5184),
	.w3(32'hbbfde44d),
	.w4(32'hbc2d80e3),
	.w5(32'hbc4432a2),
	.w6(32'hbc932dec),
	.w7(32'hbc7f61d3),
	.w8(32'hbca8dca2),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c871e),
	.w1(32'h3a83e36a),
	.w2(32'h3b94e5ff),
	.w3(32'h3bdc28eb),
	.w4(32'h38da7fb2),
	.w5(32'hbb93e917),
	.w6(32'hbc20d531),
	.w7(32'h3bbf5659),
	.w8(32'hbc0d68b9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb78937),
	.w1(32'hbcbd6845),
	.w2(32'hbc384de8),
	.w3(32'hbbebc8bf),
	.w4(32'hbb06c79d),
	.w5(32'h3bc7761e),
	.w6(32'hbc4a70d1),
	.w7(32'hbc03b06d),
	.w8(32'hbc941638),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0301c9),
	.w1(32'hbc3cb5b2),
	.w2(32'h3b860e25),
	.w3(32'hbaf9d29a),
	.w4(32'hbc11405d),
	.w5(32'hbb4eed58),
	.w6(32'hbc376a27),
	.w7(32'hbbe87080),
	.w8(32'hbbfa0f43),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabaee9),
	.w1(32'hbbbc30d5),
	.w2(32'hbaef52f2),
	.w3(32'hbc11b0d7),
	.w4(32'hbc1d1b8e),
	.w5(32'h3bed051f),
	.w6(32'hbb997b81),
	.w7(32'hbc1ff5a8),
	.w8(32'h3c04f7af),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ba4a0),
	.w1(32'hbbb8a263),
	.w2(32'h3b63a911),
	.w3(32'h3c238af0),
	.w4(32'h3c107cb4),
	.w5(32'hba584b4f),
	.w6(32'h3ac7694c),
	.w7(32'h3c5cda41),
	.w8(32'h3b1952f3),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf1e67),
	.w1(32'hbaa55cac),
	.w2(32'h3b903460),
	.w3(32'hbb28d1c3),
	.w4(32'hbbdca143),
	.w5(32'h39a94c1d),
	.w6(32'hbbb2dee5),
	.w7(32'hbb75c2b4),
	.w8(32'h3b537818),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13fdd7),
	.w1(32'hbc55bd3f),
	.w2(32'hb97defa7),
	.w3(32'hba4b603b),
	.w4(32'hbb67a949),
	.w5(32'hbc3ea046),
	.w6(32'hbb62ff43),
	.w7(32'hbac303a9),
	.w8(32'hbbbe2591),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcf55e),
	.w1(32'hbb3d1b84),
	.w2(32'hbc0d0dfd),
	.w3(32'hbbef985e),
	.w4(32'hbadd6ff9),
	.w5(32'hb86984b4),
	.w6(32'hbb656ad3),
	.w7(32'hbbf7527a),
	.w8(32'h3b82bf49),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51f663),
	.w1(32'h3b8bfc5a),
	.w2(32'h3c0db192),
	.w3(32'hbbbe124b),
	.w4(32'hbb9998c3),
	.w5(32'h3b3722af),
	.w6(32'h3b963479),
	.w7(32'h3b44bd9d),
	.w8(32'hbc5a6df7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc805628),
	.w1(32'hbc75e3e1),
	.w2(32'hbaea6f32),
	.w3(32'h3c22639d),
	.w4(32'h3c05a947),
	.w5(32'h3c12a894),
	.w6(32'hbc7558ea),
	.w7(32'h3b5aa925),
	.w8(32'h3cb6665e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8f937),
	.w1(32'h3ca2059e),
	.w2(32'h3ab102e1),
	.w3(32'hbc720e5d),
	.w4(32'hbca7be12),
	.w5(32'hbbd3b0c5),
	.w6(32'hbc6425e3),
	.w7(32'hbccbdfe8),
	.w8(32'hbbf5da06),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ef285),
	.w1(32'hbbb01b81),
	.w2(32'h3bb09ea5),
	.w3(32'hbc036a0d),
	.w4(32'h3b88e21e),
	.w5(32'h3c16adc6),
	.w6(32'hbbba8fae),
	.w7(32'hba8aed19),
	.w8(32'h3c466589),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26c0a9),
	.w1(32'h3baf8e60),
	.w2(32'hbbe481ed),
	.w3(32'hbaccd2e1),
	.w4(32'hbc567c47),
	.w5(32'h3b9b8cab),
	.w6(32'h3c2fe873),
	.w7(32'hbc3523f6),
	.w8(32'hbbabbbb4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b2583a),
	.w1(32'hbb0b841e),
	.w2(32'hbc115535),
	.w3(32'h3c466778),
	.w4(32'h3c90e8c7),
	.w5(32'hbb8589f1),
	.w6(32'hbb4202c3),
	.w7(32'h3bf9b7bd),
	.w8(32'hbbc45886),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fedb8),
	.w1(32'hbc1e895b),
	.w2(32'hb9663a4e),
	.w3(32'hbbfbcfa3),
	.w4(32'hba837ef2),
	.w5(32'h3c11911c),
	.w6(32'hbc46536d),
	.w7(32'h391dfdf8),
	.w8(32'h3c6f1247),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb63f98),
	.w1(32'h3bc72be0),
	.w2(32'hbb05ee66),
	.w3(32'h3b5a4ad1),
	.w4(32'hbc33da2f),
	.w5(32'h3c2d7214),
	.w6(32'h3cbe0186),
	.w7(32'hbc328845),
	.w8(32'hb7bcf942),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6147e6),
	.w1(32'hbbf0a5a4),
	.w2(32'h3aca4e3e),
	.w3(32'h3af30019),
	.w4(32'hbb986b70),
	.w5(32'hba9bb8a3),
	.w6(32'hbba52502),
	.w7(32'h3b253a84),
	.w8(32'h3c2f2011),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95666c),
	.w1(32'hbaf4f102),
	.w2(32'hbb98ea90),
	.w3(32'hbbf8dee2),
	.w4(32'hbc13d003),
	.w5(32'h3c4cc582),
	.w6(32'h3bfeaeb7),
	.w7(32'h382ce37a),
	.w8(32'h3c985a7c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcad17c),
	.w1(32'h3c1c9f1e),
	.w2(32'h3c67b223),
	.w3(32'h3b8fe559),
	.w4(32'h3bc84769),
	.w5(32'h3a99e368),
	.w6(32'h3c33a533),
	.w7(32'h3c506fa5),
	.w8(32'hbb013bcf),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b5aa1),
	.w1(32'h3838522f),
	.w2(32'h3bf5e295),
	.w3(32'h3bd4f064),
	.w4(32'h3c448a49),
	.w5(32'h39ab64b3),
	.w6(32'hbb25bde4),
	.w7(32'h3c0285c9),
	.w8(32'h3bc8d756),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c206d12),
	.w1(32'h3bb8237b),
	.w2(32'hbb24a8ad),
	.w3(32'hbbe12647),
	.w4(32'hbc72eef2),
	.w5(32'h3bc1db28),
	.w6(32'h3c019743),
	.w7(32'hbbdd02c1),
	.w8(32'h3bd6728b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4624ed),
	.w1(32'hbb4b7e0e),
	.w2(32'hbb49a09c),
	.w3(32'hba52ec79),
	.w4(32'h3b52485b),
	.w5(32'hba699a44),
	.w6(32'h39228edc),
	.w7(32'h3c05f0a7),
	.w8(32'hbbbca779),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79f1b5),
	.w1(32'hbb6b7bd2),
	.w2(32'hbc1dc87b),
	.w3(32'hbb27c534),
	.w4(32'hbb54c476),
	.w5(32'h3b312344),
	.w6(32'hbbe14003),
	.w7(32'hbbdd44e0),
	.w8(32'h3b649a99),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e2863),
	.w1(32'h3b460783),
	.w2(32'h3b819ea4),
	.w3(32'hbbe39c02),
	.w4(32'h3ae9e0eb),
	.w5(32'hbbd8243a),
	.w6(32'h3b7902b5),
	.w7(32'h3c18b13b),
	.w8(32'hbac80a85),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4e54),
	.w1(32'hbb39aae5),
	.w2(32'hbc4e7385),
	.w3(32'hbc50de81),
	.w4(32'hb95000c9),
	.w5(32'hbad50536),
	.w6(32'hbbceace9),
	.w7(32'hbae439b2),
	.w8(32'hbb974a7c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e3233),
	.w1(32'hbb91fe1a),
	.w2(32'hbbb9d39a),
	.w3(32'h3aa99acb),
	.w4(32'hbbaf3f35),
	.w5(32'hbb65caa1),
	.w6(32'hbc06df5e),
	.w7(32'hbb8bd625),
	.w8(32'hbba30da0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffeb17),
	.w1(32'hbc385b85),
	.w2(32'hbb0ee14f),
	.w3(32'hb98f4ab1),
	.w4(32'hbbb2b4d3),
	.w5(32'hba7c4d0a),
	.w6(32'hbbc951f3),
	.w7(32'hbb93a438),
	.w8(32'h3b39e05b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac66b22),
	.w1(32'hbb8251a3),
	.w2(32'h3c299171),
	.w3(32'hbad354d0),
	.w4(32'hbbc4816d),
	.w5(32'hbbb0b203),
	.w6(32'h3bf546bf),
	.w7(32'hbb00bc9d),
	.w8(32'hba9b3370),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a9032),
	.w1(32'hbbaca369),
	.w2(32'hbc109892),
	.w3(32'hbc05aa85),
	.w4(32'hbbc7f14c),
	.w5(32'hbc17b247),
	.w6(32'hbc26580e),
	.w7(32'h3adb94b5),
	.w8(32'h3ab1724b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1541b9),
	.w1(32'h3b6050c5),
	.w2(32'hbaa39a42),
	.w3(32'hbb9752d8),
	.w4(32'hbc2ace9a),
	.w5(32'h3c0d1c47),
	.w6(32'h3c0b3322),
	.w7(32'hbb1f7f9d),
	.w8(32'h3c2e9d8c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63b927),
	.w1(32'h3c2fd92a),
	.w2(32'h3c12ad8d),
	.w3(32'hbb1b79c0),
	.w4(32'hbb91e9ae),
	.w5(32'h3c4a35fd),
	.w6(32'h3bbd9cbe),
	.w7(32'hba426c53),
	.w8(32'hbc247c90),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba64d7),
	.w1(32'hbc463ba2),
	.w2(32'hba6986ea),
	.w3(32'hbc233205),
	.w4(32'hbc0e2b6e),
	.w5(32'hbc289258),
	.w6(32'hbd006b6a),
	.w7(32'hbbefe2a7),
	.w8(32'hbc40fbef),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c468f),
	.w1(32'h3abe214e),
	.w2(32'h3ade273c),
	.w3(32'h3b94bde9),
	.w4(32'hbba885bb),
	.w5(32'h3aa72ae1),
	.w6(32'hbb1efa38),
	.w7(32'hba9c7378),
	.w8(32'h3be101d3),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf9339),
	.w1(32'hbbcf901b),
	.w2(32'hbb0c7c14),
	.w3(32'h3b52dbbe),
	.w4(32'hbb4d8bf1),
	.w5(32'hbb90ccd6),
	.w6(32'hbba2ec3d),
	.w7(32'h3b915029),
	.w8(32'h3a20c9cd),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f0d7a),
	.w1(32'hba752e03),
	.w2(32'h3b2748e9),
	.w3(32'h39848cc2),
	.w4(32'hbb943799),
	.w5(32'hbb9b2daf),
	.w6(32'hba2dba7e),
	.w7(32'hb9f649c2),
	.w8(32'hbba4a65d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb820d7e),
	.w1(32'hbbcdbb58),
	.w2(32'hbb13ff90),
	.w3(32'h3b5ce64d),
	.w4(32'hbbf9d35a),
	.w5(32'h3afe9d82),
	.w6(32'hbc150eda),
	.w7(32'h3a005db6),
	.w8(32'hb9b3cf79),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a3b1c),
	.w1(32'hbb472d1d),
	.w2(32'hbba72a3f),
	.w3(32'hbbc84be8),
	.w4(32'hbbc17bce),
	.w5(32'hbbf4e86a),
	.w6(32'hbc2ac6be),
	.w7(32'h3a6230a2),
	.w8(32'h3b18d32b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86be99),
	.w1(32'hbc1c3de0),
	.w2(32'hbb8d2c65),
	.w3(32'hbc7b76e1),
	.w4(32'hbc455aea),
	.w5(32'h3b18d7fe),
	.w6(32'hbc038ccc),
	.w7(32'hbb421815),
	.w8(32'h3b2ac60c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b205dd7),
	.w1(32'hbb12209f),
	.w2(32'h39c446ea),
	.w3(32'h3b8c6987),
	.w4(32'h3a9041c3),
	.w5(32'hbbe9e62b),
	.w6(32'hbb43110b),
	.w7(32'h3ab30cba),
	.w8(32'hbc11425f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b7bc8),
	.w1(32'hbb816c49),
	.w2(32'hbb1ad3bf),
	.w3(32'h3b93d0a4),
	.w4(32'hbc80f875),
	.w5(32'hbbb79226),
	.w6(32'hb9fc340d),
	.w7(32'hbc40ec4e),
	.w8(32'hbaa3328b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac9972),
	.w1(32'hbb4fb01d),
	.w2(32'h3b10a048),
	.w3(32'hbbf8b378),
	.w4(32'hb94ed1ae),
	.w5(32'h3bced6a9),
	.w6(32'h3b504d25),
	.w7(32'h3bb38292),
	.w8(32'h3c793e9e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd9dfb),
	.w1(32'h3b12783a),
	.w2(32'hbbc72564),
	.w3(32'h3b7eb0a5),
	.w4(32'hbb62aea4),
	.w5(32'hbb89ee7f),
	.w6(32'h3c0e272e),
	.w7(32'hbbddc965),
	.w8(32'hbb451ff0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00db18),
	.w1(32'h3af34479),
	.w2(32'h3be4c2fa),
	.w3(32'h3acfa723),
	.w4(32'hba5390fe),
	.w5(32'h3bda85b5),
	.w6(32'hbb29c4b0),
	.w7(32'hbaaad8fa),
	.w8(32'h3b5ff9a3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac321fe),
	.w1(32'hbae41911),
	.w2(32'h38f05e20),
	.w3(32'h3bb5642b),
	.w4(32'h3bfd50de),
	.w5(32'hbbcce668),
	.w6(32'h3c431efc),
	.w7(32'h3becd9f1),
	.w8(32'hbc37665b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35a696),
	.w1(32'hbc292625),
	.w2(32'hbc08946f),
	.w3(32'h3c19d00b),
	.w4(32'h3c1fe02c),
	.w5(32'hbb87d7d3),
	.w6(32'hbba8d8e2),
	.w7(32'h3c2a25a0),
	.w8(32'hbc4cf1b1),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e0f43),
	.w1(32'hbb85db07),
	.w2(32'hbaa7a78c),
	.w3(32'hba64685c),
	.w4(32'hbba33c5e),
	.w5(32'h3c169a0c),
	.w6(32'hba0e881c),
	.w7(32'h3bb7b2c0),
	.w8(32'hba80971e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c460c),
	.w1(32'hbc457752),
	.w2(32'hbb15d922),
	.w3(32'h3cbaaba8),
	.w4(32'h3cce1f9c),
	.w5(32'hbbbcc3e3),
	.w6(32'hbad10bd0),
	.w7(32'h3c04a1cc),
	.w8(32'hbab9ea87),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd4cc7),
	.w1(32'h3a9f87d9),
	.w2(32'h3b1e7443),
	.w3(32'hbb326df4),
	.w4(32'h3acceed1),
	.w5(32'hbbf32909),
	.w6(32'h3b7e46e5),
	.w7(32'h380f5092),
	.w8(32'h39332341),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88cb91),
	.w1(32'hbbb008ba),
	.w2(32'hbc18d866),
	.w3(32'hbb960b06),
	.w4(32'hbbc04ab4),
	.w5(32'h3c624c42),
	.w6(32'hbbc1fbe1),
	.w7(32'hbc09a8a8),
	.w8(32'h3c385e49),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff2d2e),
	.w1(32'h3c232d17),
	.w2(32'h3c243f1c),
	.w3(32'h3c159ade),
	.w4(32'h3bfd0cc6),
	.w5(32'hbc0e4f40),
	.w6(32'h3c3ee3e0),
	.w7(32'h3bf7f07d),
	.w8(32'hbba3f846),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75db8d),
	.w1(32'hba9e3327),
	.w2(32'h3c0f6d22),
	.w3(32'hb9e01f1b),
	.w4(32'h3a26b9a0),
	.w5(32'h3a570568),
	.w6(32'h3c246cb4),
	.w7(32'h3c29c061),
	.w8(32'h3c16fa45),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a1cd7),
	.w1(32'h3a9a43df),
	.w2(32'hbae2e66c),
	.w3(32'h3c559614),
	.w4(32'h3c7ae7db),
	.w5(32'h3c5b6cd5),
	.w6(32'h3c435bdd),
	.w7(32'h3c7a7f9f),
	.w8(32'h39c7d214),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27dfe7),
	.w1(32'hbbfb05da),
	.w2(32'hbbae7b38),
	.w3(32'h3c82160e),
	.w4(32'h3c95feef),
	.w5(32'hba67e6a5),
	.w6(32'h3b90bdcd),
	.w7(32'h3c0805fe),
	.w8(32'hbb447b8f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24b988),
	.w1(32'h3ad8d802),
	.w2(32'hba55b76a),
	.w3(32'hbaf559d9),
	.w4(32'h3b1e1e47),
	.w5(32'hbaadce68),
	.w6(32'h3aefa133),
	.w7(32'hba834344),
	.w8(32'h3a8d3c7a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc268394),
	.w1(32'hba989dba),
	.w2(32'h3b8db435),
	.w3(32'h3b5b6207),
	.w4(32'hbb4137c0),
	.w5(32'h3c16d34b),
	.w6(32'hbc13a614),
	.w7(32'hbba415a1),
	.w8(32'h3bf5b1e3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe19af6),
	.w1(32'hbc028a13),
	.w2(32'hb9c4ef6e),
	.w3(32'hbba4a38f),
	.w4(32'h3aa531e8),
	.w5(32'h3c0a228c),
	.w6(32'hbb0222c4),
	.w7(32'hba049e81),
	.w8(32'hba58aa99),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cc46c),
	.w1(32'hbc262299),
	.w2(32'hba18e1e6),
	.w3(32'h3c1e08ae),
	.w4(32'h3c28381c),
	.w5(32'hbbab0893),
	.w6(32'hbc23474d),
	.w7(32'hba27f823),
	.w8(32'hb8be4205),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c395ff5),
	.w1(32'h3c517af0),
	.w2(32'hbbb3e25b),
	.w3(32'hbcba218c),
	.w4(32'hbc9b2198),
	.w5(32'hbb27b55c),
	.w6(32'hbb4b0f8c),
	.w7(32'hbba999b4),
	.w8(32'h3b3d5e50),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0886af),
	.w1(32'hbb359aa6),
	.w2(32'h39851e50),
	.w3(32'h3ad2ef93),
	.w4(32'h3a8dc34d),
	.w5(32'hbbb27d1b),
	.w6(32'hbb3be423),
	.w7(32'h3baccf09),
	.w8(32'h3af9b9d1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad062c8),
	.w1(32'hba1cf3ce),
	.w2(32'h39c73ba8),
	.w3(32'hbbb5a293),
	.w4(32'hbb923162),
	.w5(32'hbb6b12ac),
	.w6(32'h3b8a2fce),
	.w7(32'hbb0665fe),
	.w8(32'hbb72d64f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc368fc),
	.w1(32'h3b6d86d3),
	.w2(32'h3bfee655),
	.w3(32'h3bb085bc),
	.w4(32'h3a67fce8),
	.w5(32'h3b49e329),
	.w6(32'h3c60206a),
	.w7(32'hbb301bef),
	.w8(32'h3ba1c017),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaace721),
	.w1(32'hbc377080),
	.w2(32'h3b5c4119),
	.w3(32'h3ba40476),
	.w4(32'h3c670bbb),
	.w5(32'h3c2e66a7),
	.w6(32'h3c2ed3f1),
	.w7(32'h3c9879ae),
	.w8(32'h3c161f4a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9a232),
	.w1(32'hbc1131d7),
	.w2(32'hbae594ef),
	.w3(32'hbc2c70fa),
	.w4(32'hbc37e23d),
	.w5(32'hbc6994e6),
	.w6(32'hbba64474),
	.w7(32'hba34530f),
	.w8(32'hbc1b0c6a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ae89e),
	.w1(32'hbc96a12a),
	.w2(32'hbb192ce1),
	.w3(32'hbbed9f57),
	.w4(32'hbc1415cc),
	.w5(32'hba832a0b),
	.w6(32'hbc707c9e),
	.w7(32'hbc822bfb),
	.w8(32'hbb900f15),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71d479),
	.w1(32'hba897b03),
	.w2(32'hbbe8abb7),
	.w3(32'h3add78a0),
	.w4(32'hbc016ffa),
	.w5(32'hbc24bd18),
	.w6(32'hbc592698),
	.w7(32'hbc9bdc6d),
	.w8(32'hbc483840),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd28f8),
	.w1(32'hbbc58a9d),
	.w2(32'h3c35700c),
	.w3(32'hbb8b3bbd),
	.w4(32'h3a4869e8),
	.w5(32'h3b885524),
	.w6(32'hbb7791e9),
	.w7(32'h3b8d9850),
	.w8(32'hbbe7cf89),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22c108),
	.w1(32'hbc0624b3),
	.w2(32'hbb0fed7a),
	.w3(32'hbb158731),
	.w4(32'hbc0dda10),
	.w5(32'h3c86f206),
	.w6(32'hbb9b5d33),
	.w7(32'h3bb7be1f),
	.w8(32'h3c151494),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997b864),
	.w1(32'h3b719708),
	.w2(32'h3b12c8b5),
	.w3(32'h3c0265be),
	.w4(32'h3b9e031f),
	.w5(32'hbbe2164a),
	.w6(32'h3c2e1214),
	.w7(32'h3c1f25a4),
	.w8(32'hbb273b45),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e497c),
	.w1(32'hbbe88604),
	.w2(32'h3b186906),
	.w3(32'hbb0504d6),
	.w4(32'hbbde39ae),
	.w5(32'hba7cc9a5),
	.w6(32'hbc09fcba),
	.w7(32'hbc30a931),
	.w8(32'hba439e0a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b18381),
	.w1(32'h3a999aee),
	.w2(32'h3b1dc91d),
	.w3(32'hbaa29be3),
	.w4(32'hbb27cc2a),
	.w5(32'hba2b2915),
	.w6(32'hbb47befd),
	.w7(32'hbb1a3862),
	.w8(32'hbae6275d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a20c6),
	.w1(32'hbbbe9043),
	.w2(32'h3bf4f077),
	.w3(32'hbb957c72),
	.w4(32'hbafc006d),
	.w5(32'h3b925a48),
	.w6(32'hba826312),
	.w7(32'hbb06c997),
	.w8(32'h3b68c5bd),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4393c),
	.w1(32'hbbc5b657),
	.w2(32'hbafef0a4),
	.w3(32'hbb16d844),
	.w4(32'hbb2ccc37),
	.w5(32'hbc24886c),
	.w6(32'h3b98bedc),
	.w7(32'h392e0cd0),
	.w8(32'h3a88ebb1),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50d978),
	.w1(32'h3bd2dd82),
	.w2(32'h3bb30cf7),
	.w3(32'hbc017407),
	.w4(32'hbbf48d68),
	.w5(32'hba26d36c),
	.w6(32'h3c763f85),
	.w7(32'h3a0c75d6),
	.w8(32'h3b9e2236),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ff31d),
	.w1(32'hbc4c5a5e),
	.w2(32'hbc1dbf60),
	.w3(32'hbc3bc95b),
	.w4(32'hbbd0c505),
	.w5(32'h3a3bdbaf),
	.w6(32'h3aa4139a),
	.w7(32'h3984accb),
	.w8(32'h3ac54d4e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00be4b),
	.w1(32'hbc058809),
	.w2(32'hbb4b5006),
	.w3(32'hb9920e80),
	.w4(32'h3b03d1a6),
	.w5(32'h3b5aaae5),
	.w6(32'hbb0dc02a),
	.w7(32'h391da610),
	.w8(32'h3c12aa7d),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6ab26),
	.w1(32'h3b85a3e8),
	.w2(32'h3b484833),
	.w3(32'hba8ca777),
	.w4(32'hbaadcc58),
	.w5(32'h3bd42064),
	.w6(32'h3b96d78c),
	.w7(32'hba85701b),
	.w8(32'hba2a6d45),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba362df5),
	.w1(32'hbaaeeddc),
	.w2(32'h3ac85b8b),
	.w3(32'h3acb98da),
	.w4(32'h3bdf3ea6),
	.w5(32'hbb36f71e),
	.w6(32'hbb10daec),
	.w7(32'h3bdcdadc),
	.w8(32'h3a9aa899),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc280803),
	.w1(32'hbbc08e77),
	.w2(32'hbbd70001),
	.w3(32'hbb327127),
	.w4(32'hbb60bc1d),
	.w5(32'h3af0098a),
	.w6(32'h3b882b2a),
	.w7(32'h3a9a231e),
	.w8(32'h3b9332a1),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a246f92),
	.w1(32'hba67d789),
	.w2(32'hb980d24d),
	.w3(32'h3b7319b0),
	.w4(32'h39363861),
	.w5(32'hb972c238),
	.w6(32'h3c5d157a),
	.w7(32'h3b836a9c),
	.w8(32'hb9c7da55),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48f1b0),
	.w1(32'h3ab6ad79),
	.w2(32'h3aa274f5),
	.w3(32'h3a82044c),
	.w4(32'hbae7c5e6),
	.w5(32'h3b9a42f6),
	.w6(32'hb8992e2e),
	.w7(32'hbae5cef9),
	.w8(32'h3a1c6a17),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca17a7),
	.w1(32'hba8f0394),
	.w2(32'hb9c25e95),
	.w3(32'h3ba3ea5e),
	.w4(32'h3ba07a44),
	.w5(32'hbb1c8fbc),
	.w6(32'hb78a621d),
	.w7(32'h3b75ea4e),
	.w8(32'hbb483f96),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0d2a1),
	.w1(32'h3a1b803a),
	.w2(32'h39c5fcb8),
	.w3(32'h3b1bf33b),
	.w4(32'hbb1c7c25),
	.w5(32'hba6ab93f),
	.w6(32'hb9f17e29),
	.w7(32'h39cf6857),
	.w8(32'hbb413366),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c91f4),
	.w1(32'h3bc79199),
	.w2(32'h3c3e4a7c),
	.w3(32'hbb3c8a23),
	.w4(32'hb9dd0f67),
	.w5(32'h3c312576),
	.w6(32'hba359c90),
	.w7(32'h3bd94cd9),
	.w8(32'h3c86a5b4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47032b),
	.w1(32'h38a307af),
	.w2(32'h3b7cf225),
	.w3(32'h390d6cd4),
	.w4(32'h3b1caece),
	.w5(32'h3bc98f02),
	.w6(32'hbaf5b7db),
	.w7(32'h3bd7f270),
	.w8(32'h3c8a509c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f9f04),
	.w1(32'h3a42535e),
	.w2(32'h3bb97283),
	.w3(32'hbbaba7ca),
	.w4(32'h3b3db750),
	.w5(32'h3b9a7a77),
	.w6(32'h3d089008),
	.w7(32'h3ca1ba83),
	.w8(32'h3bdb98ce),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996ad4d),
	.w1(32'hbbbd747b),
	.w2(32'hbb0b3eb2),
	.w3(32'h3b6a4eeb),
	.w4(32'h3c10fd0a),
	.w5(32'hbb0ae67e),
	.w6(32'h3b990ec4),
	.w7(32'h3b91eae4),
	.w8(32'h3aeaeaf7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae57290),
	.w1(32'h3ba29f6b),
	.w2(32'h3bedf1e1),
	.w3(32'hb9359bba),
	.w4(32'hbb1ca5ac),
	.w5(32'h3a27fb0b),
	.w6(32'h3a4ac81e),
	.w7(32'h38af0f80),
	.w8(32'h3b429146),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b9433),
	.w1(32'h3af70df8),
	.w2(32'h3aff7de7),
	.w3(32'h3b1348d7),
	.w4(32'h3b9a34d2),
	.w5(32'h3a7e67bd),
	.w6(32'h3abde6f8),
	.w7(32'h3bac3a6e),
	.w8(32'h3a238a5c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2aa52),
	.w1(32'h3bbbed1f),
	.w2(32'hb9b26877),
	.w3(32'hba3ca106),
	.w4(32'hbbcddce4),
	.w5(32'hbac2826a),
	.w6(32'h3b50328d),
	.w7(32'hbbae5336),
	.w8(32'hbbb16036),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc094bc9),
	.w1(32'hbc23dc5f),
	.w2(32'hbb211e38),
	.w3(32'hbbb9ebfe),
	.w4(32'hbc079513),
	.w5(32'hb9875de7),
	.w6(32'hbbe8e3c1),
	.w7(32'hbbf221b3),
	.w8(32'h3b4c35d5),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ad934),
	.w1(32'hbbbff602),
	.w2(32'hbbb94591),
	.w3(32'h3ab4b93c),
	.w4(32'hba2ab2c8),
	.w5(32'h3adc0904),
	.w6(32'h387018c5),
	.w7(32'hbb6fb58d),
	.w8(32'h396a208f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0f5b2),
	.w1(32'h3be61e3e),
	.w2(32'h3bc57086),
	.w3(32'h3bba7da2),
	.w4(32'h3a9856e1),
	.w5(32'h3b09e130),
	.w6(32'hbb0aea0d),
	.w7(32'hbaf87214),
	.w8(32'h3b82bb76),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba90e77),
	.w1(32'hbb8111b5),
	.w2(32'hbbbdfe72),
	.w3(32'h39fc4efd),
	.w4(32'h3b6e4697),
	.w5(32'hbb724ed5),
	.w6(32'hbb8e10fd),
	.w7(32'hbb88c997),
	.w8(32'h3aa787a1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d8c56),
	.w1(32'h3a82395d),
	.w2(32'h399dce72),
	.w3(32'hbb953767),
	.w4(32'hbba6300b),
	.w5(32'hbb14710d),
	.w6(32'h3cfa1804),
	.w7(32'h3c4e1a29),
	.w8(32'hba93d8de),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a44ae),
	.w1(32'h3bda770d),
	.w2(32'hbafcdba1),
	.w3(32'h3c0b1b40),
	.w4(32'h3be1808e),
	.w5(32'hbbd0d8dd),
	.w6(32'hbb0c20ea),
	.w7(32'h39f31172),
	.w8(32'h3c3e90de),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5edf09),
	.w1(32'h3b9cbe9f),
	.w2(32'h3b1a0087),
	.w3(32'hbc1de6d4),
	.w4(32'hbbd2a430),
	.w5(32'h3bff0899),
	.w6(32'h3cf09f20),
	.w7(32'h3c22400d),
	.w8(32'h3c58d44a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b7213),
	.w1(32'hbc1e0612),
	.w2(32'hbb5d0b6b),
	.w3(32'hbc30730a),
	.w4(32'hbc25e3cb),
	.w5(32'h3989d3d2),
	.w6(32'h3ccdf602),
	.w7(32'h3ca40962),
	.w8(32'h3c695dec),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45d3ff),
	.w1(32'hbac701dc),
	.w2(32'hbb449c7b),
	.w3(32'h3b05d3ef),
	.w4(32'hba8ebfae),
	.w5(32'hb9b6e3d5),
	.w6(32'h3c681566),
	.w7(32'h3b5ab62a),
	.w8(32'hbaf56f59),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc041cec),
	.w1(32'hbbf4820f),
	.w2(32'hbb472171),
	.w3(32'h3bd525f9),
	.w4(32'hbb77cedf),
	.w5(32'h3bccdc5b),
	.w6(32'h3bb91757),
	.w7(32'hbb5e0c65),
	.w8(32'h3a4b8774),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule