module layer_10_featuremap_161(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acdae5),
	.w1(32'hbb8dd5fe),
	.w2(32'hbc3cab4e),
	.w3(32'h3b10355c),
	.w4(32'hb9d5cc1b),
	.w5(32'h39e0fd34),
	.w6(32'hbc5cc5f9),
	.w7(32'hbc2235dd),
	.w8(32'hbc4d1baa),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21f93a),
	.w1(32'h3b6628d0),
	.w2(32'hba909f57),
	.w3(32'hbc3fa06e),
	.w4(32'h3bf74e79),
	.w5(32'h3b1ec5e8),
	.w6(32'hba716aec),
	.w7(32'hbb5e3511),
	.w8(32'hbb62d4fb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5ebc0),
	.w1(32'h3b958f59),
	.w2(32'h3a1e22d8),
	.w3(32'h3af8db1a),
	.w4(32'h3b09406f),
	.w5(32'hbb41051b),
	.w6(32'h3ae54949),
	.w7(32'h3a997d30),
	.w8(32'h3b4801c2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b286bf1),
	.w1(32'hbc4bf5f4),
	.w2(32'hbb1b4633),
	.w3(32'h3a8821d0),
	.w4(32'hbb433d54),
	.w5(32'hbb5fcdf0),
	.w6(32'hbb423fb9),
	.w7(32'h3b2c6232),
	.w8(32'hb8cbe1ec),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf418b5),
	.w1(32'hba8e9648),
	.w2(32'hba9d8952),
	.w3(32'hbb0d96f3),
	.w4(32'hbc0d9a57),
	.w5(32'hbb6131a3),
	.w6(32'hb998c334),
	.w7(32'hbb7db1f4),
	.w8(32'hbb8280d6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78c411),
	.w1(32'h3b029c22),
	.w2(32'h3b8741a7),
	.w3(32'h3a3d6305),
	.w4(32'h3b9f9554),
	.w5(32'h3bf9e16b),
	.w6(32'h3bac9039),
	.w7(32'h3b035167),
	.w8(32'hbaafe3f5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b95a1),
	.w1(32'hbbdc94fa),
	.w2(32'hbb0fe314),
	.w3(32'h3bb93540),
	.w4(32'h3b0338a7),
	.w5(32'h3c723582),
	.w6(32'hbb9239a5),
	.w7(32'hbbd76b2e),
	.w8(32'h3bbfcad0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad492f),
	.w1(32'hbb265d74),
	.w2(32'h3c1e1781),
	.w3(32'hbc7a4c50),
	.w4(32'hbc573bcb),
	.w5(32'hbc2f1c2a),
	.w6(32'hbb9b9a53),
	.w7(32'h3b9d1786),
	.w8(32'hbb7fcc80),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c2cd8),
	.w1(32'h3ae5d926),
	.w2(32'hb981b950),
	.w3(32'hb83e8b9a),
	.w4(32'h39f3dc5c),
	.w5(32'h3a76c7ed),
	.w6(32'h3afe32fb),
	.w7(32'h3a009139),
	.w8(32'hb9e01cd2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c5fa8),
	.w1(32'h3c0ef955),
	.w2(32'h3c44dbe6),
	.w3(32'hbb9e0149),
	.w4(32'h3be2216a),
	.w5(32'h3c1ef05d),
	.w6(32'h3a2a258c),
	.w7(32'hba8c0d59),
	.w8(32'h3b2df957),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bac2bd),
	.w1(32'hbc3ecedb),
	.w2(32'hbc49f848),
	.w3(32'hba7db55e),
	.w4(32'h3a73a3e2),
	.w5(32'hbaf93db8),
	.w6(32'h3a86a679),
	.w7(32'hbb299c49),
	.w8(32'hbb0bd894),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc807aaf),
	.w1(32'hbc004131),
	.w2(32'h3bc25a46),
	.w3(32'hbbdafcd4),
	.w4(32'hbbcc3009),
	.w5(32'hbb006758),
	.w6(32'hbbcac959),
	.w7(32'h3b47b8ba),
	.w8(32'h3bd4e937),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86db81),
	.w1(32'h3a88b193),
	.w2(32'h3b936ad8),
	.w3(32'hbc5ce2da),
	.w4(32'hbb64bceb),
	.w5(32'h3b5706c7),
	.w6(32'hbbe1a1ba),
	.w7(32'hb9ec41fc),
	.w8(32'h3b4aff81),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac55805),
	.w1(32'hba2c2256),
	.w2(32'h3aaf7d55),
	.w3(32'hba839d1f),
	.w4(32'hbb8438b1),
	.w5(32'hbc4e041c),
	.w6(32'h3b7771f1),
	.w7(32'h3c778fe4),
	.w8(32'h3bad7b9f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedf8d3),
	.w1(32'hbc340d11),
	.w2(32'h3a8d8252),
	.w3(32'hbbe7a553),
	.w4(32'hbc14bdf9),
	.w5(32'hbc7ae124),
	.w6(32'hbb9344d5),
	.w7(32'hbbf58137),
	.w8(32'hbb87bb34),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3872a5),
	.w1(32'h3c849cde),
	.w2(32'h3c2f6d8e),
	.w3(32'hbc3e1b4a),
	.w4(32'h3b843847),
	.w5(32'h3bbde6e3),
	.w6(32'hb982d5ed),
	.w7(32'hbb00df70),
	.w8(32'hbb0594d0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01e4a6),
	.w1(32'h3af7f708),
	.w2(32'h39bbfdbb),
	.w3(32'h3b0d0b05),
	.w4(32'hba80d1ea),
	.w5(32'h3a3574e6),
	.w6(32'hbb48c49f),
	.w7(32'hbb590b8e),
	.w8(32'hbacdbe92),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb970dc8),
	.w1(32'h3c3c4df9),
	.w2(32'h3cba3818),
	.w3(32'hbb42aaac),
	.w4(32'h3bb82077),
	.w5(32'h3c9c50b5),
	.w6(32'hbb8eed4b),
	.w7(32'hbb3f918f),
	.w8(32'h3ba96942),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb380f01),
	.w1(32'h3b9bd234),
	.w2(32'h3c2adf10),
	.w3(32'h384933aa),
	.w4(32'h3b170439),
	.w5(32'h3c015e63),
	.w6(32'hbb58135d),
	.w7(32'h3afe0618),
	.w8(32'h3b928152),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada40f4),
	.w1(32'h39b55a18),
	.w2(32'hbacc0506),
	.w3(32'h3b0dde0d),
	.w4(32'h39919e69),
	.w5(32'h3892b6bf),
	.w6(32'h3a64169c),
	.w7(32'hb9971861),
	.w8(32'hba959f7d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1890f0),
	.w1(32'hba07ccaa),
	.w2(32'h3a432227),
	.w3(32'h38f7ec86),
	.w4(32'hbb8d5d9a),
	.w5(32'hbb87b9bf),
	.w6(32'h39d08b8e),
	.w7(32'h3999f111),
	.w8(32'h3a3b75d7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd3f47),
	.w1(32'h3b7247b2),
	.w2(32'hbc1b4145),
	.w3(32'hba0fde32),
	.w4(32'h3a29d42a),
	.w5(32'hbb862e17),
	.w6(32'h39b822d3),
	.w7(32'h39e6707f),
	.w8(32'hbb4eef39),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc058485),
	.w1(32'h3c945510),
	.w2(32'h3c683f17),
	.w3(32'hbbaf657f),
	.w4(32'hbae42414),
	.w5(32'h3b26f792),
	.w6(32'hbc1f00ac),
	.w7(32'hbbfab860),
	.w8(32'h3ba25c8f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70fa04),
	.w1(32'h3af2aa19),
	.w2(32'hb9e6905c),
	.w3(32'hbaf1a347),
	.w4(32'hbb45a6e3),
	.w5(32'hbba29821),
	.w6(32'hba98590e),
	.w7(32'h3b3b13d5),
	.w8(32'hbb00a910),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09efa4),
	.w1(32'h3b35f88e),
	.w2(32'hbc0fa8ac),
	.w3(32'h3b5d05db),
	.w4(32'h3a83a59a),
	.w5(32'hbc238ce5),
	.w6(32'h3b0c26d6),
	.w7(32'hb9aa5c95),
	.w8(32'hbb3b54b6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df2d1f),
	.w1(32'h3bdea4d1),
	.w2(32'hbb4471e8),
	.w3(32'h3af9658b),
	.w4(32'h3bdaeca4),
	.w5(32'hbaaafac4),
	.w6(32'hbae2674b),
	.w7(32'hbbd5b6f3),
	.w8(32'hba9b9f7a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba572229),
	.w1(32'hb996e13c),
	.w2(32'hbb03e182),
	.w3(32'hb9baab6f),
	.w4(32'hba3dbf6b),
	.w5(32'hb8d8817a),
	.w6(32'h3a46b0e6),
	.w7(32'hba716970),
	.w8(32'hbad1105c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a33dc),
	.w1(32'h3ca77da2),
	.w2(32'h3ad6a761),
	.w3(32'hbc4b7aa9),
	.w4(32'h3bfabab6),
	.w5(32'h3b960615),
	.w6(32'h3bae1a0b),
	.w7(32'h3c1721de),
	.w8(32'h3ae46f99),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc194e6a),
	.w1(32'hbb861c32),
	.w2(32'hbabc15ff),
	.w3(32'hbb34a946),
	.w4(32'hbb03df9f),
	.w5(32'h392f9c04),
	.w6(32'hbb79c9b5),
	.w7(32'hbb76eb71),
	.w8(32'hba0f9a7e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39890ea7),
	.w1(32'h3c137146),
	.w2(32'hbb6d371f),
	.w3(32'h3a38c935),
	.w4(32'h3baf4b2d),
	.w5(32'hbbb16a47),
	.w6(32'h3b48b036),
	.w7(32'h3c3672f4),
	.w8(32'hbb44311b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf3dce),
	.w1(32'hba832501),
	.w2(32'hba9abea8),
	.w3(32'hbb2cdefd),
	.w4(32'hbb17b98d),
	.w5(32'hbb1b5b30),
	.w6(32'h39db3471),
	.w7(32'hb8d5f578),
	.w8(32'hb978d661),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98954f6),
	.w1(32'hbae3376b),
	.w2(32'hbb26ad09),
	.w3(32'hba120bb1),
	.w4(32'hbacc8960),
	.w5(32'hbb0b7010),
	.w6(32'hba9277d2),
	.w7(32'hbb16ea2c),
	.w8(32'hba09212a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d86ed),
	.w1(32'hbb84601a),
	.w2(32'h3b148dc5),
	.w3(32'hbb532e52),
	.w4(32'hbb6fe95f),
	.w5(32'hbab13bc5),
	.w6(32'hbb5e0146),
	.w7(32'hb9d3475c),
	.w8(32'hbb01d218),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb718520),
	.w1(32'h3a7e0fbf),
	.w2(32'hbaf91bed),
	.w3(32'hba36da2f),
	.w4(32'h3c1033b8),
	.w5(32'h3bda3601),
	.w6(32'h3b4f10cd),
	.w7(32'h389c6f34),
	.w8(32'h3b38c7af),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb972b5f),
	.w1(32'h3ad54c07),
	.w2(32'h3b42b2cb),
	.w3(32'hba0db592),
	.w4(32'h3bc65ad3),
	.w5(32'h3ba42838),
	.w6(32'hbb21f208),
	.w7(32'hbc0b65bb),
	.w8(32'hbb08426e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee72c7),
	.w1(32'hbb2080e9),
	.w2(32'hba4e2a8d),
	.w3(32'h39486c2d),
	.w4(32'hbb77a63b),
	.w5(32'hbab7127b),
	.w6(32'hbb18af92),
	.w7(32'hbb272d9d),
	.w8(32'h3b2411b5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bd8e4),
	.w1(32'hbc6fcecb),
	.w2(32'h3a90045c),
	.w3(32'hbbc339af),
	.w4(32'hbc178316),
	.w5(32'hbc194f11),
	.w6(32'h3b2c835f),
	.w7(32'hbc40dd7d),
	.w8(32'hbc056d3d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaa7bc),
	.w1(32'h3b443891),
	.w2(32'hbc97428c),
	.w3(32'h3b8773c5),
	.w4(32'h3bd09e33),
	.w5(32'hbc0c2f86),
	.w6(32'h399971d5),
	.w7(32'hbb4ebf02),
	.w8(32'hbbfdf107),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfaf09a),
	.w1(32'h3c65ced3),
	.w2(32'hbb2424a1),
	.w3(32'h3ae40d3c),
	.w4(32'h3bcb6650),
	.w5(32'hbb0faf3e),
	.w6(32'h3c105620),
	.w7(32'h3bcec75b),
	.w8(32'hbaf90dd8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48f375),
	.w1(32'hba5754b5),
	.w2(32'hbb0afdd2),
	.w3(32'h394997ac),
	.w4(32'h3a1f4fdc),
	.w5(32'hbaa6935d),
	.w6(32'hbaa3b20c),
	.w7(32'hbb070fd3),
	.w8(32'hbb087c99),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeea6f0),
	.w1(32'hba56823d),
	.w2(32'h3ac3165c),
	.w3(32'h39c7b3f5),
	.w4(32'hbbcaf1f0),
	.w5(32'hbbaefa6d),
	.w6(32'hbb8324af),
	.w7(32'hba52e110),
	.w8(32'hbb0226bf),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70b044),
	.w1(32'hbb6e8a29),
	.w2(32'hbb6ee4bf),
	.w3(32'hbbe51386),
	.w4(32'h3a400955),
	.w5(32'hba801842),
	.w6(32'hbb330315),
	.w7(32'hbb7b0782),
	.w8(32'hbaaa15d1),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb24ea6),
	.w1(32'hbb0e4459),
	.w2(32'hbb7483f8),
	.w3(32'hba0f13d0),
	.w4(32'hbaaca5f5),
	.w5(32'hbb45e246),
	.w6(32'hb9e553ba),
	.w7(32'hb9c49116),
	.w8(32'h3a8f3605),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ae812),
	.w1(32'h3c7648e6),
	.w2(32'h3c8e5eb0),
	.w3(32'hbbc5e1d0),
	.w4(32'h3c64513d),
	.w5(32'h3cb89e20),
	.w6(32'hbac17384),
	.w7(32'hb98f89b5),
	.w8(32'h3c209f4e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e653b),
	.w1(32'h3b17324d),
	.w2(32'hbc4e6bf3),
	.w3(32'hbb412f66),
	.w4(32'hba1a8a30),
	.w5(32'hbc0165a5),
	.w6(32'hbb44370e),
	.w7(32'h3b566729),
	.w8(32'hbb752a77),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dd391),
	.w1(32'h3b65de79),
	.w2(32'hbbfbd16b),
	.w3(32'hbc04faea),
	.w4(32'hbc051371),
	.w5(32'hbc1a4a49),
	.w6(32'hbc0c11ce),
	.w7(32'h3a1dc734),
	.w8(32'hbbe25497),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8b866),
	.w1(32'hba29180c),
	.w2(32'h3c541717),
	.w3(32'hbba030af),
	.w4(32'hbb8251dc),
	.w5(32'hbbba6f43),
	.w6(32'hbab36a25),
	.w7(32'h3b21175f),
	.w8(32'hbb9636d0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79feec),
	.w1(32'h3a84caba),
	.w2(32'h3ca6cb41),
	.w3(32'hbc4e3dd4),
	.w4(32'h3aa2568f),
	.w5(32'h3c81fee1),
	.w6(32'hbbde3481),
	.w7(32'h3b899d41),
	.w8(32'h3c44fc30),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc336e),
	.w1(32'hbafd3a73),
	.w2(32'hbb87f1e1),
	.w3(32'h3a6a57c1),
	.w4(32'h38e29909),
	.w5(32'hbaf82dae),
	.w6(32'hbaa58019),
	.w7(32'hbaf7813f),
	.w8(32'hba91e040),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb369b1e),
	.w1(32'h39de0bf1),
	.w2(32'hbadc0896),
	.w3(32'hbaea07d0),
	.w4(32'hbb42d091),
	.w5(32'hbbb57e95),
	.w6(32'h3aeafe28),
	.w7(32'h3bc2cae4),
	.w8(32'h3a9c9815),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41a743),
	.w1(32'h3b215cab),
	.w2(32'h3a95023a),
	.w3(32'hb9995820),
	.w4(32'hba88004c),
	.w5(32'hbbd5dc7c),
	.w6(32'hba71399c),
	.w7(32'h3b00db43),
	.w8(32'hbaaa895e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cbf1c),
	.w1(32'h3af048e0),
	.w2(32'h3c0c80ca),
	.w3(32'h39e4c415),
	.w4(32'hbb091df1),
	.w5(32'hbbebc507),
	.w6(32'hbc42acf4),
	.w7(32'hbc5d62dc),
	.w8(32'hbbcd97d8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a46ec),
	.w1(32'h3ba37e0b),
	.w2(32'h3c498536),
	.w3(32'hbc1659b8),
	.w4(32'h3c0300bf),
	.w5(32'h3c6d102a),
	.w6(32'h3a7665a9),
	.w7(32'h3aad0fe9),
	.w8(32'h3b51aa24),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad5b7c),
	.w1(32'h3941d1b3),
	.w2(32'h3c8c53c0),
	.w3(32'hbad725a6),
	.w4(32'hbb32e7e5),
	.w5(32'h3c5cc97b),
	.w6(32'hbc258b0f),
	.w7(32'hbba99ab8),
	.w8(32'h3b949a7a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82e891),
	.w1(32'h3c071138),
	.w2(32'h3c2eeb63),
	.w3(32'hbab0d102),
	.w4(32'h3bcd0c87),
	.w5(32'h3bdedad9),
	.w6(32'h3a5d92bf),
	.w7(32'h39d63e6e),
	.w8(32'h3b0897f0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6318e6),
	.w1(32'hbaa88fea),
	.w2(32'hbb826c33),
	.w3(32'h3ad4501f),
	.w4(32'hbbea1ad8),
	.w5(32'hbbe694ea),
	.w6(32'h3973e8f5),
	.w7(32'h3a54e428),
	.w8(32'hba4f566a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71e2b1),
	.w1(32'h3becc1f8),
	.w2(32'h3b9fbcf9),
	.w3(32'hbbd65a76),
	.w4(32'h3ae4e192),
	.w5(32'hba7b288e),
	.w6(32'h3b5229a2),
	.w7(32'h3bbd099e),
	.w8(32'h3b8e0b02),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a5cf2),
	.w1(32'hbb9e9e1d),
	.w2(32'hbc03dcd4),
	.w3(32'hba6ef107),
	.w4(32'hbc26058c),
	.w5(32'hbc5dec32),
	.w6(32'hbc136364),
	.w7(32'hbb20760f),
	.w8(32'hbb16bf39),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99122ed),
	.w1(32'hbb4accc4),
	.w2(32'h3ae0bb37),
	.w3(32'hbb8c7bd1),
	.w4(32'h3ac10d1a),
	.w5(32'h3b652916),
	.w6(32'hbb87687a),
	.w7(32'hbba115f9),
	.w8(32'hb91094a9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab844be),
	.w1(32'h3ab5be20),
	.w2(32'h3a5b886e),
	.w3(32'hbacc4459),
	.w4(32'hba404743),
	.w5(32'h39b09b14),
	.w6(32'h3b115f50),
	.w7(32'h3b530103),
	.w8(32'h3aadabc3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba43bed),
	.w1(32'h3bc98a4b),
	.w2(32'h3ba5286a),
	.w3(32'hbacc5bef),
	.w4(32'h3b54bb21),
	.w5(32'h3b13c8d4),
	.w6(32'hbaf49c26),
	.w7(32'hba8c8813),
	.w8(32'h39faa62d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf9618),
	.w1(32'h3c244775),
	.w2(32'h3b4c651d),
	.w3(32'hbb950dbd),
	.w4(32'h3acd080e),
	.w5(32'h3ab080f4),
	.w6(32'h3aa58b16),
	.w7(32'h3c07c50e),
	.w8(32'h3b57dc3f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb238451),
	.w1(32'h39665b1c),
	.w2(32'h3a845eff),
	.w3(32'hbadd5145),
	.w4(32'h3b633e94),
	.w5(32'h3b842af1),
	.w6(32'hbb6f1db9),
	.w7(32'hbb60a80a),
	.w8(32'hbb4136fa),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a825231),
	.w1(32'h3aa1be53),
	.w2(32'h3b1a1550),
	.w3(32'h3b17f963),
	.w4(32'h3ba6d7b8),
	.w5(32'h3ba0c046),
	.w6(32'hb98ab015),
	.w7(32'hbb4dcc31),
	.w8(32'hb96d9a59),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3865aefc),
	.w1(32'h3b46ae2e),
	.w2(32'h3b2aa586),
	.w3(32'hbabf77ff),
	.w4(32'h3ab808b3),
	.w5(32'h3b5381a1),
	.w6(32'h3afb30b0),
	.w7(32'hbb5fe425),
	.w8(32'hbbb96f8f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9afee3),
	.w1(32'hbb701ac3),
	.w2(32'hbbc5bd1e),
	.w3(32'hba3827a0),
	.w4(32'hbbc418e5),
	.w5(32'hbc03b498),
	.w6(32'hbb8151ca),
	.w7(32'h3a69bacb),
	.w8(32'hbb74dda1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd07589),
	.w1(32'hba1b3975),
	.w2(32'h3caceb14),
	.w3(32'hbca6ad2a),
	.w4(32'hbac3bad9),
	.w5(32'h3c5e5d4e),
	.w6(32'hbc1f3fa3),
	.w7(32'hbb81eb39),
	.w8(32'h3bb66949),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a3e7d),
	.w1(32'h3ca48d8e),
	.w2(32'h3cc76d6d),
	.w3(32'hbc470ca1),
	.w4(32'hbbd3d220),
	.w5(32'hbad67eff),
	.w6(32'hbc62adca),
	.w7(32'h3939e164),
	.w8(32'h3b2639d8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7a8d9),
	.w1(32'h3c72b828),
	.w2(32'h3cbdf767),
	.w3(32'hbaf972e1),
	.w4(32'h3ba6633d),
	.w5(32'h3c43ef4e),
	.w6(32'h3b2d8490),
	.w7(32'h3c183189),
	.w8(32'h3c4ba0ef),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23901a),
	.w1(32'hb9b6d7d2),
	.w2(32'hbccdb514),
	.w3(32'h3b59c61f),
	.w4(32'hbc5e2aac),
	.w5(32'hbd1b4bc3),
	.w6(32'hba0c9207),
	.w7(32'h3b81b53d),
	.w8(32'hbc7fed87),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15b89a),
	.w1(32'hba64c432),
	.w2(32'h3af7dd0e),
	.w3(32'hbc234717),
	.w4(32'h3b98535e),
	.w5(32'h3bd76843),
	.w6(32'hbbb2739f),
	.w7(32'hbc16bde4),
	.w8(32'hbabbaeaa),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b172b4a),
	.w1(32'hbaa139e3),
	.w2(32'h3a01c164),
	.w3(32'h3b3f32c6),
	.w4(32'hbb0a1482),
	.w5(32'hba10a6e1),
	.w6(32'hb9596271),
	.w7(32'hb58d9cde),
	.w8(32'h3959e2ee),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe3544),
	.w1(32'h394fb747),
	.w2(32'h3a8f98f1),
	.w3(32'h3afb7707),
	.w4(32'hba8af901),
	.w5(32'hbaa6fd9a),
	.w6(32'h3a97d9d7),
	.w7(32'h3a904dbc),
	.w8(32'h3a0c86e4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a4c4b),
	.w1(32'hbaa11dc7),
	.w2(32'h3ae83176),
	.w3(32'hbaf7b1e9),
	.w4(32'hbaf177ce),
	.w5(32'hba851609),
	.w6(32'hbb26dcfb),
	.w7(32'h39d97b4d),
	.w8(32'h3b0e6897),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bd233),
	.w1(32'hb938d631),
	.w2(32'h3b4261b2),
	.w3(32'hbab985ba),
	.w4(32'h3a813409),
	.w5(32'h3a53027d),
	.w6(32'hbb5af61e),
	.w7(32'hbbc52bed),
	.w8(32'hbae8cf49),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb1b19),
	.w1(32'hbc120c0a),
	.w2(32'h3c39f9dd),
	.w3(32'hbbc4b536),
	.w4(32'hbb41be53),
	.w5(32'hbb0d77be),
	.w6(32'hbbd2080d),
	.w7(32'hbb6f8481),
	.w8(32'hbb01dda8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89ddfe),
	.w1(32'h3aa3af5e),
	.w2(32'h3c17d796),
	.w3(32'hbc2dda63),
	.w4(32'hbbfe7e11),
	.w5(32'hb9c0bc2a),
	.w6(32'hba68b043),
	.w7(32'h3c2f27aa),
	.w8(32'h3c06153e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396faf31),
	.w1(32'h3b284c3e),
	.w2(32'hbb87de7c),
	.w3(32'hbaf46c58),
	.w4(32'h3bb6edce),
	.w5(32'hbac2171a),
	.w6(32'hbba18c95),
	.w7(32'hbb81c6d9),
	.w8(32'hbac54ba2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad53b0a),
	.w1(32'h3b2418d1),
	.w2(32'h3af89ebe),
	.w3(32'h3868384b),
	.w4(32'h3bb34a86),
	.w5(32'h39c082ef),
	.w6(32'hbb55cc9f),
	.w7(32'h3aab698f),
	.w8(32'h38351224),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe70f5f),
	.w1(32'hbab3539c),
	.w2(32'h3c2f9680),
	.w3(32'hbc1511c6),
	.w4(32'hbba42c44),
	.w5(32'h3adc6d38),
	.w6(32'h3b6660a7),
	.w7(32'h3a7d8b1a),
	.w8(32'h3bf1a741),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a476597),
	.w1(32'h3ba2eb46),
	.w2(32'h3a74105e),
	.w3(32'hbadb3ff0),
	.w4(32'hba16fa7d),
	.w5(32'hbad3196a),
	.w6(32'hb929199c),
	.w7(32'hba688987),
	.w8(32'hba72e593),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb294d5b),
	.w1(32'h3b42c9c8),
	.w2(32'h3c28cf72),
	.w3(32'hbb7888af),
	.w4(32'h3ac323c2),
	.w5(32'h3c03b269),
	.w6(32'h391a61ee),
	.w7(32'hb9e55c87),
	.w8(32'h3bbb7146),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f6b6b),
	.w1(32'hbb8f4e23),
	.w2(32'hbaf586f4),
	.w3(32'hba97f414),
	.w4(32'hbae29c6f),
	.w5(32'hbad9031b),
	.w6(32'hba0c099b),
	.w7(32'h39d39294),
	.w8(32'h3b8788ba),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03ee6e),
	.w1(32'hb95bd0fb),
	.w2(32'hba5d1e3c),
	.w3(32'hba337d00),
	.w4(32'h3b63ec66),
	.w5(32'h3b5df902),
	.w6(32'hbaf8e0ad),
	.w7(32'hbb084e45),
	.w8(32'hb9d94c1b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba847097),
	.w1(32'h3aa6fa24),
	.w2(32'h391ba5de),
	.w3(32'hbb1e67c3),
	.w4(32'h3bc6638a),
	.w5(32'h3b8f7c88),
	.w6(32'hb9bbd26d),
	.w7(32'hbb40bf94),
	.w8(32'h398ec0fa),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a487688),
	.w1(32'h3b9df6fe),
	.w2(32'h3aeb0ebd),
	.w3(32'h3c021769),
	.w4(32'h3b83194f),
	.w5(32'h3af42090),
	.w6(32'h3b4093b3),
	.w7(32'h3b176585),
	.w8(32'h3b6545f6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7d150),
	.w1(32'hba17521b),
	.w2(32'hbbef8ccb),
	.w3(32'hb9b52ed1),
	.w4(32'hb970884e),
	.w5(32'hbc0734b7),
	.w6(32'hba821560),
	.w7(32'h392d4442),
	.w8(32'hbb2d206f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfaa8f),
	.w1(32'hbaaa0d5b),
	.w2(32'hba834c81),
	.w3(32'hbaea659f),
	.w4(32'hbb508a85),
	.w5(32'hbb5a6ede),
	.w6(32'h39a2f038),
	.w7(32'hb9e08362),
	.w8(32'h39f6f396),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b592d5e),
	.w1(32'h3bff0d72),
	.w2(32'h3bf64567),
	.w3(32'hbb64cb35),
	.w4(32'h3b772740),
	.w5(32'h3ae94e5b),
	.w6(32'hbb984965),
	.w7(32'hbb126505),
	.w8(32'hbb1ddc06),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbc213),
	.w1(32'h3bc2bb7c),
	.w2(32'h3c5491a9),
	.w3(32'h3a5333a5),
	.w4(32'h3aabe5ae),
	.w5(32'h3bf770e1),
	.w6(32'hbb4658c6),
	.w7(32'h3baeb89d),
	.w8(32'h3c1b21a5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fe340),
	.w1(32'h3b3a9216),
	.w2(32'hbc04de9b),
	.w3(32'h3a8875b1),
	.w4(32'h3a7d0cc6),
	.w5(32'hbb59c7c1),
	.w6(32'h3b6be6f3),
	.w7(32'hb9b593dc),
	.w8(32'hbb29d1a7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc995738),
	.w1(32'hba1667b0),
	.w2(32'h3ca19295),
	.w3(32'hbc70fa51),
	.w4(32'h3ba68aeb),
	.w5(32'h3c95da8f),
	.w6(32'hbbbab2ec),
	.w7(32'hbaa48ef1),
	.w8(32'h3c4c63a8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06d624),
	.w1(32'h3bb20990),
	.w2(32'h3b8def31),
	.w3(32'h3bb5c000),
	.w4(32'h3c3f5ec5),
	.w5(32'h3c12149b),
	.w6(32'hbb20a65e),
	.w7(32'hbbb7fb84),
	.w8(32'hbb8a544b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a9598),
	.w1(32'h3c337905),
	.w2(32'h3c8648bf),
	.w3(32'hbb3f6d76),
	.w4(32'h3a6e968c),
	.w5(32'h3bb1e4a1),
	.w6(32'hbaabf59b),
	.w7(32'h3bcae2e2),
	.w8(32'h3b986997),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b836dd5),
	.w1(32'h3c2eb6b8),
	.w2(32'h3bfe5d83),
	.w3(32'hbb80e34c),
	.w4(32'h3bbd3605),
	.w5(32'h3b14ae95),
	.w6(32'h3b2ff892),
	.w7(32'h3bb14a2e),
	.w8(32'h3b8f46b0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fc26c),
	.w1(32'hbb8c3d6d),
	.w2(32'hbc9bbe2f),
	.w3(32'h3b6c6180),
	.w4(32'h3b029ec3),
	.w5(32'h3a3bdede),
	.w6(32'hbbe6ee5f),
	.w7(32'hbc0f2687),
	.w8(32'hbc883b3d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0369b),
	.w1(32'hbb1a5ae1),
	.w2(32'hbb5e8ce2),
	.w3(32'h3b016996),
	.w4(32'hba8801ca),
	.w5(32'hbaf3eb17),
	.w6(32'hbb06eb7d),
	.w7(32'hbbc0eb75),
	.w8(32'hbaedf3f6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93d057),
	.w1(32'hba865dfd),
	.w2(32'h3c19eeb6),
	.w3(32'hbae91fe5),
	.w4(32'hba2b0737),
	.w5(32'h3c63f4de),
	.w6(32'hbc274287),
	.w7(32'hbc0d9d7e),
	.w8(32'hbb72ee1c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1718ff),
	.w1(32'hbb02c15d),
	.w2(32'h3c75cad3),
	.w3(32'hbb9c6b0e),
	.w4(32'h3b2e0397),
	.w5(32'h3ca3e401),
	.w6(32'h39771763),
	.w7(32'hbb8bcb65),
	.w8(32'h3b2af15c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fc5b3),
	.w1(32'hbaa484da),
	.w2(32'h3c00fe9d),
	.w3(32'h3c2ff88e),
	.w4(32'h3b6a126b),
	.w5(32'hbb999a68),
	.w6(32'hbc45eae8),
	.w7(32'hbc1ff4de),
	.w8(32'h3b39767e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be69f86),
	.w1(32'hbb9d181a),
	.w2(32'hbcb6cd8f),
	.w3(32'h3c033860),
	.w4(32'hbb7ead2e),
	.w5(32'hbc8c807c),
	.w6(32'hbb7f32bf),
	.w7(32'h3b072a2d),
	.w8(32'hbba2447d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c150176),
	.w1(32'hbabbbe17),
	.w2(32'hbca4a20f),
	.w3(32'h3b4ed390),
	.w4(32'hbb7acd50),
	.w5(32'hbc3a6ece),
	.w6(32'hbc31c606),
	.w7(32'hbc1d93b1),
	.w8(32'hbc850c7b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0b620),
	.w1(32'hb9ae09d1),
	.w2(32'h3b2b7932),
	.w3(32'hbb7a6b1e),
	.w4(32'hbbfe8a61),
	.w5(32'hbb8b8718),
	.w6(32'h3c21f6f3),
	.w7(32'h3c734a56),
	.w8(32'h3c3d0df9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaca31),
	.w1(32'h396efd3d),
	.w2(32'h3a8295c5),
	.w3(32'hbb1e63c0),
	.w4(32'hba91f31b),
	.w5(32'h3a49bb73),
	.w6(32'h3b05ca6b),
	.w7(32'h3b149ef6),
	.w8(32'h3af164bf),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc26cf),
	.w1(32'hbbb71330),
	.w2(32'hbc1398b2),
	.w3(32'hbb133449),
	.w4(32'hbb63c726),
	.w5(32'hbce8d963),
	.w6(32'h3b6fee2a),
	.w7(32'h3bf34b63),
	.w8(32'hbb9dce25),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa577d4),
	.w1(32'hbb24bb28),
	.w2(32'hba671b19),
	.w3(32'hbba3f65b),
	.w4(32'hbb0d6f8a),
	.w5(32'h39bdd5ef),
	.w6(32'hba168fea),
	.w7(32'hbac7fd30),
	.w8(32'h3b08b67f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c4487),
	.w1(32'h3b169cb1),
	.w2(32'h3ab5ec9f),
	.w3(32'hba50bfda),
	.w4(32'h3b0f6049),
	.w5(32'hba99ca80),
	.w6(32'h3a9836a9),
	.w7(32'h37ef567b),
	.w8(32'h3b13a2e1),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b156708),
	.w1(32'h3a0bf9d7),
	.w2(32'h39800db4),
	.w3(32'h3aad076c),
	.w4(32'hbaae6d37),
	.w5(32'hbb3513ba),
	.w6(32'h3aaf4071),
	.w7(32'hbaa71a56),
	.w8(32'h3a356ded),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc65ba6),
	.w1(32'h3abcdf5e),
	.w2(32'h3b5e3fc4),
	.w3(32'hbb8e61d2),
	.w4(32'hbb383d70),
	.w5(32'h3a6169cb),
	.w6(32'h3abc9ca3),
	.w7(32'h3c036f33),
	.w8(32'h3bbda31f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1da287),
	.w1(32'h3b42c4e9),
	.w2(32'hbbcb10e1),
	.w3(32'h38e92005),
	.w4(32'h3b140d01),
	.w5(32'hbc10d7ee),
	.w6(32'hbb416e48),
	.w7(32'h3ac4ea5d),
	.w8(32'hbb869666),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7973ce),
	.w1(32'h3c26a871),
	.w2(32'h3b97d2c4),
	.w3(32'hbbb567ee),
	.w4(32'h3bcd0952),
	.w5(32'h3afb0a46),
	.w6(32'h3ba46217),
	.w7(32'h3b40d93d),
	.w8(32'h3a43bc38),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b537e25),
	.w1(32'hb9c4ea33),
	.w2(32'hbc3fcbd3),
	.w3(32'h3a8ca038),
	.w4(32'hba75e392),
	.w5(32'hbc887c82),
	.w6(32'hbc11b27e),
	.w7(32'hbc1e7032),
	.w8(32'hbc2034e4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1bb23),
	.w1(32'h3c0a6425),
	.w2(32'h3c4901f1),
	.w3(32'hbc3afb9d),
	.w4(32'h399645f8),
	.w5(32'h3b61d05a),
	.w6(32'hbbb00916),
	.w7(32'hb8c8c6bb),
	.w8(32'hbb16baf8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb860c6f),
	.w1(32'h3c350071),
	.w2(32'h3bfce184),
	.w3(32'hbace993e),
	.w4(32'h3b896b68),
	.w5(32'hbb02ed61),
	.w6(32'hbb38a612),
	.w7(32'hba27a4a5),
	.w8(32'hbafc18d6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ee670),
	.w1(32'hbaa7c312),
	.w2(32'hbb8558b8),
	.w3(32'hbb27e44a),
	.w4(32'hbb8373ce),
	.w5(32'hbbdec038),
	.w6(32'hbb294132),
	.w7(32'h3954d992),
	.w8(32'hbb40ffa4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a90d0),
	.w1(32'hb7b04afb),
	.w2(32'hbb85e6d3),
	.w3(32'hbb53b787),
	.w4(32'hbb86c262),
	.w5(32'hbbc502bd),
	.w6(32'h3bce1c5f),
	.w7(32'h3c2507c5),
	.w8(32'h3b624f0d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0fdae),
	.w1(32'h3b13a4af),
	.w2(32'h38b66617),
	.w3(32'hbaca1986),
	.w4(32'hb8728af9),
	.w5(32'hb909be1f),
	.w6(32'h3b988ad0),
	.w7(32'h3b5f7d06),
	.w8(32'h3a5511ce),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b18459),
	.w1(32'h3ad4de8e),
	.w2(32'hb9988e33),
	.w3(32'h3ac1a64a),
	.w4(32'h3982ad50),
	.w5(32'h38f5fb62),
	.w6(32'h3b8785e3),
	.w7(32'h3b61fc0e),
	.w8(32'h3988c1e2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98202a4),
	.w1(32'hbb270653),
	.w2(32'hbbf61f68),
	.w3(32'h3ae71cca),
	.w4(32'hbbdb1f36),
	.w5(32'hbbc68ebe),
	.w6(32'hbbf8ae54),
	.w7(32'hbb64c378),
	.w8(32'hbbdc1fd1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe450b0),
	.w1(32'h3b8092ce),
	.w2(32'hb9bf0b88),
	.w3(32'hbc10eacb),
	.w4(32'hbb17949e),
	.w5(32'hbb3b69c0),
	.w6(32'hba8e1936),
	.w7(32'h3b43bb79),
	.w8(32'hb9f48e51),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e3c98),
	.w1(32'hba74d502),
	.w2(32'hbb16ee7b),
	.w3(32'h3b96ec77),
	.w4(32'h3a5f41c3),
	.w5(32'h3b200365),
	.w6(32'hba936454),
	.w7(32'h397aff13),
	.w8(32'hba664159),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64354f),
	.w1(32'hba337dd5),
	.w2(32'h3b9db338),
	.w3(32'h39cf2e6e),
	.w4(32'h3a302222),
	.w5(32'h3c045e57),
	.w6(32'hbbdb03f5),
	.w7(32'hbb9f12e1),
	.w8(32'hba917aa8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b632755),
	.w1(32'h39cf82a7),
	.w2(32'hbc526644),
	.w3(32'h3bbfbfdf),
	.w4(32'hba352656),
	.w5(32'hbc40e269),
	.w6(32'h3b62fce0),
	.w7(32'h3b8fc171),
	.w8(32'hbba98c4a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73d582),
	.w1(32'hbbfcae13),
	.w2(32'hbc8c0f61),
	.w3(32'hba05b9ac),
	.w4(32'hbbbbcd54),
	.w5(32'hbb39533d),
	.w6(32'hbc478567),
	.w7(32'hbc28550d),
	.w8(32'hbc878a04),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a7d06),
	.w1(32'hba69227c),
	.w2(32'h3baf2d9f),
	.w3(32'hbc1bbfda),
	.w4(32'h3c055f75),
	.w5(32'h3c9b1389),
	.w6(32'h3aba0f44),
	.w7(32'hbb58e269),
	.w8(32'hb9c78cb1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97f491),
	.w1(32'hbaa60a44),
	.w2(32'hba52c055),
	.w3(32'h3c2af9eb),
	.w4(32'hbb24d6b7),
	.w5(32'hbab27ace),
	.w6(32'h3a398689),
	.w7(32'hba442b9f),
	.w8(32'hb967ebfe),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e9e19),
	.w1(32'hbb86b161),
	.w2(32'hba195f46),
	.w3(32'hba0144d0),
	.w4(32'h3abd0acf),
	.w5(32'h3bbce8e7),
	.w6(32'hbb4e17d0),
	.w7(32'h3b37aa3a),
	.w8(32'hba5b5a56),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeddb78),
	.w1(32'h3bf0c803),
	.w2(32'h3c614095),
	.w3(32'hbb3ce069),
	.w4(32'hb9badd05),
	.w5(32'h3bf41981),
	.w6(32'h3b41054d),
	.w7(32'h3c4c27fc),
	.w8(32'h3c473a27),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3d52e),
	.w1(32'h3c135aa9),
	.w2(32'h3d383c36),
	.w3(32'hbc0ae63a),
	.w4(32'h3bd2b9bf),
	.w5(32'hbc4a18d5),
	.w6(32'hbb7611f7),
	.w7(32'h3bffd6c5),
	.w8(32'h3c216b3a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52175d),
	.w1(32'hb98cd0b9),
	.w2(32'hba524cb1),
	.w3(32'hbbd46ebd),
	.w4(32'hbacce714),
	.w5(32'hbc1a5c84),
	.w6(32'h3afb1569),
	.w7(32'h3c310d93),
	.w8(32'h3b11aeec),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3973495e),
	.w1(32'hbbf35d1b),
	.w2(32'hbbe63dd0),
	.w3(32'hbb9e2277),
	.w4(32'hbb80babb),
	.w5(32'h3b60db0e),
	.w6(32'hba513d5e),
	.w7(32'hb9e11f06),
	.w8(32'hbbb754be),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc420632),
	.w1(32'h3c179a93),
	.w2(32'hbc3918ea),
	.w3(32'hbb297552),
	.w4(32'hbb996440),
	.w5(32'h3a8e8021),
	.w6(32'hbbc9e401),
	.w7(32'h3b1f1f6e),
	.w8(32'hb9cf724f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92398f),
	.w1(32'h3acd7805),
	.w2(32'hbc20af99),
	.w3(32'hb9ae414a),
	.w4(32'h3bf96773),
	.w5(32'hb9bd20b7),
	.w6(32'hbbe5b17b),
	.w7(32'h3c5f2078),
	.w8(32'h3c984e4e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c555710),
	.w1(32'h3c8c18f6),
	.w2(32'hba76edec),
	.w3(32'hbbf006b1),
	.w4(32'hbbba2617),
	.w5(32'hbcefecc0),
	.w6(32'h3c9a146a),
	.w7(32'h3d0ae8a1),
	.w8(32'h3c8f43fd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e1d7d),
	.w1(32'hba1d2b28),
	.w2(32'h3c860094),
	.w3(32'hbcc6c334),
	.w4(32'h3a50b1e4),
	.w5(32'h3c029366),
	.w6(32'hbbe548f8),
	.w7(32'hbafa36f3),
	.w8(32'h3bb2c2f6),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4268c2),
	.w1(32'hbb68ef92),
	.w2(32'hbc59ad19),
	.w3(32'hbbc21548),
	.w4(32'hbb33c3fc),
	.w5(32'hba8799d2),
	.w6(32'hba887cd5),
	.w7(32'hbaa1eb31),
	.w8(32'hbb7a1946),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4ef71),
	.w1(32'hbb033206),
	.w2(32'h3b2f977b),
	.w3(32'h3a2bf9d8),
	.w4(32'hbb1763cf),
	.w5(32'hbb50c7e7),
	.w6(32'hbb57584d),
	.w7(32'h3c06e24c),
	.w8(32'h3a7198d8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95e209),
	.w1(32'hba8d9364),
	.w2(32'h3c309214),
	.w3(32'h3a3522fc),
	.w4(32'h3c025485),
	.w5(32'h3c501474),
	.w6(32'hbbf9429c),
	.w7(32'h3a069d2d),
	.w8(32'h3bdcc23f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eefb7),
	.w1(32'hbb878d11),
	.w2(32'hbcbd924f),
	.w3(32'h3afbfadc),
	.w4(32'hbb6c1271),
	.w5(32'h3b08c346),
	.w6(32'hbb39e2b5),
	.w7(32'hbbd0fbb4),
	.w8(32'hbaa7f5cf),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9db3f5),
	.w1(32'hbc50f12b),
	.w2(32'hbc0fdccf),
	.w3(32'hbbe22fbc),
	.w4(32'hbc6c7757),
	.w5(32'hb9283e29),
	.w6(32'hbcb2f19f),
	.w7(32'hbcba1d83),
	.w8(32'hbc499e88),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc469ba0),
	.w1(32'hbb4bb8e5),
	.w2(32'hbaa62bc3),
	.w3(32'hbbdbd9d2),
	.w4(32'hb98d7fcd),
	.w5(32'hb99832ae),
	.w6(32'h3a76ed71),
	.w7(32'h3b4c8d83),
	.w8(32'hbb1f1efe),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6bf42),
	.w1(32'hbb94c452),
	.w2(32'hbb9d82f6),
	.w3(32'hbaf27c63),
	.w4(32'h3c67e7cf),
	.w5(32'h3d2ab98f),
	.w6(32'hbc86205a),
	.w7(32'hbc9327ee),
	.w8(32'hbc4baf49),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb364fda),
	.w1(32'h3c30fc9f),
	.w2(32'hbcd56175),
	.w3(32'h3c632035),
	.w4(32'h3bc738d6),
	.w5(32'h3c87ae4c),
	.w6(32'hb82f6a42),
	.w7(32'h3c56ca9f),
	.w8(32'h3baaacf1),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc38b19),
	.w1(32'h3b06320d),
	.w2(32'hbb3b91e3),
	.w3(32'h3c26f632),
	.w4(32'hbb12567b),
	.w5(32'hbc1d7035),
	.w6(32'h3c0c216c),
	.w7(32'h3c7cc858),
	.w8(32'h3ab8eb38),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac99dc),
	.w1(32'hb9fafe20),
	.w2(32'hbb5d4d40),
	.w3(32'hb986caae),
	.w4(32'hbadc55d9),
	.w5(32'hbc306a59),
	.w6(32'h3bc2c984),
	.w7(32'h3aadcb6e),
	.w8(32'h3bd0e63f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba954143),
	.w1(32'hbaec3de9),
	.w2(32'h3b23bdc3),
	.w3(32'hbbe6b7b0),
	.w4(32'h3ba24bc3),
	.w5(32'hba24b745),
	.w6(32'hbabd7a11),
	.w7(32'h3b376f35),
	.w8(32'hbb146d68),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01479a),
	.w1(32'hbb5688c4),
	.w2(32'hbbf8ce41),
	.w3(32'hb9b88235),
	.w4(32'h3aa5bdac),
	.w5(32'hbc03102d),
	.w6(32'h3a21a989),
	.w7(32'hba4e855b),
	.w8(32'hbb3f191b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb579dab),
	.w1(32'h3b476f4b),
	.w2(32'h3b2b1906),
	.w3(32'hbbdb61eb),
	.w4(32'hbaab327c),
	.w5(32'hbb9c402f),
	.w6(32'hbb95475f),
	.w7(32'h3b437f69),
	.w8(32'hbb35f587),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56a13e),
	.w1(32'hba1c7ad0),
	.w2(32'hbb8644e5),
	.w3(32'hbb19c779),
	.w4(32'hbb11f268),
	.w5(32'h3a949f08),
	.w6(32'hbb3ae894),
	.w7(32'h3a943b4f),
	.w8(32'hbaa0a78f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd01a4),
	.w1(32'hbd40ce33),
	.w2(32'hbd02c92e),
	.w3(32'hbb42fd30),
	.w4(32'hbc0bc65b),
	.w5(32'hbbacc19f),
	.w6(32'hbc0da7c3),
	.w7(32'hbc045798),
	.w8(32'hbc521e51),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd73ec61),
	.w1(32'hbb0c064f),
	.w2(32'h3ac52ef7),
	.w3(32'hbc33ec67),
	.w4(32'hb90aae7a),
	.w5(32'h38440bff),
	.w6(32'hbbd6e522),
	.w7(32'hbad58c7c),
	.w8(32'hbaae7a12),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb979732),
	.w1(32'hbbbc264f),
	.w2(32'hba8cb9ce),
	.w3(32'hba3831b7),
	.w4(32'hbbb00bd5),
	.w5(32'h3c04286d),
	.w6(32'hbbcc9b19),
	.w7(32'hbb3906cb),
	.w8(32'h39dba525),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f7b82),
	.w1(32'h3cb5130d),
	.w2(32'hbb9a3ad3),
	.w3(32'hbb5645b5),
	.w4(32'h3b96971c),
	.w5(32'hbc559132),
	.w6(32'h3b6a8aab),
	.w7(32'h3c86e158),
	.w8(32'h3aa7d831),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f67bf),
	.w1(32'h3c544b4c),
	.w2(32'h3ab1c996),
	.w3(32'h3b8c3f03),
	.w4(32'h3bede30a),
	.w5(32'h3ba1f221),
	.w6(32'h3b4d5a8f),
	.w7(32'hbab1676b),
	.w8(32'h3a9bfa46),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1c5cb),
	.w1(32'hb96e7144),
	.w2(32'hbb5297fc),
	.w3(32'h3b765c3d),
	.w4(32'h3a157d09),
	.w5(32'hbaae7d32),
	.w6(32'h39cd23f4),
	.w7(32'h3b1f048a),
	.w8(32'hba9bd736),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb206bd0),
	.w1(32'hbb3dc9ce),
	.w2(32'hbb36b764),
	.w3(32'hbb22a138),
	.w4(32'hbb7d623a),
	.w5(32'hbc0a34a2),
	.w6(32'hbbaa56c6),
	.w7(32'h3cb41d40),
	.w8(32'h3c739567),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29eea1),
	.w1(32'h3b27ed8d),
	.w2(32'hbb48ad6b),
	.w3(32'h3a217d6d),
	.w4(32'hb894301f),
	.w5(32'hbb2a79ea),
	.w6(32'h3b5d98a2),
	.w7(32'h3c061a5e),
	.w8(32'h3a8dbc56),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a541d41),
	.w1(32'h3b62cb37),
	.w2(32'hbbc1e0f9),
	.w3(32'h3a20381b),
	.w4(32'h3a87dd84),
	.w5(32'hbbf99a3f),
	.w6(32'h3b4047cb),
	.w7(32'h3abe0785),
	.w8(32'h3a7fc55a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41decc),
	.w1(32'hba609753),
	.w2(32'h393ed751),
	.w3(32'hb8d2c1a1),
	.w4(32'hbab48df3),
	.w5(32'h3ab1a051),
	.w6(32'hbb770d9a),
	.w7(32'h3b075025),
	.w8(32'h3b49e0dc),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aea10a),
	.w1(32'hb9bb39a9),
	.w2(32'hbb83302d),
	.w3(32'h3a315eba),
	.w4(32'h378474cf),
	.w5(32'hbb4b505e),
	.w6(32'hb94e40a5),
	.w7(32'h3b8042c0),
	.w8(32'hba2ab5b6),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba713b5),
	.w1(32'h3b958af8),
	.w2(32'h3c038067),
	.w3(32'hbb8bd5da),
	.w4(32'h3afa5cf2),
	.w5(32'h3bff1b07),
	.w6(32'hbb8804ea),
	.w7(32'h3bb7140a),
	.w8(32'h3b8849a1),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9a49b),
	.w1(32'h3b2ec406),
	.w2(32'h3bede2fd),
	.w3(32'hbc3272dd),
	.w4(32'h3afa9648),
	.w5(32'hba151f43),
	.w6(32'h3bf49168),
	.w7(32'h39e6d4be),
	.w8(32'h3c38c096),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c7a11),
	.w1(32'h3be14dfd),
	.w2(32'hbb9a0a95),
	.w3(32'hbbab6b00),
	.w4(32'h3bc4eeb2),
	.w5(32'hbc3b6b08),
	.w6(32'h3c0d3a15),
	.w7(32'h3c80a3ee),
	.w8(32'h3af9c5fc),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a2f00),
	.w1(32'hbacb7dd7),
	.w2(32'hbb8ccf2c),
	.w3(32'h3af1af90),
	.w4(32'hbab893a3),
	.w5(32'hbafb5900),
	.w6(32'hbbd8e969),
	.w7(32'hbab60ad2),
	.w8(32'hbae39021),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb259ed9),
	.w1(32'h3a98bb31),
	.w2(32'hbc123515),
	.w3(32'hbb8ed7c7),
	.w4(32'hbbdc5439),
	.w5(32'hbc751cef),
	.w6(32'h3b9c0f49),
	.w7(32'h3ccdbbc1),
	.w8(32'h3c82daf7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ab20b),
	.w1(32'hbb0cecdb),
	.w2(32'h3b26867d),
	.w3(32'hbbd7ece8),
	.w4(32'h3aa91e7f),
	.w5(32'hbb097e2e),
	.w6(32'hbb2ec55c),
	.w7(32'hb7f00cc1),
	.w8(32'hba742289),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba959b09),
	.w1(32'hb8d0dbb8),
	.w2(32'hbbe4d9b7),
	.w3(32'hbbc782a7),
	.w4(32'hbafcb644),
	.w5(32'hbb91da78),
	.w6(32'h3b9be939),
	.w7(32'h3c0dfad0),
	.w8(32'h3b6967d8),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388cbeaa),
	.w1(32'h39edefc7),
	.w2(32'hbbccb100),
	.w3(32'h3aa074f1),
	.w4(32'h398cf111),
	.w5(32'hbbd1771d),
	.w6(32'h3a7b94d7),
	.w7(32'h3b1be4fe),
	.w8(32'h3a25c524),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953e9bc),
	.w1(32'h3b7f7088),
	.w2(32'h3c25061c),
	.w3(32'hbc344632),
	.w4(32'h3b5a63b4),
	.w5(32'h3b9e5a1e),
	.w6(32'hbc2f858b),
	.w7(32'hba503616),
	.w8(32'h3ba3eafd),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af95289),
	.w1(32'h3a2b85e5),
	.w2(32'hb90f81ba),
	.w3(32'hb9ace163),
	.w4(32'hbb8cd11d),
	.w5(32'hbb62e7f7),
	.w6(32'hbbc861e9),
	.w7(32'hbbddd5b4),
	.w8(32'hbaa2f05a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f19a4),
	.w1(32'hbab17acc),
	.w2(32'hbbca44fa),
	.w3(32'hbaa4e9f8),
	.w4(32'h392547e0),
	.w5(32'hbb7257b0),
	.w6(32'h3a9c9bda),
	.w7(32'h3b3c9ccd),
	.w8(32'hbb8304b1),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba93ea6),
	.w1(32'hbb749d01),
	.w2(32'h3c558541),
	.w3(32'hbb5c8699),
	.w4(32'h3c3d6628),
	.w5(32'h3c83565c),
	.w6(32'hbb609e56),
	.w7(32'hbb5e40d7),
	.w8(32'hba1adf40),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37c388),
	.w1(32'hbb970100),
	.w2(32'h3d429262),
	.w3(32'hbb0b7381),
	.w4(32'h3ba85a4c),
	.w5(32'h3d1892a3),
	.w6(32'hbcc326fe),
	.w7(32'hbce4931b),
	.w8(32'hbc8d324b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc372a54),
	.w1(32'hbc1101fd),
	.w2(32'h3ceab3c9),
	.w3(32'h3bb183f7),
	.w4(32'h3bebf53e),
	.w5(32'h3cbcbbe3),
	.w6(32'hbc447769),
	.w7(32'hbcbdc127),
	.w8(32'hbcc9fbde),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c8c92),
	.w1(32'h3b5049da),
	.w2(32'hbd4521a6),
	.w3(32'h3ace2be3),
	.w4(32'h3baaaaa3),
	.w5(32'h3c7b56dc),
	.w6(32'h3bd2237c),
	.w7(32'h3b89b5cf),
	.w8(32'h3c636156),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf2cc5),
	.w1(32'h39a77489),
	.w2(32'hbb7ae08a),
	.w3(32'h3ba4a7fe),
	.w4(32'hbb80b734),
	.w5(32'hbc3f0800),
	.w6(32'h3b965047),
	.w7(32'h3a35a1fa),
	.w8(32'h3b4db579),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa26717),
	.w1(32'h3be6b27a),
	.w2(32'h3b6bc032),
	.w3(32'hbaccd0fe),
	.w4(32'h3aed3c86),
	.w5(32'hbaf0564f),
	.w6(32'h3a0a3357),
	.w7(32'h3b5fc0e1),
	.w8(32'h3ace9301),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6cbd0),
	.w1(32'hbb683afd),
	.w2(32'hba910435),
	.w3(32'hbb4b25e3),
	.w4(32'hba1dbfa8),
	.w5(32'h3c3af0e6),
	.w6(32'hbb8224e1),
	.w7(32'hbb9c84b4),
	.w8(32'hbad8acd4),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d10a5),
	.w1(32'hbb0fb805),
	.w2(32'h3c7adc80),
	.w3(32'h3b19d63e),
	.w4(32'h3c6ba208),
	.w5(32'h3d4a21c2),
	.w6(32'hbc973424),
	.w7(32'hbd02a6e5),
	.w8(32'hbc951cab),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96b194),
	.w1(32'h3ba719a8),
	.w2(32'hbd0a4621),
	.w3(32'h3bf5c35f),
	.w4(32'hbc265cb8),
	.w5(32'hbc9b11ce),
	.w6(32'h3c732c67),
	.w7(32'h3c0da0b3),
	.w8(32'hbbde3cdd),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b22862),
	.w1(32'h3c2779fc),
	.w2(32'hb9dd9193),
	.w3(32'h3c01ece7),
	.w4(32'hbc44babf),
	.w5(32'hbd055fdd),
	.w6(32'h3b6e12dc),
	.w7(32'h3cad957c),
	.w8(32'hbbd199dd),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd913a5),
	.w1(32'hbb6833e7),
	.w2(32'hbc69d0c2),
	.w3(32'hbc7a5d60),
	.w4(32'hbc18fea6),
	.w5(32'hbcc6ba23),
	.w6(32'h3b705ff2),
	.w7(32'h3c892868),
	.w8(32'h3c2fcfa6),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c806201),
	.w1(32'h3977b929),
	.w2(32'hbbb6d25d),
	.w3(32'hbb2aadd0),
	.w4(32'hbb320ea1),
	.w5(32'hbc166584),
	.w6(32'h3bb4c3f0),
	.w7(32'h3c344539),
	.w8(32'h3babac74),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbf446),
	.w1(32'h3c085be1),
	.w2(32'hba0290f0),
	.w3(32'h392c3446),
	.w4(32'h3bc030c4),
	.w5(32'h3b14c00a),
	.w6(32'hbaba0725),
	.w7(32'h3bafef71),
	.w8(32'hb98af3c4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb425601),
	.w1(32'hbb929f18),
	.w2(32'h3ca21b23),
	.w3(32'h3b4c3308),
	.w4(32'hbb23fa2c),
	.w5(32'h3cbe675b),
	.w6(32'hbc11e064),
	.w7(32'hbc8a0f3d),
	.w8(32'hbc89557b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a4131),
	.w1(32'hbc17e074),
	.w2(32'hbcbef457),
	.w3(32'hbc126adb),
	.w4(32'hbb16433c),
	.w5(32'hb9c7414e),
	.w6(32'hbb88a3b1),
	.w7(32'hbc927cd5),
	.w8(32'hbc77949c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a3fe5),
	.w1(32'hbac31217),
	.w2(32'h3b14a830),
	.w3(32'hbbba5f5c),
	.w4(32'h3ae4460e),
	.w5(32'hbbb16ee7),
	.w6(32'hbb7fda48),
	.w7(32'hb9405467),
	.w8(32'hbb643c42),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f6b01),
	.w1(32'h3b520a11),
	.w2(32'h3b93a0e5),
	.w3(32'hbc1b1f61),
	.w4(32'hbb1f9025),
	.w5(32'h3b10bce0),
	.w6(32'hbba3d793),
	.w7(32'h3bfbd0ae),
	.w8(32'h3be44ebd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1070f6),
	.w1(32'h3c7011ef),
	.w2(32'hb92f1c5a),
	.w3(32'hbc43ca40),
	.w4(32'h3b2cd3f9),
	.w5(32'h3a4b4a9c),
	.w6(32'h38280367),
	.w7(32'h3b92228b),
	.w8(32'hbba1d3e3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c2ec2),
	.w1(32'hbc20b257),
	.w2(32'h3c53f432),
	.w3(32'hbba1e515),
	.w4(32'hbb53daa3),
	.w5(32'h3b7fb73e),
	.w6(32'hbb91db4b),
	.w7(32'hbb36c6b7),
	.w8(32'h3a9c8112),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1287a),
	.w1(32'h3c0f4f7d),
	.w2(32'hbc0a0ec5),
	.w3(32'h3b4b2dd4),
	.w4(32'h3aed9c9a),
	.w5(32'hbc031977),
	.w6(32'hbb42fd0f),
	.w7(32'hbc1e80af),
	.w8(32'h3ba97125),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4af07f),
	.w1(32'hbb82f8c1),
	.w2(32'h3b9189e8),
	.w3(32'hbc7d3ab9),
	.w4(32'h3be0c322),
	.w5(32'h3badf0d5),
	.w6(32'hbae9a1e4),
	.w7(32'hbaaa0d4b),
	.w8(32'hb9bc682b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33e564),
	.w1(32'h3b398dba),
	.w2(32'h3c029c49),
	.w3(32'h39bf6017),
	.w4(32'h3b1c7d5b),
	.w5(32'hbb42120e),
	.w6(32'h3b188539),
	.w7(32'h3ba6c01a),
	.w8(32'hba10e42a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32176d),
	.w1(32'h3a8c3562),
	.w2(32'hbb965c52),
	.w3(32'h39637b2d),
	.w4(32'h3ae187ac),
	.w5(32'h3c8c834b),
	.w6(32'hba4b85e9),
	.w7(32'hbc69da8a),
	.w8(32'hbb896152),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65760b),
	.w1(32'h3b79e0ba),
	.w2(32'hbb8849a4),
	.w3(32'hb8b3ccbc),
	.w4(32'hbb6e26f9),
	.w5(32'hbc0fa74c),
	.w6(32'hbb079d7e),
	.w7(32'hbaa89fe6),
	.w8(32'hbb22136e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28a63e),
	.w1(32'hbb5f10d0),
	.w2(32'hbc11a6d0),
	.w3(32'hbbae9be4),
	.w4(32'hba15ffa1),
	.w5(32'hbc25a4e2),
	.w6(32'hbb59379f),
	.w7(32'hbb1b6581),
	.w8(32'hbc17a47f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a073612),
	.w1(32'h3bbb5e50),
	.w2(32'hbba9d68d),
	.w3(32'hbaa6910f),
	.w4(32'h39921a34),
	.w5(32'hbc29388c),
	.w6(32'h3b1f8c9f),
	.w7(32'h3bfb9b31),
	.w8(32'hba4b3599),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd0dc3),
	.w1(32'hbb82ece7),
	.w2(32'h3cc0f308),
	.w3(32'hbb9fe192),
	.w4(32'h3cb21a03),
	.w5(32'h3d8b3e57),
	.w6(32'hbcce3cf3),
	.w7(32'hbd227ce2),
	.w8(32'hbce04bef),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f6da2),
	.w1(32'hb96a854c),
	.w2(32'hbb3c6c4c),
	.w3(32'h3c2d757f),
	.w4(32'hbaeeb720),
	.w5(32'hbc13ec9a),
	.w6(32'h3aa2bcf9),
	.w7(32'h3b782f51),
	.w8(32'hba918dc7),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e8156),
	.w1(32'hbb30a0a7),
	.w2(32'hbbecc46c),
	.w3(32'hbb19f696),
	.w4(32'hbae7e879),
	.w5(32'hb99ff703),
	.w6(32'hbb21750a),
	.w7(32'h3a990d98),
	.w8(32'hba54b5f4),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ad17e),
	.w1(32'h3ba6ee66),
	.w2(32'hbc11832a),
	.w3(32'h3aa93e79),
	.w4(32'h39d23623),
	.w5(32'hbbd55e2f),
	.w6(32'h3bb37981),
	.w7(32'h3c1116be),
	.w8(32'hba2cb97a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa3d76),
	.w1(32'h39ed308f),
	.w2(32'hbb9359d5),
	.w3(32'h3a3142df),
	.w4(32'hba965610),
	.w5(32'hbb3896b7),
	.w6(32'hbb986f8b),
	.w7(32'h3a19179d),
	.w8(32'hbb7e92ad),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba590fc8),
	.w1(32'h3bb19617),
	.w2(32'h3ba735f6),
	.w3(32'h3aa27c59),
	.w4(32'h3b18413d),
	.w5(32'hbaadd410),
	.w6(32'h3a9e5eeb),
	.w7(32'h3c1fb6f1),
	.w8(32'hba962507),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b8d89),
	.w1(32'h3c8bc3ba),
	.w2(32'hbc21b947),
	.w3(32'h3aa98784),
	.w4(32'h3b668261),
	.w5(32'h3d0ef8a1),
	.w6(32'hbc1b4b7c),
	.w7(32'hbc3eaf2d),
	.w8(32'h3aef272b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2e10a),
	.w1(32'hbb6c8dc2),
	.w2(32'hbb1f6a3c),
	.w3(32'hbbd4d7e1),
	.w4(32'h3aadd155),
	.w5(32'h3c45679b),
	.w6(32'hbab2cb48),
	.w7(32'h3a397967),
	.w8(32'hb9f15577),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd5e0d),
	.w1(32'h3acb0057),
	.w2(32'h3bae0b3f),
	.w3(32'h3bb2a05f),
	.w4(32'hbb809643),
	.w5(32'h3b1be958),
	.w6(32'h3a24955b),
	.w7(32'hbb5e8b85),
	.w8(32'hbb28f205),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17474e),
	.w1(32'hbb9b296f),
	.w2(32'hbc86ef89),
	.w3(32'hbb51eb7a),
	.w4(32'hbb1cd10d),
	.w5(32'hbc3711fa),
	.w6(32'h3c22b2a6),
	.w7(32'h3c10d428),
	.w8(32'hbb43a526),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb367ca2),
	.w1(32'h39c9d707),
	.w2(32'hb9122445),
	.w3(32'hbb15b499),
	.w4(32'hbb012f06),
	.w5(32'h3b3f4bbe),
	.w6(32'hbb991207),
	.w7(32'h3b6815d4),
	.w8(32'h3b6d7050),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb914c42),
	.w1(32'hb7f9e58e),
	.w2(32'hba99a445),
	.w3(32'hbaf0e67e),
	.w4(32'hbb7874c3),
	.w5(32'hbbc23d21),
	.w6(32'hbc25b40f),
	.w7(32'hbb5e0c77),
	.w8(32'hbbd52132),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f3943),
	.w1(32'h3ba5c4bb),
	.w2(32'h3b8a3f9b),
	.w3(32'hbbbbb26a),
	.w4(32'h3b954eea),
	.w5(32'hbbf2bf90),
	.w6(32'h3aa92cb4),
	.w7(32'h3b97e12c),
	.w8(32'h3b0af642),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6dd21),
	.w1(32'h3b8762ed),
	.w2(32'hbb33dff5),
	.w3(32'h3af9f24e),
	.w4(32'hbacb46d3),
	.w5(32'hbbb4ed36),
	.w6(32'h3a9b11db),
	.w7(32'h3acfbd60),
	.w8(32'hbbb770c4),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29d673),
	.w1(32'h3bbc3f48),
	.w2(32'h3ca72fa5),
	.w3(32'hbbdbb0b8),
	.w4(32'hbb599ce6),
	.w5(32'hbadf1d32),
	.w6(32'hbc27126c),
	.w7(32'hb98e477e),
	.w8(32'hb9895c28),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c15c1),
	.w1(32'h3c20e0b5),
	.w2(32'h3b98aaee),
	.w3(32'hb8bb5483),
	.w4(32'hbb91b57c),
	.w5(32'hbb47864c),
	.w6(32'hbbaaa4e4),
	.w7(32'hba8d5aee),
	.w8(32'h3c1d095f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba037e46),
	.w1(32'h3b7cba34),
	.w2(32'h3bb9799f),
	.w3(32'hbc251921),
	.w4(32'hbbf5fb74),
	.w5(32'hbbef9193),
	.w6(32'hbb329d20),
	.w7(32'hbb63a0a9),
	.w8(32'hbbd305d0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d3079),
	.w1(32'hbb31216f),
	.w2(32'h3cae3a00),
	.w3(32'hbcb350ea),
	.w4(32'h3b84afdd),
	.w5(32'h3d24a375),
	.w6(32'hbc1f28e1),
	.w7(32'hbca78de3),
	.w8(32'h3abec76a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ba6ac),
	.w1(32'h399574d1),
	.w2(32'hba9899c2),
	.w3(32'h3c11b642),
	.w4(32'hba8f9dbd),
	.w5(32'hb9833a2d),
	.w6(32'hbb55ca4f),
	.w7(32'h3a12781b),
	.w8(32'h3a976824),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391228cd),
	.w1(32'h3b197a48),
	.w2(32'hbb07b09e),
	.w3(32'hb9f0ddab),
	.w4(32'hbb50c377),
	.w5(32'hbc516120),
	.w6(32'h3b944f40),
	.w7(32'h3c45ad64),
	.w8(32'h3bcd3096),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3494ba),
	.w1(32'hbbbab837),
	.w2(32'hb9b209a0),
	.w3(32'hbba1ecd9),
	.w4(32'h39fa64df),
	.w5(32'h3bebd745),
	.w6(32'hbb8efc08),
	.w7(32'h3acd5781),
	.w8(32'h3c473f09),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a55dd),
	.w1(32'h3b9372fa),
	.w2(32'h3c1e20c5),
	.w3(32'hbb7d9606),
	.w4(32'hbade9b56),
	.w5(32'h3b6e1956),
	.w6(32'hbc125731),
	.w7(32'h3b37ae11),
	.w8(32'h3b7e9c06),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf259d3),
	.w1(32'hbc37c351),
	.w2(32'h3bc42fc7),
	.w3(32'hbb559b06),
	.w4(32'h3b763cfb),
	.w5(32'h3c7056c9),
	.w6(32'hbc8a7aa1),
	.w7(32'hbc716b26),
	.w8(32'hbc2c96da),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6ac7d),
	.w1(32'h3c0532fc),
	.w2(32'hbba928d9),
	.w3(32'hbb08281e),
	.w4(32'hbb87c129),
	.w5(32'hbd086594),
	.w6(32'h3c93dd81),
	.w7(32'h3cd14b69),
	.w8(32'h3ba9d91e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b5195),
	.w1(32'h3b95e13f),
	.w2(32'hbc3ad66f),
	.w3(32'hb8e352b0),
	.w4(32'h3bff7010),
	.w5(32'hbbebcc3a),
	.w6(32'h3b0bcc74),
	.w7(32'h3a57331b),
	.w8(32'hbb9e8294),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb934e8d7),
	.w1(32'hbb502349),
	.w2(32'hbbe50206),
	.w3(32'h3b3423c9),
	.w4(32'h39c111b9),
	.w5(32'hba49384e),
	.w6(32'hba8cff5e),
	.w7(32'hbb046ff6),
	.w8(32'hbb22eed6),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a76a3),
	.w1(32'hbc166e98),
	.w2(32'h3c6dfbf7),
	.w3(32'hb9670577),
	.w4(32'hbc0dbedf),
	.w5(32'hbcb36887),
	.w6(32'h3b3c4f66),
	.w7(32'hbaafd5eb),
	.w8(32'h3a91ceaf),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b19add),
	.w1(32'h3c047a18),
	.w2(32'h3b6fecb4),
	.w3(32'hbaf1b5c0),
	.w4(32'h399723c9),
	.w5(32'hb9a69c9f),
	.w6(32'h3ae45570),
	.w7(32'hbac370e3),
	.w8(32'h3b6b7fa5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f53e9),
	.w1(32'hba6e4d4c),
	.w2(32'hbaf310b6),
	.w3(32'hb9921c20),
	.w4(32'hbb373de0),
	.w5(32'hbc64530a),
	.w6(32'h3bba21aa),
	.w7(32'h3ccf3386),
	.w8(32'h3c5dbb3c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd0c43),
	.w1(32'h3bbc7bd5),
	.w2(32'h3bc42976),
	.w3(32'hbb96623b),
	.w4(32'h3a4674b7),
	.w5(32'hbbfa8bc2),
	.w6(32'h3a85e943),
	.w7(32'h3c012b05),
	.w8(32'h3c13e6ff),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a9436),
	.w1(32'h3b6f5e24),
	.w2(32'hbbc40e56),
	.w3(32'hbbc4952d),
	.w4(32'hbc892a00),
	.w5(32'hbd1d3259),
	.w6(32'h3c0fd7e0),
	.w7(32'h3cf28181),
	.w8(32'h3c2e2a5b),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99810fc),
	.w1(32'h3b80e548),
	.w2(32'hbc221713),
	.w3(32'hbc09cf40),
	.w4(32'hbac3bd26),
	.w5(32'h3c80f682),
	.w6(32'h3b49ff67),
	.w7(32'hbcb0d0c7),
	.w8(32'hbc21faf3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c991fab),
	.w1(32'hbbc8225b),
	.w2(32'h3ca93748),
	.w3(32'h3a92c269),
	.w4(32'hbbd90ea6),
	.w5(32'hbc9fc40c),
	.w6(32'hbb1b30af),
	.w7(32'hbb94ef75),
	.w8(32'hbc5f78fd),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d73f1),
	.w1(32'hbc4b6359),
	.w2(32'h3bb12749),
	.w3(32'hbb51f90c),
	.w4(32'hbb193ffe),
	.w5(32'h3cbaa999),
	.w6(32'hbc34e1c3),
	.w7(32'h399e576d),
	.w8(32'h3bc5a2ff),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a05f2),
	.w1(32'h39ff08d4),
	.w2(32'hbb679dd9),
	.w3(32'h3be579b7),
	.w4(32'hbb1b6c9c),
	.w5(32'h3bb682c0),
	.w6(32'hbb834fd9),
	.w7(32'h3bc12fde),
	.w8(32'h3bcc6ddd),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01c755),
	.w1(32'hbb8345ee),
	.w2(32'hbadc1fac),
	.w3(32'hba236ce6),
	.w4(32'h3a867fe2),
	.w5(32'h3c1d954a),
	.w6(32'hb9ec5479),
	.w7(32'h3b37b0f9),
	.w8(32'h3b321467),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bdd07),
	.w1(32'hbb01eecf),
	.w2(32'h3bea3f10),
	.w3(32'hb95dfdc3),
	.w4(32'h3a5cc83b),
	.w5(32'h3c129d03),
	.w6(32'hbbc657e5),
	.w7(32'h3b82cf58),
	.w8(32'h3b9498f7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba653f8a),
	.w1(32'hbc009816),
	.w2(32'hbc10609a),
	.w3(32'h3a47ed30),
	.w4(32'hb9858e26),
	.w5(32'hba25f83c),
	.w6(32'hbb7ecd60),
	.w7(32'hbb6c95f6),
	.w8(32'hba934696),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66f1de),
	.w1(32'h3a3c4c59),
	.w2(32'hbb56a0b1),
	.w3(32'hbb5eb4f3),
	.w4(32'hba6e17ec),
	.w5(32'hbb047766),
	.w6(32'hbb4c3fb0),
	.w7(32'h3a4cc36e),
	.w8(32'hba380eaf),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae254ea),
	.w1(32'hbb9660c2),
	.w2(32'h3a15bcd4),
	.w3(32'h3a28bfc2),
	.w4(32'h3af9dc9a),
	.w5(32'h3c50fe85),
	.w6(32'hbb05e9dd),
	.w7(32'hb8771464),
	.w8(32'h3acc28bd),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf2ba5),
	.w1(32'hbbf62d94),
	.w2(32'h3c7a925a),
	.w3(32'h3b8c22bf),
	.w4(32'h3bee9d55),
	.w5(32'h3d043370),
	.w6(32'hbc88577b),
	.w7(32'hbcc33c53),
	.w8(32'hbc41bc3e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcabe58),
	.w1(32'h3bca48dc),
	.w2(32'hbc70fbbc),
	.w3(32'h3b021231),
	.w4(32'hbb4dfd5f),
	.w5(32'hbc38ef77),
	.w6(32'h3c11d0b9),
	.w7(32'h3c2c59e6),
	.w8(32'hbaf86979),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74fce0),
	.w1(32'h3c33edbf),
	.w2(32'h3c3833f9),
	.w3(32'hbbd4d269),
	.w4(32'hb8795b88),
	.w5(32'h3ca925b6),
	.w6(32'hbb06d362),
	.w7(32'hbc7dff1a),
	.w8(32'h3b84b6eb),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba217c02),
	.w1(32'h3b9c4f96),
	.w2(32'hbbef2d02),
	.w3(32'h3be41e39),
	.w4(32'hbb1acc94),
	.w5(32'hbc0f2dd5),
	.w6(32'h3bd3796b),
	.w7(32'h3ca20eac),
	.w8(32'h3bd2ba37),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28b155),
	.w1(32'h3b695e64),
	.w2(32'h3c133ecb),
	.w3(32'hbbcfee1a),
	.w4(32'h3b1cc2f8),
	.w5(32'h3c9e9d3f),
	.w6(32'hbc4cc62e),
	.w7(32'hbc8b8828),
	.w8(32'hbb78849b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393cb341),
	.w1(32'hbb83e062),
	.w2(32'h3b29ba5b),
	.w3(32'h3a77ed2c),
	.w4(32'h3a882426),
	.w5(32'h3c849fe9),
	.w6(32'hbc165ae7),
	.w7(32'hbbad9ee7),
	.w8(32'h3ad63a31),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc19fe2),
	.w1(32'hbbafb63e),
	.w2(32'h3a2551dd),
	.w3(32'hbb549108),
	.w4(32'h3b10d9dc),
	.w5(32'h3c8b1ca0),
	.w6(32'hbafcd88f),
	.w7(32'h3b15e157),
	.w8(32'h3b650dad),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf452ef),
	.w1(32'hbb1cb8a3),
	.w2(32'hbbbbdacc),
	.w3(32'h3bd3708c),
	.w4(32'hbb5d2bd4),
	.w5(32'hbb511f5f),
	.w6(32'h3b10c560),
	.w7(32'h3bc80846),
	.w8(32'h3b3101e6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacb771),
	.w1(32'hba898c43),
	.w2(32'hbbb8cfe4),
	.w3(32'hbb463dd6),
	.w4(32'hbb3b1885),
	.w5(32'hbc03c38b),
	.w6(32'h3bbae903),
	.w7(32'h3c5881ac),
	.w8(32'h3bf6e16b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03020b),
	.w1(32'hbcfb9b95),
	.w2(32'hbbb6d6b5),
	.w3(32'hbbeef879),
	.w4(32'hb9e9216d),
	.w5(32'h3c0de39e),
	.w6(32'h3af80fa2),
	.w7(32'h3c85fe2b),
	.w8(32'h3865220a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1a7565),
	.w1(32'hbb7fa3df),
	.w2(32'hba707fc7),
	.w3(32'hbbb69bc2),
	.w4(32'hbacdf13d),
	.w5(32'h3b973984),
	.w6(32'hbb07b07e),
	.w7(32'hbc4057f0),
	.w8(32'hbbfdf074),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bfc90),
	.w1(32'h39f3d3ef),
	.w2(32'h3816b7b8),
	.w3(32'hbad291b0),
	.w4(32'hbc07bc0c),
	.w5(32'hbbe49f77),
	.w6(32'hbbe21e56),
	.w7(32'h3be71b6d),
	.w8(32'h3aa0117a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3953905d),
	.w1(32'h3c10364e),
	.w2(32'hba929e04),
	.w3(32'hbc0ab110),
	.w4(32'hbb9a7567),
	.w5(32'hbc91dd6e),
	.w6(32'h3b556a75),
	.w7(32'h3bd3e0b0),
	.w8(32'hbbf6d544),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc566e88),
	.w1(32'hbb3e9088),
	.w2(32'hbb8b3a28),
	.w3(32'hbc4927dd),
	.w4(32'hbb4345ea),
	.w5(32'hbb02af11),
	.w6(32'h3a17e7c7),
	.w7(32'h3ab607cd),
	.w8(32'hb95474c3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4d17f),
	.w1(32'hbc73b1d8),
	.w2(32'h3cfe6e38),
	.w3(32'hba972ea1),
	.w4(32'hbbc49000),
	.w5(32'h3b89b9e1),
	.w6(32'hbbc68908),
	.w7(32'h3b9d0080),
	.w8(32'h3863a25e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc454463),
	.w1(32'h3c007f5e),
	.w2(32'h3be84293),
	.w3(32'h39d79138),
	.w4(32'hbc389cbb),
	.w5(32'hbd3a7eba),
	.w6(32'h3c5a2194),
	.w7(32'h3d0ebff2),
	.w8(32'h3c4602c0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e24b8),
	.w1(32'h3c8c1547),
	.w2(32'h3c11c665),
	.w3(32'hbd02d03e),
	.w4(32'h3c180661),
	.w5(32'h3c0bd670),
	.w6(32'hbb776db2),
	.w7(32'h3ba907a2),
	.w8(32'h3b6123a3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaacb56),
	.w1(32'hba4d96b6),
	.w2(32'hbb02e045),
	.w3(32'h389121c6),
	.w4(32'hb9b6e9e8),
	.w5(32'hbabda53f),
	.w6(32'h3a2f5134),
	.w7(32'hba9dffe5),
	.w8(32'hb951c51c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9ad2e),
	.w1(32'h3b3ff384),
	.w2(32'hbb4a9369),
	.w3(32'hbab784f3),
	.w4(32'hbb311df5),
	.w5(32'hbbf6d568),
	.w6(32'hbb24de44),
	.w7(32'hba7be29c),
	.w8(32'hbb6c6ce6),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule