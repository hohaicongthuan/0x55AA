module layer_10_featuremap_362(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6dfc5),
	.w1(32'hbbaedce7),
	.w2(32'hbb02a7e5),
	.w3(32'hbb9e51af),
	.w4(32'hbad91eaa),
	.w5(32'h3b9b5d07),
	.w6(32'hbbbea544),
	.w7(32'hbb084513),
	.w8(32'h3b989cc1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6cfce),
	.w1(32'h3b6ea37c),
	.w2(32'h3c54985c),
	.w3(32'hb8a2e245),
	.w4(32'h3b15524f),
	.w5(32'hbbccc1f9),
	.w6(32'hbb6881a7),
	.w7(32'h3b9b4910),
	.w8(32'hbbb2d3f7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08e8cc),
	.w1(32'h3984352a),
	.w2(32'hbb085c3f),
	.w3(32'hbb74db6e),
	.w4(32'hbbe7e9ea),
	.w5(32'h385fe3e8),
	.w6(32'hbc2096c6),
	.w7(32'hbbae1c4b),
	.w8(32'h3a8d8402),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a522b05),
	.w1(32'h3ac4a70b),
	.w2(32'h3af6d952),
	.w3(32'h3a86f65e),
	.w4(32'hba6ae46c),
	.w5(32'hbba0ac44),
	.w6(32'h3b8806b8),
	.w7(32'h3aa1ec8d),
	.w8(32'hbaed506e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58d1f7),
	.w1(32'h3bb1d50b),
	.w2(32'h3b6fe6ba),
	.w3(32'h3ad3be22),
	.w4(32'h3acc38fd),
	.w5(32'hbb7bbac0),
	.w6(32'h3ba48317),
	.w7(32'h3af186e2),
	.w8(32'hbb65994e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9385a2),
	.w1(32'hbb6708af),
	.w2(32'hbb3eaf38),
	.w3(32'hbb8ca95c),
	.w4(32'hbb68e86a),
	.w5(32'hbb90ed16),
	.w6(32'hbb5bf2a2),
	.w7(32'hbb78ad78),
	.w8(32'hbb803571),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb608a90),
	.w1(32'hbb6fa94b),
	.w2(32'hbbce03ef),
	.w3(32'hbbae255a),
	.w4(32'hbb963eb6),
	.w5(32'hbc041130),
	.w6(32'hbb6f31eb),
	.w7(32'hbb77337a),
	.w8(32'hbbdf2d14),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0d4e8),
	.w1(32'hbbff5315),
	.w2(32'hbc11eace),
	.w3(32'hbb82d625),
	.w4(32'hba421764),
	.w5(32'hbbf70837),
	.w6(32'hbb8c80e9),
	.w7(32'hba9c4bb4),
	.w8(32'hbbf5a9c3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c4b14),
	.w1(32'hbb99bc98),
	.w2(32'hbb99971b),
	.w3(32'hbbc65c39),
	.w4(32'hbb8a57c7),
	.w5(32'hbaaadf26),
	.w6(32'hbbbfe435),
	.w7(32'hbba78498),
	.w8(32'hbb49c336),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc359326),
	.w1(32'hbb0e87eb),
	.w2(32'hbb9bc7ce),
	.w3(32'hbbeba1b8),
	.w4(32'hbb217239),
	.w5(32'hbb8f79a9),
	.w6(32'hbbbb86fa),
	.w7(32'h3ab83224),
	.w8(32'hba66fc0f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd374a),
	.w1(32'hbb1f0aad),
	.w2(32'hbb516f76),
	.w3(32'hbb186322),
	.w4(32'hbb24ba7e),
	.w5(32'h39caa184),
	.w6(32'hbb37f47d),
	.w7(32'hbb60f34b),
	.w8(32'hbb037f51),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d0f0b),
	.w1(32'h3b503059),
	.w2(32'hbbb9a9dc),
	.w3(32'h3b62954f),
	.w4(32'hbad62c44),
	.w5(32'h3a417347),
	.w6(32'hbc370247),
	.w7(32'hbb56f208),
	.w8(32'h3aa88a1d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03d8db),
	.w1(32'hbb2212ff),
	.w2(32'hbba65176),
	.w3(32'h3a6c27eb),
	.w4(32'h3bf36ad5),
	.w5(32'hbbb788e0),
	.w6(32'h3b25e5cf),
	.w7(32'h3c36edea),
	.w8(32'hbb2b1463),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36ecd8),
	.w1(32'hba9f0660),
	.w2(32'h3ba3e388),
	.w3(32'hbb0a47cd),
	.w4(32'h399b5223),
	.w5(32'h38c8929f),
	.w6(32'h3b0436cc),
	.w7(32'h3bd963ca),
	.w8(32'hba92231a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a47ed),
	.w1(32'hbacc61ba),
	.w2(32'hbb2f2f26),
	.w3(32'hbb89a910),
	.w4(32'hbb0bff58),
	.w5(32'h3a334ee3),
	.w6(32'hbaeaadb6),
	.w7(32'h38de5aa3),
	.w8(32'h3aaf2d94),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd41bfb),
	.w1(32'hbb5798dc),
	.w2(32'h3a6d5696),
	.w3(32'hbbf305c8),
	.w4(32'h3a689c31),
	.w5(32'hbbb1c423),
	.w6(32'hbb6d8853),
	.w7(32'h3aefde2c),
	.w8(32'hbb2aaf0f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e49c8),
	.w1(32'hbb48eb46),
	.w2(32'hbb153598),
	.w3(32'hbbb27383),
	.w4(32'hbb80ef7d),
	.w5(32'hbbb0c27a),
	.w6(32'hbb8c4b5e),
	.w7(32'hbb6fdeba),
	.w8(32'hbb5f3d10),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7621e),
	.w1(32'hbbc5bed2),
	.w2(32'hbbe1c01a),
	.w3(32'hbaf721ee),
	.w4(32'hbb2e8006),
	.w5(32'hbba11f1c),
	.w6(32'hbb7716e8),
	.w7(32'hb96a7435),
	.w8(32'hbb21fd19),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26bd0c),
	.w1(32'hbb5a732a),
	.w2(32'hbba76539),
	.w3(32'hba94e1e7),
	.w4(32'hbb01915f),
	.w5(32'hb9b3886f),
	.w6(32'hbafc6643),
	.w7(32'hbbe54511),
	.w8(32'hb83e9785),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cada4),
	.w1(32'h3b62cb6c),
	.w2(32'h3ba3cfc0),
	.w3(32'h3a262a63),
	.w4(32'hb8afda4e),
	.w5(32'h3a752c93),
	.w6(32'h3bee3c17),
	.w7(32'h39b362b7),
	.w8(32'hb9ccb856),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5b52e),
	.w1(32'hbaff80fd),
	.w2(32'h3bcb6de9),
	.w3(32'h3ad3f714),
	.w4(32'h3b41fdc8),
	.w5(32'h3a538d73),
	.w6(32'h3b84bc67),
	.w7(32'h3bc1947a),
	.w8(32'h3a6dc78e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33e77d),
	.w1(32'hba6cb2ff),
	.w2(32'hbb88cd03),
	.w3(32'h3a6d1fc7),
	.w4(32'hbac52891),
	.w5(32'hbb077dc5),
	.w6(32'h3b211c9f),
	.w7(32'hbaeda34a),
	.w8(32'hbaef8d4f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3df0aa),
	.w1(32'hbb694274),
	.w2(32'hbac373a8),
	.w3(32'hbc6886e5),
	.w4(32'hbac1b822),
	.w5(32'hbb2bf6a7),
	.w6(32'hbc939bd0),
	.w7(32'hbb7b66e9),
	.w8(32'hbbe49110),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf70d81),
	.w1(32'hbbdcc9a0),
	.w2(32'hbbb6245b),
	.w3(32'hbbd3c556),
	.w4(32'hbb21812b),
	.w5(32'hbaf77438),
	.w6(32'hbc0211ef),
	.w7(32'h3992c19a),
	.w8(32'h3b3655ee),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d507a),
	.w1(32'hbad0e4fd),
	.w2(32'hbb97c67f),
	.w3(32'hbb811ab7),
	.w4(32'hba874ad8),
	.w5(32'hbae65cec),
	.w6(32'hbc23f085),
	.w7(32'hbb5e2b39),
	.w8(32'hbab075a9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7bec1),
	.w1(32'h39e59602),
	.w2(32'hb9b8ff0c),
	.w3(32'hbb944549),
	.w4(32'hbb011fd0),
	.w5(32'hb81c18c2),
	.w6(32'hb71e7c15),
	.w7(32'hbb230ef4),
	.w8(32'h3a540557),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3fcc1),
	.w1(32'hbb1346ad),
	.w2(32'hbaca4e3c),
	.w3(32'hbb24ffb0),
	.w4(32'hbb33a548),
	.w5(32'hbb50f2e7),
	.w6(32'hba79bcb8),
	.w7(32'hbae18e68),
	.w8(32'hbba42661),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8abb2),
	.w1(32'hbbc546e2),
	.w2(32'hbb338940),
	.w3(32'hbbbbe599),
	.w4(32'hbb6400ab),
	.w5(32'hbacdbaf9),
	.w6(32'hbbcc0e66),
	.w7(32'hbb951386),
	.w8(32'h3adc5598),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eb94b),
	.w1(32'hbae2f149),
	.w2(32'h3af113ed),
	.w3(32'hbb8eebda),
	.w4(32'hbb8c0ffc),
	.w5(32'hbb6faf26),
	.w6(32'hba1072ec),
	.w7(32'hbb1fe53b),
	.w8(32'hbbb9b3bc),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18ddb9),
	.w1(32'h3b8d5d68),
	.w2(32'h3b18d9d3),
	.w3(32'hbb80dda2),
	.w4(32'hbb34cb44),
	.w5(32'hba9d7836),
	.w6(32'hbb07faa2),
	.w7(32'h3aaf6207),
	.w8(32'hbc16ac87),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75bfde),
	.w1(32'hbbd1862a),
	.w2(32'hbbcacd69),
	.w3(32'hba80a2a4),
	.w4(32'hbb4dbcb0),
	.w5(32'h3a9d0264),
	.w6(32'hbc6e23d6),
	.w7(32'hbc4a1258),
	.w8(32'h3adab9f5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b2661),
	.w1(32'h3acf658f),
	.w2(32'hba8c8cb2),
	.w3(32'hbb27a0df),
	.w4(32'hba7298df),
	.w5(32'hbb398a50),
	.w6(32'hbb479f08),
	.w7(32'hbb1af55c),
	.w8(32'hbb45ab50),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77ee3d),
	.w1(32'hbb40e3d7),
	.w2(32'hbbc75fe8),
	.w3(32'hbbb7d43e),
	.w4(32'hbb10a9f4),
	.w5(32'hbc180864),
	.w6(32'hbc4f7bcf),
	.w7(32'hbbab44fd),
	.w8(32'hbb71d53b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc240ad),
	.w1(32'hbb46c45c),
	.w2(32'hb9dddcff),
	.w3(32'hbbce3e77),
	.w4(32'hba02b74c),
	.w5(32'h3b1f778e),
	.w6(32'hbbc8d660),
	.w7(32'hbb98a6c5),
	.w8(32'h3a958fc4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5eed38),
	.w1(32'hb82a4005),
	.w2(32'h3a3bc269),
	.w3(32'hbb113741),
	.w4(32'hba57fff7),
	.w5(32'hbb213ab6),
	.w6(32'h3a560a9a),
	.w7(32'hbb08aae4),
	.w8(32'h38ac5e12),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bda74),
	.w1(32'hbb0a1440),
	.w2(32'hbbb12b55),
	.w3(32'hbb29622c),
	.w4(32'hb8d0f414),
	.w5(32'hbb06e794),
	.w6(32'hbb4795cd),
	.w7(32'hbaf2aea1),
	.w8(32'h39d1f24d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1ab56),
	.w1(32'hbb7275a5),
	.w2(32'h3b0501a4),
	.w3(32'hbbdc07e5),
	.w4(32'hbb7df433),
	.w5(32'hbb4891a6),
	.w6(32'hbc1205a3),
	.w7(32'hbc17e883),
	.w8(32'hbb3b1e74),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5afd2d),
	.w1(32'hbbbdb695),
	.w2(32'hbb634072),
	.w3(32'hbc1b00c1),
	.w4(32'hbbbfc497),
	.w5(32'hbbcc21f1),
	.w6(32'hbbf4ce99),
	.w7(32'hbbeddb14),
	.w8(32'hbb749d39),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7eb134),
	.w1(32'hbaf724f3),
	.w2(32'h3b0e7dd6),
	.w3(32'hbb530041),
	.w4(32'hbc105ae1),
	.w5(32'h3bcdd950),
	.w6(32'hbb9c91c8),
	.w7(32'hbc0b3c2b),
	.w8(32'h3a563983),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dea16),
	.w1(32'hbb0e3a70),
	.w2(32'hbba0df45),
	.w3(32'h3c1800af),
	.w4(32'h39a7e725),
	.w5(32'hbb1aa0f5),
	.w6(32'h3c482f41),
	.w7(32'h3afeab9c),
	.w8(32'hbaf6bcc1),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40f5d8),
	.w1(32'hba07762d),
	.w2(32'h3a8b08f8),
	.w3(32'hbb867432),
	.w4(32'hbb2366dd),
	.w5(32'hbb472287),
	.w6(32'hbbeefb9a),
	.w7(32'h3ac02e4d),
	.w8(32'hbb4d0304),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff42b8),
	.w1(32'h38e30a17),
	.w2(32'hba8f5157),
	.w3(32'hba37813c),
	.w4(32'hbaee24d4),
	.w5(32'h3b80f47f),
	.w6(32'h3b1d66d6),
	.w7(32'hb9566a87),
	.w8(32'h3beed088),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990e57e),
	.w1(32'hbbe96b53),
	.w2(32'hbad68f8d),
	.w3(32'hb9db553e),
	.w4(32'h3b16c108),
	.w5(32'hbb8e7229),
	.w6(32'h396b4b31),
	.w7(32'hbb500d93),
	.w8(32'h39b191b8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf5f4f),
	.w1(32'hbbd14de3),
	.w2(32'hbb3ccef7),
	.w3(32'hbc88909f),
	.w4(32'hbbf0a844),
	.w5(32'h3a2ca023),
	.w6(32'hbc3a31f1),
	.w7(32'hbb44037f),
	.w8(32'hbb460da1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd3f07),
	.w1(32'h3abfec75),
	.w2(32'hbb41ea39),
	.w3(32'hbbe780d9),
	.w4(32'hbab34233),
	.w5(32'hbbb9d54b),
	.w6(32'hbbea50b4),
	.w7(32'hb8c9235d),
	.w8(32'hbbaa1acd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d9615),
	.w1(32'hbbb91daa),
	.w2(32'hbc09eaf1),
	.w3(32'hbc1abf45),
	.w4(32'hbbb3892d),
	.w5(32'hbb6cebcb),
	.w6(32'hbbf0e018),
	.w7(32'hbaea0603),
	.w8(32'hbaf6475d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd63b37),
	.w1(32'h3a154d63),
	.w2(32'h3ac6b20a),
	.w3(32'hbb9880a6),
	.w4(32'hbb454379),
	.w5(32'h39af229c),
	.w6(32'hbafef65c),
	.w7(32'h3992bc9b),
	.w8(32'h3aeb95b9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9613818),
	.w1(32'hbc0346f4),
	.w2(32'hbc3c990d),
	.w3(32'h38774a30),
	.w4(32'hbba6f6ef),
	.w5(32'hbb28b7eb),
	.w6(32'hbb9d1601),
	.w7(32'hbb258446),
	.w8(32'hbab6f5b2),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f7be2),
	.w1(32'hba713fb8),
	.w2(32'h3a41b2d9),
	.w3(32'h3b324e86),
	.w4(32'h3b3c8d3a),
	.w5(32'h3ac9c438),
	.w6(32'h3ac1a94c),
	.w7(32'h3b429ede),
	.w8(32'h3b081115),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b6cea),
	.w1(32'h3b053bcd),
	.w2(32'hba983d0b),
	.w3(32'h3af87fa3),
	.w4(32'h3aae8e02),
	.w5(32'h3b9e7d8d),
	.w6(32'h3bbb5dc9),
	.w7(32'h3a9754ac),
	.w8(32'h3ab86419),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08bce5),
	.w1(32'h3ad25c0e),
	.w2(32'hba479f0a),
	.w3(32'hba157e82),
	.w4(32'hbaa72d07),
	.w5(32'hbb7f3869),
	.w6(32'hbb865bb7),
	.w7(32'hbbad5ca2),
	.w8(32'hbb43c89d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5822f5),
	.w1(32'hbc19caa6),
	.w2(32'hbbf9893c),
	.w3(32'hbc343c3b),
	.w4(32'hbb8a0e65),
	.w5(32'hbbc21ae5),
	.w6(32'hbb80d35a),
	.w7(32'hbba27187),
	.w8(32'hbba31773),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15774f),
	.w1(32'hb999fc9b),
	.w2(32'hbba4f164),
	.w3(32'hbb7b2879),
	.w4(32'hbb9e267c),
	.w5(32'hbbb403af),
	.w6(32'hbc0fbfa8),
	.w7(32'hbb3a2faf),
	.w8(32'hbba48837),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6126a),
	.w1(32'hbc0d500a),
	.w2(32'hbc3376fc),
	.w3(32'hbc12684b),
	.w4(32'hbb9e84a8),
	.w5(32'hbb967b79),
	.w6(32'hbbf06fe6),
	.w7(32'hbb4707d7),
	.w8(32'hbb4479a7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba339253),
	.w1(32'h3b251790),
	.w2(32'h3b881862),
	.w3(32'h3842d0aa),
	.w4(32'h3aef37bb),
	.w5(32'hb9adcc8b),
	.w6(32'h3b08c165),
	.w7(32'h394a6f99),
	.w8(32'h3b0e830f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25a76c),
	.w1(32'h3b8bc729),
	.w2(32'h3ababbb5),
	.w3(32'hbbc899e6),
	.w4(32'hbb415612),
	.w5(32'h3a39af09),
	.w6(32'hb9832de5),
	.w7(32'hbb512128),
	.w8(32'h3a9b884f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87ed7c3),
	.w1(32'h392389ee),
	.w2(32'h3a8885c7),
	.w3(32'hbb2c660b),
	.w4(32'hb961de09),
	.w5(32'hbb055cfc),
	.w6(32'h38ac2c73),
	.w7(32'h3b0f7cd3),
	.w8(32'hbb42d75f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb145b2e),
	.w1(32'hbac17e93),
	.w2(32'h3ba6d8fe),
	.w3(32'h382de550),
	.w4(32'h3b0a8b1c),
	.w5(32'hb98ef9ba),
	.w6(32'h3aaa54c7),
	.w7(32'h3b6d7c1e),
	.w8(32'h39b2dd9c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e80bd),
	.w1(32'h3a768421),
	.w2(32'hbaf14554),
	.w3(32'hbac6ad20),
	.w4(32'hbaba2895),
	.w5(32'hbaa534fa),
	.w6(32'h3aeaf4d2),
	.w7(32'hbb0788b3),
	.w8(32'h3aac6837),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b056b),
	.w1(32'hb7fdbcbd),
	.w2(32'hbb454759),
	.w3(32'h3bbdbdda),
	.w4(32'h3bdf9c09),
	.w5(32'hbaea20ff),
	.w6(32'hbb2617ea),
	.w7(32'hba6b4549),
	.w8(32'hbad9c8be),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ed8f6),
	.w1(32'hba86921f),
	.w2(32'hbab27eca),
	.w3(32'hb997324b),
	.w4(32'hbaa3fc9b),
	.w5(32'hbb6d5f27),
	.w6(32'h3b58f71a),
	.w7(32'h3b5bf776),
	.w8(32'hbb1a527f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4aef59),
	.w1(32'hbac5a1a6),
	.w2(32'h3b1db365),
	.w3(32'hbbccbe00),
	.w4(32'hbb54e253),
	.w5(32'h3a57ef01),
	.w6(32'hbb0ba5b5),
	.w7(32'hb9a4de40),
	.w8(32'h3a06f2da),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ca16e),
	.w1(32'h3bcbd25a),
	.w2(32'h3b72a807),
	.w3(32'h3b8e053a),
	.w4(32'h3aacbd65),
	.w5(32'h3ab342e5),
	.w6(32'h3b2f56de),
	.w7(32'hbb00916a),
	.w8(32'h3a1c0b69),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e2712),
	.w1(32'hbab14e2c),
	.w2(32'h39c9d82b),
	.w3(32'hbb8f6e79),
	.w4(32'hbb11d322),
	.w5(32'h3a12ee8c),
	.w6(32'hbb22d27f),
	.w7(32'h3a2ff9d4),
	.w8(32'h3b2743d6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bf076),
	.w1(32'h3b6a8782),
	.w2(32'h3b899653),
	.w3(32'h38f06c56),
	.w4(32'h3b691047),
	.w5(32'h3b0986d6),
	.w6(32'h3b93a953),
	.w7(32'h39a8d7bc),
	.w8(32'h3aaac574),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9402ec),
	.w1(32'h3b7fe6c9),
	.w2(32'h3a39d2eb),
	.w3(32'h3a81576c),
	.w4(32'hb9e8ac61),
	.w5(32'hbb9909bb),
	.w6(32'hbb4cfcac),
	.w7(32'hbb273bce),
	.w8(32'hbb548fd4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8edf61),
	.w1(32'hbb67155f),
	.w2(32'hbb4af614),
	.w3(32'hbb038aba),
	.w4(32'hbb3126f9),
	.w5(32'hbbae9dfe),
	.w6(32'hbb307f21),
	.w7(32'hbb0cf89b),
	.w8(32'hbb45e06c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a2fbe),
	.w1(32'hbc10db92),
	.w2(32'hbc27add7),
	.w3(32'hbc0f9d40),
	.w4(32'hbbc31866),
	.w5(32'hbb89d01a),
	.w6(32'hbc1056d3),
	.w7(32'hbada4e1e),
	.w8(32'hb874b5d5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e2d97),
	.w1(32'hbb2c7787),
	.w2(32'hbb64d86c),
	.w3(32'hba154dd4),
	.w4(32'h3b82286a),
	.w5(32'hbaa16ddf),
	.w6(32'h3aaf33c7),
	.w7(32'h3af06777),
	.w8(32'h3ad4c41e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb752596),
	.w1(32'hbb1f3d09),
	.w2(32'hbbef3381),
	.w3(32'hbb281008),
	.w4(32'h3bdff2dd),
	.w5(32'h3bf79a3b),
	.w6(32'h3b82661b),
	.w7(32'h3b4c084d),
	.w8(32'h3bcaf165),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32b595),
	.w1(32'hbb59f004),
	.w2(32'hbac451b7),
	.w3(32'hbaba64fe),
	.w4(32'hbb3d0b4d),
	.w5(32'hbb56b35d),
	.w6(32'hb9c8c242),
	.w7(32'hbb71da88),
	.w8(32'hba1ed8a2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803942),
	.w1(32'hbb02505a),
	.w2(32'hbb8bed97),
	.w3(32'h3a132cc7),
	.w4(32'hba9d656c),
	.w5(32'hba86ce3f),
	.w6(32'hbabb5616),
	.w7(32'hbb9c48ca),
	.w8(32'h3b113165),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb21877),
	.w1(32'hbafcc0d0),
	.w2(32'hba8b7e7c),
	.w3(32'hbacb3cbd),
	.w4(32'hbb6a5e9d),
	.w5(32'h3b2eebf7),
	.w6(32'hbab13038),
	.w7(32'hbb51c76c),
	.w8(32'h3b4aa640),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8dcbe),
	.w1(32'h3a82b22d),
	.w2(32'h3bb706b5),
	.w3(32'h3ba2c02f),
	.w4(32'h3ba5ddac),
	.w5(32'hbb87cac5),
	.w6(32'h3b1713b7),
	.w7(32'hb8d7c9a2),
	.w8(32'hba7755bd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb430e66),
	.w1(32'hbb7d1988),
	.w2(32'h38931ffe),
	.w3(32'hbad5a30f),
	.w4(32'hbac66aaf),
	.w5(32'h3a0509c7),
	.w6(32'hbacce36d),
	.w7(32'hba4c24b9),
	.w8(32'h39a4636d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57dae0),
	.w1(32'hbb4c6798),
	.w2(32'hbbb17ae3),
	.w3(32'h3bd6c8d9),
	.w4(32'h3b4e1cce),
	.w5(32'hbbc1fe18),
	.w6(32'hbb1dfb69),
	.w7(32'hba821ff5),
	.w8(32'hbbc6841d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5dc35),
	.w1(32'hbab7cea2),
	.w2(32'hbb20dafb),
	.w3(32'hbc0ce652),
	.w4(32'hbb5397ac),
	.w5(32'hbbb30a04),
	.w6(32'hbc42cda0),
	.w7(32'hb8a96739),
	.w8(32'hbad8ea34),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cb511),
	.w1(32'hbb82f02b),
	.w2(32'hbbb75ccd),
	.w3(32'hbbf11845),
	.w4(32'hbb4a7955),
	.w5(32'hbbbf1806),
	.w6(32'hbbb9d68d),
	.w7(32'hbb247678),
	.w8(32'hbb481322),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21c35b),
	.w1(32'hbbe0d35f),
	.w2(32'hbc411abe),
	.w3(32'hb94f6ce1),
	.w4(32'hba9f90ca),
	.w5(32'hbbd4ea1a),
	.w6(32'hbbb961cc),
	.w7(32'h3a18635c),
	.w8(32'hbb8d73b8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd534a1),
	.w1(32'hbba5463e),
	.w2(32'hbbb17b15),
	.w3(32'hbbe96d80),
	.w4(32'hbb9ce121),
	.w5(32'h3bf34851),
	.w6(32'hbbf571bd),
	.w7(32'hbb57ccdd),
	.w8(32'h3b9b6e54),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00fc23),
	.w1(32'h3a70c71a),
	.w2(32'hbbd79551),
	.w3(32'h3c0d3a38),
	.w4(32'h3c1cb1f6),
	.w5(32'h3960ff40),
	.w6(32'h3ace88e6),
	.w7(32'h3b8cf02f),
	.w8(32'h3b0c9b15),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab22e58),
	.w1(32'hbb6f86e0),
	.w2(32'hbbbecc42),
	.w3(32'h3b8cb755),
	.w4(32'h3bcffa7a),
	.w5(32'hbb1349b8),
	.w6(32'hbb0e477b),
	.w7(32'hbb3a58ca),
	.w8(32'hbb592831),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58ca15),
	.w1(32'hbb4edd05),
	.w2(32'hbb86c10e),
	.w3(32'hba716a5e),
	.w4(32'hba4e76ba),
	.w5(32'h3a8d2ad9),
	.w6(32'hbba4a115),
	.w7(32'hbb7cd88f),
	.w8(32'hb8788ca4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05dc7a),
	.w1(32'hb9e674d6),
	.w2(32'hbba2d25b),
	.w3(32'h3ae4e4ce),
	.w4(32'hbbc1876a),
	.w5(32'h3af33835),
	.w6(32'hba99837a),
	.w7(32'h3a597a5a),
	.w8(32'h3aa1c652),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac87e29),
	.w1(32'hbb60d0cc),
	.w2(32'hbb46437c),
	.w3(32'h39742019),
	.w4(32'h3acfefa5),
	.w5(32'hbb189229),
	.w6(32'hbb656003),
	.w7(32'hbb156a7d),
	.w8(32'hba291fa3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e5db2),
	.w1(32'h3a2550d8),
	.w2(32'hba4c9995),
	.w3(32'hba6f7f90),
	.w4(32'hbaa92bf0),
	.w5(32'hbbebe3a2),
	.w6(32'hba989511),
	.w7(32'hba30831f),
	.w8(32'hbbf3a5f5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbdaa7),
	.w1(32'hbbc17baa),
	.w2(32'hbbb39065),
	.w3(32'hbc0e2fcc),
	.w4(32'hbb8a8746),
	.w5(32'hba1e10c1),
	.w6(32'hbc0f200f),
	.w7(32'hbb97cca9),
	.w8(32'hbb7bf089),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3e4d2),
	.w1(32'h3b5f9a43),
	.w2(32'h3ba5c46e),
	.w3(32'h3a816b82),
	.w4(32'hb9e9985d),
	.w5(32'hbb991135),
	.w6(32'hbb04b377),
	.w7(32'hbb839529),
	.w8(32'hbbaa2515),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef2284),
	.w1(32'hbbca8f24),
	.w2(32'hbbfa2b3e),
	.w3(32'hbc0251b2),
	.w4(32'hbb99d008),
	.w5(32'hba2f04be),
	.w6(32'hbbebd893),
	.w7(32'hbb8ec9df),
	.w8(32'hbb5cb633),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31fdf5),
	.w1(32'hbb432c42),
	.w2(32'hbbc30560),
	.w3(32'hbc0510aa),
	.w4(32'hbbc122c0),
	.w5(32'hbb51b20d),
	.w6(32'hbbcdc85d),
	.w7(32'hba2416d3),
	.w8(32'hbbd37932),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe54406),
	.w1(32'hba68def2),
	.w2(32'h3bc67ccb),
	.w3(32'hbb412abc),
	.w4(32'hba060d1f),
	.w5(32'hba60cd7c),
	.w6(32'hb9bcb128),
	.w7(32'h3b82e2d5),
	.w8(32'hbb808f6f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7555a),
	.w1(32'h3955febc),
	.w2(32'h3b808eb4),
	.w3(32'hbb6eba90),
	.w4(32'hbaacf59b),
	.w5(32'hb8e6483f),
	.w6(32'hbb271f11),
	.w7(32'h3b81d050),
	.w8(32'h3a51faaf),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54508a),
	.w1(32'h3a9509c5),
	.w2(32'h3b685c93),
	.w3(32'hbbec824b),
	.w4(32'h3989307f),
	.w5(32'hb7d717f0),
	.w6(32'hbb047d1f),
	.w7(32'h3b8a6065),
	.w8(32'h3ad08d36),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0f23),
	.w1(32'h3b27f303),
	.w2(32'h3bdace3b),
	.w3(32'hbb80f8ae),
	.w4(32'h3b2cd7bd),
	.w5(32'hbaf9f66c),
	.w6(32'hbb335cf9),
	.w7(32'h3c0170c7),
	.w8(32'h3adfba92),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1a0a6),
	.w1(32'hbb13dcc9),
	.w2(32'hbb8649ad),
	.w3(32'h399fe332),
	.w4(32'h3b21ab52),
	.w5(32'hbb50ac54),
	.w6(32'hb9cb097e),
	.w7(32'hba66f42c),
	.w8(32'hbacd72c2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7ecf3),
	.w1(32'hbbf51937),
	.w2(32'hbc0c5508),
	.w3(32'hbbac13e3),
	.w4(32'hbbb485be),
	.w5(32'h3c19aa4a),
	.w6(32'hbb13858a),
	.w7(32'hbba5f46d),
	.w8(32'h3c1ceaca),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0826e2),
	.w1(32'h3b60bc64),
	.w2(32'h3b868a48),
	.w3(32'h3c941e8b),
	.w4(32'h3c0f2f76),
	.w5(32'hbb82a920),
	.w6(32'h3be1b0c2),
	.w7(32'h3c0df728),
	.w8(32'hbbb20b21),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc48c70),
	.w1(32'hba0be7a8),
	.w2(32'hbbe5b7d1),
	.w3(32'hbc47a267),
	.w4(32'hbbddc99d),
	.w5(32'h3ae20d1c),
	.w6(32'hbc6847bf),
	.w7(32'hbb170560),
	.w8(32'hbb1db709),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae13831),
	.w1(32'hbb4fc463),
	.w2(32'hba56b4a1),
	.w3(32'hbb099c5e),
	.w4(32'h3b24edc4),
	.w5(32'hbb4d341e),
	.w6(32'hbbcb8ae1),
	.w7(32'hbab8a39b),
	.w8(32'hbb4b9e72),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85d66d),
	.w1(32'hbc0b1a0d),
	.w2(32'hbc3f3e18),
	.w3(32'hbaf8a184),
	.w4(32'hbb5ff8e5),
	.w5(32'h393e1eea),
	.w6(32'hbb522a46),
	.w7(32'hba4754f7),
	.w8(32'hbc1d352c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b0a85),
	.w1(32'hbaf3a08e),
	.w2(32'hbb44c3f9),
	.w3(32'hbc25d090),
	.w4(32'h3af7300f),
	.w5(32'hba68caba),
	.w6(32'hbc8dc32f),
	.w7(32'hbbaf2733),
	.w8(32'h3a9b8676),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f4123),
	.w1(32'hbb52f651),
	.w2(32'hbc36cd1a),
	.w3(32'h3aa92029),
	.w4(32'h3bcd95c0),
	.w5(32'hbb21e017),
	.w6(32'h3cca78cd),
	.w7(32'h3b998752),
	.w8(32'h3c29dec2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80355f),
	.w1(32'h3c82aeb5),
	.w2(32'hbb87ef22),
	.w3(32'h3b73a3d9),
	.w4(32'h3c939852),
	.w5(32'h3bc24cb1),
	.w6(32'h3cd2bd32),
	.w7(32'h3c7daa14),
	.w8(32'hba79ac0d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb231bb0),
	.w1(32'hb9cc9fca),
	.w2(32'hbb85b35c),
	.w3(32'h3aa2927f),
	.w4(32'h38e28a07),
	.w5(32'hbb5368be),
	.w6(32'hbb10716d),
	.w7(32'h3a9d865b),
	.w8(32'h3ab96e48),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b379c),
	.w1(32'hbba1270a),
	.w2(32'hbbc68e87),
	.w3(32'hbbf90f6d),
	.w4(32'h3a0d1cb6),
	.w5(32'hbad3694e),
	.w6(32'h3b7a9c22),
	.w7(32'h3ba37013),
	.w8(32'hbbae6159),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90cabf),
	.w1(32'hb8ccf3e2),
	.w2(32'hba404a38),
	.w3(32'h3bba4b0d),
	.w4(32'h3b73434c),
	.w5(32'h3a9be20e),
	.w6(32'h3a8ef888),
	.w7(32'h3b634058),
	.w8(32'h3b1aa4a3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c2c6ab),
	.w1(32'hbb800b45),
	.w2(32'hbb5903d2),
	.w3(32'h3abbd10f),
	.w4(32'h3b80d04c),
	.w5(32'hbb3a6eed),
	.w6(32'h3c59172b),
	.w7(32'h3b735b49),
	.w8(32'hb8d0027e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbd5d9),
	.w1(32'hb8d99ce8),
	.w2(32'hbb6fd2be),
	.w3(32'hbb873bb3),
	.w4(32'hbb1e2840),
	.w5(32'h3a3e0e2e),
	.w6(32'h3acdca2f),
	.w7(32'hbb333263),
	.w8(32'hbbaa894d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a2cc5),
	.w1(32'h39c11b0f),
	.w2(32'h3c02aab5),
	.w3(32'hbc215e70),
	.w4(32'h3b496a68),
	.w5(32'h3ba16ea9),
	.w6(32'hbc8481f9),
	.w7(32'h3ab2f930),
	.w8(32'h3b76232b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf2300),
	.w1(32'h3883dd33),
	.w2(32'h3b49c9eb),
	.w3(32'hbbff302d),
	.w4(32'hbb024f4a),
	.w5(32'h3aa21960),
	.w6(32'hbc027852),
	.w7(32'h3b19e81d),
	.w8(32'hbac23288),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb998dab),
	.w1(32'hbb091a84),
	.w2(32'h3aad0209),
	.w3(32'hbb75efd5),
	.w4(32'hb9de6569),
	.w5(32'h3b640fe2),
	.w6(32'hbbbff631),
	.w7(32'hba62ab33),
	.w8(32'hbc27dac3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09ed2a),
	.w1(32'h3b1806ea),
	.w2(32'h3cb64e53),
	.w3(32'hbc80478c),
	.w4(32'hbc589d32),
	.w5(32'h3b37d383),
	.w6(32'hbbf40242),
	.w7(32'hbb61c7f3),
	.w8(32'h3abbdba9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b121e92),
	.w1(32'hbb62a299),
	.w2(32'hba1c80a8),
	.w3(32'hb9f1a479),
	.w4(32'h39c0a294),
	.w5(32'h3a230a76),
	.w6(32'hbb1a6af8),
	.w7(32'hbabd5599),
	.w8(32'h3b0abac5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8355fb),
	.w1(32'h3d0337b0),
	.w2(32'h3ca99b57),
	.w3(32'hbbab4137),
	.w4(32'h3b8b4520),
	.w5(32'hbbdc4cb2),
	.w6(32'h3c250a82),
	.w7(32'h3c418445),
	.w8(32'hbb270716),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85e391),
	.w1(32'h3a4bc41f),
	.w2(32'hbb57a45d),
	.w3(32'hbb80e505),
	.w4(32'h3b25c4f4),
	.w5(32'h3bee3585),
	.w6(32'hbbbe8137),
	.w7(32'h3b95e2aa),
	.w8(32'hbb25f3aa),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc2dc8),
	.w1(32'hbb8323f1),
	.w2(32'h3bc1c43f),
	.w3(32'hbbafadde),
	.w4(32'hbc1c9f94),
	.w5(32'h3b18a53a),
	.w6(32'hb9833df5),
	.w7(32'hbba7707d),
	.w8(32'h3a9604f8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70e34d),
	.w1(32'hb8e080c9),
	.w2(32'hbaae492a),
	.w3(32'h3b373efd),
	.w4(32'h3b73ed6b),
	.w5(32'h3ac4b694),
	.w6(32'hbac32478),
	.w7(32'h38f8d887),
	.w8(32'h3a67e8cb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a6929),
	.w1(32'hbb83850b),
	.w2(32'h3a871888),
	.w3(32'hbc12bf1c),
	.w4(32'hbc10512d),
	.w5(32'hbb417275),
	.w6(32'h3aa2de1a),
	.w7(32'hbbaa0e12),
	.w8(32'hbaedd5b0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30da81),
	.w1(32'h3ab4aba5),
	.w2(32'h3b94af0a),
	.w3(32'hbb7a2c28),
	.w4(32'hbb997f76),
	.w5(32'h3a36a895),
	.w6(32'hbb2f1ac2),
	.w7(32'hbb4dab26),
	.w8(32'h3a7b78b6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0ceda),
	.w1(32'h3b0abbde),
	.w2(32'hbc09b3fb),
	.w3(32'hbc0aa51b),
	.w4(32'h3a0cfa4c),
	.w5(32'h3c27a9a2),
	.w6(32'hbb6aeef7),
	.w7(32'h3b59808a),
	.w8(32'hbbc95ad4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395323e2),
	.w1(32'hbb682969),
	.w2(32'h3c31121a),
	.w3(32'hbc20c92a),
	.w4(32'hbb951d37),
	.w5(32'h3b720eb3),
	.w6(32'hbbeaeee9),
	.w7(32'hba902a57),
	.w8(32'h39e29df0),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a4c55),
	.w1(32'hbb8f6013),
	.w2(32'hbb90bba0),
	.w3(32'h3b1e7684),
	.w4(32'hba6e9808),
	.w5(32'h3bc31bcd),
	.w6(32'h3b875eee),
	.w7(32'hb95ac2e6),
	.w8(32'hbb31836c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba000a9),
	.w1(32'hbb9a0a57),
	.w2(32'h3aaf5005),
	.w3(32'h3c37e4c2),
	.w4(32'h3be72644),
	.w5(32'h3a7b668f),
	.w6(32'hbaa42727),
	.w7(32'hbc0a4a02),
	.w8(32'hbb9b7e5f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bd1e8),
	.w1(32'hbbcc2e1f),
	.w2(32'hbb384b25),
	.w3(32'h3a57bbf9),
	.w4(32'h3913b7c0),
	.w5(32'hbae9779e),
	.w6(32'h3a3b9a46),
	.w7(32'hbb29ed73),
	.w8(32'h3a877726),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29eabe),
	.w1(32'hb91d99d5),
	.w2(32'h3a8b2c29),
	.w3(32'h39875f7e),
	.w4(32'hbb5222b1),
	.w5(32'h3c60c3a5),
	.w6(32'h3b016d2f),
	.w7(32'hbae5b97f),
	.w8(32'h3ccbb3c9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf141ef),
	.w1(32'h3c847cd7),
	.w2(32'h3cdb5932),
	.w3(32'hbb7ffcfc),
	.w4(32'hbc1f3fd1),
	.w5(32'hbb7a8a9b),
	.w6(32'h3cdab6d7),
	.w7(32'h3c7c2613),
	.w8(32'hba0a3398),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e2d73),
	.w1(32'hbaad644e),
	.w2(32'hbb94375a),
	.w3(32'hbb13cb74),
	.w4(32'h3a914594),
	.w5(32'h39178c53),
	.w6(32'h3b2280c4),
	.w7(32'h3a9f486d),
	.w8(32'h39971f5d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d2003),
	.w1(32'h3c18193d),
	.w2(32'h3bb92a61),
	.w3(32'hbc27fdeb),
	.w4(32'hbc6b98d1),
	.w5(32'hbb3b81a5),
	.w6(32'hbbb783d9),
	.w7(32'hb8d9b4db),
	.w8(32'h39fb070d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2b897),
	.w1(32'h3b6ec86e),
	.w2(32'h3a33c089),
	.w3(32'hbb755d0b),
	.w4(32'h39b483fd),
	.w5(32'hbb956f20),
	.w6(32'hba77f5c3),
	.w7(32'hbb1667ff),
	.w8(32'hbbacc218),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f1b0c),
	.w1(32'h3b3d60de),
	.w2(32'hbaf863e6),
	.w3(32'hba8217af),
	.w4(32'h3a276bbd),
	.w5(32'hbb9e77f9),
	.w6(32'h3b5cfa9b),
	.w7(32'h395c5093),
	.w8(32'hbb931334),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc0576),
	.w1(32'hbbbb4242),
	.w2(32'hbbceaa15),
	.w3(32'hbbdcf190),
	.w4(32'hbbb69a55),
	.w5(32'h3b781ed8),
	.w6(32'h3c4f791c),
	.w7(32'hbbc74b36),
	.w8(32'h3b56f454),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7c87b),
	.w1(32'hbabbfd61),
	.w2(32'hbb9674e5),
	.w3(32'h3b50f9f3),
	.w4(32'h3b523334),
	.w5(32'hbb943827),
	.w6(32'h3b6a9de9),
	.w7(32'h3aaa2a83),
	.w8(32'hbb4d6d10),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc465a70),
	.w1(32'hbc5da717),
	.w2(32'hbbb197ed),
	.w3(32'hbc41a9ea),
	.w4(32'hbbf9e701),
	.w5(32'hbab0d35c),
	.w6(32'h39c164e3),
	.w7(32'hbb6a64f0),
	.w8(32'h38b93094),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aa59d),
	.w1(32'h39e96da3),
	.w2(32'hba0c7e1d),
	.w3(32'hbb780a51),
	.w4(32'hbb5b5375),
	.w5(32'hb8b4840e),
	.w6(32'hb99d9fe7),
	.w7(32'hbb37b9c6),
	.w8(32'hbaf1d052),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe37eca),
	.w1(32'hb95350ca),
	.w2(32'hbbcf41f0),
	.w3(32'h3b7716cb),
	.w4(32'h3b76c384),
	.w5(32'hbbb0f68a),
	.w6(32'h3b5b00d4),
	.w7(32'h3b6ebfed),
	.w8(32'hbb92a689),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08a764),
	.w1(32'hbb18a0c2),
	.w2(32'hbaa11317),
	.w3(32'hbbdd9e69),
	.w4(32'h3b327dc1),
	.w5(32'h3b755e8f),
	.w6(32'hbc1f220e),
	.w7(32'hbb10b5d4),
	.w8(32'h3afe6130),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd08e41),
	.w1(32'hbbabc5b2),
	.w2(32'hbb8b585b),
	.w3(32'hbbc3564e),
	.w4(32'hbb789904),
	.w5(32'hbb3a502f),
	.w6(32'hbbb8539b),
	.w7(32'hbb015bbb),
	.w8(32'hbb6ce62f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b9029),
	.w1(32'hb9e86ce3),
	.w2(32'hbb9dd994),
	.w3(32'hbb4c1809),
	.w4(32'hbab872e2),
	.w5(32'hbbb0dd11),
	.w6(32'hb9649990),
	.w7(32'hba1b0528),
	.w8(32'hbb20cfb4),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb031ee9),
	.w1(32'h398fc0b1),
	.w2(32'hba83f8b6),
	.w3(32'hbb32a86b),
	.w4(32'hbb2bbadc),
	.w5(32'h3b349f28),
	.w6(32'h3a9d88fa),
	.w7(32'hbb89c01f),
	.w8(32'hbb79bb35),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6de6ec),
	.w1(32'h3b34d1d3),
	.w2(32'hbad6a4e3),
	.w3(32'hba1c94bb),
	.w4(32'h3b9b7254),
	.w5(32'h3b775ed4),
	.w6(32'hba96ca27),
	.w7(32'h3c118a83),
	.w8(32'h3b92599f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16a7bd),
	.w1(32'hbbd3b252),
	.w2(32'h393e4beb),
	.w3(32'hb91b31d5),
	.w4(32'h3b657b7e),
	.w5(32'hbbf0070e),
	.w6(32'hb9a34ac0),
	.w7(32'h3bb30c0e),
	.w8(32'hbc351ae2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f4f1f),
	.w1(32'hbc01def9),
	.w2(32'h3c60e306),
	.w3(32'hbcd5edcd),
	.w4(32'hbc8fca0a),
	.w5(32'h3bd468ef),
	.w6(32'hbc9fd7bc),
	.w7(32'hbc23c678),
	.w8(32'hbb2a00b5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1675e),
	.w1(32'h3aee3f3d),
	.w2(32'h3b8a1865),
	.w3(32'h38f05c71),
	.w4(32'hba4a7eda),
	.w5(32'hbaeddad3),
	.w6(32'hbb1d8554),
	.w7(32'h3ae0f65c),
	.w8(32'h39f70c75),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba565160),
	.w1(32'hbb425a8e),
	.w2(32'hbb8c47fd),
	.w3(32'hbaeaea43),
	.w4(32'hba95685d),
	.w5(32'hbb807533),
	.w6(32'h3b1eb0b0),
	.w7(32'h3aeb0d0d),
	.w8(32'hba8e4fb0),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e052d),
	.w1(32'hbb087f0d),
	.w2(32'h3b2c136b),
	.w3(32'hbba29355),
	.w4(32'h3a8ea85b),
	.w5(32'h3b16aef9),
	.w6(32'hba211f02),
	.w7(32'h3a9e969c),
	.w8(32'h3a5eff0b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e88a2),
	.w1(32'hbc01cb07),
	.w2(32'hbbcccd95),
	.w3(32'h3b077fee),
	.w4(32'h3b4f66e2),
	.w5(32'hbb356ae7),
	.w6(32'h3a7908ab),
	.w7(32'h3ae3d92c),
	.w8(32'hbb3cb9d1),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc371691),
	.w1(32'hbb4b12ce),
	.w2(32'hba8203f4),
	.w3(32'hbc06299a),
	.w4(32'hbb1b7ed2),
	.w5(32'h3c5cd7c9),
	.w6(32'hbc07dcec),
	.w7(32'hbabc74a8),
	.w8(32'h3bb86461),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc814a90),
	.w1(32'hba2c1458),
	.w2(32'h3c7d2eb2),
	.w3(32'hbb8986ea),
	.w4(32'hbc4985b2),
	.w5(32'hbb8dda69),
	.w6(32'h3bd7d524),
	.w7(32'h3be9c05b),
	.w8(32'hbb23ae5c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e61e1),
	.w1(32'hbb34761d),
	.w2(32'hbb26b0b5),
	.w3(32'hbb2645c4),
	.w4(32'h39f5aed3),
	.w5(32'h3b3bf8d4),
	.w6(32'hb9dc5514),
	.w7(32'h3a887e3e),
	.w8(32'h3b41eaa3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998d5d5),
	.w1(32'h3b36f415),
	.w2(32'h3a46ef39),
	.w3(32'h3aa8c3c7),
	.w4(32'h3be5da12),
	.w5(32'hbbaf31e3),
	.w6(32'hbb3759ca),
	.w7(32'h3c079e14),
	.w8(32'h3b8f22d1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb6a829),
	.w1(32'h3d0f64ef),
	.w2(32'h3c59ba32),
	.w3(32'hbb6d8bd4),
	.w4(32'h3c80cdce),
	.w5(32'hbb3bed25),
	.w6(32'h3cc5bfbb),
	.w7(32'h3cb0ef5a),
	.w8(32'hbaa0bb0f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfda8cc),
	.w1(32'hbb77f5b3),
	.w2(32'hb90328f9),
	.w3(32'hba85622f),
	.w4(32'h3a8f8a55),
	.w5(32'h3c0e026d),
	.w6(32'h3b1d4246),
	.w7(32'h3b963931),
	.w8(32'hbba86a81),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba48116),
	.w1(32'hbbf626cb),
	.w2(32'hbb6fea24),
	.w3(32'hbabe1a98),
	.w4(32'hbbb4d0b6),
	.w5(32'h3b9674f6),
	.w6(32'h3af9a782),
	.w7(32'hbb9ffdff),
	.w8(32'h3b952e44),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba611982),
	.w1(32'hbb477d62),
	.w2(32'hbab8a1f0),
	.w3(32'hb98c23bc),
	.w4(32'h3b05a2d0),
	.w5(32'hbabbb6e3),
	.w6(32'h3b409dd6),
	.w7(32'h3ae85ec9),
	.w8(32'hbbc09852),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb601e5f),
	.w1(32'hbb707cdd),
	.w2(32'h3a0a3b3f),
	.w3(32'hbba42b12),
	.w4(32'h3ab129c0),
	.w5(32'h3a60fdd2),
	.w6(32'hbbb941a9),
	.w7(32'h3aef0a05),
	.w8(32'h3a509690),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b01611),
	.w1(32'h3aae654d),
	.w2(32'h3ba472b8),
	.w3(32'hbc3a07e9),
	.w4(32'hbb0a6d4d),
	.w5(32'h3b2f6bdb),
	.w6(32'hbc0c2837),
	.w7(32'h383b97dc),
	.w8(32'h3974a788),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce03d3b),
	.w1(32'hbca388d7),
	.w2(32'h3aef28c0),
	.w3(32'hbc6dd902),
	.w4(32'hbcdad722),
	.w5(32'h3b0d88af),
	.w6(32'hbb2d0539),
	.w7(32'hbb811879),
	.w8(32'hbb131a74),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadab47f),
	.w1(32'hbc05ca7b),
	.w2(32'hbc0c01e3),
	.w3(32'hbb1a7369),
	.w4(32'hbbd65226),
	.w5(32'hbb242eba),
	.w6(32'h3b0e2ff8),
	.w7(32'hbc2b998c),
	.w8(32'hbab3c6dc),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabb00e),
	.w1(32'hbaf9f991),
	.w2(32'hba0eb686),
	.w3(32'h3a3fbb95),
	.w4(32'h3aa5ef02),
	.w5(32'hbba2a340),
	.w6(32'h3bf21e14),
	.w7(32'hb8ab5954),
	.w8(32'h3a22e216),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d3719),
	.w1(32'hbbdf301d),
	.w2(32'h3a7f610c),
	.w3(32'hbb3be9c5),
	.w4(32'hba5d044e),
	.w5(32'hbb892c47),
	.w6(32'hb75cc144),
	.w7(32'hbbc1f25d),
	.w8(32'hb9cbcef9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba22cf9),
	.w1(32'h3b83fd0c),
	.w2(32'hb87d6a2d),
	.w3(32'hbb9bfae1),
	.w4(32'hbababdd7),
	.w5(32'h3b800d95),
	.w6(32'hbaed1d37),
	.w7(32'hba66eb2c),
	.w8(32'h3aaa69fa),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6a7d0),
	.w1(32'hbc2eda5b),
	.w2(32'hbbd6e378),
	.w3(32'h39def4ed),
	.w4(32'h3b893977),
	.w5(32'hbb8396db),
	.w6(32'h3b3a87ea),
	.w7(32'h3a06aa2b),
	.w8(32'hbc0eccf6),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bdaeb),
	.w1(32'h3c1be986),
	.w2(32'h3bf03c49),
	.w3(32'hbbe49c2c),
	.w4(32'h3c1e1e72),
	.w5(32'hbb8b88c5),
	.w6(32'hbc6cba34),
	.w7(32'hbbf0877b),
	.w8(32'hbb885bd6),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc63f8f),
	.w1(32'hbbb05af3),
	.w2(32'hbb8214db),
	.w3(32'hbc4468b6),
	.w4(32'hbb72d2ac),
	.w5(32'hbb592496),
	.w6(32'hbb0b00b3),
	.w7(32'hb9c0b9db),
	.w8(32'hbb3b36fb),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebf093),
	.w1(32'hbb63dd08),
	.w2(32'hbb0e30f4),
	.w3(32'h3b2c1a30),
	.w4(32'hbb5f418c),
	.w5(32'h3b3ac9aa),
	.w6(32'hba8cda8d),
	.w7(32'hbb847e02),
	.w8(32'hbab2c833),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1288a),
	.w1(32'hbacde5db),
	.w2(32'hb9c9e44f),
	.w3(32'hba1e4b61),
	.w4(32'h3a362975),
	.w5(32'h3b146764),
	.w6(32'h3997ec72),
	.w7(32'hbaf4b805),
	.w8(32'hba994c22),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab74f53),
	.w1(32'hbb1a6a9a),
	.w2(32'hb94cf150),
	.w3(32'h3bf53658),
	.w4(32'h3c0884fb),
	.w5(32'hba475bdb),
	.w6(32'h3b84d5fc),
	.w7(32'h38c27cc0),
	.w8(32'hbbc63626),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b6da2),
	.w1(32'h3ba2738a),
	.w2(32'h3b3bafa7),
	.w3(32'hbbc261a6),
	.w4(32'hbb705cf1),
	.w5(32'hbbfde4b7),
	.w6(32'hbc4877dc),
	.w7(32'hbb856cb3),
	.w8(32'hbc1944fa),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33a5de),
	.w1(32'hbb9d1e90),
	.w2(32'hbbd7819a),
	.w3(32'hbb19f2da),
	.w4(32'h3bbcf3c4),
	.w5(32'hba807e67),
	.w6(32'hbbfd0120),
	.w7(32'h3aba02e2),
	.w8(32'hb942817c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ee7b3),
	.w1(32'hbbc55214),
	.w2(32'hbbd3ea8e),
	.w3(32'hbac8c7f2),
	.w4(32'h39ee6785),
	.w5(32'h3aa01228),
	.w6(32'h3b187d2b),
	.w7(32'hba4f0513),
	.w8(32'hba33324c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe74970),
	.w1(32'h3b1d9794),
	.w2(32'hb8aecb77),
	.w3(32'h3b1f440e),
	.w4(32'h3ba5cd34),
	.w5(32'hbb9d20e3),
	.w6(32'hbb6eb780),
	.w7(32'h3b505775),
	.w8(32'hbb1cc614),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bd9be),
	.w1(32'hbae13e82),
	.w2(32'hba344bd1),
	.w3(32'hbbf85a53),
	.w4(32'hbab56589),
	.w5(32'h3b63f1fc),
	.w6(32'h3acab0b5),
	.w7(32'h3aeb3ad9),
	.w8(32'hba42709a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ce85e),
	.w1(32'hbc18c86e),
	.w2(32'hbc5d3b68),
	.w3(32'h3b489ca5),
	.w4(32'hba8ead67),
	.w5(32'hbb2b3321),
	.w6(32'h3b06717d),
	.w7(32'h3b98f088),
	.w8(32'h39c5915e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14ef97),
	.w1(32'hbc0b9056),
	.w2(32'hbb85a936),
	.w3(32'hbb624eb3),
	.w4(32'h3a957d97),
	.w5(32'h3b0422fb),
	.w6(32'hb9158dad),
	.w7(32'h3bb81a77),
	.w8(32'h3a8b7d1b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb946e94),
	.w1(32'hbbafc745),
	.w2(32'hbbb9aa06),
	.w3(32'hbbf0cf95),
	.w4(32'hba1c2e40),
	.w5(32'h3adceec4),
	.w6(32'hbb1f26cc),
	.w7(32'h3bd2fdb0),
	.w8(32'h3b4bee64),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4aee0),
	.w1(32'hbad783aa),
	.w2(32'h3b1dc078),
	.w3(32'h3b57ad06),
	.w4(32'h3b4d84a2),
	.w5(32'hba8ff164),
	.w6(32'hbb6b3079),
	.w7(32'h3a9be727),
	.w8(32'hbaa2977c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32185a),
	.w1(32'hbb84a286),
	.w2(32'hbb7151cd),
	.w3(32'hba3d1aa5),
	.w4(32'h3a6c0cfb),
	.w5(32'h3ab2bc1f),
	.w6(32'hbb0afdeb),
	.w7(32'h39ef83f9),
	.w8(32'h3ac9f10d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff7813),
	.w1(32'hba09a9cd),
	.w2(32'hbb217e42),
	.w3(32'h3ac1f2f3),
	.w4(32'h3b6b61a1),
	.w5(32'h3c4bc4f6),
	.w6(32'hb996489b),
	.w7(32'h3ac5c2c5),
	.w8(32'h3c01a3f3),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3df2f4),
	.w1(32'hbbee3f65),
	.w2(32'h3c255377),
	.w3(32'hbb881489),
	.w4(32'hbbf7912a),
	.w5(32'hbb2611cb),
	.w6(32'hbb68ea33),
	.w7(32'h3acf382a),
	.w8(32'hb905f321),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d2e8b),
	.w1(32'hbab51b46),
	.w2(32'h3a4de3a1),
	.w3(32'hbaa71352),
	.w4(32'h3af9a73f),
	.w5(32'hbbca829e),
	.w6(32'h3b743f49),
	.w7(32'h3a0df1fc),
	.w8(32'hbc23e63b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc939465),
	.w1(32'hbcb709fc),
	.w2(32'hbc9e397d),
	.w3(32'hbc05cd09),
	.w4(32'hbc125c26),
	.w5(32'h3ac04913),
	.w6(32'hbbed7474),
	.w7(32'hbc5c3020),
	.w8(32'hbbdd0869),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81ce78),
	.w1(32'hbb088f15),
	.w2(32'hbc08adfa),
	.w3(32'hbb94d1ce),
	.w4(32'hbb0b8c80),
	.w5(32'hbb46bd7c),
	.w6(32'hbb7ccac4),
	.w7(32'h3ab55f31),
	.w8(32'hbba777e7),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc544d7b),
	.w1(32'hbb85426c),
	.w2(32'h3acc3ec4),
	.w3(32'hbbc1739d),
	.w4(32'hbc51c5d6),
	.w5(32'hbbb7ac00),
	.w6(32'hbb371cbc),
	.w7(32'hbc0c8375),
	.w8(32'hbc08b30b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46ab9a),
	.w1(32'hbbf4dcc1),
	.w2(32'hbbae5248),
	.w3(32'hbbb9fdb4),
	.w4(32'hbb876cfc),
	.w5(32'hbb33eef0),
	.w6(32'hbbe45da5),
	.w7(32'hbbfe365a),
	.w8(32'hbbae439b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98aa795),
	.w1(32'hbb3308c9),
	.w2(32'hbaf312d0),
	.w3(32'hbaee78e1),
	.w4(32'h3b924060),
	.w5(32'hba9bb746),
	.w6(32'hbc45f3bf),
	.w7(32'hbb0be440),
	.w8(32'hbbd31d58),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd376a9),
	.w1(32'hbb61d957),
	.w2(32'hba509261),
	.w3(32'hbbe086bf),
	.w4(32'hbbd97c3a),
	.w5(32'h3b134f7b),
	.w6(32'hbb1e06df),
	.w7(32'hbc16a69c),
	.w8(32'h3aaeac54),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc06e4),
	.w1(32'hbb6b6486),
	.w2(32'hbba11510),
	.w3(32'h3aa76361),
	.w4(32'h3acd1561),
	.w5(32'hbc1844c6),
	.w6(32'h3a27eb2c),
	.w7(32'h3a42f617),
	.w8(32'h38d3d242),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d5dbf),
	.w1(32'hbbd339ba),
	.w2(32'hbc181bd8),
	.w3(32'hbc2ee17b),
	.w4(32'h3b32d601),
	.w5(32'hba961246),
	.w6(32'h3af2acc6),
	.w7(32'h3c4fbdbc),
	.w8(32'h3b813bf3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc87543),
	.w1(32'hbb52ca1c),
	.w2(32'h3b920fde),
	.w3(32'hbb638f81),
	.w4(32'h3a638ada),
	.w5(32'hbad8bcbc),
	.w6(32'hbbcf3531),
	.w7(32'hbb32d7f1),
	.w8(32'hbb8ad319),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1edd9),
	.w1(32'hbb886b6d),
	.w2(32'hbba8265c),
	.w3(32'hbb3f33ba),
	.w4(32'h3ac3c1cf),
	.w5(32'hb9335c51),
	.w6(32'h3b841305),
	.w7(32'h3b3c8c28),
	.w8(32'hbc274c0e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05175d),
	.w1(32'hbba47aeb),
	.w2(32'h3b6c6d13),
	.w3(32'hbb8768f2),
	.w4(32'hbab5f8ad),
	.w5(32'hbc10131d),
	.w6(32'hbb92cac6),
	.w7(32'hbc173e8d),
	.w8(32'hbc40cd31),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd44461),
	.w1(32'h3b73f9b4),
	.w2(32'h3af444d9),
	.w3(32'hbb715e5f),
	.w4(32'h3c2ecbd6),
	.w5(32'hbc1f2883),
	.w6(32'hbbd11f28),
	.w7(32'h3b1177a8),
	.w8(32'hbc4b6fa2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfc80e),
	.w1(32'hbbd587c2),
	.w2(32'hbc6d8913),
	.w3(32'hbc33afff),
	.w4(32'hbc0f0f05),
	.w5(32'hbbc84c58),
	.w6(32'hbc6f7efa),
	.w7(32'hbc9b1f41),
	.w8(32'hbb194561),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6e6f4),
	.w1(32'h3743295a),
	.w2(32'hbb8443a1),
	.w3(32'h3b1de03d),
	.w4(32'hbac918cb),
	.w5(32'h3acc4556),
	.w6(32'h3c39d158),
	.w7(32'hbadbe907),
	.w8(32'hbb1a2274),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafa1e2),
	.w1(32'hbbac814d),
	.w2(32'hbbce1d6e),
	.w3(32'hb90e2d27),
	.w4(32'h3abfabf6),
	.w5(32'hbb918adc),
	.w6(32'hbb5f844c),
	.w7(32'hbb5cabbc),
	.w8(32'h39fe916d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9c837),
	.w1(32'hbc2e072d),
	.w2(32'hba8db32f),
	.w3(32'hbbc11b53),
	.w4(32'hbb5e1d4f),
	.w5(32'hbc1a3bd0),
	.w6(32'hbba96979),
	.w7(32'h3c15971a),
	.w8(32'hbc33e6e5),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc212972),
	.w1(32'hbc30d3a3),
	.w2(32'hbc42b10f),
	.w3(32'hbc0bdcb1),
	.w4(32'hbbd3887c),
	.w5(32'h3b8e9b4b),
	.w6(32'hbc1b12ca),
	.w7(32'hbc2e6c91),
	.w8(32'hbb88c4af),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ad92c),
	.w1(32'hbab64f6b),
	.w2(32'hb9e07a69),
	.w3(32'hbb811f0e),
	.w4(32'h3b820de3),
	.w5(32'hbad23fbf),
	.w6(32'hbc11c67a),
	.w7(32'h3c037e9e),
	.w8(32'hbae00b78),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a891d13),
	.w1(32'h3b762786),
	.w2(32'hba10af68),
	.w3(32'hbb4507c4),
	.w4(32'h3b3e961c),
	.w5(32'h3b0878e9),
	.w6(32'hbb90203c),
	.w7(32'h3b3d0596),
	.w8(32'h3b547b6e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afaccb9),
	.w1(32'hbad70125),
	.w2(32'h399c4591),
	.w3(32'hba82bf87),
	.w4(32'h3a829318),
	.w5(32'h3b048b04),
	.w6(32'h3b52621d),
	.w7(32'h3aa8cacc),
	.w8(32'h3b7ec159),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cd142),
	.w1(32'hbb33fc53),
	.w2(32'hbb70fb96),
	.w3(32'hbb49d75f),
	.w4(32'hb91ee31b),
	.w5(32'hbb48021b),
	.w6(32'h3b1f3fc0),
	.w7(32'hba6f98e9),
	.w8(32'hbba61fd1),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7e040),
	.w1(32'hbb425dd3),
	.w2(32'hb9a73235),
	.w3(32'hbb3d46bc),
	.w4(32'hba15b732),
	.w5(32'h3933bb29),
	.w6(32'hbb0495e4),
	.w7(32'hbb597154),
	.w8(32'hb905b238),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6230b3),
	.w1(32'h3a90c553),
	.w2(32'h3b8006d8),
	.w3(32'hbaf0c185),
	.w4(32'h3a898e69),
	.w5(32'h3b7c5729),
	.w6(32'hbb3578e4),
	.w7(32'hba6fbd3f),
	.w8(32'h3b6c8af7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fe387),
	.w1(32'h3a12b9bf),
	.w2(32'h3b285951),
	.w3(32'h3b1eaecb),
	.w4(32'h3bb7a0d2),
	.w5(32'hbba8184e),
	.w6(32'h3b0519b0),
	.w7(32'h3b31b49f),
	.w8(32'h3bcd9952),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4286b7),
	.w1(32'h3cb3032a),
	.w2(32'h3ab97688),
	.w3(32'h3b84722b),
	.w4(32'h3c5c3654),
	.w5(32'h3bd1dddb),
	.w6(32'h3ce6e6d3),
	.w7(32'h3c8a6693),
	.w8(32'h3ad8de4c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb109a29),
	.w1(32'hbab31d24),
	.w2(32'h3a386bca),
	.w3(32'h3a7d7138),
	.w4(32'h3b84076d),
	.w5(32'h3a4c8d8c),
	.w6(32'h3b755864),
	.w7(32'h3bc77427),
	.w8(32'hbaaa0149),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11bf9b),
	.w1(32'hbb521b27),
	.w2(32'h3b52d8e3),
	.w3(32'hbbd0f477),
	.w4(32'hb8257510),
	.w5(32'h3b013e6c),
	.w6(32'hbc1e3d72),
	.w7(32'hbad6d5b2),
	.w8(32'h3abddc54),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba638bbc),
	.w1(32'h389bf92a),
	.w2(32'hba39c53d),
	.w3(32'hbb7ce7eb),
	.w4(32'hb9bb25ee),
	.w5(32'hbbc9e90a),
	.w6(32'hbad2a61e),
	.w7(32'h3ab37a88),
	.w8(32'hbb051386),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b9931),
	.w1(32'h3a951b86),
	.w2(32'hbbd48a86),
	.w3(32'hbaffd17c),
	.w4(32'h3a311f62),
	.w5(32'h3b79b08d),
	.w6(32'hbbbd47b0),
	.w7(32'hbadc0d55),
	.w8(32'hb8af5818),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bb1c7),
	.w1(32'hbac25cb6),
	.w2(32'h3a42fb78),
	.w3(32'h3b953b1e),
	.w4(32'h3b9d0740),
	.w5(32'hbc1a89eb),
	.w6(32'hba476633),
	.w7(32'h3ae98020),
	.w8(32'hbb1e6af5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14d659),
	.w1(32'h3bebb969),
	.w2(32'hbc610faf),
	.w3(32'hbb3671f1),
	.w4(32'h3c191ce7),
	.w5(32'hbb5b32ad),
	.w6(32'h3cbef455),
	.w7(32'hbb0c0739),
	.w8(32'h3b2fe24d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb462d8e),
	.w1(32'hbba9707f),
	.w2(32'h3b0acfa0),
	.w3(32'hbb03a620),
	.w4(32'hbbc2658d),
	.w5(32'hbc1b73b2),
	.w6(32'h3af26370),
	.w7(32'hbaed037c),
	.w8(32'h3a09f851),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c578171),
	.w1(32'h3cbdb7dc),
	.w2(32'h39c6f811),
	.w3(32'hbc5abf1d),
	.w4(32'h3bd6edb6),
	.w5(32'hbc138b38),
	.w6(32'h3cb28e7a),
	.w7(32'h3c626012),
	.w8(32'hbacb05a2),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba442ba),
	.w1(32'hbb155b00),
	.w2(32'hbbac9c59),
	.w3(32'hbba7cbae),
	.w4(32'hbb1679d3),
	.w5(32'h3be1fd65),
	.w6(32'h3a87ec38),
	.w7(32'hbafa32c9),
	.w8(32'hbb52d56f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01e3fb),
	.w1(32'hbbea090f),
	.w2(32'hbbebe074),
	.w3(32'hbb9f32c7),
	.w4(32'hbb8f1c0c),
	.w5(32'h3be95c40),
	.w6(32'hbbd61f06),
	.w7(32'hbb899973),
	.w8(32'h3cf8f7fb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc68acd),
	.w1(32'h3c297d63),
	.w2(32'h3c530ef3),
	.w3(32'h3c1a5fec),
	.w4(32'h3b959b0d),
	.w5(32'h389368f0),
	.w6(32'h3d4269a3),
	.w7(32'h3cd8733f),
	.w8(32'h3a199afb),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8980fda),
	.w1(32'h3a70ed7f),
	.w2(32'h3b8ab274),
	.w3(32'hbb445b18),
	.w4(32'hbb32c169),
	.w5(32'h3b82a09a),
	.w6(32'hba01bbf0),
	.w7(32'h3b20fc08),
	.w8(32'h3b504512),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf5b6b),
	.w1(32'hbba1ad26),
	.w2(32'hbbcadd28),
	.w3(32'h3c3f5404),
	.w4(32'h3b2ad418),
	.w5(32'h3b432ba8),
	.w6(32'h3b9ff9ed),
	.w7(32'hbb7828bf),
	.w8(32'hba5a2677),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf41bb7),
	.w1(32'hbbbce19c),
	.w2(32'hbbc9a80e),
	.w3(32'hb9c19b2b),
	.w4(32'h3b3fe4c7),
	.w5(32'hbb29421c),
	.w6(32'h3b2ddae2),
	.w7(32'h3c05356f),
	.w8(32'h3b34c641),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba08536),
	.w1(32'hbc190004),
	.w2(32'hbc254b18),
	.w3(32'h3b407180),
	.w4(32'hbbb253e9),
	.w5(32'hb9d65d62),
	.w6(32'h3b92dba0),
	.w7(32'hbbf1d579),
	.w8(32'hbaf807c7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eca32),
	.w1(32'hbbd8aa43),
	.w2(32'hbbb6e036),
	.w3(32'hb8d4ec61),
	.w4(32'hbac3f93b),
	.w5(32'hbab8eeb1),
	.w6(32'h3b4aad57),
	.w7(32'h3adb6528),
	.w8(32'hbb0e4d8d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e64d0),
	.w1(32'hbb6e6f2a),
	.w2(32'h3b3bef77),
	.w3(32'hbbeff07d),
	.w4(32'hbbd29f9e),
	.w5(32'h3b4584ce),
	.w6(32'hbbe0539f),
	.w7(32'hbbe5a978),
	.w8(32'h3aa527e7),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397acb29),
	.w1(32'hbadaab5b),
	.w2(32'hbad5bd58),
	.w3(32'h3b2aa540),
	.w4(32'hba04418b),
	.w5(32'h3b856d38),
	.w6(32'h3b00c380),
	.w7(32'hb9ce2ce5),
	.w8(32'hbb2a77de),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac31b69),
	.w1(32'hbba51cb5),
	.w2(32'hbab67d02),
	.w3(32'h3c02c224),
	.w4(32'h3b25ad35),
	.w5(32'hba745351),
	.w6(32'h3b30bed5),
	.w7(32'hbae7b2bc),
	.w8(32'hb875b391),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fe527),
	.w1(32'h3969f0e7),
	.w2(32'h3a85889d),
	.w3(32'hbba0a4e4),
	.w4(32'hbb3e5f15),
	.w5(32'hbb97100c),
	.w6(32'hbbcf9ba0),
	.w7(32'h3ab26249),
	.w8(32'hbb43c85c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa01fe8),
	.w1(32'h39d410bc),
	.w2(32'hbc0070d1),
	.w3(32'h3b9d4cfc),
	.w4(32'h3b96f7cb),
	.w5(32'hb9c2bf0b),
	.w6(32'h3b7fcc40),
	.w7(32'h3aa750cf),
	.w8(32'hba1f2e18),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba947882),
	.w1(32'hba8e5449),
	.w2(32'hba9f799b),
	.w3(32'hba29a090),
	.w4(32'hba25bf06),
	.w5(32'hb9743ba6),
	.w6(32'hba89d98c),
	.w7(32'hba5b5762),
	.w8(32'hbac3666d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aa3ca),
	.w1(32'hbae5203c),
	.w2(32'hba51b52b),
	.w3(32'hbb6c0764),
	.w4(32'hb90c1a27),
	.w5(32'h3a10c3cf),
	.w6(32'hbbadf2ea),
	.w7(32'h3a377373),
	.w8(32'h3b5269ce),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02e452),
	.w1(32'h39c13edd),
	.w2(32'h3a74ffac),
	.w3(32'hbad7205f),
	.w4(32'h3b0bcf03),
	.w5(32'h3b1d74e5),
	.w6(32'hbb1d51d0),
	.w7(32'h3a8d500e),
	.w8(32'h388caa08),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaa53d),
	.w1(32'hbacb4ee9),
	.w2(32'hba6c3711),
	.w3(32'hba29c339),
	.w4(32'hba4bfd30),
	.w5(32'h389e876b),
	.w6(32'hba96b52b),
	.w7(32'hbad8ac34),
	.w8(32'hb99fadf0),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b2925),
	.w1(32'hbae1bf34),
	.w2(32'hbb7e8dc8),
	.w3(32'hba506997),
	.w4(32'h3a0c07bb),
	.w5(32'hbb842af3),
	.w6(32'hba0ab012),
	.w7(32'h3aee01d2),
	.w8(32'hbb44dc93),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a70c2),
	.w1(32'hbb507adc),
	.w2(32'hbb5e0865),
	.w3(32'hbb1bd007),
	.w4(32'hbace6a80),
	.w5(32'hbb195c51),
	.w6(32'hbaf8d3d6),
	.w7(32'h3a20c6c0),
	.w8(32'h398e133a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6698ed),
	.w1(32'hba5c2e6f),
	.w2(32'hba22dc52),
	.w3(32'hba6bb98b),
	.w4(32'hba946fcd),
	.w5(32'hb936e696),
	.w6(32'h3862709a),
	.w7(32'hbaf031ec),
	.w8(32'hb9c851d8),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01fe09),
	.w1(32'hba782c50),
	.w2(32'hbb09b4d5),
	.w3(32'hbad76a99),
	.w4(32'hba47e07f),
	.w5(32'hbaea595c),
	.w6(32'hba8bbbf8),
	.w7(32'h39ac1c29),
	.w8(32'hbabb0227),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f0730),
	.w1(32'h394a9881),
	.w2(32'h395fe1b0),
	.w3(32'hba655b28),
	.w4(32'hba4a15df),
	.w5(32'h3a6c3d18),
	.w6(32'hba39851a),
	.w7(32'hb9d52f7e),
	.w8(32'h3a436a6d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d589c),
	.w1(32'hb89284f8),
	.w2(32'h393f8a12),
	.w3(32'h389f9d5e),
	.w4(32'h38194145),
	.w5(32'hba8b2c7d),
	.w6(32'hb7024f5b),
	.w7(32'hba17334b),
	.w8(32'hbaa7442a),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a4b6),
	.w1(32'hbaa83d51),
	.w2(32'hbb0b479d),
	.w3(32'hba9088c5),
	.w4(32'hbad24d5d),
	.w5(32'h3a0a54f9),
	.w6(32'hba426ec9),
	.w7(32'hba9fd63f),
	.w8(32'h39a3fe36),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3530cf),
	.w1(32'h3a139fb1),
	.w2(32'h3a6b32e0),
	.w3(32'h38884b82),
	.w4(32'h39ea3099),
	.w5(32'h3a39bafd),
	.w6(32'h39a98175),
	.w7(32'h3a8307f9),
	.w8(32'hb90c0f7c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb446ea5),
	.w1(32'hbabda6cf),
	.w2(32'hb9227af3),
	.w3(32'hbacd88a2),
	.w4(32'hb8cdde8d),
	.w5(32'h3a028644),
	.w6(32'hbafbaac3),
	.w7(32'hb964a9f6),
	.w8(32'hba13fbed),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba185c8),
	.w1(32'hbad71e20),
	.w2(32'hbb8ffdf2),
	.w3(32'hbb74c5d6),
	.w4(32'hb9bbdc6e),
	.w5(32'hba57617d),
	.w6(32'hbb9fd2c9),
	.w7(32'h3ac759e1),
	.w8(32'h3acc60a8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb774894),
	.w1(32'h3a15e34b),
	.w2(32'hbb1d5811),
	.w3(32'hbb11c7ca),
	.w4(32'h3ad1eba4),
	.w5(32'hbb03661b),
	.w6(32'hb9966d7f),
	.w7(32'h3ba52c10),
	.w8(32'h3a4cb1b8),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d65a5),
	.w1(32'hba01f66a),
	.w2(32'hbb674aa5),
	.w3(32'hbaafa621),
	.w4(32'hb97ec7c2),
	.w5(32'hba8aa153),
	.w6(32'hbb0bdca5),
	.w7(32'h3a45e3b4),
	.w8(32'hb825db3c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1deae3),
	.w1(32'h381c6015),
	.w2(32'hba846fd1),
	.w3(32'h3a91ca91),
	.w4(32'h377f6428),
	.w5(32'h392f5b63),
	.w6(32'hba020e67),
	.w7(32'hba619e50),
	.w8(32'hbae069b9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba742657),
	.w1(32'hba899db9),
	.w2(32'hba40ac1f),
	.w3(32'hba2aebf9),
	.w4(32'hb9d1af4b),
	.w5(32'h3a412b65),
	.w6(32'hbb16bc83),
	.w7(32'hba97c7e5),
	.w8(32'h3a77de0f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ebe00),
	.w1(32'h3a23ae75),
	.w2(32'h3a804611),
	.w3(32'h39c6a105),
	.w4(32'h399aac0e),
	.w5(32'hbac6d788),
	.w6(32'h3a29c58a),
	.w7(32'h3a7e8dee),
	.w8(32'h3a175945),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d6432),
	.w1(32'h3aad23a7),
	.w2(32'h3a9eaf3f),
	.w3(32'hb9aebe29),
	.w4(32'hb96222a0),
	.w5(32'hb9d6532b),
	.w6(32'h3a737ae0),
	.w7(32'hbacf75cb),
	.w8(32'hba3591b5),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ac5aa),
	.w1(32'hbb118f97),
	.w2(32'hbaa91023),
	.w3(32'hbaffe4b7),
	.w4(32'hb9cbdb35),
	.w5(32'hbac7593f),
	.w6(32'hbb10a5ae),
	.w7(32'h3a7de7fd),
	.w8(32'hbac6ff7d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb411741),
	.w1(32'hbb2f9320),
	.w2(32'hbae86447),
	.w3(32'hbb13b8a7),
	.w4(32'hbb099545),
	.w5(32'h3aad2d86),
	.w6(32'hbaefccfa),
	.w7(32'hba655f3b),
	.w8(32'h3a11cf16),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e65402),
	.w1(32'hbac11d7b),
	.w2(32'hb9faae86),
	.w3(32'h39a59c75),
	.w4(32'hba465e13),
	.w5(32'hba873f65),
	.w6(32'hb9ad6008),
	.w7(32'hbaabe1ff),
	.w8(32'hbad44598),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b577d),
	.w1(32'hbab39e64),
	.w2(32'hba87255d),
	.w3(32'hba810c49),
	.w4(32'hb89ceb63),
	.w5(32'hba3a6120),
	.w6(32'hba898945),
	.w7(32'hbaad619f),
	.w8(32'hb9e9103d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b49064),
	.w1(32'h3924fb09),
	.w2(32'h39dd7f39),
	.w3(32'hba80d15b),
	.w4(32'hbac100fc),
	.w5(32'hba65e9c9),
	.w6(32'h3aa01255),
	.w7(32'h3a43776f),
	.w8(32'hb9bc8a0d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10917e),
	.w1(32'hbb06d148),
	.w2(32'hbaed9bc7),
	.w3(32'hbaa31a02),
	.w4(32'hb9a476a3),
	.w5(32'hba775d43),
	.w6(32'hba580307),
	.w7(32'hb9b5730e),
	.w8(32'hba97af54),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38942d82),
	.w1(32'h3998d477),
	.w2(32'h3a1e0fd8),
	.w3(32'hb927e0b7),
	.w4(32'hb9c1a903),
	.w5(32'hb9ed04fc),
	.w6(32'h39c0033d),
	.w7(32'hb96ac811),
	.w8(32'h39b5a4b4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae65d73),
	.w1(32'hb8be58e2),
	.w2(32'hbb2c74e1),
	.w3(32'hb9cd44dc),
	.w4(32'h3ab05a48),
	.w5(32'h39633426),
	.w6(32'hbac64431),
	.w7(32'h39a60583),
	.w8(32'h39c1e5e1),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d44aba),
	.w1(32'hba200ceb),
	.w2(32'h39194cdc),
	.w3(32'hb9babe32),
	.w4(32'h394053ef),
	.w5(32'h3a5dcab4),
	.w6(32'hb99ce398),
	.w7(32'h398aae2b),
	.w8(32'h3a8d36ef),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2d2dc),
	.w1(32'hba1ecdb4),
	.w2(32'h39d88433),
	.w3(32'hbb527a22),
	.w4(32'hbb148432),
	.w5(32'hb7a153cf),
	.w6(32'hbaa1280d),
	.w7(32'h3b0394a3),
	.w8(32'h3ae3c285),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule