module layer_8_featuremap_12(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe03367),
	.w1(32'h3bc9effb),
	.w2(32'h3c197ca2),
	.w3(32'hbc6c684a),
	.w4(32'h3bc283b7),
	.w5(32'h3b827749),
	.w6(32'hbc5c9dac),
	.w7(32'h3b886061),
	.w8(32'h3b0bdd7f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45dd3c),
	.w1(32'h3c59776e),
	.w2(32'h3bbbdc27),
	.w3(32'h3c51c646),
	.w4(32'h3c4c9f84),
	.w5(32'h3b8614bf),
	.w6(32'h3c3a1439),
	.w7(32'h3c2b1a24),
	.w8(32'h3b6a6f6a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e319d),
	.w1(32'h3bfa908e),
	.w2(32'h3c094dc1),
	.w3(32'h3c3500f9),
	.w4(32'h3c8971a6),
	.w5(32'h3c944b15),
	.w6(32'h3c1b76bb),
	.w7(32'h3c0465be),
	.w8(32'h3bfc94c6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8000f),
	.w1(32'hbcf4ff51),
	.w2(32'hbd285981),
	.w3(32'hba34d03d),
	.w4(32'hbd2b9217),
	.w5(32'hbd8429b7),
	.w6(32'hbc2a62c3),
	.w7(32'hbcd2bd22),
	.w8(32'hbd28e34f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce1079e),
	.w1(32'h3bf4a851),
	.w2(32'h3be16e84),
	.w3(32'hbd2c996d),
	.w4(32'h3c10546a),
	.w5(32'h3bffead3),
	.w6(32'hbcdacbb4),
	.w7(32'h3baff951),
	.w8(32'h3b1a6a92),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3fd12),
	.w1(32'hbae8f806),
	.w2(32'hb9b6443b),
	.w3(32'h3c21501d),
	.w4(32'hbb04289a),
	.w5(32'hbc99c268),
	.w6(32'h3c09e9b8),
	.w7(32'hbb0b296d),
	.w8(32'hbc259282),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e6e57),
	.w1(32'hbc52a8f7),
	.w2(32'h3b79ce1e),
	.w3(32'hbc14fdc9),
	.w4(32'hbbe92040),
	.w5(32'h3c4d9abc),
	.w6(32'h3b8230f6),
	.w7(32'hbc164236),
	.w8(32'h3c05e9e5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d41ab),
	.w1(32'h3bb8a480),
	.w2(32'h3bb89aac),
	.w3(32'h3c6418a8),
	.w4(32'h3c1ac2c5),
	.w5(32'h3c7411d7),
	.w6(32'h3c3b51c0),
	.w7(32'hbb80f4b4),
	.w8(32'hba70588d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e92fc),
	.w1(32'h3bb848e7),
	.w2(32'hbb24b08d),
	.w3(32'h3c1c84e0),
	.w4(32'h3a471d91),
	.w5(32'hbba18bb2),
	.w6(32'h3b428932),
	.w7(32'hbbbf59f3),
	.w8(32'hbc399509),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8da674),
	.w1(32'h3a9b77c8),
	.w2(32'hbb8a8728),
	.w3(32'hbabf1164),
	.w4(32'h3aefa3d9),
	.w5(32'h3c5f67ec),
	.w6(32'hb9e78516),
	.w7(32'h3c8cfa90),
	.w8(32'hb92000f1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4d7bc),
	.w1(32'hbcc5b1f2),
	.w2(32'hbb1d326b),
	.w3(32'h3ad83464),
	.w4(32'hbbf76b66),
	.w5(32'hb997e8f3),
	.w6(32'h3bda7470),
	.w7(32'hbca5fc67),
	.w8(32'hbbca7513),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb818010),
	.w1(32'hbb04973e),
	.w2(32'h3bb55748),
	.w3(32'hba913a54),
	.w4(32'hbaed51f3),
	.w5(32'h3c4d159e),
	.w6(32'h3914fb6e),
	.w7(32'h3beee001),
	.w8(32'h3c1ada29),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ea722),
	.w1(32'hbc4a01f0),
	.w2(32'h3cf2a58d),
	.w3(32'h3be3a1c2),
	.w4(32'hbbe923b1),
	.w5(32'h3c296c9b),
	.w6(32'h3cb1161d),
	.w7(32'hbc258999),
	.w8(32'hbb401950),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1db41),
	.w1(32'hbc244ee7),
	.w2(32'h3917b962),
	.w3(32'hb961daeb),
	.w4(32'hbbab48ab),
	.w5(32'h3b74a7f3),
	.w6(32'h3c8c7888),
	.w7(32'hbb8ca526),
	.w8(32'h3bb8321b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a4626),
	.w1(32'hbc317868),
	.w2(32'h3af52329),
	.w3(32'h3bd31860),
	.w4(32'hbb9ec8e4),
	.w5(32'h3c2f9b42),
	.w6(32'h3bec4799),
	.w7(32'hbbdb6a38),
	.w8(32'h3bdad37f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb331589),
	.w1(32'hba10c8f7),
	.w2(32'hbbb687bf),
	.w3(32'h3b495ac8),
	.w4(32'h3c529639),
	.w5(32'h3c0519e6),
	.w6(32'h3a682ead),
	.w7(32'hbbb99519),
	.w8(32'hbc05dabd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb865519),
	.w1(32'hbbb5c494),
	.w2(32'h3c8333ef),
	.w3(32'h3c2d4ffb),
	.w4(32'h3c94e7cb),
	.w5(32'hbc9b047a),
	.w6(32'hbac6bd6d),
	.w7(32'hbb877715),
	.w8(32'hbc46b77b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e850ba),
	.w1(32'h3c209895),
	.w2(32'h3b9f8757),
	.w3(32'h3bd19281),
	.w4(32'h3c1343a6),
	.w5(32'h3c07ca6c),
	.w6(32'h3bd7ea17),
	.w7(32'h3c1056e5),
	.w8(32'h3ba8b294),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e6170),
	.w1(32'hbcf81bfb),
	.w2(32'hb9c50f21),
	.w3(32'h3bb76f1f),
	.w4(32'hbc48ea00),
	.w5(32'h3c236337),
	.w6(32'h3ca2455c),
	.w7(32'hbbcbc4da),
	.w8(32'h3bd4cfa4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c1fc5),
	.w1(32'hbcf6c7e8),
	.w2(32'hbc99b913),
	.w3(32'h3b3e216b),
	.w4(32'hbcc6ceb5),
	.w5(32'hbc85d5a7),
	.w6(32'h3c866ed5),
	.w7(32'hbc1ff5ed),
	.w8(32'hba3938db),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd4c8f),
	.w1(32'hbd01ce99),
	.w2(32'h3b15f2df),
	.w3(32'h3c26addb),
	.w4(32'hbcab1887),
	.w5(32'h3c10ece8),
	.w6(32'h3c5d8be9),
	.w7(32'hbcb882fd),
	.w8(32'h3c172ce3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd9c9),
	.w1(32'hbab92712),
	.w2(32'hbb92a958),
	.w3(32'h3bec7720),
	.w4(32'hbc3bdfd5),
	.w5(32'h3cdd438a),
	.w6(32'h3ba4a641),
	.w7(32'h3c16641d),
	.w8(32'h3c0897c3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e277d),
	.w1(32'hbcd5bcbd),
	.w2(32'h3c0881e5),
	.w3(32'h3cc17e37),
	.w4(32'hbbfd2768),
	.w5(32'h3b73c2c5),
	.w6(32'h3c52f5d2),
	.w7(32'hbce52354),
	.w8(32'h3ca14478),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5987c),
	.w1(32'hbcdd08f8),
	.w2(32'hbb80f99c),
	.w3(32'h3c8b27f8),
	.w4(32'hbc8cc724),
	.w5(32'h3c11dde2),
	.w6(32'h3bf12fb2),
	.w7(32'hbcbd88dd),
	.w8(32'h3b397eb7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8cb0f),
	.w1(32'h3c856617),
	.w2(32'h3ccaf857),
	.w3(32'h3bfc0b13),
	.w4(32'h3ca219ca),
	.w5(32'h3d1002b8),
	.w6(32'h3be82751),
	.w7(32'h3c95d030),
	.w8(32'h3cae14f3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc20f2),
	.w1(32'h3ba67cb9),
	.w2(32'hbb2ad197),
	.w3(32'h3ce0e251),
	.w4(32'h393da723),
	.w5(32'hbc7e3174),
	.w6(32'h3ce85622),
	.w7(32'h3b979dcf),
	.w8(32'hbbb4f509),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b517427),
	.w1(32'hbc5d760d),
	.w2(32'h3c36eea7),
	.w3(32'hbb0759b9),
	.w4(32'hbb8fc16e),
	.w5(32'h3cd30728),
	.w6(32'h3a7a9e59),
	.w7(32'hbc6ee6e3),
	.w8(32'h3c8dc564),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0262f6),
	.w1(32'hbdb1ef17),
	.w2(32'hbdd2e184),
	.w3(32'hbcd6ec46),
	.w4(32'hbb922582),
	.w5(32'hbdae52f9),
	.w6(32'hbd896fc9),
	.w7(32'hbd80cf71),
	.w8(32'hbd6551e5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9df2f),
	.w1(32'h3b3d00e2),
	.w2(32'hbb889a92),
	.w3(32'hbca1d439),
	.w4(32'h3b2eb71a),
	.w5(32'hbc3adac4),
	.w6(32'hbbaed5e3),
	.w7(32'hbad2ae4d),
	.w8(32'hbc2b92e6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3433ba),
	.w1(32'h3b2aca2b),
	.w2(32'h3b856d66),
	.w3(32'hb9a307b4),
	.w4(32'h3b9d517b),
	.w5(32'h3b7a42ec),
	.w6(32'hbb809515),
	.w7(32'h3b09bf29),
	.w8(32'hbb2531de),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922da14),
	.w1(32'hbcda2e03),
	.w2(32'hbccad7e1),
	.w3(32'h39995c58),
	.w4(32'hbcfcc87a),
	.w5(32'hbcdd9aec),
	.w6(32'hbb38dd31),
	.w7(32'hbc8ee867),
	.w8(32'hbcb3ddf6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b874c),
	.w1(32'hbc0d50c6),
	.w2(32'h3bc0e2d4),
	.w3(32'hbd06d6c6),
	.w4(32'hbaaab1d4),
	.w5(32'h3c4dacde),
	.w6(32'hbc9bff4e),
	.w7(32'hbbd51e10),
	.w8(32'h3bc0dc18),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc214e0),
	.w1(32'hbb307668),
	.w2(32'hb91399f2),
	.w3(32'h3b06c35c),
	.w4(32'hbadbab1b),
	.w5(32'h3a1e10ca),
	.w6(32'hbb85f596),
	.w7(32'hbab8e0bb),
	.w8(32'h3ae50250),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb157ff7),
	.w1(32'hba5f372b),
	.w2(32'h3b62c7d3),
	.w3(32'h3a6847a7),
	.w4(32'h3b71b73d),
	.w5(32'h3bf67941),
	.w6(32'hbada9cad),
	.w7(32'hbb0fb602),
	.w8(32'hbc2cba7a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c877109),
	.w1(32'h3b4c3bff),
	.w2(32'h3b81bf73),
	.w3(32'h3b950611),
	.w4(32'h3bffd26e),
	.w5(32'h35e52a79),
	.w6(32'h399c9695),
	.w7(32'h3c12887a),
	.w8(32'h3bd405bd),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f3166),
	.w1(32'hbc28fa85),
	.w2(32'hbc694240),
	.w3(32'hbafc7071),
	.w4(32'hbad50f0d),
	.w5(32'hbc2b431f),
	.w6(32'hbad03f2c),
	.w7(32'h3b8e6d11),
	.w8(32'hbc52c43c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd56a1b),
	.w1(32'hbcfd28cd),
	.w2(32'hbb5697cc),
	.w3(32'hbad2ccea),
	.w4(32'hbb5a0b01),
	.w5(32'h3ca06dcf),
	.w6(32'h3bea4531),
	.w7(32'hbc3364bb),
	.w8(32'h3c335658),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb499be3),
	.w1(32'h39b7040e),
	.w2(32'h3c0c0c56),
	.w3(32'h3a943cfa),
	.w4(32'h3c0345e5),
	.w5(32'h3bcd3f68),
	.w6(32'h3bf3f71a),
	.w7(32'h3c3b4a15),
	.w8(32'hba45cfed),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65ca5a),
	.w1(32'hbacfd0c5),
	.w2(32'hbc4a1f9f),
	.w3(32'h3b2914bf),
	.w4(32'hbb804ddc),
	.w5(32'hbc94b26b),
	.w6(32'h3c258faa),
	.w7(32'hbc5a16da),
	.w8(32'hbc9cf8e8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb711560),
	.w1(32'h3c6804c5),
	.w2(32'h3c020ae1),
	.w3(32'h3ab67f48),
	.w4(32'h3c804b63),
	.w5(32'h3bb43baa),
	.w6(32'hbc5e822f),
	.w7(32'h3c99f618),
	.w8(32'h3beca0ee),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf52da),
	.w1(32'h3baf6876),
	.w2(32'h3c803804),
	.w3(32'h3c5263d4),
	.w4(32'h3c031f54),
	.w5(32'h3c56bafc),
	.w6(32'h3b0f971e),
	.w7(32'hbc58b05a),
	.w8(32'hbb40c6fd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fe239),
	.w1(32'hbc6b5331),
	.w2(32'h38d2db3a),
	.w3(32'h3bdcd031),
	.w4(32'hbbf3efd8),
	.w5(32'h3b7dcb93),
	.w6(32'h3c81a855),
	.w7(32'hbb978810),
	.w8(32'h3c241f3a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86347d),
	.w1(32'h3c5139b7),
	.w2(32'h3b3864cc),
	.w3(32'h3bac76be),
	.w4(32'h3c031efb),
	.w5(32'hbaec2230),
	.w6(32'h3bba1791),
	.w7(32'h3c15ac27),
	.w8(32'h3ab7c66a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba38558),
	.w1(32'hbc69008c),
	.w2(32'hbcabf864),
	.w3(32'h3aa5013f),
	.w4(32'hbcbaf62e),
	.w5(32'hbceb3cf9),
	.w6(32'hb91f36c8),
	.w7(32'hbc812991),
	.w8(32'hbcc74f82),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc425d16),
	.w1(32'hbc94b7ed),
	.w2(32'h3be5c8f8),
	.w3(32'hbbcb3912),
	.w4(32'hbbcdab6d),
	.w5(32'h3acbaf7a),
	.w6(32'hbb9e8117),
	.w7(32'hba4249f8),
	.w8(32'h3c61d421),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba67242),
	.w1(32'hbc327f0f),
	.w2(32'h3af24e81),
	.w3(32'hbbe24c68),
	.w4(32'hbc1f764a),
	.w5(32'h3c5bd300),
	.w6(32'h3c6878d4),
	.w7(32'hbbdcc881),
	.w8(32'h3c9cfd05),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1a97f),
	.w1(32'hbc704d0d),
	.w2(32'hbbaf1382),
	.w3(32'h3c0f9136),
	.w4(32'hbc0e634d),
	.w5(32'hb993141f),
	.w6(32'h3b3cb260),
	.w7(32'hbb695d73),
	.w8(32'hbc2e4416),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e8d1d),
	.w1(32'hbc950a8d),
	.w2(32'hbc3cf78c),
	.w3(32'h3c069819),
	.w4(32'hbc3e5de8),
	.w5(32'hbb126cc8),
	.w6(32'h3c74b3c4),
	.w7(32'hbbbbc761),
	.w8(32'hbb8eb83a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b314f),
	.w1(32'h3b42f80b),
	.w2(32'hbbbbb8ee),
	.w3(32'hbc4947d0),
	.w4(32'hbab69a84),
	.w5(32'hbb526dac),
	.w6(32'hbcd7ec4b),
	.w7(32'h3b7d16d6),
	.w8(32'h3898d3d1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c83a2),
	.w1(32'hbb6c7dda),
	.w2(32'h3d94b616),
	.w3(32'h3b49e642),
	.w4(32'h3dbf3e77),
	.w5(32'hbe81fa48),
	.w6(32'h3b42dce4),
	.w7(32'hbe13f16b),
	.w8(32'h3e3e8c5b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8b4abb),
	.w1(32'h3c0d0edb),
	.w2(32'h3c4d6038),
	.w3(32'h3e2e5601),
	.w4(32'h3acbb9f9),
	.w5(32'h3c7046ef),
	.w6(32'hbd2fcf61),
	.w7(32'hba83d343),
	.w8(32'h3c0aa5fc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb35b2d),
	.w1(32'hbc1f2460),
	.w2(32'hbc7a681d),
	.w3(32'hbb6e0c6d),
	.w4(32'hbc5f32ea),
	.w5(32'hbc9dd53d),
	.w6(32'h3b3b5cb4),
	.w7(32'h3bbfb41e),
	.w8(32'hbb9d961b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43810d),
	.w1(32'hbc82fc11),
	.w2(32'hbb2140aa),
	.w3(32'hbb5fa26c),
	.w4(32'hbbc9db7c),
	.w5(32'h3c8a9c90),
	.w6(32'hbb2ce45e),
	.w7(32'hbbdf7cf9),
	.w8(32'hba4b3397),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba38c2e),
	.w1(32'hbbcd6a39),
	.w2(32'h3a3ad7aa),
	.w3(32'h3b6f2974),
	.w4(32'hbc468adc),
	.w5(32'h3c0b73cd),
	.w6(32'h3b200500),
	.w7(32'hbb7c4eb6),
	.w8(32'h3d085d7c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b523793),
	.w1(32'hbb2a76a5),
	.w2(32'hbca4435d),
	.w3(32'h3c876703),
	.w4(32'hbc7a003e),
	.w5(32'hb92e4cdf),
	.w6(32'hbc68852e),
	.w7(32'hbb75d9b6),
	.w8(32'h3c58373c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc468f5a),
	.w1(32'hbb0bad52),
	.w2(32'hbc4b826d),
	.w3(32'h3cbceaf3),
	.w4(32'h3b20d029),
	.w5(32'hbc028be3),
	.w6(32'h3aa0b4fc),
	.w7(32'hb9684efc),
	.w8(32'hbbc4e76a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cc2e9),
	.w1(32'hbbeaef27),
	.w2(32'h3b6c6bdd),
	.w3(32'hba9d5a8e),
	.w4(32'hba9a31e2),
	.w5(32'h3c18be17),
	.w6(32'hb9c2c4f4),
	.w7(32'h3ad227c2),
	.w8(32'h3c1c8cdf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda49db),
	.w1(32'h3befa383),
	.w2(32'h3ad5797d),
	.w3(32'h3bcbf23f),
	.w4(32'hba81859b),
	.w5(32'hbbda8a82),
	.w6(32'h3c59325c),
	.w7(32'h3a92cf01),
	.w8(32'hbc11b2a5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65484b),
	.w1(32'hbb225639),
	.w2(32'hbc22049c),
	.w3(32'hbc3205df),
	.w4(32'hbb64eded),
	.w5(32'hbc0591c7),
	.w6(32'hbb906b48),
	.w7(32'hbb6ec30c),
	.w8(32'hbc1f73a6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a40c8d),
	.w1(32'hbb83d73a),
	.w2(32'h3c9bc92d),
	.w3(32'hbba33f29),
	.w4(32'h3c125d2f),
	.w5(32'h3b59f897),
	.w6(32'hbc08189c),
	.w7(32'hbbb91d99),
	.w8(32'h3c8cdcd3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1857f),
	.w1(32'h3b327359),
	.w2(32'h3b43d5cc),
	.w3(32'h3a84eaef),
	.w4(32'h3c9ff6d5),
	.w5(32'h3c858eb3),
	.w6(32'h3c796c52),
	.w7(32'h3c2c6b13),
	.w8(32'h3c43d5cd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb479699),
	.w1(32'hbc0799e8),
	.w2(32'h3be4696a),
	.w3(32'h3c84afe7),
	.w4(32'h3b119c91),
	.w5(32'hbbd3773a),
	.w6(32'hbb9078cf),
	.w7(32'hbbd9f19b),
	.w8(32'hbc1b1793),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389dd22f),
	.w1(32'h39faacd3),
	.w2(32'hbc4a8eb1),
	.w3(32'hbc0f5c77),
	.w4(32'hbbbec73c),
	.w5(32'hbc81adae),
	.w6(32'h3bcb36ca),
	.w7(32'h3b43bb26),
	.w8(32'hbbc501f7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e3837),
	.w1(32'hbc911707),
	.w2(32'hbc0150fb),
	.w3(32'h3a1d5e8e),
	.w4(32'hbcd772f9),
	.w5(32'h3d187f5f),
	.w6(32'h3bf758d8),
	.w7(32'h3c0e90aa),
	.w8(32'hbc3d89c0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c959a73),
	.w1(32'h3ac87e1b),
	.w2(32'h3c36647e),
	.w3(32'hbbd8db65),
	.w4(32'h3a10fa55),
	.w5(32'h3c713e3f),
	.w6(32'h3c1d90fb),
	.w7(32'hbb80b11f),
	.w8(32'h3c274ca2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21ba79),
	.w1(32'hba84f99b),
	.w2(32'hbb19aa61),
	.w3(32'h39ff0fee),
	.w4(32'hba99c4ea),
	.w5(32'hbb5327a7),
	.w6(32'hbb3dc0e1),
	.w7(32'h39c5dede),
	.w8(32'hbae5f468),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87f404),
	.w1(32'h3c194121),
	.w2(32'h3aff073c),
	.w3(32'h3c1c312f),
	.w4(32'h3c34c7ba),
	.w5(32'h399905c1),
	.w6(32'h3bd97be2),
	.w7(32'h3c22f806),
	.w8(32'h3b1ec74d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d233e),
	.w1(32'hbc7937be),
	.w2(32'hbb8b6763),
	.w3(32'hb8bc8fce),
	.w4(32'hbc7530fc),
	.w5(32'hbbafbd7b),
	.w6(32'hba835c02),
	.w7(32'hbc05ca6b),
	.w8(32'h3be7a640),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07e79f),
	.w1(32'hbb33709e),
	.w2(32'h3be1441f),
	.w3(32'h3c39c302),
	.w4(32'hb92f7557),
	.w5(32'h3c553f14),
	.w6(32'h3c5a19e3),
	.w7(32'hbb8c9143),
	.w8(32'h3bf3eeb5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985428a),
	.w1(32'hbc93d8f1),
	.w2(32'hbc309e89),
	.w3(32'h3b5870d7),
	.w4(32'h3c3bd918),
	.w5(32'hbc160612),
	.w6(32'hbb0545aa),
	.w7(32'h3c3b9656),
	.w8(32'h3c22421b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dd889),
	.w1(32'hbb6c0f32),
	.w2(32'hbbe45973),
	.w3(32'hbc23e0b7),
	.w4(32'h3b990bc5),
	.w5(32'h3b4b3304),
	.w6(32'h3ccd406b),
	.w7(32'h3bd5f119),
	.w8(32'h3b7c631c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc019fbe),
	.w1(32'hbb53f6e0),
	.w2(32'hbc91a621),
	.w3(32'h3a6e28e6),
	.w4(32'hbbd5b16b),
	.w5(32'h3b98b1e3),
	.w6(32'h3896561c),
	.w7(32'hbbb009b0),
	.w8(32'hbcc2b720),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27d586),
	.w1(32'h3a6bd5d5),
	.w2(32'h3b0bdaba),
	.w3(32'h3bfaa338),
	.w4(32'hbb9a0d64),
	.w5(32'hbb9634c7),
	.w6(32'hba609a40),
	.w7(32'hbbac4d6b),
	.w8(32'hbbb1f633),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d9828),
	.w1(32'h3c062369),
	.w2(32'h3c90a82a),
	.w3(32'h3bc0fe95),
	.w4(32'h3c54ed5e),
	.w5(32'hba84a3ab),
	.w6(32'h3b6b56df),
	.w7(32'h3bae12bf),
	.w8(32'h3c02df4d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01273e),
	.w1(32'h3ae689c2),
	.w2(32'h3b97e349),
	.w3(32'hbb071b90),
	.w4(32'hbc007674),
	.w5(32'hbb81d295),
	.w6(32'h3c91e477),
	.w7(32'hbc833bc5),
	.w8(32'hbc62f0e0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e039e),
	.w1(32'h3cde2b7d),
	.w2(32'h3ca27d5b),
	.w3(32'h3bb3609d),
	.w4(32'hbbde4ad0),
	.w5(32'h3af93b56),
	.w6(32'hbbff4474),
	.w7(32'hbc14ff5f),
	.w8(32'hbccfd76e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baea2d6),
	.w1(32'hbc78c2f2),
	.w2(32'h39a6324f),
	.w3(32'h3c6ec75c),
	.w4(32'hbc8c9a38),
	.w5(32'hbcd21220),
	.w6(32'hbcc4d0f2),
	.w7(32'h3cdc0f25),
	.w8(32'hbc14ac75),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c175c39),
	.w1(32'hbb9529bc),
	.w2(32'hbc26d987),
	.w3(32'hbc15a30e),
	.w4(32'h3b307049),
	.w5(32'hbc13e7de),
	.w6(32'hbcdb6417),
	.w7(32'hbbe42e15),
	.w8(32'h3a3b6bc8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c2763),
	.w1(32'hbb88a858),
	.w2(32'hba6bc100),
	.w3(32'hbbfacc51),
	.w4(32'hb9674ebc),
	.w5(32'h3a1b73d5),
	.w6(32'h3c466a7f),
	.w7(32'h3c23fa45),
	.w8(32'h3beb651c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa29ba),
	.w1(32'hbb3e3f97),
	.w2(32'hb94774db),
	.w3(32'h3c03906f),
	.w4(32'h3c1a652d),
	.w5(32'h3b8171ed),
	.w6(32'h3a5ae9c2),
	.w7(32'h3c1af564),
	.w8(32'h3c145fb1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc0d1e),
	.w1(32'h3a932885),
	.w2(32'h3bce1b9f),
	.w3(32'h3a6d7a91),
	.w4(32'hbc71401f),
	.w5(32'hbcdf80e3),
	.w6(32'h3c319f20),
	.w7(32'hbceaac6f),
	.w8(32'hbd2a05a2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fc202),
	.w1(32'hba0ca8d8),
	.w2(32'h39eca563),
	.w3(32'hbc5e600f),
	.w4(32'h3b216016),
	.w5(32'h3a5b9431),
	.w6(32'hbd04d1d9),
	.w7(32'h3ac0370c),
	.w8(32'h3b375975),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c060451),
	.w1(32'h3a8d10d9),
	.w2(32'h3a800a0c),
	.w3(32'h3bba7292),
	.w4(32'hbc44fd7c),
	.w5(32'h399667cc),
	.w6(32'h3c070878),
	.w7(32'hbd00598e),
	.w8(32'hbd5df425),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bc9d7),
	.w1(32'h3963cffc),
	.w2(32'hba4206ea),
	.w3(32'h3c5c8d54),
	.w4(32'hba4b75b1),
	.w5(32'hbc225ac6),
	.w6(32'hbcdab1c4),
	.w7(32'h3b8507a3),
	.w8(32'hbb5cdec7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25174c),
	.w1(32'hbae39033),
	.w2(32'hbbd858ee),
	.w3(32'h3c8180ff),
	.w4(32'h3b9403b8),
	.w5(32'hbc48bbf3),
	.w6(32'h3b69aa7d),
	.w7(32'hbb8f9ecf),
	.w8(32'hbb9e7eea),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17f4e6),
	.w1(32'hbaf0d9af),
	.w2(32'hbc2b8234),
	.w3(32'h3b96ab73),
	.w4(32'hbc860b90),
	.w5(32'hbd32a207),
	.w6(32'h3c1f8e1c),
	.w7(32'h390a4ef1),
	.w8(32'hbc319e45),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac15192),
	.w1(32'hbc7ea275),
	.w2(32'hbc2258d2),
	.w3(32'hbd5b4eb9),
	.w4(32'h3c4376fe),
	.w5(32'hbc952a7a),
	.w6(32'hbc045b74),
	.w7(32'h3cf58a31),
	.w8(32'h3d0d148a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cd9bb),
	.w1(32'hbac53751),
	.w2(32'hbb5ee128),
	.w3(32'hbc880fb0),
	.w4(32'h3b722744),
	.w5(32'hba6c9b30),
	.w6(32'hbb86ea59),
	.w7(32'h3c1d7dff),
	.w8(32'h3b4e55ba),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb724787),
	.w1(32'h3c6d6862),
	.w2(32'h3c9366ce),
	.w3(32'hbb5fcc25),
	.w4(32'h3ab46b29),
	.w5(32'hbc5fa970),
	.w6(32'hbb890ffa),
	.w7(32'hbb8a5118),
	.w8(32'hbcd1d815),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b92d8),
	.w1(32'hba5921aa),
	.w2(32'hbb4d239d),
	.w3(32'h3bf38603),
	.w4(32'h3bb69d27),
	.w5(32'hbbbc0644),
	.w6(32'hbc8ed142),
	.w7(32'h3cb806ad),
	.w8(32'h3bf4fe4a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba7b71),
	.w1(32'h3b2d9138),
	.w2(32'hba8db2b2),
	.w3(32'hbaf22de9),
	.w4(32'h39978307),
	.w5(32'hbb806b34),
	.w6(32'hbbdb0cab),
	.w7(32'hbb4bf1c1),
	.w8(32'hbc18f432),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7f97e),
	.w1(32'hbc2673a6),
	.w2(32'hbc4890e5),
	.w3(32'h3bb89409),
	.w4(32'h3c9e8e6f),
	.w5(32'h3a2b5b6a),
	.w6(32'hba8e8d8f),
	.w7(32'hb90f56a0),
	.w8(32'h3cd6c31f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6847a),
	.w1(32'h3c1848a6),
	.w2(32'h3c895e38),
	.w3(32'hbc690707),
	.w4(32'hba446bdf),
	.w5(32'h3c4e0682),
	.w6(32'h3cfba172),
	.w7(32'h3c69f42c),
	.w8(32'h3bb611a4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c998cdf),
	.w1(32'h3a6324b1),
	.w2(32'hbb1ed30f),
	.w3(32'h3c971e8c),
	.w4(32'hb9d786f0),
	.w5(32'hbb840afc),
	.w6(32'h3b96cb52),
	.w7(32'h3b3b4491),
	.w8(32'h3a74319b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab13ab5),
	.w1(32'h3ca1f516),
	.w2(32'h3c91fed0),
	.w3(32'hb887e305),
	.w4(32'hbb9460a7),
	.w5(32'hbc3c6100),
	.w6(32'h3bb20824),
	.w7(32'h3c1aa7e4),
	.w8(32'hba355ab7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b7aaf),
	.w1(32'hbbaf3831),
	.w2(32'hbbd41470),
	.w3(32'hba9a7d4a),
	.w4(32'h3a6f7482),
	.w5(32'hbbcf006f),
	.w6(32'hbc1ca448),
	.w7(32'h3ac233c0),
	.w8(32'hbabe228d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c056caf),
	.w1(32'h3ba8483a),
	.w2(32'h3ab36cfd),
	.w3(32'h3c051a80),
	.w4(32'h3bb2d15d),
	.w5(32'hb9e6c60d),
	.w6(32'h3c1d6a42),
	.w7(32'h3b20e96e),
	.w8(32'hbab6e1eb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b5bab),
	.w1(32'h3bb029a4),
	.w2(32'h3a67950c),
	.w3(32'hbb056ec3),
	.w4(32'h3c765a6b),
	.w5(32'hbba8feff),
	.w6(32'hba3c1b78),
	.w7(32'h3c63de66),
	.w8(32'h3c74d130),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a6665),
	.w1(32'h3a3cd71f),
	.w2(32'hb972ab4f),
	.w3(32'hbb929437),
	.w4(32'hbadde743),
	.w5(32'hbb4bba17),
	.w6(32'hbbaf4bd3),
	.w7(32'h3b598a05),
	.w8(32'h3a8186fa),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b148a),
	.w1(32'hbc46e992),
	.w2(32'hbb18592f),
	.w3(32'hbb3a7174),
	.w4(32'hbc2f361d),
	.w5(32'hbc830b1b),
	.w6(32'h3b233f82),
	.w7(32'hbb48ec1d),
	.w8(32'hbc5ca705),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb234ee3),
	.w1(32'h3b975ccb),
	.w2(32'h3c93871e),
	.w3(32'hbc133be2),
	.w4(32'h3c478d66),
	.w5(32'h3c491ae1),
	.w6(32'hbcabd647),
	.w7(32'hbc868c5a),
	.w8(32'hbd234cf4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c746301),
	.w1(32'h3af851c0),
	.w2(32'h3b1bbe83),
	.w3(32'h3cd78360),
	.w4(32'h3b00236e),
	.w5(32'h3c2e1679),
	.w6(32'hbcda0551),
	.w7(32'h3c8d64cb),
	.w8(32'h3c8e98ae),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15d2cc),
	.w1(32'hbcc0a83a),
	.w2(32'hbc8cd750),
	.w3(32'h3b282068),
	.w4(32'hbc6557aa),
	.w5(32'hbd13d9ee),
	.w6(32'h3cf90920),
	.w7(32'h3d13ea5f),
	.w8(32'h3d1439ab),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabce43a),
	.w1(32'h3a96736c),
	.w2(32'h3a0c91da),
	.w3(32'hbd0514c0),
	.w4(32'h3b4e0415),
	.w5(32'h3b3a50fa),
	.w6(32'h3ce02640),
	.w7(32'hbb29de43),
	.w8(32'hbb88907a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb801e60e),
	.w1(32'hbbb37a29),
	.w2(32'hbaa43c84),
	.w3(32'hbae32526),
	.w4(32'h3c1e16ee),
	.w5(32'h3ba052e2),
	.w6(32'hbc2e7ebf),
	.w7(32'h3c0ffec5),
	.w8(32'h3c2bcc44),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84cf04),
	.w1(32'hbb6c3c7d),
	.w2(32'hbc1786f7),
	.w3(32'h3bc0360f),
	.w4(32'h3a5a41ef),
	.w5(32'hbbb77d33),
	.w6(32'h3c670a19),
	.w7(32'hbb9af2ee),
	.w8(32'hbaf4a015),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1601a),
	.w1(32'h3a0918a8),
	.w2(32'hbab83658),
	.w3(32'h3ae0a9ad),
	.w4(32'hbace4eef),
	.w5(32'hbb949c5b),
	.w6(32'h3aefdd10),
	.w7(32'hbb5b3984),
	.w8(32'hbb93169a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b164be3),
	.w1(32'hbcc58dc1),
	.w2(32'hbcfea3de),
	.w3(32'h3a830c12),
	.w4(32'h3c8a181f),
	.w5(32'hbc45aeb8),
	.w6(32'h3b8a4577),
	.w7(32'h3d061f25),
	.w8(32'h3d36ee46),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86374e),
	.w1(32'hbb92f350),
	.w2(32'h3b2e3693),
	.w3(32'hbd08b561),
	.w4(32'hbbd61acd),
	.w5(32'hbca0fd2e),
	.w6(32'h3d164b80),
	.w7(32'h3a138fac),
	.w8(32'hbb29eb51),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5892d1),
	.w1(32'h3c727fe0),
	.w2(32'hbc0e56a7),
	.w3(32'h3a250817),
	.w4(32'hbc37f65e),
	.w5(32'h3c0e43de),
	.w6(32'h3c618f1e),
	.w7(32'hbd01e59a),
	.w8(32'hbd036ec1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7728f3),
	.w1(32'h3c562900),
	.w2(32'h3c4a3655),
	.w3(32'h3d072900),
	.w4(32'hbca065b3),
	.w5(32'hbc83428c),
	.w6(32'hbc1306fa),
	.w7(32'hbc4376a6),
	.w8(32'hbccbfe2f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac431f6),
	.w1(32'hba9c1ac0),
	.w2(32'hbc5b6944),
	.w3(32'h391bec56),
	.w4(32'h3bce832f),
	.w5(32'h3b9af111),
	.w6(32'hbcc78bfb),
	.w7(32'h3caea75f),
	.w8(32'h3c037594),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f2090),
	.w1(32'h3bb87304),
	.w2(32'h3c09e95a),
	.w3(32'hbc22cee5),
	.w4(32'h3aeae928),
	.w5(32'h3bc8114a),
	.w6(32'hbc0381de),
	.w7(32'h3c161281),
	.w8(32'h3bf44ee5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba057f43),
	.w1(32'h3bd6bc41),
	.w2(32'h3b952523),
	.w3(32'hbabd9f37),
	.w4(32'h3b0b9612),
	.w5(32'h3c2de6a9),
	.w6(32'hbb30d49f),
	.w7(32'hbbd035ad),
	.w8(32'hbc01b0e4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36c782),
	.w1(32'h3ade7c3a),
	.w2(32'hbadf47f4),
	.w3(32'h3c597ed2),
	.w4(32'h3a893417),
	.w5(32'h3ba6ce05),
	.w6(32'h3a56f022),
	.w7(32'hba3f8fd3),
	.w8(32'hbbf3c600),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f2aef),
	.w1(32'h3b519e42),
	.w2(32'h3aee114a),
	.w3(32'h3c16a53e),
	.w4(32'h3b1f05e1),
	.w5(32'h3aa3ce63),
	.w6(32'h3b12393b),
	.w7(32'h374a3701),
	.w8(32'h3ada8618),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada94c0),
	.w1(32'hbc1ea0a4),
	.w2(32'h3b9286d5),
	.w3(32'hb871ae51),
	.w4(32'hbb8ac5fa),
	.w5(32'hbc3ac883),
	.w6(32'h39c220a7),
	.w7(32'h3b608f2c),
	.w8(32'hbbfa1fb8),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d07ea),
	.w1(32'h3c1dd221),
	.w2(32'h3bb4f63a),
	.w3(32'hbbe988bf),
	.w4(32'hbce3a552),
	.w5(32'h3a6a8016),
	.w6(32'hbab45181),
	.w7(32'h3cd8d196),
	.w8(32'h3c370471),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36e599),
	.w1(32'h3c019ace),
	.w2(32'h3cb56683),
	.w3(32'h3c90436b),
	.w4(32'hbc3827c5),
	.w5(32'hbcf40b9a),
	.w6(32'hbcd7ded8),
	.w7(32'hbbed02b8),
	.w8(32'hbc8fd71f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd20dc9),
	.w1(32'hb9ed1f35),
	.w2(32'hba79d5d2),
	.w3(32'hbc0cf39f),
	.w4(32'h39c25ca2),
	.w5(32'hba83b024),
	.w6(32'hbc8e14cb),
	.w7(32'hbae95d63),
	.w8(32'h39b44432),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8039f5),
	.w1(32'h3b141650),
	.w2(32'h3b9e0463),
	.w3(32'h395d9250),
	.w4(32'hbbd98cf5),
	.w5(32'h3b03c3fc),
	.w6(32'h3ba220a4),
	.w7(32'hbb1208b0),
	.w8(32'hbc470485),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dc5ea),
	.w1(32'hbba76469),
	.w2(32'hbc02608b),
	.w3(32'h3b10e8cb),
	.w4(32'hbc24e30a),
	.w5(32'hbc1d5d08),
	.w6(32'hbc078e63),
	.w7(32'hbc26729c),
	.w8(32'hbc3aaa46),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7015b3),
	.w1(32'hbae64608),
	.w2(32'h3ab5cc68),
	.w3(32'hbaa9b4bf),
	.w4(32'hbb077c74),
	.w5(32'hba8cb3d3),
	.w6(32'hbbcde6a9),
	.w7(32'h3a2cbea2),
	.w8(32'h3a364e53),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6540a),
	.w1(32'h3c8f666b),
	.w2(32'h3d1d07c7),
	.w3(32'h3b8034ea),
	.w4(32'hbcad6478),
	.w5(32'hbbca1731),
	.w6(32'h3b8af6cd),
	.w7(32'hbd34d90b),
	.w8(32'hbd8b228e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c989f02),
	.w1(32'h3b4edc62),
	.w2(32'h3b3a9cdf),
	.w3(32'h3cb403f9),
	.w4(32'hbab08e7e),
	.w5(32'hbbb9bd51),
	.w6(32'hbc8d86e0),
	.w7(32'h3b9245c9),
	.w8(32'h3bc3fe48),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7ed14),
	.w1(32'h3c839fbc),
	.w2(32'h3c1e7b68),
	.w3(32'hbb669d13),
	.w4(32'hba8184b9),
	.w5(32'hbbc22a72),
	.w6(32'h3ca85978),
	.w7(32'hbc694d7c),
	.w8(32'hbcbcdf38),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8949db),
	.w1(32'h3beda018),
	.w2(32'h3c309ac7),
	.w3(32'h3c8f26d0),
	.w4(32'h3b9ba444),
	.w5(32'h3bc1c8cc),
	.w6(32'hbcb47c94),
	.w7(32'h3b7e323c),
	.w8(32'h3b521b42),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c415f88),
	.w1(32'hbbb9ea76),
	.w2(32'h3b5235b8),
	.w3(32'h3bc2135c),
	.w4(32'h3c7af040),
	.w5(32'h3c7bc52b),
	.w6(32'h3b6f01cb),
	.w7(32'hbd11b19d),
	.w8(32'h3abf3cde),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule