module layer_10_featuremap_146(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3854154b),
	.w1(32'h39e8edaa),
	.w2(32'h3aba0274),
	.w3(32'h38a833f8),
	.w4(32'hb637e885),
	.w5(32'h3a65b251),
	.w6(32'h3a02bd15),
	.w7(32'h3a513280),
	.w8(32'h399c1f40),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5055a),
	.w1(32'hba0c5b62),
	.w2(32'hb936a206),
	.w3(32'h39c315bb),
	.w4(32'hb9ea7da7),
	.w5(32'hb9374dbd),
	.w6(32'hb9d7d054),
	.w7(32'hb9375776),
	.w8(32'hb93f2b5b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af1b56),
	.w1(32'hb9be5385),
	.w2(32'hb928b02d),
	.w3(32'hb9555144),
	.w4(32'hb9aa0811),
	.w5(32'hb9b62afe),
	.w6(32'hb98fdcdd),
	.w7(32'hb98f939e),
	.w8(32'hb9a59f2e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96dff5c),
	.w1(32'hba016867),
	.w2(32'hba7f0b79),
	.w3(32'hb9c5d806),
	.w4(32'h39dd6c34),
	.w5(32'hb89c6ac3),
	.w6(32'hb9b31a1b),
	.w7(32'hba3b9673),
	.w8(32'hb9e768fe),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387c6f51),
	.w1(32'h379dad0c),
	.w2(32'h3a04958e),
	.w3(32'hb9001da9),
	.w4(32'h39ad477f),
	.w5(32'h39f10f79),
	.w6(32'h37d1eaa8),
	.w7(32'h38fe084b),
	.w8(32'h39a18149),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39065fe1),
	.w1(32'h395fbdbb),
	.w2(32'h3971ff71),
	.w3(32'h39dd6f05),
	.w4(32'h39979cbd),
	.w5(32'h38c4598a),
	.w6(32'h39172ff2),
	.w7(32'h391f6a25),
	.w8(32'h3973ccb3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b2720),
	.w1(32'hba770907),
	.w2(32'hb9c9b1a0),
	.w3(32'h39a64b6b),
	.w4(32'hba269140),
	.w5(32'hb9d4e087),
	.w6(32'hba30b70d),
	.w7(32'hb9b6db83),
	.w8(32'hb9aa1120),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfc6e9),
	.w1(32'h3a4ede9e),
	.w2(32'h3a2ba970),
	.w3(32'hb958c9de),
	.w4(32'h3a6165fb),
	.w5(32'h39d154de),
	.w6(32'h39d82323),
	.w7(32'h3a1ecd49),
	.w8(32'h3a2a0cbe),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8d65f),
	.w1(32'h35c09477),
	.w2(32'hb8f58f51),
	.w3(32'h398d4068),
	.w4(32'hb7dfa7ac),
	.w5(32'hb979a947),
	.w6(32'hb67ff3f6),
	.w7(32'hb9b5d781),
	.w8(32'hb92eb06a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383f45ae),
	.w1(32'hb90c71e8),
	.w2(32'hb8a8c464),
	.w3(32'h39020a9f),
	.w4(32'hb8d5c78c),
	.w5(32'hb815b5bd),
	.w6(32'hb8dfa790),
	.w7(32'hb730bc9d),
	.w8(32'hb847fcb6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5cb2e),
	.w1(32'h3a202fd2),
	.w2(32'h39a715a1),
	.w3(32'hb992a1b9),
	.w4(32'h39bcf108),
	.w5(32'h39f0f81e),
	.w6(32'h39f50a84),
	.w7(32'h39a814b0),
	.w8(32'h3998c532),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f86954),
	.w1(32'h3925cba4),
	.w2(32'hb9e063c1),
	.w3(32'h39c84721),
	.w4(32'h3a2d130b),
	.w5(32'h39af1007),
	.w6(32'h3947a9a7),
	.w7(32'h389871ef),
	.w8(32'h39d3973a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a828ad6),
	.w1(32'h3a0a9443),
	.w2(32'h3a1b4a4c),
	.w3(32'h3a42f780),
	.w4(32'h3a0af952),
	.w5(32'h3a166f4e),
	.w6(32'hb85b0005),
	.w7(32'h3930e122),
	.w8(32'h390c682b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391ebb05),
	.w1(32'h3a81fdc6),
	.w2(32'h3a28248b),
	.w3(32'h38a2503e),
	.w4(32'h3a3b7225),
	.w5(32'h39b3708e),
	.w6(32'h3a5f5895),
	.w7(32'h39d1ba76),
	.w8(32'h3a3a6c8a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a251447),
	.w1(32'h3a540a77),
	.w2(32'h3a7b1740),
	.w3(32'h39a95432),
	.w4(32'h3ad2ab36),
	.w5(32'h3aad7470),
	.w6(32'h3988ae35),
	.w7(32'h39d65e4e),
	.w8(32'h39b0a5fc),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c030b),
	.w1(32'h399adc3c),
	.w2(32'h39f0e863),
	.w3(32'h3a4b4901),
	.w4(32'h39636c05),
	.w5(32'h3989e0d6),
	.w6(32'h38482e25),
	.w7(32'h382de371),
	.w8(32'h38a2cc68),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88e369f),
	.w1(32'hb81ffa41),
	.w2(32'h3854b77c),
	.w3(32'h38dc1426),
	.w4(32'hb80b9198),
	.w5(32'hb9e21625),
	.w6(32'hb8616248),
	.w7(32'hb97f9b4e),
	.w8(32'h388588c9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8de6432),
	.w1(32'hba3b55dc),
	.w2(32'hb9495621),
	.w3(32'hb962f686),
	.w4(32'hba041ed9),
	.w5(32'hb99350c3),
	.w6(32'hba459679),
	.w7(32'hba12fa98),
	.w8(32'hba16e262),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fc2a9),
	.w1(32'hb9c098a5),
	.w2(32'hb9320157),
	.w3(32'hba3e0d70),
	.w4(32'hb9a9d019),
	.w5(32'hb95f661e),
	.w6(32'hba0ce0e1),
	.w7(32'hb9a9b621),
	.w8(32'hb9a5f551),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe0c79),
	.w1(32'h3975afc3),
	.w2(32'h392cc34b),
	.w3(32'hb9b7ddca),
	.w4(32'h3929a0d6),
	.w5(32'h368048b4),
	.w6(32'h390f8ced),
	.w7(32'hb83b9c69),
	.w8(32'h38565b80),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb773c880),
	.w1(32'h38b40ae5),
	.w2(32'h38f46fb3),
	.w3(32'h38fb0d57),
	.w4(32'h372fb5cb),
	.w5(32'hb8fd5dad),
	.w6(32'hb93ccc70),
	.w7(32'hb9427fc9),
	.w8(32'hb90a284c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35afb70b),
	.w1(32'h398d3312),
	.w2(32'h386020a6),
	.w3(32'hb8fc9d97),
	.w4(32'h39c9c5e9),
	.w5(32'h39ccae85),
	.w6(32'h3a349dd2),
	.w7(32'h3a41c789),
	.w8(32'h3a23fe0b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390bd540),
	.w1(32'h3934435f),
	.w2(32'h39a1012c),
	.w3(32'hb9a30c11),
	.w4(32'hb803c384),
	.w5(32'hb8724772),
	.w6(32'h38b4a1c0),
	.w7(32'h3909444c),
	.w8(32'h39e403a7),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ddb09),
	.w1(32'h3a0b645d),
	.w2(32'h3a0a788d),
	.w3(32'h39dc1985),
	.w4(32'h39c99ebe),
	.w5(32'h39bf0a28),
	.w6(32'h391044a4),
	.w7(32'h36741df6),
	.w8(32'h39afad45),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b8ca5),
	.w1(32'hb94ccc9e),
	.w2(32'h37fc3440),
	.w3(32'h38851cb6),
	.w4(32'h392c891d),
	.w5(32'h39a9dcd8),
	.w6(32'hb9ebf85f),
	.w7(32'hb97e69fe),
	.w8(32'hb93eb5c7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91fb363),
	.w1(32'h39f59219),
	.w2(32'h390e064c),
	.w3(32'h38cb8221),
	.w4(32'h3a2a7b9b),
	.w5(32'h394ebca1),
	.w6(32'h3a1fba21),
	.w7(32'h3a0f687e),
	.w8(32'h3a15a796),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39891ad8),
	.w1(32'h39cf2375),
	.w2(32'h3999ed85),
	.w3(32'h39776d4b),
	.w4(32'h39add286),
	.w5(32'h3917ad35),
	.w6(32'h3986a8ca),
	.w7(32'h3901b502),
	.w8(32'h39213e71),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fa71e),
	.w1(32'h3a175a5d),
	.w2(32'h3960e472),
	.w3(32'hb9a69469),
	.w4(32'h3a606b6f),
	.w5(32'h3a48cbab),
	.w6(32'hba161ba8),
	.w7(32'h3a08e51f),
	.w8(32'hb888bb0f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c6a47),
	.w1(32'h392ec79b),
	.w2(32'hba0e8707),
	.w3(32'h3972a008),
	.w4(32'h389c298c),
	.w5(32'hba2a2a8e),
	.w6(32'h399fb517),
	.w7(32'hba3579f2),
	.w8(32'hb98773db),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a4b69),
	.w1(32'hb973a1bd),
	.w2(32'hb83b62b1),
	.w3(32'hb9ddda4a),
	.w4(32'hb9d2b6f9),
	.w5(32'hb939d9c6),
	.w6(32'hba1bf50a),
	.w7(32'hba00f32c),
	.w8(32'hba315401),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1dde7d),
	.w1(32'h395a7433),
	.w2(32'h39403f37),
	.w3(32'hba54310d),
	.w4(32'h3933bf64),
	.w5(32'h37d21551),
	.w6(32'hb627dc75),
	.w7(32'hb7d74a57),
	.w8(32'h38836ea8),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39529c58),
	.w1(32'h3951cacb),
	.w2(32'h3967f3aa),
	.w3(32'h3827715d),
	.w4(32'h39254d5a),
	.w5(32'h38263feb),
	.w6(32'h38819c86),
	.w7(32'h38a431e8),
	.w8(32'h38909b69),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396fe306),
	.w1(32'h39afc524),
	.w2(32'h3a914003),
	.w3(32'h388e7a06),
	.w4(32'h39d74ff5),
	.w5(32'h3a519241),
	.w6(32'h3a03a8ec),
	.w7(32'h399272df),
	.w8(32'h39a535d2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37996095),
	.w1(32'hb95ff4f0),
	.w2(32'h39cce104),
	.w3(32'h397d9079),
	.w4(32'hb9f47041),
	.w5(32'h3895e1e0),
	.w6(32'hb987bbf9),
	.w7(32'hb90af962),
	.w8(32'hb93ee46e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91889c6),
	.w1(32'hba6ac07a),
	.w2(32'hba3095f3),
	.w3(32'h3965f5ef),
	.w4(32'hba4a7b5c),
	.w5(32'hba249858),
	.w6(32'hba5327f0),
	.w7(32'hb9fa3e95),
	.w8(32'hba11b6e0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d0475),
	.w1(32'h39d0fff4),
	.w2(32'h3a0500a1),
	.w3(32'hb9f5c759),
	.w4(32'h3a1cf3e1),
	.w5(32'h39c75afe),
	.w6(32'h3808c2eb),
	.w7(32'h39255045),
	.w8(32'h3981845b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7335b4),
	.w1(32'hba1ad1af),
	.w2(32'h39a8cb5f),
	.w3(32'h39e3ba61),
	.w4(32'hb98b4fd9),
	.w5(32'h38b08e20),
	.w6(32'hb9031cfe),
	.w7(32'hb98ee01e),
	.w8(32'h38ae481f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bd755),
	.w1(32'hba449855),
	.w2(32'hb99195c4),
	.w3(32'hba65d680),
	.w4(32'hba62745f),
	.w5(32'hba1ce89e),
	.w6(32'hba9558e8),
	.w7(32'hb9f6ba04),
	.w8(32'hba0f50b5),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ba81b),
	.w1(32'h3987aa86),
	.w2(32'hb9aa0c49),
	.w3(32'hbaae498c),
	.w4(32'h39088814),
	.w5(32'hb97290e0),
	.w6(32'hb9ea684c),
	.w7(32'h381a2c91),
	.w8(32'hb932d64f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b96caf),
	.w1(32'hba0e2446),
	.w2(32'hb99681b1),
	.w3(32'hb82566df),
	.w4(32'hb9fcdc0a),
	.w5(32'hb9b192b1),
	.w6(32'hb9d94a26),
	.w7(32'hb991474f),
	.w8(32'hb9738c0f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8ea58),
	.w1(32'hb9a1f5e6),
	.w2(32'h3903cd7d),
	.w3(32'hb939427c),
	.w4(32'hba02d8ab),
	.w5(32'hb980e105),
	.w6(32'hb95460f9),
	.w7(32'hb9961bd3),
	.w8(32'hba51ef69),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba010319),
	.w1(32'hb7cfbc8b),
	.w2(32'hb91326c0),
	.w3(32'hba49a644),
	.w4(32'h3947b4ff),
	.w5(32'h38beda4c),
	.w6(32'hb89b98cf),
	.w7(32'h393053d7),
	.w8(32'hb89bc166),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ccbec1),
	.w1(32'hb7a27e42),
	.w2(32'h391b0b82),
	.w3(32'h3903c7dd),
	.w4(32'hb9187476),
	.w5(32'hb8288690),
	.w6(32'hb89754e2),
	.w7(32'hb820a1c8),
	.w8(32'h38855523),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39768cdb),
	.w1(32'h38a38b4e),
	.w2(32'h3790182e),
	.w3(32'h399124aa),
	.w4(32'h383b0fd0),
	.w5(32'hb745fce4),
	.w6(32'h397f16e0),
	.w7(32'h3716c9c4),
	.w8(32'h382cb074),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2aa71),
	.w1(32'h39ccadca),
	.w2(32'h3a0c6380),
	.w3(32'hba1516f5),
	.w4(32'hb933fd93),
	.w5(32'h38fc6f7c),
	.w6(32'h394406b0),
	.w7(32'hb8558255),
	.w8(32'hb8d56cff),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fef4e7),
	.w1(32'hb89795b8),
	.w2(32'hb917902f),
	.w3(32'hb9df3777),
	.w4(32'hb9398f3d),
	.w5(32'hb940ada0),
	.w6(32'hb9c175a4),
	.w7(32'hb9781964),
	.w8(32'hb95f42ff),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb3d2a),
	.w1(32'h38cad5a0),
	.w2(32'hba5e4286),
	.w3(32'hba4539a7),
	.w4(32'h3aa7ab18),
	.w5(32'h3a39b27b),
	.w6(32'hb524d000),
	.w7(32'hb9b0b224),
	.w8(32'hb6db5c7c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efb6c3),
	.w1(32'h398863cd),
	.w2(32'h389afada),
	.w3(32'h3a1586b9),
	.w4(32'h39c4b070),
	.w5(32'hb90cb311),
	.w6(32'h39860d9a),
	.w7(32'hb9fc7408),
	.w8(32'h3891310e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8087d1d),
	.w1(32'h3960334d),
	.w2(32'h39a5211d),
	.w3(32'hb8ebb3a8),
	.w4(32'h391d1902),
	.w5(32'h38ab2d10),
	.w6(32'h392e091b),
	.w7(32'h391469a4),
	.w8(32'h3963cc0d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3970778d),
	.w1(32'h39f4aee8),
	.w2(32'h399a6a2f),
	.w3(32'h39088db1),
	.w4(32'h39c9b41e),
	.w5(32'h396d2999),
	.w6(32'h39c7a902),
	.w7(32'h3938973d),
	.w8(32'h39a667b5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c23923),
	.w1(32'hb923f21f),
	.w2(32'hb9789c53),
	.w3(32'h399a9b93),
	.w4(32'hb8cbac7a),
	.w5(32'hb989924a),
	.w6(32'hb780a233),
	.w7(32'h37c823b6),
	.w8(32'hb91575bb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a50eed),
	.w1(32'h3a428552),
	.w2(32'h36f0a218),
	.w3(32'hb947d3a1),
	.w4(32'h3a590bca),
	.w5(32'h3aae54d1),
	.w6(32'h3a3a3490),
	.w7(32'h3a3ba361),
	.w8(32'h3a35a694),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389d56f4),
	.w1(32'h39808c0c),
	.w2(32'h39c3fac6),
	.w3(32'h3a623405),
	.w4(32'h3a0e387c),
	.w5(32'h39c4550e),
	.w6(32'h3926df52),
	.w7(32'h38ace5d7),
	.w8(32'h38c51be8),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c29204),
	.w1(32'h379e2987),
	.w2(32'h39c44b5e),
	.w3(32'h39cc2326),
	.w4(32'h3a197e20),
	.w5(32'h3a3b0ce8),
	.w6(32'hb976cee1),
	.w7(32'hb99e9afe),
	.w8(32'h39e0b551),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374afc7b),
	.w1(32'hb957af43),
	.w2(32'hb8d7b5fd),
	.w3(32'h39c0ad14),
	.w4(32'hb745d21f),
	.w5(32'hb89b61ec),
	.w6(32'hb985964f),
	.w7(32'hb92ea62e),
	.w8(32'h389b7e86),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8496426),
	.w1(32'h3985c10c),
	.w2(32'h39a164ff),
	.w3(32'hb910cd6f),
	.w4(32'h398c92ff),
	.w5(32'h38cabb27),
	.w6(32'h397e5d3a),
	.w7(32'hb90b9278),
	.w8(32'hb9813c83),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3887cb6b),
	.w1(32'h393c0a5e),
	.w2(32'h39cb9719),
	.w3(32'hb9288c45),
	.w4(32'h3941527e),
	.w5(32'h393a6459),
	.w6(32'h394cc1df),
	.w7(32'h398dec97),
	.w8(32'h388c3b91),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38368177),
	.w1(32'h397d5dd0),
	.w2(32'h3a32b6ee),
	.w3(32'hb92bbe5b),
	.w4(32'h39a790c7),
	.w5(32'h3a1efe1f),
	.w6(32'h39470eb2),
	.w7(32'h3a00c8e6),
	.w8(32'h3a1d0d6f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f710ea),
	.w1(32'hba4549bb),
	.w2(32'hb9f58aff),
	.w3(32'h39ebe7c2),
	.w4(32'hba305057),
	.w5(32'hb9d2de32),
	.w6(32'hba193ee2),
	.w7(32'hb9a337c8),
	.w8(32'hb9f90aab),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9df78),
	.w1(32'h39038ac9),
	.w2(32'hb787e8fd),
	.w3(32'hb9c50b05),
	.w4(32'h39096083),
	.w5(32'hb882f350),
	.w6(32'h39100036),
	.w7(32'hb85aaa9a),
	.w8(32'h3840b0db),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f11fa2),
	.w1(32'hb9fc84c2),
	.w2(32'hb99aa475),
	.w3(32'h3910b030),
	.w4(32'hb9e82282),
	.w5(32'hb98813f4),
	.w6(32'hb9f4ae82),
	.w7(32'hb999887c),
	.w8(32'hb930d923),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebd611),
	.w1(32'h3a498327),
	.w2(32'h3a013019),
	.w3(32'hb97fadff),
	.w4(32'h39b2a9b9),
	.w5(32'h399962f2),
	.w6(32'h39c5a5ea),
	.w7(32'h391f1283),
	.w8(32'h39cd3934),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991d716),
	.w1(32'h3969d3db),
	.w2(32'h3ac8eee0),
	.w3(32'h39088a2d),
	.w4(32'hba16e5e2),
	.w5(32'h3a14f64d),
	.w6(32'h3a43a9c0),
	.w7(32'h397cb93e),
	.w8(32'h379b277e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ecc07a),
	.w1(32'hb99d59ae),
	.w2(32'hb9ce3f12),
	.w3(32'h398e274a),
	.w4(32'hb95ce35b),
	.w5(32'hb99d7601),
	.w6(32'h382f7425),
	.w7(32'hb87168c2),
	.w8(32'hb8da70c9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c45f1),
	.w1(32'hb98b0fc9),
	.w2(32'hb9852135),
	.w3(32'hb98ef72d),
	.w4(32'hb9ac4841),
	.w5(32'hb9371cce),
	.w6(32'hb8242506),
	.w7(32'hb8b901aa),
	.w8(32'hb89f23cc),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9113687),
	.w1(32'h391070ec),
	.w2(32'h3951945f),
	.w3(32'hb946dd27),
	.w4(32'h38b4ba24),
	.w5(32'h39c8ecb1),
	.w6(32'h3917ddf3),
	.w7(32'h391fbf5b),
	.w8(32'h39092ef3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39971a99),
	.w1(32'hb960b179),
	.w2(32'h3985274c),
	.w3(32'h399042f5),
	.w4(32'hb99ef494),
	.w5(32'h38c2efaa),
	.w6(32'h39a00af4),
	.w7(32'h38ae9a4c),
	.w8(32'hb9a26b79),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d31c7f),
	.w1(32'hb74e4460),
	.w2(32'h39597c25),
	.w3(32'hb9da677c),
	.w4(32'h381acf2d),
	.w5(32'h38be2c9c),
	.w6(32'hb9829440),
	.w7(32'hb9956ebe),
	.w8(32'hb91ac427),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8006f05),
	.w1(32'hb7bae222),
	.w2(32'h39db3644),
	.w3(32'hb9446640),
	.w4(32'h391c0140),
	.w5(32'h3994806c),
	.w6(32'hb995dcc4),
	.w7(32'hb99ea114),
	.w8(32'hb91a644d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba009c48),
	.w1(32'h37ce6c2d),
	.w2(32'h3a0e2c53),
	.w3(32'hba03e496),
	.w4(32'hb800619e),
	.w5(32'h39c021c4),
	.w6(32'hb9ee439a),
	.w7(32'h394680d9),
	.w8(32'h399580a0),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a90253),
	.w1(32'hba34345a),
	.w2(32'hb9b9b4f5),
	.w3(32'h39637b6c),
	.w4(32'hba27f51a),
	.w5(32'hba079233),
	.w6(32'hba17f442),
	.w7(32'hb9ae577c),
	.w8(32'hba0061c4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e26918),
	.w1(32'h38e913e3),
	.w2(32'h3867e7f2),
	.w3(32'hba1c686a),
	.w4(32'h3921faba),
	.w5(32'hb7d9b060),
	.w6(32'h3761cb4c),
	.w7(32'hb8818feb),
	.w8(32'hb810259c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38667235),
	.w1(32'h37db7a00),
	.w2(32'hb8b4312b),
	.w3(32'hb58885b2),
	.w4(32'h38341ce6),
	.w5(32'hb9046311),
	.w6(32'h38072058),
	.w7(32'hb91e4f2c),
	.w8(32'hb894f9e7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3885853b),
	.w1(32'h39bc16c2),
	.w2(32'h39b66616),
	.w3(32'h389d30ec),
	.w4(32'h39ae8db9),
	.w5(32'h38dcd117),
	.w6(32'h39121280),
	.w7(32'h390db557),
	.w8(32'h389011ec),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39871db7),
	.w1(32'hb9e38d39),
	.w2(32'hb9e11d3b),
	.w3(32'h38e415de),
	.w4(32'hb994294c),
	.w5(32'hb8b9e18d),
	.w6(32'hb9c48461),
	.w7(32'hb98420dd),
	.w8(32'hb975191f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a4585),
	.w1(32'h3a1154c1),
	.w2(32'hba58405d),
	.w3(32'hb8af8596),
	.w4(32'h3ab6741d),
	.w5(32'h3acb4acd),
	.w6(32'h39d4c8de),
	.w7(32'h3982741c),
	.w8(32'h3a2ed1fe),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67f6b8),
	.w1(32'h3a4be725),
	.w2(32'h3a20c5d1),
	.w3(32'h3a899961),
	.w4(32'h3a209acc),
	.w5(32'h39cb3ba0),
	.w6(32'h39fd0d31),
	.w7(32'h390915f2),
	.w8(32'h3a26e594),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08c701),
	.w1(32'hba036845),
	.w2(32'h390c802e),
	.w3(32'h39c00380),
	.w4(32'hba2f0459),
	.w5(32'hb8f4ceff),
	.w6(32'hba14e16b),
	.w7(32'hb9cf780b),
	.w8(32'hb9a25ac2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c18b56),
	.w1(32'h39b4c1fc),
	.w2(32'h39b64150),
	.w3(32'hb938f39c),
	.w4(32'h39e420d9),
	.w5(32'h39bc307e),
	.w6(32'h39d437d0),
	.w7(32'h39851f3c),
	.w8(32'h3a5e53d7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1542c3),
	.w1(32'h39760c46),
	.w2(32'h394849b3),
	.w3(32'h3a0d428d),
	.w4(32'h39374e6c),
	.w5(32'h3824cc3e),
	.w6(32'h3951e111),
	.w7(32'h389ef767),
	.w8(32'h3951e0dc),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993a6f2),
	.w1(32'hb6d026f6),
	.w2(32'h3925a86e),
	.w3(32'h38b95534),
	.w4(32'hb93cb6ed),
	.w5(32'hb8e13154),
	.w6(32'h389a4f2f),
	.w7(32'hb955fab7),
	.w8(32'hb953f4c0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h355e8745),
	.w1(32'hba2b50a0),
	.w2(32'hba046ef5),
	.w3(32'hb8cf1296),
	.w4(32'hb993d015),
	.w5(32'hb9303043),
	.w6(32'hba16b103),
	.w7(32'hb9ee0037),
	.w8(32'hb999e499),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e68d1a),
	.w1(32'hb91eac85),
	.w2(32'hb7c6d559),
	.w3(32'hb93c56a7),
	.w4(32'h3885168d),
	.w5(32'hb841716a),
	.w6(32'hb8cd1cdf),
	.w7(32'hb9498b7d),
	.w8(32'hb9658c45),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b36278),
	.w1(32'hba1a4949),
	.w2(32'hb9c60c83),
	.w3(32'hb811f1f4),
	.w4(32'hba0c3da0),
	.w5(32'hb9aebbcd),
	.w6(32'hb9e49f8c),
	.w7(32'hb9ae0569),
	.w8(32'hb97e5700),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a40ac),
	.w1(32'hb9632235),
	.w2(32'hb8df7cbf),
	.w3(32'hb9310fce),
	.w4(32'hb95930e8),
	.w5(32'hb9dca999),
	.w6(32'hb8e40ac9),
	.w7(32'hb9a71934),
	.w8(32'h39605362),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3957455b),
	.w1(32'h3881764a),
	.w2(32'h396fc232),
	.w3(32'hb8e264be),
	.w4(32'h3889b694),
	.w5(32'h391870a5),
	.w6(32'h37e779fa),
	.w7(32'h38b07d03),
	.w8(32'hb826874a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cefb15),
	.w1(32'h39948e2d),
	.w2(32'h3809a347),
	.w3(32'hb9994eed),
	.w4(32'h398394fb),
	.w5(32'h398af7c3),
	.w6(32'h38d266ec),
	.w7(32'hb8ec3b2c),
	.w8(32'h374638f9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953ceea),
	.w1(32'h38ab35b1),
	.w2(32'h38cc4c6c),
	.w3(32'h3892a4cf),
	.w4(32'h37e06d2e),
	.w5(32'hb88c741c),
	.w6(32'hb8ba8417),
	.w7(32'hb8f09498),
	.w8(32'hb8ab894a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380edc39),
	.w1(32'hb99bc235),
	.w2(32'hb93e4b64),
	.w3(32'hb8c72baf),
	.w4(32'hb91aa70c),
	.w5(32'hb92322e3),
	.w6(32'hba06301d),
	.w7(32'hb93b896e),
	.w8(32'hb93734ae),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99bf7c0),
	.w1(32'h38ca4931),
	.w2(32'h39c2f818),
	.w3(32'hb9adf202),
	.w4(32'h390a14b2),
	.w5(32'h3997b267),
	.w6(32'hb9a56392),
	.w7(32'hb8f19c06),
	.w8(32'h3993b9ff),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eda432),
	.w1(32'h39296575),
	.w2(32'h37aba843),
	.w3(32'hb998e610),
	.w4(32'h38da6f17),
	.w5(32'hb7194918),
	.w6(32'hb992e773),
	.w7(32'hb8df4986),
	.w8(32'hb839d293),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393bbb19),
	.w1(32'hb962d5e8),
	.w2(32'h392d5e00),
	.w3(32'h3842499b),
	.w4(32'hb9d2eb4a),
	.w5(32'hb9c210fe),
	.w6(32'hb8fb6f8f),
	.w7(32'hb840547a),
	.w8(32'hb861aef1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a18f6),
	.w1(32'hb9255053),
	.w2(32'hb8142f0b),
	.w3(32'hba2c7195),
	.w4(32'h36ba760e),
	.w5(32'h37e85ba7),
	.w6(32'hb9826571),
	.w7(32'hb92e340b),
	.w8(32'hb8a3f49f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f0d481),
	.w1(32'h396957bb),
	.w2(32'h39238dff),
	.w3(32'hb913fa6c),
	.w4(32'hb923c6c1),
	.w5(32'hb969e5b9),
	.w6(32'h393dc982),
	.w7(32'hb9731f61),
	.w8(32'hb7be7220),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e8399b),
	.w1(32'hb990f742),
	.w2(32'h37f671c8),
	.w3(32'hb9152047),
	.w4(32'hb98d8e80),
	.w5(32'hb97967d0),
	.w6(32'hb90edb7c),
	.w7(32'hb91cc4e5),
	.w8(32'hb8f0920c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c0d48),
	.w1(32'h37dd9cb6),
	.w2(32'hb947dac0),
	.w3(32'hb9ff7cff),
	.w4(32'h39c77621),
	.w5(32'h39c9b407),
	.w6(32'hb9b75a79),
	.w7(32'h38b81af3),
	.w8(32'h3a0c3860),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ff5b7),
	.w1(32'hb9ef20b8),
	.w2(32'hb8f636e4),
	.w3(32'h3990404f),
	.w4(32'hba07d37b),
	.w5(32'hb9f5e1c3),
	.w6(32'hb92a1683),
	.w7(32'h38a492db),
	.w8(32'h3a19a04e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5597ca),
	.w1(32'h39a8c0b6),
	.w2(32'h3a2ac87d),
	.w3(32'h3a79b050),
	.w4(32'h382f0bff),
	.w5(32'h39d33869),
	.w6(32'h395f7e53),
	.w7(32'h3979c875),
	.w8(32'hb8bee08d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ed9a11),
	.w1(32'hba1ead15),
	.w2(32'hb9f5b91c),
	.w3(32'h370ad12b),
	.w4(32'hba0d1bac),
	.w5(32'hba0b7759),
	.w6(32'hb9fcd855),
	.w7(32'hb9e5733c),
	.w8(32'hb9bcc7cb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e2fcc),
	.w1(32'h37eba2d8),
	.w2(32'h3a2c3d96),
	.w3(32'hb84f3efc),
	.w4(32'h3a12748e),
	.w5(32'h3a3e7932),
	.w6(32'hb9521f68),
	.w7(32'h37eeae65),
	.w8(32'h39abe8b1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd44a0),
	.w1(32'hb9cfb507),
	.w2(32'h3a4ee055),
	.w3(32'hb99bf033),
	.w4(32'hb9df02a4),
	.w5(32'h391653fe),
	.w6(32'hb86a5d3d),
	.w7(32'h3a0ee1bc),
	.w8(32'hb88bc3a3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88dbd27),
	.w1(32'hb8a3b726),
	.w2(32'hb9a4ce07),
	.w3(32'h39148329),
	.w4(32'h39e360ce),
	.w5(32'h3a2e0c17),
	.w6(32'hb9beb58c),
	.w7(32'h39b87bd1),
	.w8(32'h3a5c1f12),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7151e7),
	.w1(32'h3a9cbfbe),
	.w2(32'h3a609b83),
	.w3(32'h3a2404a3),
	.w4(32'h3a722cf1),
	.w5(32'h3a08df39),
	.w6(32'h3a847dda),
	.w7(32'h39a4fd1c),
	.w8(32'h3a850a15),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32d085),
	.w1(32'h39456c52),
	.w2(32'h3900b86e),
	.w3(32'h3a01ff0f),
	.w4(32'h39802b7a),
	.w5(32'h3826b00d),
	.w6(32'h38eab9e8),
	.w7(32'h38145e3a),
	.w8(32'h38bd1480),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29d4ef),
	.w1(32'h3a2f516c),
	.w2(32'h3a42cb05),
	.w3(32'h38b58716),
	.w4(32'h3a0661b5),
	.w5(32'h3a5ed1d2),
	.w6(32'h3a677086),
	.w7(32'h39ea664c),
	.w8(32'h3a42577a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0beafd),
	.w1(32'h398499bc),
	.w2(32'h39952eea),
	.w3(32'h3a01d814),
	.w4(32'h3992b830),
	.w5(32'h395207ec),
	.w6(32'h3964de7f),
	.w7(32'h38da8620),
	.w8(32'h39830614),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72b2fe3),
	.w1(32'hb9d94345),
	.w2(32'hb973d1cd),
	.w3(32'h3884d68b),
	.w4(32'hb9ffa9da),
	.w5(32'hb9a6a171),
	.w6(32'hb98b0956),
	.w7(32'hb995f7de),
	.w8(32'hb9d40faa),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94cc368),
	.w1(32'h398ac84f),
	.w2(32'h399df2fa),
	.w3(32'hb99f1b2f),
	.w4(32'h38f5b5bc),
	.w5(32'h36245c5e),
	.w6(32'hb8f308fc),
	.w7(32'hb87b83cb),
	.w8(32'hb80f224f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a12c80),
	.w1(32'h3a47af7e),
	.w2(32'h39f3c44b),
	.w3(32'h3807d021),
	.w4(32'h3a242941),
	.w5(32'h39ae7310),
	.w6(32'h3a0acfc0),
	.w7(32'h39819280),
	.w8(32'h39ecd40f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a429a),
	.w1(32'hb8cb20d0),
	.w2(32'hb95250e7),
	.w3(32'h392f8420),
	.w4(32'hb909660b),
	.w5(32'hb7bd85a9),
	.w6(32'hb798955b),
	.w7(32'hb9509338),
	.w8(32'hb9651b71),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84c0564),
	.w1(32'h39bc4096),
	.w2(32'hb94487af),
	.w3(32'hb98965a4),
	.w4(32'h398a1939),
	.w5(32'hb895de6f),
	.w6(32'hb6188631),
	.w7(32'h3750b078),
	.w8(32'hb999daa6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e060ff),
	.w1(32'h3a157ba8),
	.w2(32'h3a426815),
	.w3(32'h384f14c3),
	.w4(32'hb94fbff4),
	.w5(32'h3a3d16dc),
	.w6(32'h3a2d9c7a),
	.w7(32'h394c9d34),
	.w8(32'h3991d4a8),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c80e69),
	.w1(32'hb8c323f5),
	.w2(32'hb8c66cb7),
	.w3(32'h3947d6f5),
	.w4(32'h39812d67),
	.w5(32'h38844b09),
	.w6(32'hb9f887ab),
	.w7(32'hb9a09c8c),
	.w8(32'hb97dbc72),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80f09e4),
	.w1(32'hb7b14ed6),
	.w2(32'h398a0a3f),
	.w3(32'h38c9c573),
	.w4(32'hb9169b1b),
	.w5(32'h38c44d73),
	.w6(32'hb9140ac8),
	.w7(32'h3975a6de),
	.w8(32'h3891583b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6899f1e),
	.w1(32'h39cbe3bd),
	.w2(32'h3a24f31b),
	.w3(32'hb7cc6c3d),
	.w4(32'h39c04c0e),
	.w5(32'h39f8227e),
	.w6(32'h38d9209d),
	.w7(32'hb8b054ef),
	.w8(32'h392cab2a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c7200),
	.w1(32'h3a5c56a1),
	.w2(32'h39c39774),
	.w3(32'h39774151),
	.w4(32'h3a328e0d),
	.w5(32'h395e6a09),
	.w6(32'h3a4ed5e7),
	.w7(32'h39987d95),
	.w8(32'h3a12e82f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09dba4),
	.w1(32'h39b7bdb2),
	.w2(32'h394b8d62),
	.w3(32'h39c81afa),
	.w4(32'h39539076),
	.w5(32'h3843ec91),
	.w6(32'h398a8cb8),
	.w7(32'h38c95cff),
	.w8(32'h39832774),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5c8eb),
	.w1(32'h39cdd735),
	.w2(32'h391ea602),
	.w3(32'h39002d81),
	.w4(32'h39a1a005),
	.w5(32'h388dea49),
	.w6(32'h397b1b73),
	.w7(32'h380b4dbd),
	.w8(32'h39685ad4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a283a9),
	.w1(32'h3a06f899),
	.w2(32'h39b1f025),
	.w3(32'h392eca32),
	.w4(32'h39c90a90),
	.w5(32'h3a12ad01),
	.w6(32'h39a2eebc),
	.w7(32'h39a8edb4),
	.w8(32'h39648591),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38d88b),
	.w1(32'hba189946),
	.w2(32'hb9960cb6),
	.w3(32'h3916c8da),
	.w4(32'hba2b3b6a),
	.w5(32'hba11bbd3),
	.w6(32'hba2caf5d),
	.w7(32'hba02c563),
	.w8(32'hb9ffe7a3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30d030),
	.w1(32'h39bf817c),
	.w2(32'h399d16ce),
	.w3(32'hba0fe501),
	.w4(32'h39da2083),
	.w5(32'hb7d9d0f3),
	.w6(32'h396c77ac),
	.w7(32'h38ff898d),
	.w8(32'h3942653f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1b6ad),
	.w1(32'h3989e760),
	.w2(32'h39fadd16),
	.w3(32'h391a2d7a),
	.w4(32'h39632a76),
	.w5(32'h38c93382),
	.w6(32'h3921e38b),
	.w7(32'h3975cbbf),
	.w8(32'h391f65a2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9783e3c),
	.w1(32'h398a98e7),
	.w2(32'h39327ead),
	.w3(32'hb89159ad),
	.w4(32'h39a899a1),
	.w5(32'h390ed1d4),
	.w6(32'h38808910),
	.w7(32'h395f8fa4),
	.w8(32'h39d466dd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398abc92),
	.w1(32'hb923ed9f),
	.w2(32'hba58f4bd),
	.w3(32'h3959874e),
	.w4(32'hb999fde2),
	.w5(32'hb81b8f20),
	.w6(32'hb98c68c7),
	.w7(32'h387cd8ac),
	.w8(32'hb7217a33),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bde59c),
	.w1(32'hb8a33656),
	.w2(32'hb8a13bec),
	.w3(32'hb939326b),
	.w4(32'h3999793c),
	.w5(32'h38ceecac),
	.w6(32'hb8ffbaaf),
	.w7(32'hb95a8bce),
	.w8(32'hb7e37fff),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc19cf),
	.w1(32'h39ecd3c6),
	.w2(32'h392a41b4),
	.w3(32'h3986d544),
	.w4(32'h39a8bc28),
	.w5(32'hb86e8324),
	.w6(32'h393d8872),
	.w7(32'hb91400e4),
	.w8(32'hb77ab792),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393722ae),
	.w1(32'h3853daac),
	.w2(32'hb68fdfc3),
	.w3(32'h385329ae),
	.w4(32'h383195c0),
	.w5(32'hb6405193),
	.w6(32'h387436a1),
	.w7(32'h37a911b6),
	.w8(32'h37cf6597),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94bf1ab),
	.w1(32'h38f3a144),
	.w2(32'h38f220b7),
	.w3(32'h39615054),
	.w4(32'h39aaa0b3),
	.w5(32'h38e14e30),
	.w6(32'hba0e54ce),
	.w7(32'hb9898509),
	.w8(32'h38d0ea9e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b0cbfc),
	.w1(32'h39926dfe),
	.w2(32'h39ca9fbf),
	.w3(32'h38f67059),
	.w4(32'h39454433),
	.w5(32'h399b008b),
	.w6(32'hb7f05424),
	.w7(32'h38f049e4),
	.w8(32'h3868f108),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb628ab38),
	.w1(32'hb6b05c29),
	.w2(32'hb57c109a),
	.w3(32'hb86207a2),
	.w4(32'hb8029860),
	.w5(32'hb76e96c3),
	.w6(32'hb5ad3768),
	.w7(32'hb5fa7e15),
	.w8(32'h370f93cf),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dd0a71),
	.w1(32'h37f3a6e8),
	.w2(32'h387dee09),
	.w3(32'h3826bfec),
	.w4(32'h3787bacf),
	.w5(32'hb7bdf554),
	.w6(32'hb85bbc35),
	.w7(32'h37496124),
	.w8(32'h381d732f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360fe391),
	.w1(32'h375b88c4),
	.w2(32'h37d97f43),
	.w3(32'hb7e31d0e),
	.w4(32'h37bc7039),
	.w5(32'h38ad233a),
	.w6(32'h386baa41),
	.w7(32'h38d7c2cf),
	.w8(32'h39085b2d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb828b7d3),
	.w1(32'h38abcb13),
	.w2(32'h3882e8a8),
	.w3(32'hb7b0cf1d),
	.w4(32'h3883ba36),
	.w5(32'h38bf5185),
	.w6(32'h37cb6970),
	.w7(32'hb6ab82ff),
	.w8(32'h3912c97a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a83b7b),
	.w1(32'h398cce14),
	.w2(32'h39d46f57),
	.w3(32'hb851e38c),
	.w4(32'h38ee4224),
	.w5(32'h3991f58e),
	.w6(32'h38a14b48),
	.w7(32'h395bef9b),
	.w8(32'h39b8f698),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382a7b87),
	.w1(32'h391d54be),
	.w2(32'h3988f24e),
	.w3(32'h38c51c7a),
	.w4(32'h395b3248),
	.w5(32'h3981f95c),
	.w6(32'h36dd3f1c),
	.w7(32'h380f2c96),
	.w8(32'h394c35fe),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9398c18),
	.w1(32'h37841bbe),
	.w2(32'h3639e440),
	.w3(32'hb946108a),
	.w4(32'hb7411858),
	.w5(32'h385f74d5),
	.w6(32'hb8afec0d),
	.w7(32'h365b6867),
	.w8(32'h388398e7),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39092f54),
	.w1(32'h396caed1),
	.w2(32'h392c27e1),
	.w3(32'h39160489),
	.w4(32'h391d89eb),
	.w5(32'h38f9cb0e),
	.w6(32'h388f04ac),
	.w7(32'h38ecd63f),
	.w8(32'h3898cd94),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38abdc56),
	.w1(32'h3946e582),
	.w2(32'h39a40592),
	.w3(32'h38782b1c),
	.w4(32'h3910e4a2),
	.w5(32'h3983817f),
	.w6(32'hb691ee58),
	.w7(32'h38646b85),
	.w8(32'h38e8ca53),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ae1c59),
	.w1(32'h38f5a768),
	.w2(32'h38e545df),
	.w3(32'hb84aed7b),
	.w4(32'h38b51219),
	.w5(32'h38814919),
	.w6(32'hb919f31a),
	.w7(32'h36db8f2d),
	.w8(32'h383009fe),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38613d18),
	.w1(32'h38634298),
	.w2(32'h38a81262),
	.w3(32'h37c0549e),
	.w4(32'h38758d39),
	.w5(32'h38ee595a),
	.w6(32'h38e71a61),
	.w7(32'h38f58966),
	.w8(32'h39065ecd),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76a7636),
	.w1(32'h38862b83),
	.w2(32'h38b71db2),
	.w3(32'h383844b4),
	.w4(32'h382ed30a),
	.w5(32'h38858e1e),
	.w6(32'hb79490cc),
	.w7(32'hb64ee232),
	.w8(32'h37f4d428),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba720a53),
	.w1(32'h38c9203b),
	.w2(32'hb5fcd3b8),
	.w3(32'hba32eb99),
	.w4(32'h39183b72),
	.w5(32'h391ae780),
	.w6(32'hba2eea48),
	.w7(32'h392d22bc),
	.w8(32'h3923321c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dce758),
	.w1(32'hb784344c),
	.w2(32'hb829cd40),
	.w3(32'hb77bfdc5),
	.w4(32'h389884bd),
	.w5(32'h38bae47c),
	.w6(32'hb759ab3f),
	.w7(32'h3774d209),
	.w8(32'h39014a6c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ddd598),
	.w1(32'h371eac0c),
	.w2(32'hb446b351),
	.w3(32'h3889ec7d),
	.w4(32'h3758da89),
	.w5(32'h3767d082),
	.w6(32'h373991e4),
	.w7(32'h36e7c9b3),
	.w8(32'h34997e9a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77a5258),
	.w1(32'h37986df8),
	.w2(32'h3737dd30),
	.w3(32'hb5964649),
	.w4(32'h365a67c3),
	.w5(32'hb746cac4),
	.w6(32'h378b8f50),
	.w7(32'h37601df9),
	.w8(32'hb74ca0ca),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a8dbc),
	.w1(32'h389c495b),
	.w2(32'h38a7975a),
	.w3(32'h36888e5d),
	.w4(32'h382fa478),
	.w5(32'h3878e737),
	.w6(32'h38146c40),
	.w7(32'h3875b177),
	.w8(32'h38529a64),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb864492b),
	.w1(32'h3889001d),
	.w2(32'h38b9b5eb),
	.w3(32'hb941f812),
	.w4(32'h36e4b478),
	.w5(32'h3862a4ff),
	.w6(32'hb8f5e65e),
	.w7(32'h374cd42c),
	.w8(32'h38b38c5e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ce81e),
	.w1(32'h39a0ebf9),
	.w2(32'h39c17e6a),
	.w3(32'h39508b70),
	.w4(32'h399611e2),
	.w5(32'h399b7870),
	.w6(32'h369562c9),
	.w7(32'h38f04ae6),
	.w8(32'h38c4346d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71caaa8),
	.w1(32'h379814aa),
	.w2(32'hb74ca86d),
	.w3(32'h349e3e93),
	.w4(32'h37866967),
	.w5(32'hb76bd9a8),
	.w6(32'h37fd9361),
	.w7(32'hb60e0a68),
	.w8(32'h36b1f8c9),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39057b9b),
	.w1(32'h39a09939),
	.w2(32'h39b833bd),
	.w3(32'h38a5a3d3),
	.w4(32'h393393a2),
	.w5(32'h3962d582),
	.w6(32'hb74d473e),
	.w7(32'h389ad68e),
	.w8(32'h3890815d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6667b),
	.w1(32'h3949b1f6),
	.w2(32'h38e56326),
	.w3(32'hb889d4a1),
	.w4(32'h38d46806),
	.w5(32'h3881414a),
	.w6(32'h37f2b273),
	.w7(32'hb8143a85),
	.w8(32'h37346a61),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900be80),
	.w1(32'h38a64660),
	.w2(32'h394a5750),
	.w3(32'h380e11cd),
	.w4(32'h38bb97ad),
	.w5(32'h39041822),
	.w6(32'h378235b8),
	.w7(32'hb7b64c0c),
	.w8(32'h392d862c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2862f),
	.w1(32'h39884369),
	.w2(32'h39459bd8),
	.w3(32'hb9e6ae71),
	.w4(32'h392b1262),
	.w5(32'h39642a84),
	.w6(32'hb91304a5),
	.w7(32'h394ec81c),
	.w8(32'h3889ac62),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89707f1),
	.w1(32'hb8788470),
	.w2(32'hb6bac01b),
	.w3(32'hb8ab43ca),
	.w4(32'hb84562fc),
	.w5(32'hb65bffa1),
	.w6(32'h37cf8f83),
	.w7(32'h3826ccde),
	.w8(32'h38ae0d66),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83231db),
	.w1(32'hb4281515),
	.w2(32'hb76b687f),
	.w3(32'hb7add26c),
	.w4(32'h36eaacca),
	.w5(32'hb70fe2fc),
	.w6(32'h37b0008b),
	.w7(32'h376802ca),
	.w8(32'hb5517cae),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93cf19c),
	.w1(32'hb871353c),
	.w2(32'hb78d09a1),
	.w3(32'hb94a28f9),
	.w4(32'hb893bf8d),
	.w5(32'hb7aa310f),
	.w6(32'hb92737e1),
	.w7(32'hb823a854),
	.w8(32'hb82d5b47),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c1550b),
	.w1(32'h3914676f),
	.w2(32'h390ed678),
	.w3(32'hb8af86e0),
	.w4(32'hb777d4ab),
	.w5(32'h386356bf),
	.w6(32'h38160a37),
	.w7(32'h367500d5),
	.w8(32'h38af7716),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9422efd),
	.w1(32'hb8595010),
	.w2(32'hb7afc3e2),
	.w3(32'hb936ae4e),
	.w4(32'hb8205fd5),
	.w5(32'hb785fff9),
	.w6(32'hb804b225),
	.w7(32'h37952cbb),
	.w8(32'hb71533b4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7db787f),
	.w1(32'h368b3a74),
	.w2(32'h37a5f0b5),
	.w3(32'hb89d45b2),
	.w4(32'h37bff9c4),
	.w5(32'h387c6e10),
	.w6(32'hb7c8eeda),
	.w7(32'hb7a6087a),
	.w8(32'h38521c80),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378aa6cb),
	.w1(32'h379e9f47),
	.w2(32'h34d1af30),
	.w3(32'h373ad16f),
	.w4(32'h35376a22),
	.w5(32'hb76afc43),
	.w6(32'h381e97a7),
	.w7(32'h37a44662),
	.w8(32'h37825b50),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d368bd),
	.w1(32'h38fdb0ee),
	.w2(32'h393efa73),
	.w3(32'hb6ee280f),
	.w4(32'h3807d7a9),
	.w5(32'h38fbfef8),
	.w6(32'hb844a328),
	.w7(32'h3897f00a),
	.w8(32'h377c9cb0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e3f268),
	.w1(32'h375520d3),
	.w2(32'hb813e913),
	.w3(32'hb80a25d6),
	.w4(32'h37da0899),
	.w5(32'hb771edc3),
	.w6(32'hb6eb5042),
	.w7(32'hb83d832c),
	.w8(32'hb895db82),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dd5eb),
	.w1(32'h38457bf6),
	.w2(32'h3848a294),
	.w3(32'hb93b6d3a),
	.w4(32'h38ac6f98),
	.w5(32'h38e4974e),
	.w6(32'hb9026110),
	.w7(32'h38840176),
	.w8(32'h388f567f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb797bd88),
	.w1(32'h37623e5f),
	.w2(32'hb6c59004),
	.w3(32'hb794f1d3),
	.w4(32'h37883006),
	.w5(32'hb6831b3c),
	.w6(32'h37a97e97),
	.w7(32'h37330ddf),
	.w8(32'h3722fd18),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92cf1e7),
	.w1(32'hb82fee22),
	.w2(32'h365751de),
	.w3(32'h37d900a3),
	.w4(32'h3912b798),
	.w5(32'h392b045e),
	.w6(32'hb900a5be),
	.w7(32'h376b6198),
	.w8(32'h38c2192e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb748931f),
	.w1(32'h37007c78),
	.w2(32'h3659f767),
	.w3(32'hb5f7c95e),
	.w4(32'h35b14d07),
	.w5(32'hb6c4ada0),
	.w6(32'h36e1c603),
	.w7(32'h35d4420a),
	.w8(32'hb543e6c7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3d4af29),
	.w1(32'h35f2e7d3),
	.w2(32'hb76fdd6e),
	.w3(32'hb680a359),
	.w4(32'h36f68c7d),
	.w5(32'hb708cc11),
	.w6(32'h36b8c92b),
	.w7(32'hb63205e0),
	.w8(32'hb703884b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fb386c),
	.w1(32'hb7f84d18),
	.w2(32'h37f42c9f),
	.w3(32'hb92af56d),
	.w4(32'hb89b08a0),
	.w5(32'hb77b3dca),
	.w6(32'hb890cf0e),
	.w7(32'hb7dc3737),
	.w8(32'h386fcce2),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d2309c),
	.w1(32'h37c4534f),
	.w2(32'h39201a5c),
	.w3(32'h38aecb5c),
	.w4(32'h39a1d67f),
	.w5(32'h398f11bf),
	.w6(32'hb939f9f2),
	.w7(32'hb8eecbaf),
	.w8(32'hb604479c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b80ec7),
	.w1(32'hb87dc992),
	.w2(32'hb8856922),
	.w3(32'hb8b9d9a1),
	.w4(32'hb7c8598a),
	.w5(32'hb7c6125f),
	.w6(32'hb5c3f7ce),
	.w7(32'h36f8aa1b),
	.w8(32'hb5c64952),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90467cf),
	.w1(32'h38612bd5),
	.w2(32'h38b767e8),
	.w3(32'hb8b7973e),
	.w4(32'h38900b2f),
	.w5(32'h38edff94),
	.w6(32'hb7f6816f),
	.w7(32'h384841ef),
	.w8(32'h38a2cfe4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a6ed66),
	.w1(32'h392cede7),
	.w2(32'h38efff8b),
	.w3(32'hb8ae143b),
	.w4(32'h38aef327),
	.w5(32'h38c206af),
	.w6(32'hb7252b6a),
	.w7(32'h38695bf8),
	.w8(32'h37eae788),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930882f),
	.w1(32'h39d4dfd2),
	.w2(32'h3a0c1c2f),
	.w3(32'h39675e6d),
	.w4(32'h398ab373),
	.w5(32'h39c1df7c),
	.w6(32'h38cac696),
	.w7(32'hb6bb3b0d),
	.w8(32'h38972e2b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a75048),
	.w1(32'h39135f17),
	.w2(32'h3971d56e),
	.w3(32'hb89fb42b),
	.w4(32'h37125034),
	.w5(32'h38bbd368),
	.w6(32'hb7d238bc),
	.w7(32'hb8311eb4),
	.w8(32'h38c0a3a4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dd6268),
	.w1(32'h390bd8e1),
	.w2(32'h397b0050),
	.w3(32'h38e802da),
	.w4(32'h39788497),
	.w5(32'h39b1cbdc),
	.w6(32'h38895d42),
	.w7(32'h38c7edea),
	.w8(32'h393f13e7),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8955fb6),
	.w1(32'h3836175a),
	.w2(32'h378f757b),
	.w3(32'h383a6957),
	.w4(32'h38052b52),
	.w5(32'hb6423851),
	.w6(32'h38589c7a),
	.w7(32'h37bc34ac),
	.w8(32'hb82cd899),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90bd343),
	.w1(32'h38909a2a),
	.w2(32'h390c6607),
	.w3(32'hb92e335c),
	.w4(32'h37213820),
	.w5(32'h38d44d1c),
	.w6(32'h3864e56f),
	.w7(32'h3887e141),
	.w8(32'h391bc7b6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362d2d39),
	.w1(32'h36b457f4),
	.w2(32'hb68bcbe8),
	.w3(32'h3580f5c2),
	.w4(32'h3692a4f4),
	.w5(32'hb68f0a1b),
	.w6(32'h36cfa541),
	.w7(32'hb6fb4f31),
	.w8(32'hb67ada39),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3853df60),
	.w1(32'h37d4d482),
	.w2(32'h3879c40d),
	.w3(32'h38602ef5),
	.w4(32'h3877eefe),
	.w5(32'h38118f26),
	.w6(32'h38910fba),
	.w7(32'h3816a33b),
	.w8(32'h382d1062),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c3a3ac),
	.w1(32'hb8c94713),
	.w2(32'h3824720f),
	.w3(32'hb887b04a),
	.w4(32'hb6beb11e),
	.w5(32'h38da670d),
	.w6(32'hb83fdcef),
	.w7(32'h38e7255f),
	.w8(32'h353a7cec),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c01e6e),
	.w1(32'h38f6b93d),
	.w2(32'h3905dee8),
	.w3(32'h38d56ed8),
	.w4(32'h380b08b5),
	.w5(32'h38d60d0d),
	.w6(32'h391e1d9c),
	.w7(32'h38c54e98),
	.w8(32'h393f4f2f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f26554),
	.w1(32'h376c9b84),
	.w2(32'hb85522a5),
	.w3(32'hb7a62e43),
	.w4(32'h37e03956),
	.w5(32'hb837aedf),
	.w6(32'h3693176b),
	.w7(32'hb806fcb2),
	.w8(32'h37402dfc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363f9f76),
	.w1(32'h37ad2ef5),
	.w2(32'h37c64558),
	.w3(32'hb5ecaa6d),
	.w4(32'h37723b4e),
	.w5(32'h37517835),
	.w6(32'h37a8919c),
	.w7(32'h37e256b0),
	.w8(32'h37a733c2),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d9100),
	.w1(32'h38c4c070),
	.w2(32'hb689d7a1),
	.w3(32'hb8c3b588),
	.w4(32'h388a9a1a),
	.w5(32'hb750bc63),
	.w6(32'hb8c3585d),
	.w7(32'hb8662990),
	.w8(32'hb804bc61),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39402a27),
	.w1(32'h38c9c4f3),
	.w2(32'h39654eb2),
	.w3(32'h37ea2fa3),
	.w4(32'hb826567b),
	.w5(32'h3932e839),
	.w6(32'h368be6a4),
	.w7(32'hb956f7df),
	.w8(32'h3924e1c6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39878aaa),
	.w1(32'h3906f374),
	.w2(32'h3923ea4d),
	.w3(32'h3901c90a),
	.w4(32'h3904438b),
	.w5(32'h39104e02),
	.w6(32'h3874bffd),
	.w7(32'h38909ca9),
	.w8(32'h38d63589),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8166912),
	.w1(32'hb5a9f60e),
	.w2(32'hb650f12f),
	.w3(32'hb79217cf),
	.w4(32'hb7841900),
	.w5(32'h37ad047c),
	.w6(32'hb789cb22),
	.w7(32'h36f5e213),
	.w8(32'h38299c32),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6001f),
	.w1(32'h3a1526e6),
	.w2(32'h3a514062),
	.w3(32'h39f5319a),
	.w4(32'h3a1dbae8),
	.w5(32'h3a23a3af),
	.w6(32'h38a72926),
	.w7(32'h38e3f519),
	.w8(32'h392b8319),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a1951),
	.w1(32'h39a7d477),
	.w2(32'h39ce7dd2),
	.w3(32'hb9b3d82e),
	.w4(32'h390222f3),
	.w5(32'h397b5531),
	.w6(32'hb8ec853e),
	.w7(32'h39052775),
	.w8(32'h3852dacf),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72d7109),
	.w1(32'hb781d437),
	.w2(32'h38288f8f),
	.w3(32'h37055aa3),
	.w4(32'hb7f45516),
	.w5(32'h37e9434a),
	.w6(32'hb76ed129),
	.w7(32'h3816859c),
	.w8(32'hb765c6f4),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37539a18),
	.w1(32'hb84da537),
	.w2(32'h37facfc5),
	.w3(32'hb68b2820),
	.w4(32'hb800a96a),
	.w5(32'h37f9ba69),
	.w6(32'hb82df005),
	.w7(32'h37b054b5),
	.w8(32'hb8969a7d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86ab3b7),
	.w1(32'h37121e76),
	.w2(32'h36f6ca58),
	.w3(32'hb83685d2),
	.w4(32'h370d025e),
	.w5(32'h36ddf682),
	.w6(32'h36fa114a),
	.w7(32'h3705d3a8),
	.w8(32'hb70cda4f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76f8d6b),
	.w1(32'h377680cf),
	.w2(32'h3778d660),
	.w3(32'hb7347600),
	.w4(32'h375eb3c1),
	.w5(32'h376e539d),
	.w6(32'h37527cf2),
	.w7(32'h376a187b),
	.w8(32'h3734009e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b1541b),
	.w1(32'hb7af060a),
	.w2(32'hb7d68674),
	.w3(32'h3870e4e1),
	.w4(32'h38bc2267),
	.w5(32'h38041216),
	.w6(32'hb8af79d7),
	.w7(32'h3744cdef),
	.w8(32'h3872e43e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381825ea),
	.w1(32'h38cef7cc),
	.w2(32'h3922c513),
	.w3(32'hb8208bf8),
	.w4(32'h388082ee),
	.w5(32'h391c3a8f),
	.w6(32'hb8a98c8c),
	.w7(32'hb80761fd),
	.w8(32'h37d0a64d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389fe22e),
	.w1(32'h39af3b5d),
	.w2(32'h3998b7d5),
	.w3(32'hb72de78f),
	.w4(32'h396bbc06),
	.w5(32'h3938391c),
	.w6(32'h38ea6086),
	.w7(32'h38cfa319),
	.w8(32'h38a6ea97),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cd378b),
	.w1(32'hb67beb17),
	.w2(32'hb78579eb),
	.w3(32'hb8f95d48),
	.w4(32'hb63bb112),
	.w5(32'hb6cc684e),
	.w6(32'hb868fcb5),
	.w7(32'hb813ff12),
	.w8(32'hb77eeca4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39310b4e),
	.w1(32'h3988ab9a),
	.w2(32'h396580bb),
	.w3(32'h39158acf),
	.w4(32'h3981ab32),
	.w5(32'h394f68cc),
	.w6(32'h385a259d),
	.w7(32'h376c53a0),
	.w8(32'h38905ef5),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39365648),
	.w1(32'h38f47f1a),
	.w2(32'h39152608),
	.w3(32'h38a77890),
	.w4(32'h38cd09a5),
	.w5(32'h39436acf),
	.w6(32'h36c21911),
	.w7(32'h38482f0b),
	.w8(32'h3837ae99),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73e297a),
	.w1(32'h3739ea0a),
	.w2(32'hb753dd0d),
	.w3(32'hb727b2b7),
	.w4(32'h3722e43a),
	.w5(32'hb75ba6b7),
	.w6(32'h371b2dc9),
	.w7(32'hb740f89c),
	.w8(32'h35d26ac1),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3883e0f7),
	.w1(32'h3799e402),
	.w2(32'h38c5088b),
	.w3(32'h38be6fd9),
	.w4(32'h38476b17),
	.w5(32'h3932050e),
	.w6(32'h38a16dea),
	.w7(32'h38b91dbb),
	.w8(32'h38a784b0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7199e28),
	.w1(32'h37805be9),
	.w2(32'hb69d9dbc),
	.w3(32'hb6315933),
	.w4(32'h377f27cd),
	.w5(32'hb6ee3101),
	.w6(32'h37c098ef),
	.w7(32'h3733dcc3),
	.w8(32'h376381fb),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383cc18e),
	.w1(32'h389f1345),
	.w2(32'h395e84f1),
	.w3(32'hb7bdfd76),
	.w4(32'h388af709),
	.w5(32'h39595f5e),
	.w6(32'hb822e2e4),
	.w7(32'h37e62397),
	.w8(32'h38f780ec),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88df599),
	.w1(32'h37362d90),
	.w2(32'h38ecb64a),
	.w3(32'hb934a8a4),
	.w4(32'hb61a9b1d),
	.w5(32'h38e77597),
	.w6(32'hb8927627),
	.w7(32'h38cda0a4),
	.w8(32'h38a0628a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8941503),
	.w1(32'h38dc943c),
	.w2(32'h39109dfd),
	.w3(32'hb86f1795),
	.w4(32'hb6a7510a),
	.w5(32'h3885351f),
	.w6(32'hb8938328),
	.w7(32'hb89aed36),
	.w8(32'h379734fb),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8179133),
	.w1(32'hb8728ae1),
	.w2(32'hb7bcef2e),
	.w3(32'hb849c15a),
	.w4(32'hb872ead0),
	.w5(32'hb7fca1d4),
	.w6(32'hb81d2076),
	.w7(32'hb710ba2f),
	.w8(32'hb82e9391),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9182a8b),
	.w1(32'h39379d7a),
	.w2(32'h3985115d),
	.w3(32'hb96a373b),
	.w4(32'hb7407e5e),
	.w5(32'h39140115),
	.w6(32'hb85baf65),
	.w7(32'h38b51fef),
	.w8(32'h39408f68),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d37c0e),
	.w1(32'h390058b4),
	.w2(32'h391138b3),
	.w3(32'h35cb6955),
	.w4(32'h39081983),
	.w5(32'h392388fc),
	.w6(32'h384c85be),
	.w7(32'h386fae72),
	.w8(32'h390de34e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39991e6a),
	.w1(32'h39f5046f),
	.w2(32'h39ccdec8),
	.w3(32'h3950b577),
	.w4(32'h39bbe3ec),
	.w5(32'h3992af53),
	.w6(32'h38f6a914),
	.w7(32'h383ff850),
	.w8(32'h36f88e2f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85f9757),
	.w1(32'hb73b07df),
	.w2(32'hb70672ce),
	.w3(32'hb8969759),
	.w4(32'hb776a7be),
	.w5(32'hb7566035),
	.w6(32'hb7171565),
	.w7(32'hb679bedb),
	.w8(32'h3600fcfe),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c1fb81),
	.w1(32'hb6aeff35),
	.w2(32'hb673de83),
	.w3(32'hb7b4641a),
	.w4(32'hb738e163),
	.w5(32'h35f51fd1),
	.w6(32'h36e6cabe),
	.w7(32'h36f5be6d),
	.w8(32'h370c90ab),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3909b8f4),
	.w1(32'h38ec0199),
	.w2(32'h38dac0d5),
	.w3(32'h3838a280),
	.w4(32'h38e247e4),
	.w5(32'h381739be),
	.w6(32'hb9de3eb3),
	.w7(32'hb948498b),
	.w8(32'hb8b3e72c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7dc4b),
	.w1(32'h385c5f04),
	.w2(32'h38e6100c),
	.w3(32'h37fbfbc4),
	.w4(32'h3975f085),
	.w5(32'h39948039),
	.w6(32'hb90205e7),
	.w7(32'hb92e0c2c),
	.w8(32'hb6f6ad8e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a93ba8),
	.w1(32'h395293bd),
	.w2(32'h3986c2b9),
	.w3(32'hb82900a4),
	.w4(32'h389409e2),
	.w5(32'h390a01c0),
	.w6(32'hb8cf7515),
	.w7(32'hb818c6dc),
	.w8(32'h3877d24b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3741007a),
	.w1(32'hb78a5613),
	.w2(32'h38a60609),
	.w3(32'h37198616),
	.w4(32'h391b7f13),
	.w5(32'h38c5382a),
	.w6(32'h398a0cb0),
	.w7(32'h393f04c3),
	.w8(32'h393bcad5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7aeb073),
	.w1(32'h35b4eff3),
	.w2(32'h37a7f50f),
	.w3(32'h38327901),
	.w4(32'h37c526a9),
	.w5(32'h37b59f9d),
	.w6(32'h37cdb88e),
	.w7(32'hb6aa03ab),
	.w8(32'h37962c57),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3829e573),
	.w1(32'h381bfa49),
	.w2(32'h3829d3e3),
	.w3(32'h37ac8bd0),
	.w4(32'h379ee698),
	.w5(32'h37e6c145),
	.w6(32'h3661773d),
	.w7(32'h35ad8838),
	.w8(32'h3651ce8f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388808ab),
	.w1(32'hb68e6858),
	.w2(32'h39442c38),
	.w3(32'h39c3eb85),
	.w4(32'h39f11380),
	.w5(32'h39d57561),
	.w6(32'hb8e7340f),
	.w7(32'h391e2fb0),
	.w8(32'h396d4306),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fa3f39),
	.w1(32'h39a8075d),
	.w2(32'h39f9917d),
	.w3(32'h3940d1c2),
	.w4(32'h39b2b42a),
	.w5(32'h39cb4697),
	.w6(32'hb7a4c676),
	.w7(32'h37b9660a),
	.w8(32'h38d91749),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fcacc2),
	.w1(32'hb88272ea),
	.w2(32'h39121c4d),
	.w3(32'h378d210b),
	.w4(32'h37b7900f),
	.w5(32'h39405164),
	.w6(32'hb8e38a1f),
	.w7(32'hb8ff46bc),
	.w8(32'h391010f9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988eb99),
	.w1(32'hb876f57d),
	.w2(32'hb6a0c68d),
	.w3(32'hb960bd9b),
	.w4(32'hb8312940),
	.w5(32'h38337a8a),
	.w6(32'hb93fb5f1),
	.w7(32'hb6459dc1),
	.w8(32'h375899f0),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0cc3b),
	.w1(32'h3972310a),
	.w2(32'h3951ffbe),
	.w3(32'hb92cee20),
	.w4(32'h38c3eaa6),
	.w5(32'h38989f46),
	.w6(32'h37b5ecff),
	.w7(32'h3812b67e),
	.w8(32'h38d801b2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8389951),
	.w1(32'h3754c189),
	.w2(32'h378ddf2d),
	.w3(32'hb877b8a8),
	.w4(32'hb54d0121),
	.w5(32'h36977298),
	.w6(32'h3702790d),
	.w7(32'h36f5e2ae),
	.w8(32'h369849d7),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37281fab),
	.w1(32'h380c08fe),
	.w2(32'h36cc2ea2),
	.w3(32'h35df79f8),
	.w4(32'hb526d3ba),
	.w5(32'hb8367a1c),
	.w6(32'hb5d35a94),
	.w7(32'hb7e89de5),
	.w8(32'hb5c54672),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86f747c),
	.w1(32'hb78fdb9e),
	.w2(32'hb8f8cf4b),
	.w3(32'hb81628cd),
	.w4(32'h38211b92),
	.w5(32'hb898fb2b),
	.w6(32'hb74ec2f5),
	.w7(32'hb7335e6b),
	.w8(32'hb88ba90f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8320f96),
	.w1(32'hb780b3aa),
	.w2(32'h37924b97),
	.w3(32'hb838d466),
	.w4(32'hb71c2fac),
	.w5(32'h37e9bc16),
	.w6(32'hb7201428),
	.w7(32'h37be6b83),
	.w8(32'hb82795d0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3604926e),
	.w1(32'h37cfef8e),
	.w2(32'h3820480a),
	.w3(32'h384637c4),
	.w4(32'h385f69be),
	.w5(32'h38767818),
	.w6(32'hb6e2751c),
	.w7(32'h381822ee),
	.w8(32'h385a755f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7efc620),
	.w1(32'h36dade2d),
	.w2(32'h394cd391),
	.w3(32'h38cc43ef),
	.w4(32'h3907afe1),
	.w5(32'h395a7538),
	.w6(32'hb92bcad0),
	.w7(32'hb8da5a3f),
	.w8(32'h375cd7ec),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b42c71),
	.w1(32'h38e148b2),
	.w2(32'hb80b8d23),
	.w3(32'hb867f729),
	.w4(32'h38b22e5a),
	.w5(32'hb7c562e2),
	.w6(32'hb7f9eab2),
	.w7(32'hb8bf3c9f),
	.w8(32'h36eb24f8),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb702f8ac),
	.w1(32'h38b6020d),
	.w2(32'h37d7494b),
	.w3(32'hb7b0c6c5),
	.w4(32'h384e3fa2),
	.w5(32'hb8394177),
	.w6(32'h378c6b2b),
	.w7(32'hb8109d27),
	.w8(32'h37cee394),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0210f9),
	.w1(32'hb903cdb9),
	.w2(32'h39ec3ab9),
	.w3(32'h39547ee1),
	.w4(32'h392759fc),
	.w5(32'h39c5e16c),
	.w6(32'h3823d887),
	.w7(32'hb881fa89),
	.w8(32'h3966695c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ef85b6),
	.w1(32'h3895bd5f),
	.w2(32'h38fd1767),
	.w3(32'h381b7a5a),
	.w4(32'h38fd9a99),
	.w5(32'h38c6e53c),
	.w6(32'h3654a443),
	.w7(32'h3788d32c),
	.w8(32'h386233a5),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370b24aa),
	.w1(32'h3787dc98),
	.w2(32'hb65416b7),
	.w3(32'h370e75ae),
	.w4(32'h3788a20e),
	.w5(32'hb68c615d),
	.w6(32'h3744bcd1),
	.w7(32'hb717ec6e),
	.w8(32'hb62a004e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75bf513),
	.w1(32'h37db97c9),
	.w2(32'h38b0983b),
	.w3(32'hb7f09b70),
	.w4(32'h385d55d6),
	.w5(32'h38f64ebf),
	.w6(32'hb8c45554),
	.w7(32'hb75896ae),
	.w8(32'h384cc4bf),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cac726),
	.w1(32'h3799fc5d),
	.w2(32'h37bca042),
	.w3(32'h34419893),
	.w4(32'h35c99cc0),
	.w5(32'h36dbd354),
	.w6(32'h36eabffe),
	.w7(32'h3702c7c6),
	.w8(32'h352b2f32),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378dfaa2),
	.w1(32'h37cd95a8),
	.w2(32'h370ab14d),
	.w3(32'h377ad6db),
	.w4(32'h37aa7978),
	.w5(32'h368e6852),
	.w6(32'h37e1134b),
	.w7(32'h3688c89b),
	.w8(32'h37792832),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3724ea4d),
	.w1(32'h378c145a),
	.w2(32'hb6d20764),
	.w3(32'h3623bc41),
	.w4(32'h3781ea27),
	.w5(32'hb729277c),
	.w6(32'h37317e1d),
	.w7(32'hb76a68b1),
	.w8(32'hb6a86dfd),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3409f4d9),
	.w1(32'hb768d450),
	.w2(32'h3752b857),
	.w3(32'hb6aaf0ed),
	.w4(32'hb72b95dd),
	.w5(32'h3791ff5a),
	.w6(32'hb7c43a1f),
	.w7(32'h350901e9),
	.w8(32'hb7b0ac00),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b671c4),
	.w1(32'hb860720f),
	.w2(32'hb8929194),
	.w3(32'hb847bebb),
	.w4(32'hb7c8c5ee),
	.w5(32'hb6e81275),
	.w6(32'hb7e61a13),
	.w7(32'hb7cb6093),
	.w8(32'hb7f84e2e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c5ff9f),
	.w1(32'h3913093a),
	.w2(32'h39ac1474),
	.w3(32'h37ec7ff0),
	.w4(32'h390ed784),
	.w5(32'h3999f27c),
	.w6(32'h390eaddb),
	.w7(32'h390ea500),
	.w8(32'h3907d2e3),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37809393),
	.w1(32'h38e92a01),
	.w2(32'h392c1bfd),
	.w3(32'h370514a1),
	.w4(32'h388b2c17),
	.w5(32'h3918c820),
	.w6(32'hb81429dc),
	.w7(32'h370cce3f),
	.w8(32'h3850a56c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb776f1fb),
	.w1(32'h395625ce),
	.w2(32'h395baedb),
	.w3(32'h38fdb89c),
	.w4(32'h3966dcb0),
	.w5(32'h3957e029),
	.w6(32'h389e397d),
	.w7(32'h38e613eb),
	.w8(32'h38b738b1),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b5bee7),
	.w1(32'hb780560c),
	.w2(32'h355dbf83),
	.w3(32'hb6b20b8e),
	.w4(32'hb7fd19cc),
	.w5(32'hb7516021),
	.w6(32'hb6823c5d),
	.w7(32'hb5e8da9a),
	.w8(32'hb7925301),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79f6e79),
	.w1(32'h37ea0b81),
	.w2(32'hb797a248),
	.w3(32'hb7ca18c2),
	.w4(32'h37c585fe),
	.w5(32'hb7a4468a),
	.w6(32'h37629556),
	.w7(32'hb7b2a0e9),
	.w8(32'hb717d92b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36374d6b),
	.w1(32'h371d5c8a),
	.w2(32'hb7158877),
	.w3(32'hb66871eb),
	.w4(32'h3730b6b5),
	.w5(32'hb707e22c),
	.w6(32'h36bb38f6),
	.w7(32'hb74befee),
	.w8(32'hb5a171f6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368e65f3),
	.w1(32'h37412a75),
	.w2(32'hb6f8658b),
	.w3(32'h368a0e94),
	.w4(32'h37509591),
	.w5(32'hb705ddb1),
	.w6(32'h36f69154),
	.w7(32'hb725cd39),
	.w8(32'hb617570d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7eeb8db),
	.w1(32'h392bc968),
	.w2(32'h3988ad05),
	.w3(32'hb78d8a38),
	.w4(32'h3733bf1d),
	.w5(32'h38b583c8),
	.w6(32'hb58151cd),
	.w7(32'hb7addc29),
	.w8(32'h382f3129),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3772debc),
	.w1(32'h377ca74b),
	.w2(32'hb7b61906),
	.w3(32'hb84e5f70),
	.w4(32'h375db6b3),
	.w5(32'hb7b94456),
	.w6(32'h3712aea0),
	.w7(32'hb7a4cf5d),
	.w8(32'hb7335c47),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d2928e),
	.w1(32'hb6a9370c),
	.w2(32'hb8551baf),
	.w3(32'hb81c0d9c),
	.w4(32'h37384d8d),
	.w5(32'hb805591f),
	.w6(32'h378f2ff5),
	.w7(32'hb1a23794),
	.w8(32'h37a4d7d8),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bfdf5c),
	.w1(32'h38adf0f6),
	.w2(32'h38b44385),
	.w3(32'h387e771a),
	.w4(32'h386164af),
	.w5(32'h38ca3163),
	.w6(32'h385c2de8),
	.w7(32'h3899f111),
	.w8(32'h3867dc87),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7103e5f),
	.w1(32'h368d3c87),
	.w2(32'hb6ce2358),
	.w3(32'hb692f14e),
	.w4(32'h3551dc73),
	.w5(32'hb73071b5),
	.w6(32'h362b9390),
	.w7(32'hb7140b41),
	.w8(32'hb6e40200),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38813e7d),
	.w1(32'h3908384d),
	.w2(32'h390ca8d7),
	.w3(32'h387882b0),
	.w4(32'h38a0ebb2),
	.w5(32'h381ca0ed),
	.w6(32'h37dea6c5),
	.w7(32'hb6037b69),
	.w8(32'hb82d3e06),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3861854b),
	.w1(32'h341a14ca),
	.w2(32'hb83d00bf),
	.w3(32'hb78eb585),
	.w4(32'h37a349cf),
	.w5(32'hb7ee0f1a),
	.w6(32'h382046cf),
	.w7(32'hb6df9281),
	.w8(32'h36b39d62),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c905cf),
	.w1(32'h39a15d34),
	.w2(32'h3993f3a7),
	.w3(32'hb88af2d7),
	.w4(32'h38ab601e),
	.w5(32'h38f9cc38),
	.w6(32'h3996f2f4),
	.w7(32'h3991f51d),
	.w8(32'h399f8fd2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368b63cc),
	.w1(32'hb818f050),
	.w2(32'hb853e81a),
	.w3(32'h375264fb),
	.w4(32'hb91bca75),
	.w5(32'h36554912),
	.w6(32'hb99b131e),
	.w7(32'hb9e45b6f),
	.w8(32'hb8101ed8),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37780d88),
	.w1(32'hb9bb8ce2),
	.w2(32'hb9f98287),
	.w3(32'h38929ab2),
	.w4(32'hb9aa666d),
	.w5(32'hb8929616),
	.w6(32'hba00e5ce),
	.w7(32'hb9b9b5d0),
	.w8(32'hb90da4fb),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule