module layer_8_featuremap_66(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbab8e),
	.w1(32'hbc6fec35),
	.w2(32'hbc90969d),
	.w3(32'h3cbc49ac),
	.w4(32'h3ca7aac8),
	.w5(32'hba3a2ba6),
	.w6(32'hba39ff1e),
	.w7(32'hb9873a05),
	.w8(32'hbb3b969d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b065cd7),
	.w1(32'hb93bc8e7),
	.w2(32'h39680e72),
	.w3(32'h3bdd1fde),
	.w4(32'h3c48741c),
	.w5(32'h3bbff246),
	.w6(32'hbc64e089),
	.w7(32'hbc0cdd73),
	.w8(32'hbbe6b4a2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0583e),
	.w1(32'h3bbcad1e),
	.w2(32'h3bd25f29),
	.w3(32'h3c3b94e1),
	.w4(32'h3c8ef1ab),
	.w5(32'h3c3c4ef7),
	.w6(32'hbc0e9394),
	.w7(32'hbb8fa3ce),
	.w8(32'h3bbff60e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fe471),
	.w1(32'hbc49a89e),
	.w2(32'hbbfb7f73),
	.w3(32'hbc4b0758),
	.w4(32'hbcb50ce9),
	.w5(32'hbce2c73c),
	.w6(32'h3b9a8478),
	.w7(32'h39ba4d6e),
	.w8(32'hbc7bf577),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad42726),
	.w1(32'h3bb3b659),
	.w2(32'h3b728ae7),
	.w3(32'h3c4e6978),
	.w4(32'h3cee3c34),
	.w5(32'h3cb261a6),
	.w6(32'hbca0b270),
	.w7(32'hbc4d236d),
	.w8(32'hbcbc9aaa),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9eda4c),
	.w1(32'h3c5d518f),
	.w2(32'h3c43cc95),
	.w3(32'h3d2573ae),
	.w4(32'h3dabb6c4),
	.w5(32'h3d3e1f38),
	.w6(32'hbd34b622),
	.w7(32'hbce13240),
	.w8(32'h3a65ca1b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5ee54),
	.w1(32'h3a4eb688),
	.w2(32'h3aa37c06),
	.w3(32'h3bd8e12e),
	.w4(32'h3c561919),
	.w5(32'h3c07c3f5),
	.w6(32'hbc345a79),
	.w7(32'hbbe330d9),
	.w8(32'hbc8a40b1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49dd39),
	.w1(32'hbb8183eb),
	.w2(32'hbbddceb3),
	.w3(32'h3c259702),
	.w4(32'h3c8e7a66),
	.w5(32'h3b4a7f27),
	.w6(32'hbc7d1c2e),
	.w7(32'hbc8535ce),
	.w8(32'hbc40ca6b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8c191),
	.w1(32'h3c0bc2b5),
	.w2(32'h3c16ec34),
	.w3(32'h3c7b97ae),
	.w4(32'h3cd77932),
	.w5(32'h3c99bec9),
	.w6(32'hbc544e2f),
	.w7(32'hbbefa76e),
	.w8(32'hbc1a45e2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fb1b2),
	.w1(32'hbc041901),
	.w2(32'hbcb0618a),
	.w3(32'h3bf4804d),
	.w4(32'h3bc36003),
	.w5(32'hbadca50d),
	.w6(32'h3bd25de7),
	.w7(32'hbbbbdee1),
	.w8(32'hbcda79d3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0410af),
	.w1(32'hbc55c080),
	.w2(32'h3b4ea918),
	.w3(32'h3c63def5),
	.w4(32'h3ca214a7),
	.w5(32'h3bc65341),
	.w6(32'hbc1faeab),
	.w7(32'hbb8894a3),
	.w8(32'hbab29c8d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bc07a),
	.w1(32'hbc6d9626),
	.w2(32'hbc9bd719),
	.w3(32'h3c4c004a),
	.w4(32'h3c8a91c4),
	.w5(32'h3abeebbc),
	.w6(32'hbb3bbfc9),
	.w7(32'h3c0fec0e),
	.w8(32'h3bf065cb),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf69f71),
	.w1(32'h3b630cd6),
	.w2(32'hb8ec9138),
	.w3(32'h3bc13e00),
	.w4(32'h3ca1eb40),
	.w5(32'h3c719e82),
	.w6(32'hbc51c5a9),
	.w7(32'hbbf0e08b),
	.w8(32'hbccd35c8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a131b94),
	.w1(32'h3b8d7f28),
	.w2(32'hbbd324e4),
	.w3(32'h3d504d12),
	.w4(32'h3db2750a),
	.w5(32'h3d48091c),
	.w6(32'hbd2d235d),
	.w7(32'hbd0a7b09),
	.w8(32'hbc5d1e04),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b571bfd),
	.w1(32'h3b9ea422),
	.w2(32'hb964a0a0),
	.w3(32'h3ce613b2),
	.w4(32'h3d353ecf),
	.w5(32'h3cd52194),
	.w6(32'hbcc99329),
	.w7(32'hbc84a5b7),
	.w8(32'hbbebe0aa),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafded5),
	.w1(32'hba07b007),
	.w2(32'hbb927423),
	.w3(32'h3c3cb2ae),
	.w4(32'h3c80d9d0),
	.w5(32'h3a6c7bc8),
	.w6(32'hbc357615),
	.w7(32'hbbe60d33),
	.w8(32'hbb8b3f75),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79b3a4),
	.w1(32'hbb16e7d7),
	.w2(32'hbbfb14ec),
	.w3(32'h3ca57e32),
	.w4(32'h3b4127cd),
	.w5(32'h3c2c64ef),
	.w6(32'hbc3b838d),
	.w7(32'hbc9ca566),
	.w8(32'hbc801fa4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d940d),
	.w1(32'hbc576b8f),
	.w2(32'hbc903300),
	.w3(32'h3beea310),
	.w4(32'h3c781048),
	.w5(32'h3bd34ab7),
	.w6(32'hbc04d974),
	.w7(32'h3a420283),
	.w8(32'hbbd3a26d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e9f7f),
	.w1(32'hbd88fa59),
	.w2(32'hbd86d414),
	.w3(32'h3d5f7341),
	.w4(32'h3d231800),
	.w5(32'hbcc44dc9),
	.w6(32'h3ceda813),
	.w7(32'h3c84a918),
	.w8(32'h3bce45fb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc122938),
	.w1(32'hbcf7ee45),
	.w2(32'hbca49612),
	.w3(32'h3cae3446),
	.w4(32'h3c75c162),
	.w5(32'h3cc71213),
	.w6(32'hbcc39834),
	.w7(32'hbcc37dab),
	.w8(32'hbc1b114e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21428a),
	.w1(32'h3b982901),
	.w2(32'hbace5c6a),
	.w3(32'h3c187347),
	.w4(32'h3cb8450a),
	.w5(32'h3c1853e3),
	.w6(32'hbc1f5978),
	.w7(32'h3c0da59a),
	.w8(32'hbbf109df),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab12d2),
	.w1(32'h3c1fd3ef),
	.w2(32'h3c169e74),
	.w3(32'h3c8a28ee),
	.w4(32'h3d092500),
	.w5(32'h3ccdce3b),
	.w6(32'hbd029f97),
	.w7(32'hbcb9b3f2),
	.w8(32'h3d0ea091),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10dd54),
	.w1(32'hbd0744e1),
	.w2(32'hbd5e4a80),
	.w3(32'hbbd61b07),
	.w4(32'hbd8e789f),
	.w5(32'hbdaa5267),
	.w6(32'h3dd19926),
	.w7(32'h3d611c1d),
	.w8(32'hbc96056f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7d868),
	.w1(32'h3bc13ed2),
	.w2(32'h3a3a8ee1),
	.w3(32'h3c909764),
	.w4(32'h3cd93c3e),
	.w5(32'h3c453419),
	.w6(32'hbcc8b959),
	.w7(32'hbca5477a),
	.w8(32'hbcb93761),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d72c7),
	.w1(32'hbc22dcd9),
	.w2(32'h3783c98c),
	.w3(32'h3cd3fe9c),
	.w4(32'h3ccd987f),
	.w5(32'h3d0e1511),
	.w6(32'hbd022a83),
	.w7(32'hbce6bd35),
	.w8(32'h3d10e163),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fdf6b),
	.w1(32'hbc38e4e8),
	.w2(32'hbce02fa3),
	.w3(32'hbce23144),
	.w4(32'hbd5042ed),
	.w5(32'hbd4556b2),
	.w6(32'h3da58b08),
	.w7(32'h3d5e2f38),
	.w8(32'h3d24ae07),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fc11e),
	.w1(32'hbb76b9e1),
	.w2(32'hbc2b0864),
	.w3(32'hbd06998a),
	.w4(32'hbd453e60),
	.w5(32'hbd10bae1),
	.w6(32'h3d4dd967),
	.w7(32'h3cf959ed),
	.w8(32'hbbe6310e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd39e55d),
	.w1(32'hbdb0ab14),
	.w2(32'hbd7b0edf),
	.w3(32'h3d174729),
	.w4(32'hbd04c5f5),
	.w5(32'hbd408882),
	.w6(32'h3dd9dde2),
	.w7(32'h3df283e4),
	.w8(32'hbccf3a7f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ed3a3f),
	.w1(32'hbb896cee),
	.w2(32'hbc8fa383),
	.w3(32'h3cc06110),
	.w4(32'h3d0e0c45),
	.w5(32'hbc90eea1),
	.w6(32'hbb637c8a),
	.w7(32'h3c3fa56b),
	.w8(32'h39b688ed),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac710d5),
	.w1(32'hbb050f35),
	.w2(32'hb9ba7c9b),
	.w3(32'h3b8a5a0b),
	.w4(32'h3bfb9ca7),
	.w5(32'h3b8e8c5b),
	.w6(32'hbc2db137),
	.w7(32'hbbde92b9),
	.w8(32'hb9b3a89d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3599f7),
	.w1(32'hbca9ac7a),
	.w2(32'hbd011138),
	.w3(32'h3c0c86b9),
	.w4(32'h3bd3af54),
	.w5(32'hbc02456a),
	.w6(32'hbbd29cac),
	.w7(32'hbc513d8e),
	.w8(32'hbcf8d218),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f948d),
	.w1(32'hbba2aae8),
	.w2(32'hbabc84d9),
	.w3(32'h3c994608),
	.w4(32'h3c9070cc),
	.w5(32'h3cfb6aaa),
	.w6(32'hbd11a137),
	.w7(32'hbd09d13b),
	.w8(32'h3c17d807),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac07b98),
	.w1(32'hbb089e59),
	.w2(32'hbc9e7832),
	.w3(32'hbc4276a5),
	.w4(32'hbc99bd1c),
	.w5(32'hbcbdbfd6),
	.w6(32'h3b0231a7),
	.w7(32'h3bb7865d),
	.w8(32'hbc71d814),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75c294),
	.w1(32'hbc9f1ab8),
	.w2(32'hbc87e9c7),
	.w3(32'h3adf75b8),
	.w4(32'h3b01b474),
	.w5(32'hbb45f918),
	.w6(32'hbb5b2dd2),
	.w7(32'hbc8a1211),
	.w8(32'hbccc5ccf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb3201),
	.w1(32'h3c39a0c6),
	.w2(32'hb9c71f8d),
	.w3(32'h3d32ffbd),
	.w4(32'h3da70a97),
	.w5(32'h3d51bf6c),
	.w6(32'hbd6e5835),
	.w7(32'hbd460c5b),
	.w8(32'hbca9a58f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abab390),
	.w1(32'hbc0e9eb1),
	.w2(32'hbcdb8f1d),
	.w3(32'h3cc3812f),
	.w4(32'h3cefe199),
	.w5(32'hb9c72a90),
	.w6(32'hbc594496),
	.w7(32'hbc0dc91d),
	.w8(32'hbca7d624),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2a33f),
	.w1(32'hb82653f1),
	.w2(32'h3bd24c95),
	.w3(32'h3cd1365a),
	.w4(32'h3cd5f326),
	.w5(32'h3ceb5de0),
	.w6(32'hbcc5c9b3),
	.w7(32'hbc69ce47),
	.w8(32'hbc453444),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adee729),
	.w1(32'h3a274fc4),
	.w2(32'h3b5a0589),
	.w3(32'h3c49ba7c),
	.w4(32'h3c8ef6c1),
	.w5(32'h3c5a83d2),
	.w6(32'hbc6611af),
	.w7(32'hbc0fac8f),
	.w8(32'hbc896021),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1be5a),
	.w1(32'h3c201aeb),
	.w2(32'h392fbb89),
	.w3(32'h3d39e597),
	.w4(32'h3d968017),
	.w5(32'h3d30f498),
	.w6(32'hbd286a9b),
	.w7(32'hbcc888e3),
	.w8(32'hbc2ba3b3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e07ff),
	.w1(32'hbafa1668),
	.w2(32'h3ab4b542),
	.w3(32'h3c141e4e),
	.w4(32'h3ba190f5),
	.w5(32'h3c61036f),
	.w6(32'hbc30faa0),
	.w7(32'hbc32ea74),
	.w8(32'h3c743689),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf610e4),
	.w1(32'hbc9474da),
	.w2(32'hbc328a82),
	.w3(32'hbc51da10),
	.w4(32'hbcbe38ec),
	.w5(32'hbbae1195),
	.w6(32'h3d6d711f),
	.w7(32'h3d80afac),
	.w8(32'h3d2b499a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5eee86),
	.w1(32'hbbae4a02),
	.w2(32'hbbf558fc),
	.w3(32'h3a9b62b8),
	.w4(32'hbc01cbdd),
	.w5(32'hbc57e895),
	.w6(32'h3b706c22),
	.w7(32'h3ae048c6),
	.w8(32'hbc8908ee),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebf5bf),
	.w1(32'h3b41cb02),
	.w2(32'h3b8f5566),
	.w3(32'h3c10b3d5),
	.w4(32'h3c73ec17),
	.w5(32'hbc167a38),
	.w6(32'hbc9b0e70),
	.w7(32'h3b53cf46),
	.w8(32'h3bbc9648),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3438f),
	.w1(32'hbb0745f2),
	.w2(32'hb9ecc58f),
	.w3(32'hbbc44416),
	.w4(32'hbc62b92a),
	.w5(32'hbc3b9700),
	.w6(32'h3c9d6ee3),
	.w7(32'h3c67f8f5),
	.w8(32'h3c752f91),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a2b65),
	.w1(32'hbcb3ca1d),
	.w2(32'hbc9548be),
	.w3(32'hb8f1aeba),
	.w4(32'hbcbae3d5),
	.w5(32'hbcfeb55e),
	.w6(32'h3cdc02bc),
	.w7(32'h3c91fa77),
	.w8(32'h3a249958),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e788e),
	.w1(32'hbc8f7f30),
	.w2(32'hbcb1ccd7),
	.w3(32'h3be777a2),
	.w4(32'hbc0cac11),
	.w5(32'hbc9070cb),
	.w6(32'hbb6066d8),
	.w7(32'hbbbd8cba),
	.w8(32'hbc5b6064),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d0e8a),
	.w1(32'hbab10f92),
	.w2(32'hbbaaadac),
	.w3(32'hba0a72f6),
	.w4(32'hbba5dc37),
	.w5(32'hbc29399a),
	.w6(32'hbb1a0568),
	.w7(32'h3b92b1de),
	.w8(32'h3b095b29),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f7f98),
	.w1(32'hbbe774cc),
	.w2(32'hbcb100fc),
	.w3(32'h3c11a740),
	.w4(32'hbc1f0d37),
	.w5(32'hbcd6e4a8),
	.w6(32'h3c35164a),
	.w7(32'hbb9ed32c),
	.w8(32'hbce16587),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe99287),
	.w1(32'h3aa71dd1),
	.w2(32'hbb7cdb7c),
	.w3(32'h3cde138a),
	.w4(32'h3d3805d2),
	.w5(32'h3cedb367),
	.w6(32'hbcbe2fba),
	.w7(32'hbc5a24ac),
	.w8(32'h3c19cb1c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3804faa8),
	.w1(32'hbc405dfa),
	.w2(32'hbc522d60),
	.w3(32'hbbab7707),
	.w4(32'hbc8c9830),
	.w5(32'hbccd678b),
	.w6(32'h3ca9c69f),
	.w7(32'h3c89bfc3),
	.w8(32'h3bfd0168),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cf1aa),
	.w1(32'h3b93cae7),
	.w2(32'h3b010375),
	.w3(32'hbbf2f583),
	.w4(32'h3b22a8f3),
	.w5(32'h3c031b7d),
	.w6(32'hbb2b1200),
	.w7(32'h3c1fda1e),
	.w8(32'h3cd8b059),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc868e43),
	.w1(32'hbcc4e1fb),
	.w2(32'hbbcef954),
	.w3(32'hbc84e4c3),
	.w4(32'hbd5ce232),
	.w5(32'hbd485c44),
	.w6(32'h3d4b2568),
	.w7(32'h3cfb5a61),
	.w8(32'hb9950a24),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cd5e8),
	.w1(32'hbb25a10f),
	.w2(32'h3bced1f5),
	.w3(32'hbaee66b7),
	.w4(32'h3a9d8b19),
	.w5(32'h3b3f367f),
	.w6(32'hbb0adfe0),
	.w7(32'h3bfee254),
	.w8(32'hbc795287),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e103a),
	.w1(32'hbc13e690),
	.w2(32'hbce1bf73),
	.w3(32'h3c984666),
	.w4(32'h3cd83ed8),
	.w5(32'h3c894f06),
	.w6(32'hbca534fc),
	.w7(32'hbccfff7c),
	.w8(32'hbc91b3de),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11c818),
	.w1(32'h3b969ec7),
	.w2(32'h3c2a16f7),
	.w3(32'h3c49084a),
	.w4(32'hbb98edda),
	.w5(32'hb97f279e),
	.w6(32'hb7c2842d),
	.w7(32'h3c4b11a6),
	.w8(32'h3a94a5c8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca967cf),
	.w1(32'hbcaa4e91),
	.w2(32'hbd816b65),
	.w3(32'h3c2fff8f),
	.w4(32'h3bb578af),
	.w5(32'hbcca440d),
	.w6(32'h3c35482b),
	.w7(32'hbc0e0db8),
	.w8(32'hbc5de8af),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b393c4d),
	.w1(32'hb8f6465a),
	.w2(32'hbb175ca4),
	.w3(32'hbb7dd0d0),
	.w4(32'hbbb603b6),
	.w5(32'hbadfda6c),
	.w6(32'h3bb8f237),
	.w7(32'hba02853c),
	.w8(32'hbc000af2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16847f),
	.w1(32'hbc953329),
	.w2(32'hbb91693c),
	.w3(32'hbb9b2f62),
	.w4(32'hbc7b29ef),
	.w5(32'hbcd4550e),
	.w6(32'h3c121d7e),
	.w7(32'h3c148d46),
	.w8(32'h3c5c5f07),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2deb1e),
	.w1(32'hbc00837c),
	.w2(32'hbc891e11),
	.w3(32'hbb24c27d),
	.w4(32'hbbd164eb),
	.w5(32'hbc82c90c),
	.w6(32'h3ce27608),
	.w7(32'h3c9a9699),
	.w8(32'hbbe6e6f5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd385cf),
	.w1(32'hbbec7e9f),
	.w2(32'hbb0ccef4),
	.w3(32'hbbaa8459),
	.w4(32'hbbd31c9f),
	.w5(32'hbb319526),
	.w6(32'hbc9076a3),
	.w7(32'hbb246e89),
	.w8(32'h3be06d24),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5f317),
	.w1(32'hb9431131),
	.w2(32'h3aee7b2a),
	.w3(32'h3c01ecdf),
	.w4(32'h3b3af5d7),
	.w5(32'h3bcd189f),
	.w6(32'hbb639817),
	.w7(32'hbaa41573),
	.w8(32'hbbf1ac17),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb300689),
	.w1(32'hbba70172),
	.w2(32'hbbfb4744),
	.w3(32'hbb35f200),
	.w4(32'hbbde53fa),
	.w5(32'hbb3a5ee9),
	.w6(32'hbba823d2),
	.w7(32'hbbdcff5e),
	.w8(32'h3c2b83c7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2eba44),
	.w1(32'hbcc1ed10),
	.w2(32'hbcdbce32),
	.w3(32'hbc2c590e),
	.w4(32'hbc99a5fe),
	.w5(32'hbc8f405e),
	.w6(32'h3d0c4be0),
	.w7(32'h3ce795b1),
	.w8(32'h3c1f08a5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83291c),
	.w1(32'h3bd7080d),
	.w2(32'h3a9e6048),
	.w3(32'hbc0b6a7f),
	.w4(32'hbc8555ff),
	.w5(32'hbc8b1466),
	.w6(32'hbc0ae45b),
	.w7(32'hbb004fe0),
	.w8(32'h3b339983),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c991d),
	.w1(32'h3b2f2d57),
	.w2(32'h3709fdd4),
	.w3(32'hbb1718e8),
	.w4(32'hbbdfa347),
	.w5(32'hbb94330a),
	.w6(32'h3c080975),
	.w7(32'h3b4f46b3),
	.w8(32'h3bb16ea8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e0636e),
	.w1(32'hbbaf87ce),
	.w2(32'hbb9e531a),
	.w3(32'hba00421e),
	.w4(32'hbbbafa6b),
	.w5(32'hbbe5ccb4),
	.w6(32'h3c387467),
	.w7(32'h3c132754),
	.w8(32'h3b972e7f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15b43e),
	.w1(32'h3b9476d7),
	.w2(32'h3bb594a5),
	.w3(32'hbba814f9),
	.w4(32'hbb6efa0f),
	.w5(32'hba6d4a80),
	.w6(32'h3c0fe3af),
	.w7(32'h3c170d6e),
	.w8(32'h3a26fe9f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ada06),
	.w1(32'hbc3947bb),
	.w2(32'hbcc7bbaf),
	.w3(32'h3c007de8),
	.w4(32'h3bedb977),
	.w5(32'h3bad106e),
	.w6(32'h3ac85c81),
	.w7(32'hb9f1f903),
	.w8(32'h3c3ac2d4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af59915),
	.w1(32'hb93f8dcc),
	.w2(32'hba879fcd),
	.w3(32'hbb864c3a),
	.w4(32'hbc155a26),
	.w5(32'hbbe30b72),
	.w6(32'h3c111257),
	.w7(32'h3b64c7ba),
	.w8(32'h3d47f8e7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20d354),
	.w1(32'hbc0fbb80),
	.w2(32'hbc61ade6),
	.w3(32'hbd18227a),
	.w4(32'hbd57eb1b),
	.w5(32'hbd83e1e0),
	.w6(32'h3da4a4a4),
	.w7(32'h3d87eb66),
	.w8(32'h3c1771d6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c258e9),
	.w1(32'hbaaf26fe),
	.w2(32'hbb1e4ba2),
	.w3(32'hbb66d0c1),
	.w4(32'hbbfdf642),
	.w5(32'hbb9cc41f),
	.w6(32'h3b824d6b),
	.w7(32'h39e736f1),
	.w8(32'h3bbeef0c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c219189),
	.w1(32'h3b129a1b),
	.w2(32'hbabec70f),
	.w3(32'h3b1c5926),
	.w4(32'hbc0ed170),
	.w5(32'hbc03e41d),
	.w6(32'h3c704509),
	.w7(32'h3bfb86b5),
	.w8(32'h3c049549),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa05075),
	.w1(32'hbadb3e76),
	.w2(32'hbabedc32),
	.w3(32'hbb83e351),
	.w4(32'hbc2c3ab7),
	.w5(32'hbbcd4bde),
	.w6(32'h3bdac0bd),
	.w7(32'h3b50e593),
	.w8(32'hbaa83f51),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3881e8),
	.w1(32'hbccbd997),
	.w2(32'hbcd222ec),
	.w3(32'hbbbc3916),
	.w4(32'hbbaa358e),
	.w5(32'hbb4a0bdf),
	.w6(32'hbbcf010d),
	.w7(32'hba8164bd),
	.w8(32'hbab015c0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bfd6a),
	.w1(32'hbb9c2124),
	.w2(32'hbba577dd),
	.w3(32'hbbc420ff),
	.w4(32'hbc438a1d),
	.w5(32'hbc241cb8),
	.w6(32'h3a932a10),
	.w7(32'hbb0a1c58),
	.w8(32'h3b80b305),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f1e25),
	.w1(32'hbb2ed598),
	.w2(32'hbb77db0c),
	.w3(32'hbba38511),
	.w4(32'hbc27abc7),
	.w5(32'hbc2e48a8),
	.w6(32'h3c5bf120),
	.w7(32'h3c0bdb70),
	.w8(32'h39cd04ac),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae73cc4),
	.w1(32'hbb899f1e),
	.w2(32'hbb74aa32),
	.w3(32'hbba6d427),
	.w4(32'hbc227118),
	.w5(32'hbbcd5f2d),
	.w6(32'h3a32b6b7),
	.w7(32'hbaaf8ea3),
	.w8(32'h3d652e39),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39df27),
	.w1(32'hbcaef80d),
	.w2(32'hbcdfb551),
	.w3(32'hbcdfcffe),
	.w4(32'hbd438d67),
	.w5(32'hbd501eef),
	.w6(32'h3dd23699),
	.w7(32'h3d953842),
	.w8(32'h3d3a1de0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88e91b),
	.w1(32'hbc8b8acb),
	.w2(32'hbd18aafb),
	.w3(32'hbc9d0440),
	.w4(32'hbd28c34f),
	.w5(32'hbd34bdd5),
	.w6(32'h3d139c92),
	.w7(32'h3bcee161),
	.w8(32'hbc585330),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979aad0),
	.w1(32'hb8eec2f0),
	.w2(32'h3ad3fe5a),
	.w3(32'hba922805),
	.w4(32'hbb1e3748),
	.w5(32'h3aa9d2be),
	.w6(32'h3ba4057f),
	.w7(32'h3b2d65dc),
	.w8(32'h3b77a88f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfe154),
	.w1(32'h3b0de3da),
	.w2(32'hbb2d1c2d),
	.w3(32'hbbc3e66a),
	.w4(32'h3b23f02d),
	.w5(32'hbb874aec),
	.w6(32'h3beff88e),
	.w7(32'h3be303c3),
	.w8(32'hbab278c2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7bd88),
	.w1(32'hbb7d8a9a),
	.w2(32'h3c35511e),
	.w3(32'h3a5032b4),
	.w4(32'hbc2ad1cc),
	.w5(32'hbbc53954),
	.w6(32'hbb411644),
	.w7(32'hbbd1c83e),
	.w8(32'h3a95deb9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf75b4),
	.w1(32'hbc13e399),
	.w2(32'hbbca1d6d),
	.w3(32'h3bbc4754),
	.w4(32'hbbac463c),
	.w5(32'hbbbacaaf),
	.w6(32'h3cff31bf),
	.w7(32'h3ce7325e),
	.w8(32'h3ca0dc66),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1dec19),
	.w1(32'hbcc034bb),
	.w2(32'hbd1012a5),
	.w3(32'hbd44146f),
	.w4(32'hbce3605b),
	.w5(32'hbbbf9d02),
	.w6(32'h3c0c70ba),
	.w7(32'h3cd77aef),
	.w8(32'h3c693980),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57c149),
	.w1(32'hbcb76f5f),
	.w2(32'hbcb004ae),
	.w3(32'h3ceb317c),
	.w4(32'h3c66abc7),
	.w5(32'h39fb6833),
	.w6(32'h3c811006),
	.w7(32'h3c8d8c7f),
	.w8(32'h3d0cca74),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cf354),
	.w1(32'hbc8f3c6f),
	.w2(32'h3a770e52),
	.w3(32'hbbaf7a38),
	.w4(32'hbcdc9987),
	.w5(32'hbcafbaf0),
	.w6(32'h3cb99372),
	.w7(32'h3c0a9055),
	.w8(32'hbcfabbd2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2800b7),
	.w1(32'h3b12c7b3),
	.w2(32'hbba7e70c),
	.w3(32'h3d0a9de0),
	.w4(32'h3d6d7a51),
	.w5(32'h3d1edcf8),
	.w6(32'hbd057904),
	.w7(32'hbcbbb033),
	.w8(32'h3b56c542),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c598d),
	.w1(32'h3b0c60b7),
	.w2(32'h39d6b271),
	.w3(32'hbb1442c9),
	.w4(32'hbbd0bf88),
	.w5(32'h3a910308),
	.w6(32'h3bfebd20),
	.w7(32'h3abc0536),
	.w8(32'hbc1558da),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb183827),
	.w1(32'hba2be08a),
	.w2(32'hbada972e),
	.w3(32'hbaa84024),
	.w4(32'h3c0e4571),
	.w5(32'h3a5b47a5),
	.w6(32'hbc7a7f43),
	.w7(32'hbbbe92ea),
	.w8(32'hbceaf149),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6911a),
	.w1(32'h3b5831ec),
	.w2(32'hbba30a5c),
	.w3(32'h3d0933c2),
	.w4(32'h3d5a8898),
	.w5(32'h3d0d3910),
	.w6(32'hbcdae2eb),
	.w7(32'hbca1f2c5),
	.w8(32'hbcc715b8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84bc51),
	.w1(32'hbc08d463),
	.w2(32'hbc1770bc),
	.w3(32'h3cc394d6),
	.w4(32'h3d265b71),
	.w5(32'h3ce5d481),
	.w6(32'hbcc48bdf),
	.w7(32'hbc82de86),
	.w8(32'hbc968690),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2250ac),
	.w1(32'h3aad254a),
	.w2(32'hbb1678bd),
	.w3(32'h3c67bec8),
	.w4(32'h3cbbc3c3),
	.w5(32'h3c4bcd4a),
	.w6(32'hbc935303),
	.w7(32'hbc7b9842),
	.w8(32'h3c102b6b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac61ac),
	.w1(32'h3c520bd3),
	.w2(32'h3ccbf583),
	.w3(32'hbc2884fb),
	.w4(32'hbbaa77bd),
	.w5(32'h3c5999df),
	.w6(32'hbba9bb61),
	.w7(32'hbc3a2e9b),
	.w8(32'h3c0682cb),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a871d38),
	.w1(32'hbbb9182a),
	.w2(32'hbbdb02fd),
	.w3(32'h3b05ed1c),
	.w4(32'hbbbf84dd),
	.w5(32'hbc021e72),
	.w6(32'h3c74eeb7),
	.w7(32'h3c3ad78d),
	.w8(32'hbc645f24),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad22747),
	.w1(32'hbc028d2e),
	.w2(32'hbc74e07a),
	.w3(32'hbc2e88ab),
	.w4(32'hbc26148d),
	.w5(32'hbc52c4fc),
	.w6(32'hbc8794e1),
	.w7(32'hbca2b307),
	.w8(32'hbd0449bc),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac583c2),
	.w1(32'h3aa2bd3a),
	.w2(32'hbc1b1cea),
	.w3(32'h3ce9abb2),
	.w4(32'h3cfe77c6),
	.w5(32'h3c0bae03),
	.w6(32'hbcce3261),
	.w7(32'hbc68e424),
	.w8(32'hbca26830),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c1329),
	.w1(32'hbc7a5a7f),
	.w2(32'hbc843ca9),
	.w3(32'h3b1f80bb),
	.w4(32'h3ae6d778),
	.w5(32'h3b0990d7),
	.w6(32'h3c4f4189),
	.w7(32'h3a6060f5),
	.w8(32'h3c442e30),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a66bfb),
	.w1(32'h3af3c411),
	.w2(32'hbb708696),
	.w3(32'hbc3fcea3),
	.w4(32'hbc6e956a),
	.w5(32'hbc576786),
	.w6(32'hbacb6ea0),
	.w7(32'hba99dd87),
	.w8(32'h3d48346b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf32743),
	.w1(32'hbb934a46),
	.w2(32'hbc570905),
	.w3(32'hbd08222f),
	.w4(32'hbd371d02),
	.w5(32'hbd133940),
	.w6(32'h3d88cc69),
	.w7(32'h3d243270),
	.w8(32'h3b89bd00),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38943386),
	.w1(32'h3a0753ed),
	.w2(32'h3a5a0023),
	.w3(32'hbb7c0192),
	.w4(32'hbc097328),
	.w5(32'hbabf28d2),
	.w6(32'h3c05f926),
	.w7(32'h3b617bb3),
	.w8(32'hbc6b59cc),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb902fda),
	.w1(32'hbb47035f),
	.w2(32'hbb12bfb3),
	.w3(32'h3bc2656d),
	.w4(32'h3c58aca1),
	.w5(32'h3b12bfcb),
	.w6(32'hbc9878ae),
	.w7(32'hbbf4cd51),
	.w8(32'h3bb3ab5f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61392b),
	.w1(32'h3a2b7bda),
	.w2(32'h3a982343),
	.w3(32'hbb430405),
	.w4(32'hbbe3efac),
	.w5(32'hbba6cc05),
	.w6(32'h3bb5bc3f),
	.w7(32'h3b0bc18b),
	.w8(32'h3d22f382),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc553d2),
	.w1(32'hbbbaaafc),
	.w2(32'hbc327ff5),
	.w3(32'hbd0dab9c),
	.w4(32'hbd56b87c),
	.w5(32'hbd160697),
	.w6(32'h3d8061b0),
	.w7(32'h3d04faff),
	.w8(32'hbca3ba0f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe4605),
	.w1(32'h3ab2e724),
	.w2(32'h3c119161),
	.w3(32'h3c1488b7),
	.w4(32'h3ca00fef),
	.w5(32'h3cb43190),
	.w6(32'hbcd5fcc3),
	.w7(32'hbcea4365),
	.w8(32'hbcacf6c5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac043a9),
	.w1(32'h3b96a7e0),
	.w2(32'h3aa91ff7),
	.w3(32'h3c404064),
	.w4(32'h3cba257f),
	.w5(32'h3c7c2f3d),
	.w6(32'hbca758e1),
	.w7(32'hbc817bfb),
	.w8(32'hbbd8aa0d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf143fc),
	.w1(32'hbc665970),
	.w2(32'hbc0c7cdb),
	.w3(32'hbbb6fe72),
	.w4(32'hbc5979cb),
	.w5(32'hbc9cf15c),
	.w6(32'h3bdfee59),
	.w7(32'h3c17be92),
	.w8(32'hbb80695c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5dc8f0),
	.w1(32'hbb28d29a),
	.w2(32'h39db3c2e),
	.w3(32'h3ab29ca8),
	.w4(32'h3a8384d7),
	.w5(32'hbaaefddf),
	.w6(32'h3b917e67),
	.w7(32'h3a2d1621),
	.w8(32'hba528bae),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4c8c5),
	.w1(32'h3bc58ae9),
	.w2(32'h3bbdc8aa),
	.w3(32'hbbf151aa),
	.w4(32'hbb34291a),
	.w5(32'hbacd4ab9),
	.w6(32'hbbdbc20c),
	.w7(32'hbb841d35),
	.w8(32'hbb738057),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b93ba),
	.w1(32'h3a9bdee3),
	.w2(32'h3ae8a9fe),
	.w3(32'hbbbb7917),
	.w4(32'hbb6c506e),
	.w5(32'hb97ccebc),
	.w6(32'hbbc85d98),
	.w7(32'hbbbada3c),
	.w8(32'hba2101e3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe34a0),
	.w1(32'h3ac56569),
	.w2(32'h3bd77799),
	.w3(32'h3b7a7bad),
	.w4(32'h3b988ebf),
	.w5(32'h3be32c78),
	.w6(32'h3bec1122),
	.w7(32'h3b9bf1d9),
	.w8(32'hba3fae98),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81b8a4),
	.w1(32'h3a0dd892),
	.w2(32'hbc5345ff),
	.w3(32'h3aebba18),
	.w4(32'h3c0fcb7d),
	.w5(32'hb7867e00),
	.w6(32'hbbebc645),
	.w7(32'h3b00f40a),
	.w8(32'h3be4d1fc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd84dcd),
	.w1(32'hbb2575e7),
	.w2(32'h3a47bad2),
	.w3(32'hbbb80f10),
	.w4(32'h3aecaa50),
	.w5(32'h3b9fdfc6),
	.w6(32'h3afe447e),
	.w7(32'h3b3ee130),
	.w8(32'h3b143e13),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60bfc1),
	.w1(32'h3bd9d5c8),
	.w2(32'h3c05248a),
	.w3(32'hbb57fbb8),
	.w4(32'h39b310f8),
	.w5(32'h3b06eb19),
	.w6(32'hbc1bd6d6),
	.w7(32'hbbba0e5b),
	.w8(32'hbb9b225a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba288500),
	.w1(32'h3aa80367),
	.w2(32'h3b1a14e4),
	.w3(32'hbb234dcd),
	.w4(32'hb9a5e648),
	.w5(32'h3b6dfd24),
	.w6(32'h38c35277),
	.w7(32'h3b038a99),
	.w8(32'hba916cbb),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78c72b),
	.w1(32'hba4cf7df),
	.w2(32'hbb2d75d4),
	.w3(32'h3b205561),
	.w4(32'hbb1ea53b),
	.w5(32'hbbba5d60),
	.w6(32'h3aaed169),
	.w7(32'h3a724b64),
	.w8(32'hbc185df4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20a300),
	.w1(32'hbb1b2844),
	.w2(32'h3b263a96),
	.w3(32'hba97d37c),
	.w4(32'hbb159bfe),
	.w5(32'hb994e228),
	.w6(32'hbab35e5a),
	.w7(32'h3b2ea7c5),
	.w8(32'hbb3c55bf),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6020c0),
	.w1(32'h3ae491c5),
	.w2(32'hbbf3215a),
	.w3(32'h3949be54),
	.w4(32'h3b8ace28),
	.w5(32'hbc0530c3),
	.w6(32'hba8cc063),
	.w7(32'hbb7bd8ec),
	.w8(32'hbaa71cb7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b047d17),
	.w1(32'hbb6ba2f9),
	.w2(32'hbc1b9e07),
	.w3(32'h3ad5ae15),
	.w4(32'hbb2400c1),
	.w5(32'hbc2ed380),
	.w6(32'h3c4e9a48),
	.w7(32'h3c485bcb),
	.w8(32'h3c174478),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e21d34),
	.w1(32'hba7b5f29),
	.w2(32'hbc0c9704),
	.w3(32'hba7c2c2d),
	.w4(32'h3b411c0e),
	.w5(32'hbbb99ad5),
	.w6(32'hba33cec3),
	.w7(32'hbbfedb24),
	.w8(32'hbb575e54),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c0486),
	.w1(32'hbb9672e0),
	.w2(32'hbba16928),
	.w3(32'hba7fa731),
	.w4(32'hbb523b54),
	.w5(32'hbb540810),
	.w6(32'hbb92e1a2),
	.w7(32'hbb3144db),
	.w8(32'hbae19744),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09cc8e),
	.w1(32'h3a83bd0a),
	.w2(32'hbb914da8),
	.w3(32'hbad8f5d4),
	.w4(32'hbc6c00f8),
	.w5(32'hbc27d874),
	.w6(32'hbbd47bcc),
	.w7(32'hbc5501a5),
	.w8(32'hbc6a05af),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc086a59),
	.w1(32'hbbfef02d),
	.w2(32'hbc0a91b4),
	.w3(32'h3b0840e1),
	.w4(32'h3a8d7ec6),
	.w5(32'h3a540fea),
	.w6(32'h3bd54801),
	.w7(32'hbb29b095),
	.w8(32'h3bcb5c92),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39500c0e),
	.w1(32'hb909561d),
	.w2(32'h3b1cdff3),
	.w3(32'h3a5d8809),
	.w4(32'h3a1c2ff2),
	.w5(32'h3b3ce120),
	.w6(32'h3ad97bcb),
	.w7(32'h3b80271d),
	.w8(32'hbb87a7a9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb751468),
	.w1(32'hbb5fbefb),
	.w2(32'hbb594fbe),
	.w3(32'hbbc38b0f),
	.w4(32'hbbaa5980),
	.w5(32'hbbb48198),
	.w6(32'hbbea0043),
	.w7(32'hbbd34e35),
	.w8(32'h3b9934eb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39984004),
	.w1(32'hbb6fb340),
	.w2(32'h3b2011a2),
	.w3(32'h3bbce6e1),
	.w4(32'h3bd6661a),
	.w5(32'h3b548216),
	.w6(32'h3b1f699d),
	.w7(32'h3a549d46),
	.w8(32'h3b6bc1b4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf74ff),
	.w1(32'h3bef16f2),
	.w2(32'h3aa4f730),
	.w3(32'hbb0e0626),
	.w4(32'h3b948381),
	.w5(32'h3b19f04e),
	.w6(32'hbb435ac1),
	.w7(32'h3b1e7d14),
	.w8(32'hbb0a7ffa),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25e609),
	.w1(32'hbb9a717d),
	.w2(32'hbbcfa622),
	.w3(32'h3b41959e),
	.w4(32'h3896d307),
	.w5(32'hb9facc6e),
	.w6(32'h3b5b19a0),
	.w7(32'h3ba3ef18),
	.w8(32'hbb3fcfe5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9cbe5),
	.w1(32'hbb71d758),
	.w2(32'hbc0310a6),
	.w3(32'h3bb9afa1),
	.w4(32'h3aba668d),
	.w5(32'hbc828a1b),
	.w6(32'h3afe1a38),
	.w7(32'hbb1b59f0),
	.w8(32'hbc474d05),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule