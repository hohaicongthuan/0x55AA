module layer_10_featuremap_266(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad113fe),
	.w1(32'hbc12c3bd),
	.w2(32'hbb759e08),
	.w3(32'hbc028341),
	.w4(32'hbbbb0474),
	.w5(32'h3b040098),
	.w6(32'hbc218a01),
	.w7(32'hbbe8e452),
	.w8(32'h37ed6762),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81c476),
	.w1(32'hbac38e08),
	.w2(32'hbb3414f3),
	.w3(32'h3bb9c2a4),
	.w4(32'hb98893be),
	.w5(32'hbc1348f6),
	.w6(32'h3ac680d4),
	.w7(32'hbb813760),
	.w8(32'hbc45fb99),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e0de6),
	.w1(32'h3c1b7958),
	.w2(32'h3b79e676),
	.w3(32'h3bef0eac),
	.w4(32'h3b87ccf9),
	.w5(32'h39a97ecb),
	.w6(32'h3c13ef65),
	.w7(32'h3c6d7bf7),
	.w8(32'hbb6f0882),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabaf88),
	.w1(32'hbb928476),
	.w2(32'hbb1bf45b),
	.w3(32'h3a1db11e),
	.w4(32'h3a940050),
	.w5(32'hbb9e8e6c),
	.w6(32'hbaf3c61a),
	.w7(32'hb9eeb755),
	.w8(32'hbb48a168),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6d49f),
	.w1(32'h3b356776),
	.w2(32'hbb0e5913),
	.w3(32'hbb04a292),
	.w4(32'hbb0c6c2a),
	.w5(32'h39c5503f),
	.w6(32'h3c0aa4f8),
	.w7(32'hba5a299c),
	.w8(32'h3a8092d3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb099390),
	.w1(32'hbb0b99c6),
	.w2(32'h39c198cd),
	.w3(32'h3a6bca70),
	.w4(32'h3b3b5ee5),
	.w5(32'h3b28ec2f),
	.w6(32'h390b8d65),
	.w7(32'h3b858207),
	.w8(32'h3a1eba0f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb925865),
	.w1(32'h3b80b671),
	.w2(32'hbb3931bf),
	.w3(32'h3bf8eb23),
	.w4(32'hbb938d80),
	.w5(32'hbc7116ec),
	.w6(32'h3c3001bc),
	.w7(32'hb9bb77d4),
	.w8(32'hbc3b5d64),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82e00d),
	.w1(32'hbc7ae76c),
	.w2(32'h3b8f4059),
	.w3(32'hbc20efb9),
	.w4(32'hbc248634),
	.w5(32'h3bd668be),
	.w6(32'hbb2b860c),
	.w7(32'h39950e20),
	.w8(32'h39ceab0b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5bf55),
	.w1(32'h3a04bc17),
	.w2(32'h3a1d439e),
	.w3(32'h3ada4b07),
	.w4(32'h39827ba0),
	.w5(32'h3a00889f),
	.w6(32'hba161d90),
	.w7(32'hba51b2a7),
	.w8(32'h3aab6c57),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca576e),
	.w1(32'hbb0782e2),
	.w2(32'h3b0d49e5),
	.w3(32'hbc120857),
	.w4(32'hbb4456fb),
	.w5(32'h3a9a5fce),
	.w6(32'hbbbce8f4),
	.w7(32'hb8ffef80),
	.w8(32'h3bc4a426),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3391a),
	.w1(32'hbb9716ab),
	.w2(32'h3b21cfb3),
	.w3(32'hbb4f1128),
	.w4(32'hba2a3ae0),
	.w5(32'hbb22df2b),
	.w6(32'hb9b09f07),
	.w7(32'h3b0d4921),
	.w8(32'h3c744b83),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04d976),
	.w1(32'h3b63c4b8),
	.w2(32'h3c70ff43),
	.w3(32'h3bafc15e),
	.w4(32'hb9f4ff7d),
	.w5(32'hbbbe9651),
	.w6(32'h3ac7201a),
	.w7(32'h3b365234),
	.w8(32'hb9d719ea),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7fb7d),
	.w1(32'h3c02a05e),
	.w2(32'h3b203f2e),
	.w3(32'h3a0569cb),
	.w4(32'hbb96550c),
	.w5(32'hbc461e44),
	.w6(32'h3c106928),
	.w7(32'h3b41326c),
	.w8(32'hbbd0659c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d9165),
	.w1(32'hbc435df3),
	.w2(32'h3a0363f6),
	.w3(32'hbc44ba5e),
	.w4(32'h3c2de478),
	.w5(32'hbbb52a36),
	.w6(32'h3acf9911),
	.w7(32'h3b2de594),
	.w8(32'hbb6521c2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3db73),
	.w1(32'h3b932533),
	.w2(32'h3bae7ab5),
	.w3(32'hbb22a803),
	.w4(32'h3a518588),
	.w5(32'hba68d908),
	.w6(32'hbb3bc158),
	.w7(32'hbaf14973),
	.w8(32'h3abd4388),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf23e4d),
	.w1(32'hbc1c381e),
	.w2(32'hbc01de4a),
	.w3(32'hbc207db4),
	.w4(32'hbba663b2),
	.w5(32'hbb1741cd),
	.w6(32'hbba2f1b0),
	.w7(32'hbc0877c7),
	.w8(32'h3986a619),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813c79),
	.w1(32'h3bd3aeba),
	.w2(32'h3b5b3394),
	.w3(32'h3b86f987),
	.w4(32'h3b3320df),
	.w5(32'hbb744236),
	.w6(32'h3b4484db),
	.w7(32'h3ac0d781),
	.w8(32'hbb213b27),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde10e4),
	.w1(32'h3a80e522),
	.w2(32'hbac95964),
	.w3(32'h39be5ea9),
	.w4(32'hbb59b070),
	.w5(32'hbc30705b),
	.w6(32'h3aa7d263),
	.w7(32'h3bf0c685),
	.w8(32'hbb7c86d6),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47b82e),
	.w1(32'hbb079fb9),
	.w2(32'h3b200219),
	.w3(32'hbb8e3d4b),
	.w4(32'hbb7ff047),
	.w5(32'h3cb474ef),
	.w6(32'hbbb2961e),
	.w7(32'h3bd1190b),
	.w8(32'h3cce71b5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc195d5),
	.w1(32'h3c287895),
	.w2(32'h3c4aba17),
	.w3(32'h3bd50002),
	.w4(32'h3a9be273),
	.w5(32'hbbe3b60d),
	.w6(32'h3c34831c),
	.w7(32'h3c73bf0e),
	.w8(32'hbc1a107d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaad0ea),
	.w1(32'hbba6ae46),
	.w2(32'hbb0b21e5),
	.w3(32'h3a6e2178),
	.w4(32'h3b1e5168),
	.w5(32'h3b251205),
	.w6(32'h3c1df89c),
	.w7(32'hba47f72d),
	.w8(32'hba9b296e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbc810),
	.w1(32'hba7341f8),
	.w2(32'h3b02e2e7),
	.w3(32'h3a8ce885),
	.w4(32'h3b73f2ee),
	.w5(32'h3a4f228d),
	.w6(32'hbb87e2f8),
	.w7(32'h3a10b123),
	.w8(32'h3b3f8236),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98012e8),
	.w1(32'h3b99d218),
	.w2(32'h3a84da48),
	.w3(32'h38c48b65),
	.w4(32'hbb5c55f7),
	.w5(32'hbc79ba80),
	.w6(32'h3c0c4a8c),
	.w7(32'hbb393666),
	.w8(32'hbbd3c912),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1388cc),
	.w1(32'hbbe3abc6),
	.w2(32'h3a4a5f12),
	.w3(32'hbbecd96a),
	.w4(32'hbb8c43d2),
	.w5(32'h39a3f322),
	.w6(32'h3a06a7ed),
	.w7(32'h3b792336),
	.w8(32'h3aa7ca41),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7daff1),
	.w1(32'hbae77324),
	.w2(32'hba3f4806),
	.w3(32'h3c6ebe54),
	.w4(32'hbb7a4aaf),
	.w5(32'h3bab10b9),
	.w6(32'h3c005394),
	.w7(32'h3b32aad6),
	.w8(32'h3b02bbd7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d5f84),
	.w1(32'hbb428220),
	.w2(32'h3b49cd2f),
	.w3(32'hbb061655),
	.w4(32'h3a0b161f),
	.w5(32'h3789214e),
	.w6(32'hbc21d260),
	.w7(32'hb9a23124),
	.w8(32'hbb7c47ad),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabf164),
	.w1(32'h3c4b5168),
	.w2(32'h3a50bd9c),
	.w3(32'h3c1de70d),
	.w4(32'hba7cbf16),
	.w5(32'h3b0a35cd),
	.w6(32'h3c21e976),
	.w7(32'hbaa676e1),
	.w8(32'h3aace817),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b570f85),
	.w1(32'hba76a573),
	.w2(32'hbbf36e3b),
	.w3(32'h3ae127f1),
	.w4(32'hbc10f63b),
	.w5(32'hbc6fdc38),
	.w6(32'h3b340455),
	.w7(32'hbc2368f2),
	.w8(32'hbc02121a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c047be4),
	.w1(32'hbc581d68),
	.w2(32'hbc42c5f0),
	.w3(32'hbc1b5d79),
	.w4(32'h3c0f7ac9),
	.w5(32'h3ab4a94e),
	.w6(32'hbbf6c7aa),
	.w7(32'hbc1e18e2),
	.w8(32'h3b2b11a1),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab33be6),
	.w1(32'h3c6fa7c3),
	.w2(32'h3c3a4a87),
	.w3(32'hbbb7895d),
	.w4(32'hbb4a10ec),
	.w5(32'hbba9ba6d),
	.w6(32'hba47e053),
	.w7(32'h3b2065ce),
	.w8(32'hbb1578a6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c344b),
	.w1(32'hbbb50503),
	.w2(32'hbb0a4404),
	.w3(32'h3b7e837a),
	.w4(32'hba8ada91),
	.w5(32'hbbb62d75),
	.w6(32'hba23a56e),
	.w7(32'h3b8358d2),
	.w8(32'h3baec634),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968f267),
	.w1(32'h3bef8bbf),
	.w2(32'h3bfbab0b),
	.w3(32'hbbfcfc16),
	.w4(32'hbb472af4),
	.w5(32'h3c0342e1),
	.w6(32'h3ba168c0),
	.w7(32'hbb465a20),
	.w8(32'h3d01baa2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca713cc),
	.w1(32'hbc4dbb6e),
	.w2(32'h3b235b69),
	.w3(32'h3b1ca22c),
	.w4(32'h3b190eaf),
	.w5(32'hbbf00a42),
	.w6(32'hbb7932d8),
	.w7(32'h3b733224),
	.w8(32'h3a98e0cd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb178c1e),
	.w1(32'hbbb7b00d),
	.w2(32'hbc2242d8),
	.w3(32'hbb2ee970),
	.w4(32'h3a802e3a),
	.w5(32'hbb07fc01),
	.w6(32'hbc3ba47a),
	.w7(32'hba44e2ed),
	.w8(32'hbbf54f29),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b1d93),
	.w1(32'hbb14ff87),
	.w2(32'hbc15463e),
	.w3(32'hbb701410),
	.w4(32'hbbf9d69e),
	.w5(32'hbc0080ad),
	.w6(32'h3b4012e8),
	.w7(32'hbc3a39c8),
	.w8(32'hbc20a1f4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae81c65),
	.w1(32'h3b82e81c),
	.w2(32'h3b8437eb),
	.w3(32'h3c36e4b0),
	.w4(32'h3b575bd7),
	.w5(32'hbacfc499),
	.w6(32'h3c320264),
	.w7(32'h3ba1af54),
	.w8(32'h3b0426ea),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02fcd9),
	.w1(32'hbb903032),
	.w2(32'h3c7077b6),
	.w3(32'h3c51906e),
	.w4(32'h3c98cf96),
	.w5(32'hbbeba6bc),
	.w6(32'h3b604a4b),
	.w7(32'h3be9cdf4),
	.w8(32'hbc71ecae),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba90808),
	.w1(32'hbbd4e224),
	.w2(32'h3b39311e),
	.w3(32'hbb4a0736),
	.w4(32'h39be1ebf),
	.w5(32'h3a5ec5ff),
	.w6(32'hbc2cb2f9),
	.w7(32'hbc11f91d),
	.w8(32'hbc0a545f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfebdf),
	.w1(32'hbb81d74f),
	.w2(32'h39f82523),
	.w3(32'h3c1693d0),
	.w4(32'hbae19112),
	.w5(32'h3a9b6e3f),
	.w6(32'h3bc49926),
	.w7(32'hbb1d4b56),
	.w8(32'hbc036111),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398302f8),
	.w1(32'h3a103f30),
	.w2(32'h39d650a9),
	.w3(32'h3b359304),
	.w4(32'h3ba45764),
	.w5(32'h3b6162d3),
	.w6(32'h39184a72),
	.w7(32'h3b523851),
	.w8(32'h3c6adb0a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c480714),
	.w1(32'hbb7ffe98),
	.w2(32'h3bbfb94b),
	.w3(32'hbb28f022),
	.w4(32'h3c96fec1),
	.w5(32'h3b1c79aa),
	.w6(32'hbb145d70),
	.w7(32'h3c907953),
	.w8(32'h38f9ed49),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cb1a2),
	.w1(32'hbb11de88),
	.w2(32'h3b26e3a0),
	.w3(32'hbaedd8ec),
	.w4(32'h3b48d3c8),
	.w5(32'h3a9c5555),
	.w6(32'hbb8ba4c9),
	.w7(32'h3b492acd),
	.w8(32'hbb439cf0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9eff9),
	.w1(32'hbc3db2ff),
	.w2(32'hbbea9376),
	.w3(32'hbbdcea06),
	.w4(32'hbadc3878),
	.w5(32'hbc2753cb),
	.w6(32'hbbde790a),
	.w7(32'hba56cc21),
	.w8(32'hb9c06024),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91e7ee),
	.w1(32'h3b9d2a9e),
	.w2(32'hbbe27616),
	.w3(32'hbbabcc23),
	.w4(32'h3aa4d9ff),
	.w5(32'hbbcae9cb),
	.w6(32'h3b23c8dd),
	.w7(32'h3b81fbe7),
	.w8(32'h3a8ff1a3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4243ef),
	.w1(32'hb883aa99),
	.w2(32'hbb6b8730),
	.w3(32'hbb41b610),
	.w4(32'h3b27558d),
	.w5(32'h3c01c3a3),
	.w6(32'hba4d6796),
	.w7(32'h3b216935),
	.w8(32'h3af14301),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4be4e9),
	.w1(32'h3ad5e90a),
	.w2(32'h3c075256),
	.w3(32'h3bdf3bd4),
	.w4(32'h3b5f59d5),
	.w5(32'h3ae5b060),
	.w6(32'h3b6c32f8),
	.w7(32'h3bc1f78d),
	.w8(32'h3a86e08f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c8a39),
	.w1(32'h3b76cd20),
	.w2(32'hbaddd290),
	.w3(32'h3a8e722a),
	.w4(32'hba86e598),
	.w5(32'hb9c1b0d0),
	.w6(32'h392469b2),
	.w7(32'hba2d84e4),
	.w8(32'hbabb0e8d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab19e3),
	.w1(32'hbb5798d2),
	.w2(32'hbb60dbd8),
	.w3(32'hbb08a258),
	.w4(32'hbb3dca6d),
	.w5(32'hbbda54fb),
	.w6(32'hbb5c0f90),
	.w7(32'hba54942e),
	.w8(32'h3b24d0ab),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e119aa),
	.w1(32'hbae00b76),
	.w2(32'hbb94b39b),
	.w3(32'h3b2a1be1),
	.w4(32'h3ade3b60),
	.w5(32'hbb0a7952),
	.w6(32'hbb70c0d8),
	.w7(32'hba02ff68),
	.w8(32'hbb7908e6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb432390),
	.w1(32'hba9f5b9c),
	.w2(32'hbae308ad),
	.w3(32'hbae6931c),
	.w4(32'h3b388891),
	.w5(32'hbc16c82e),
	.w6(32'hbbf09c6a),
	.w7(32'hbb1ce7a1),
	.w8(32'hbc64c981),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17193c),
	.w1(32'h3c756f05),
	.w2(32'hba857232),
	.w3(32'h3ccf1da8),
	.w4(32'hb9b98f4d),
	.w5(32'h3b30bb78),
	.w6(32'h3cea0b37),
	.w7(32'hbb4b0a2a),
	.w8(32'hba1f982f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ba39d),
	.w1(32'h3afa3256),
	.w2(32'h3b9b59c7),
	.w3(32'hba8890da),
	.w4(32'hbb5d6a71),
	.w5(32'hbbdcb6c1),
	.w6(32'h3c6a8590),
	.w7(32'h3c0aa69b),
	.w8(32'h3a8baefe),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc2225),
	.w1(32'hbc807beb),
	.w2(32'hbb0afee8),
	.w3(32'hbc439b38),
	.w4(32'hb959cd08),
	.w5(32'hbb99f83c),
	.w6(32'hbc6a3487),
	.w7(32'hbafd159a),
	.w8(32'hbb524ce9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1fd9d),
	.w1(32'hbabae670),
	.w2(32'h3b18773e),
	.w3(32'hbb0bb195),
	.w4(32'h3ba472c9),
	.w5(32'h3d0158ad),
	.w6(32'h3c78568b),
	.w7(32'hbad1dbac),
	.w8(32'h3d1fb6e9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd0d17),
	.w1(32'h3c800df1),
	.w2(32'h3c39b3c6),
	.w3(32'h3bd58e65),
	.w4(32'h3b7a0ac9),
	.w5(32'hbbba24ea),
	.w6(32'h3ca7ebf7),
	.w7(32'h3c34a1a0),
	.w8(32'hbc603db3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d24a3),
	.w1(32'hbc784fbe),
	.w2(32'hbbdf9bbd),
	.w3(32'h3b080b58),
	.w4(32'h3b5e4a90),
	.w5(32'h3b116434),
	.w6(32'hbc178a68),
	.w7(32'hbb562fae),
	.w8(32'h3c5c5ea4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93b34b),
	.w1(32'hbb950f25),
	.w2(32'h3b2cce3d),
	.w3(32'h3bfc0a04),
	.w4(32'h3c979c7a),
	.w5(32'hbb460831),
	.w6(32'hbb9de1e0),
	.w7(32'h3c748b87),
	.w8(32'hbafc7136),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9a59c),
	.w1(32'h3c11ab84),
	.w2(32'h3c03ae9b),
	.w3(32'h3c0c9482),
	.w4(32'h388aced5),
	.w5(32'hbaa99c83),
	.w6(32'h3cb3dc1e),
	.w7(32'h3b553f44),
	.w8(32'hbae68d94),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc1883),
	.w1(32'hba1a4f6c),
	.w2(32'hbae5b610),
	.w3(32'hbb06708c),
	.w4(32'hbb0a1a5b),
	.w5(32'hbb5bba60),
	.w6(32'hbbcc57f5),
	.w7(32'hbba05084),
	.w8(32'hbc2dd8c9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac29b3b),
	.w1(32'hbb8cb9a9),
	.w2(32'h3b44edcf),
	.w3(32'hbbb9f118),
	.w4(32'hb8925ce5),
	.w5(32'h3b8e1601),
	.w6(32'hbc3a93e6),
	.w7(32'hba14696d),
	.w8(32'hba932885),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8049a),
	.w1(32'hbb2eebaf),
	.w2(32'hbafb982c),
	.w3(32'hba5d3cf0),
	.w4(32'hbb13b0eb),
	.w5(32'hba7cde96),
	.w6(32'h3aff3333),
	.w7(32'h3b69de0c),
	.w8(32'h3bec2916),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba16ff2),
	.w1(32'h3b2d04d7),
	.w2(32'hbbcbe7b4),
	.w3(32'hba66f1c9),
	.w4(32'hbb0ca59a),
	.w5(32'h3b6e76a5),
	.w6(32'h3add4e96),
	.w7(32'hbb3468c5),
	.w8(32'hbaa43183),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc386902),
	.w1(32'h3ae52f9e),
	.w2(32'h397b42ed),
	.w3(32'hbb9f1dd4),
	.w4(32'hbbe798d8),
	.w5(32'hbb77b434),
	.w6(32'h3c22ca8f),
	.w7(32'hbb07a57b),
	.w8(32'hbaef000d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18d086),
	.w1(32'hbc1eff1d),
	.w2(32'hbc32c1e5),
	.w3(32'hbbdd0f80),
	.w4(32'h3be73c53),
	.w5(32'h3c3317f0),
	.w6(32'h38c8c28f),
	.w7(32'hbbb8cca2),
	.w8(32'h3c505514),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc722767),
	.w1(32'h3c8c93cf),
	.w2(32'hb7a32640),
	.w3(32'h3c24ff43),
	.w4(32'h3b8b2920),
	.w5(32'h3c63b0ac),
	.w6(32'h3d02bf97),
	.w7(32'h3abffc9c),
	.w8(32'h3d176cc6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb916711),
	.w1(32'h3c4c3789),
	.w2(32'h3c6505a7),
	.w3(32'hbbb5ddfd),
	.w4(32'h3c36c9c5),
	.w5(32'hbc042ab2),
	.w6(32'h3c5ae521),
	.w7(32'h3c86f9ae),
	.w8(32'hbc15b8b8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d552b),
	.w1(32'h3ba98741),
	.w2(32'h3c0df54e),
	.w3(32'hbb72d924),
	.w4(32'hbac046a5),
	.w5(32'h3a3f70f0),
	.w6(32'h3b8ccb1c),
	.w7(32'h3ad1a476),
	.w8(32'h3b3dc56f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e432b),
	.w1(32'h3a840928),
	.w2(32'h3a50515d),
	.w3(32'h3c9baf30),
	.w4(32'h3c0ceb63),
	.w5(32'h3c639e4c),
	.w6(32'h3c7a3579),
	.w7(32'h3b86d00c),
	.w8(32'h3d0eb7f7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c760acd),
	.w1(32'h3d02dd8a),
	.w2(32'hbc4ac480),
	.w3(32'h3cc4a6ac),
	.w4(32'hbaf641a2),
	.w5(32'hbb110cfc),
	.w6(32'h3cae5cf3),
	.w7(32'hbbc70d9f),
	.w8(32'h3a83b85f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb074c),
	.w1(32'hbae4411e),
	.w2(32'hba5d16d9),
	.w3(32'hbc1d7f2c),
	.w4(32'hbb2964a4),
	.w5(32'h3b091757),
	.w6(32'hbcaa2b00),
	.w7(32'hbb932569),
	.w8(32'hbc18d5ac),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80d57d),
	.w1(32'h3985a516),
	.w2(32'hbb0d151e),
	.w3(32'h3a956ac6),
	.w4(32'h37e2a7cc),
	.w5(32'h3b00f1c3),
	.w6(32'hb9dcdf7b),
	.w7(32'h38028c29),
	.w8(32'hbb1f8d16),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4fe3d),
	.w1(32'h3a7a91af),
	.w2(32'h3bdb8e0b),
	.w3(32'h3a8349e4),
	.w4(32'h3a252c58),
	.w5(32'hbbed83f4),
	.w6(32'h3b163e1d),
	.w7(32'h39737692),
	.w8(32'hba1ae57e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e42f2),
	.w1(32'hbaa41c7d),
	.w2(32'h3a6a5e11),
	.w3(32'hba5a9a19),
	.w4(32'hbbbc2e51),
	.w5(32'h3bba5935),
	.w6(32'hba87d4bb),
	.w7(32'hbba5a2f0),
	.w8(32'h3bc57756),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8c1ca),
	.w1(32'hbb3e1df3),
	.w2(32'hbb6da2b7),
	.w3(32'h3bdd0418),
	.w4(32'h3bc387f9),
	.w5(32'hbba4275d),
	.w6(32'hbbc403c6),
	.w7(32'h3c09e02f),
	.w8(32'hbb093021),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae01c9),
	.w1(32'hbbcadfa5),
	.w2(32'hba67b666),
	.w3(32'hbab1c213),
	.w4(32'h3a2fb39c),
	.w5(32'hbc2735fc),
	.w6(32'hba79be24),
	.w7(32'h3aea0d22),
	.w8(32'hbc2ad016),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b4904),
	.w1(32'hbb41449f),
	.w2(32'h3b22850f),
	.w3(32'h3b746da6),
	.w4(32'h3b39cedf),
	.w5(32'hbbcc67d4),
	.w6(32'h3b87517b),
	.w7(32'h3bb2b62d),
	.w8(32'hbb395977),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2b98c),
	.w1(32'hbc490f7c),
	.w2(32'hbb221e0c),
	.w3(32'hbc7e889f),
	.w4(32'h3a222019),
	.w5(32'hbc0cf325),
	.w6(32'hbc7d01f1),
	.w7(32'h3b40d61f),
	.w8(32'hbae61cc0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81d0a4),
	.w1(32'hb8eb8e3a),
	.w2(32'h3ad32fe2),
	.w3(32'hbba1eabb),
	.w4(32'h3b26c393),
	.w5(32'hbaaafe8f),
	.w6(32'h3c07f0a4),
	.w7(32'h3b77457a),
	.w8(32'hbae81b6b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2fa4e),
	.w1(32'hbb6eb88a),
	.w2(32'hbae31222),
	.w3(32'hbb41a214),
	.w4(32'hbb60f691),
	.w5(32'hb9b1be15),
	.w6(32'hbb8717f2),
	.w7(32'hba84aac0),
	.w8(32'h3acff745),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3eea27),
	.w1(32'h3b567d42),
	.w2(32'h3bea5762),
	.w3(32'h3bf4eeee),
	.w4(32'h3badecba),
	.w5(32'hb9d3dbee),
	.w6(32'h3b80c132),
	.w7(32'h3b2f4f2c),
	.w8(32'hbba17d24),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0f849),
	.w1(32'h3b393841),
	.w2(32'h3ad61952),
	.w3(32'hbbb9b137),
	.w4(32'h3ba874fc),
	.w5(32'hbbca9892),
	.w6(32'hbbaecbc6),
	.w7(32'h3ad96833),
	.w8(32'hbb2f0680),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba254b),
	.w1(32'hbb882dfd),
	.w2(32'hbb91a310),
	.w3(32'hbb8ebd04),
	.w4(32'h381f82df),
	.w5(32'hbc3c7976),
	.w6(32'hbc07b8e8),
	.w7(32'h3b228237),
	.w8(32'hbb867fa8),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa25337),
	.w1(32'h3c089979),
	.w2(32'hbb301bd6),
	.w3(32'h3bc35445),
	.w4(32'hbb7d1fd2),
	.w5(32'hbb2f50fb),
	.w6(32'h3c738d4a),
	.w7(32'h39896fb0),
	.w8(32'hbbfafd9d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1749e0),
	.w1(32'hbb3edd75),
	.w2(32'h3ab01c5b),
	.w3(32'hbb787f2d),
	.w4(32'hbb569bf4),
	.w5(32'hbbba6e65),
	.w6(32'hbb43e9aa),
	.w7(32'h3ac16c64),
	.w8(32'hbc1d69f2),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba571aa),
	.w1(32'hb9f64cc6),
	.w2(32'hbb26d320),
	.w3(32'h3b9ea82f),
	.w4(32'hbb4b3219),
	.w5(32'hba8b6368),
	.w6(32'h3ac68249),
	.w7(32'hbae473f3),
	.w8(32'h3b6c14f4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d5e36),
	.w1(32'h3b4380a0),
	.w2(32'h39b10a71),
	.w3(32'h3a8b2019),
	.w4(32'hba9e894f),
	.w5(32'hbc02f019),
	.w6(32'h3b2487a2),
	.w7(32'h3aa0963c),
	.w8(32'hbc596007),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5efecb),
	.w1(32'h3c676de7),
	.w2(32'hba04dbee),
	.w3(32'h3b8f175f),
	.w4(32'hbbcf035e),
	.w5(32'h3b97a070),
	.w6(32'h3c0e18c8),
	.w7(32'hbae41574),
	.w8(32'h3c2f0fba),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17e315),
	.w1(32'hbb34b6ff),
	.w2(32'hbc55a534),
	.w3(32'hbb8a05b0),
	.w4(32'hbae4a504),
	.w5(32'h387738eb),
	.w6(32'h3bc2261c),
	.w7(32'hbb297adf),
	.w8(32'hba7fa04f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2aef41),
	.w1(32'h3b7b90ea),
	.w2(32'h3b592050),
	.w3(32'h3b4946e2),
	.w4(32'h3be0ee3f),
	.w5(32'hbb742870),
	.w6(32'h3af13983),
	.w7(32'h3b165c82),
	.w8(32'hbba9cfce),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c5fd0),
	.w1(32'hbc4f960d),
	.w2(32'h3b4e8ffe),
	.w3(32'hbc566255),
	.w4(32'hbb24b87a),
	.w5(32'hb95b2f97),
	.w6(32'hbb37b230),
	.w7(32'h3b7f02a3),
	.w8(32'h3b997ac9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd78947),
	.w1(32'hbacb56ba),
	.w2(32'h3801983a),
	.w3(32'h3bab05b4),
	.w4(32'hbbb3436b),
	.w5(32'h3ba15205),
	.w6(32'h3bc68012),
	.w7(32'hbb9cb195),
	.w8(32'h3c933073),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45abdd),
	.w1(32'h3814b7a4),
	.w2(32'h3bf2e61b),
	.w3(32'hbbaa68d8),
	.w4(32'h3b9e2517),
	.w5(32'hbc55d19a),
	.w6(32'hb90d9529),
	.w7(32'h3a734483),
	.w8(32'hbc059304),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3dda5d),
	.w1(32'hbb94b1e0),
	.w2(32'h3a7b60cc),
	.w3(32'hbb755efb),
	.w4(32'hba1745bd),
	.w5(32'hbb98f7e7),
	.w6(32'hbb177f4c),
	.w7(32'hbc0f7512),
	.w8(32'hbbf44f70),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba01e38),
	.w1(32'h3ccf19b4),
	.w2(32'h3a9e904a),
	.w3(32'h3c574c9b),
	.w4(32'hbb474a13),
	.w5(32'h3a151949),
	.w6(32'h3cbd4d28),
	.w7(32'hba04ce27),
	.w8(32'h3bab4410),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c1b7f),
	.w1(32'hbb91f6d1),
	.w2(32'h393b7fd0),
	.w3(32'hbba87d2d),
	.w4(32'hbb879184),
	.w5(32'hbbf02e20),
	.w6(32'hbc045041),
	.w7(32'hbbb60469),
	.w8(32'hbac0ab17),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4416a3),
	.w1(32'hbb59574b),
	.w2(32'h3bd1ceac),
	.w3(32'hbc00da40),
	.w4(32'hbbffebb8),
	.w5(32'hb9ccabdd),
	.w6(32'hbbaa74ee),
	.w7(32'hbaeae82b),
	.w8(32'hbbc1ddd0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd50dd),
	.w1(32'hbbe10c6d),
	.w2(32'hbb4cfa5c),
	.w3(32'h3c1256d8),
	.w4(32'hba3a4c5c),
	.w5(32'hbcac1fe4),
	.w6(32'h3b2a8ece),
	.w7(32'h3b53439a),
	.w8(32'hbca438e9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81df4b),
	.w1(32'hbc2fb0e6),
	.w2(32'hbb099254),
	.w3(32'hbc5ca932),
	.w4(32'h3bfc9cfa),
	.w5(32'hbac9fdf8),
	.w6(32'hbb784ef1),
	.w7(32'h3c077136),
	.w8(32'h3a78e629),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20a323),
	.w1(32'h3a9c152c),
	.w2(32'h3ba9396c),
	.w3(32'h3b954e1c),
	.w4(32'h3b11e068),
	.w5(32'hb97571f4),
	.w6(32'h3af2244c),
	.w7(32'h3a1c0a53),
	.w8(32'hba9d0e46),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac8137),
	.w1(32'hbb898a8d),
	.w2(32'h3b09335f),
	.w3(32'h3ba268f9),
	.w4(32'h3c34026d),
	.w5(32'hbb976815),
	.w6(32'h3b10f8a7),
	.w7(32'h3ba55834),
	.w8(32'hb9a10b00),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71eb8f),
	.w1(32'h385a3b3e),
	.w2(32'h3c14bc87),
	.w3(32'hbba1e9bf),
	.w4(32'hbae0c08f),
	.w5(32'h3be19c53),
	.w6(32'hbc1c9e83),
	.w7(32'hbbc9313b),
	.w8(32'h3a6403ff),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8d6fd),
	.w1(32'hb9820cb3),
	.w2(32'h3abe66c7),
	.w3(32'h3a85f892),
	.w4(32'h3a4ed391),
	.w5(32'h3b403c2a),
	.w6(32'hba144166),
	.w7(32'hbace1eb7),
	.w8(32'h3a97e58a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac66ef),
	.w1(32'h3b255e60),
	.w2(32'h3c220337),
	.w3(32'h3b8ed6c2),
	.w4(32'h3bd2db8c),
	.w5(32'hbb52c119),
	.w6(32'h3b842726),
	.w7(32'h3b5e4f83),
	.w8(32'h3ad28c7e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd44dd),
	.w1(32'h3ab03486),
	.w2(32'hbaaa9a5b),
	.w3(32'h3a2cf156),
	.w4(32'hb9973daf),
	.w5(32'hb9a30ead),
	.w6(32'h3ab00897),
	.w7(32'h3a8b8dfc),
	.w8(32'hbb2786a6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9049d5),
	.w1(32'hbb969191),
	.w2(32'h3c2f1b2d),
	.w3(32'h3b7fedb3),
	.w4(32'h3c3c404e),
	.w5(32'hba86d8e4),
	.w6(32'h3b3d27e9),
	.w7(32'h3c0c9800),
	.w8(32'hba72376e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb089f6d),
	.w1(32'hbacd66c5),
	.w2(32'hbaa389d5),
	.w3(32'hbb2cfdab),
	.w4(32'h3a7096a2),
	.w5(32'h3a350174),
	.w6(32'h3ab1a6a6),
	.w7(32'h3a434655),
	.w8(32'h39a986a5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a829ac8),
	.w1(32'h39d962e3),
	.w2(32'h3a597b3c),
	.w3(32'h3ad31941),
	.w4(32'h3ab16dab),
	.w5(32'hb9d208b7),
	.w6(32'h3b383380),
	.w7(32'h37ace48a),
	.w8(32'hb7bb9646),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9697634),
	.w1(32'hb8e42a55),
	.w2(32'hb91d2944),
	.w3(32'hb80e39de),
	.w4(32'h38f6c37a),
	.w5(32'h3a03d79e),
	.w6(32'h3a5bb270),
	.w7(32'hb9b15835),
	.w8(32'hba22d5cf),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb332b5d),
	.w1(32'h3a77abd6),
	.w2(32'hb96e0d92),
	.w3(32'hbb0b3250),
	.w4(32'hba87459c),
	.w5(32'hbb044032),
	.w6(32'h3805ba88),
	.w7(32'h3b06cf33),
	.w8(32'h3adfb537),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa07494),
	.w1(32'h3b473980),
	.w2(32'h3b2a467b),
	.w3(32'hbae51a5d),
	.w4(32'hb9c449bc),
	.w5(32'h3ae360d5),
	.w6(32'hb990b1c1),
	.w7(32'h3a88a66f),
	.w8(32'h3b807721),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cb0bd),
	.w1(32'h3911b220),
	.w2(32'h3b05533c),
	.w3(32'h3b0e8704),
	.w4(32'hb86605c3),
	.w5(32'h3ad0ae63),
	.w6(32'hba0ea328),
	.w7(32'hbb94b893),
	.w8(32'h3a27c31b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a702a9a),
	.w1(32'h3b11e86a),
	.w2(32'h3b12a940),
	.w3(32'h39a74b26),
	.w4(32'h39b853e9),
	.w5(32'hba42fb46),
	.w6(32'hb80cc43a),
	.w7(32'hba7f3d47),
	.w8(32'hbab1501d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f94dd),
	.w1(32'h3a80aff8),
	.w2(32'h3aba0f22),
	.w3(32'h3a1768bd),
	.w4(32'h3a885eb3),
	.w5(32'h3acd4099),
	.w6(32'hb9e79839),
	.w7(32'h3aedd6f9),
	.w8(32'h3b9129d3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce1b32),
	.w1(32'h3b6c350f),
	.w2(32'h3b5089f2),
	.w3(32'hbb851684),
	.w4(32'hbb1126f8),
	.w5(32'hb9a82779),
	.w6(32'hb90f5b79),
	.w7(32'hba88b415),
	.w8(32'hbaf08705),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bc0d7),
	.w1(32'hb9dcacba),
	.w2(32'h3aacc612),
	.w3(32'hbb18d8b6),
	.w4(32'h3a08e0b7),
	.w5(32'h3b8c2831),
	.w6(32'hbaed07be),
	.w7(32'hba4764a6),
	.w8(32'h3b69e6ed),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39428d05),
	.w1(32'h3aa99bc9),
	.w2(32'h3a5eb299),
	.w3(32'h3a73a329),
	.w4(32'h3a156f28),
	.w5(32'hbb0ef259),
	.w6(32'h3ab9ebd5),
	.w7(32'h3a4d315a),
	.w8(32'hba5fb551),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1a161),
	.w1(32'hbadcf998),
	.w2(32'hbb078380),
	.w3(32'hbb3312bb),
	.w4(32'hbb1020d1),
	.w5(32'h3adbef1e),
	.w6(32'hbad3abc9),
	.w7(32'hbae41885),
	.w8(32'hbae8475e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37963671),
	.w1(32'hba97ee6d),
	.w2(32'h3a99f503),
	.w3(32'h3aae4936),
	.w4(32'h3a341e9d),
	.w5(32'h3a3cec8d),
	.w6(32'hba59b9b3),
	.w7(32'h3a000528),
	.w8(32'h3893663d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2754a4),
	.w1(32'h3ab1dca6),
	.w2(32'h3ad6859e),
	.w3(32'h39e0dee5),
	.w4(32'hb8e03f5f),
	.w5(32'hbafec723),
	.w6(32'h3a7bc383),
	.w7(32'h3a7168bc),
	.w8(32'hbb227609),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba95caf),
	.w1(32'hbb699b8b),
	.w2(32'hba48d3a4),
	.w3(32'hbba9f0a0),
	.w4(32'hba95ff4c),
	.w5(32'h3b2b158b),
	.w6(32'hbba94a21),
	.w7(32'hbb0e9858),
	.w8(32'h3ad3c41e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f8bed),
	.w1(32'h3b66ebf1),
	.w2(32'h3b05fbfb),
	.w3(32'h37e77e09),
	.w4(32'hb98c95db),
	.w5(32'hbad3cec9),
	.w6(32'h3a69831f),
	.w7(32'h3afea40e),
	.w8(32'hbae218d7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5030c7),
	.w1(32'hba9f4901),
	.w2(32'h3ac801f2),
	.w3(32'hba1ade7b),
	.w4(32'h3a44e8be),
	.w5(32'h3a507274),
	.w6(32'hbacdd80f),
	.w7(32'h3aa39e1c),
	.w8(32'h3b3db330),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b582471),
	.w1(32'h3b32d7f7),
	.w2(32'h3b2bfc05),
	.w3(32'hbab3afde),
	.w4(32'hb9e8a2b1),
	.w5(32'hbafc7f6c),
	.w6(32'h3b0f2404),
	.w7(32'hb9e0acaf),
	.w8(32'hbb9068ec),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69120a),
	.w1(32'hba439eed),
	.w2(32'hbaa6175a),
	.w3(32'hbaa4b0f7),
	.w4(32'hb9b6f302),
	.w5(32'h3adb28fb),
	.w6(32'hbad7b1bd),
	.w7(32'hba85dd29),
	.w8(32'h3a28aec9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e56e4),
	.w1(32'h3b944bba),
	.w2(32'h3b0b23a7),
	.w3(32'h3ac4d488),
	.w4(32'h39d05e4c),
	.w5(32'h3ad554b5),
	.w6(32'h3acf6836),
	.w7(32'h38e17543),
	.w8(32'h390ebdb5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38405fca),
	.w1(32'hb80d6186),
	.w2(32'h3a78a67f),
	.w3(32'h3aef01e2),
	.w4(32'h3b12cd4c),
	.w5(32'hba5948c6),
	.w6(32'h3a31bba1),
	.w7(32'h3aad5401),
	.w8(32'hb842f492),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba045d67),
	.w1(32'hb9e357f4),
	.w2(32'h3875730f),
	.w3(32'hb9fd3059),
	.w4(32'hba827189),
	.w5(32'hb81eea5e),
	.w6(32'h3ac62eaf),
	.w7(32'h3a9f4e6f),
	.w8(32'h39973867),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c57e7),
	.w1(32'h3a4a73eb),
	.w2(32'hbafda64b),
	.w3(32'h3b479c76),
	.w4(32'hbb1528a7),
	.w5(32'hbba8af01),
	.w6(32'h3b207087),
	.w7(32'h3b5d464d),
	.w8(32'h3b90056a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8420d9),
	.w1(32'h3b60979f),
	.w2(32'h3ab69cb0),
	.w3(32'hbb7f8044),
	.w4(32'hbb4fc5dd),
	.w5(32'h3b214d60),
	.w6(32'hb9ba2da4),
	.w7(32'h3ad7bb2f),
	.w8(32'h3b72a9f5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e6c6f1),
	.w1(32'h3ad96d31),
	.w2(32'h3aba9422),
	.w3(32'h3af87268),
	.w4(32'h3a5c38fc),
	.w5(32'h3b0c3c1a),
	.w6(32'h3b4ff3bf),
	.w7(32'h3ab4b6d6),
	.w8(32'h3b3c3963),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394dd26a),
	.w1(32'hb986fe9d),
	.w2(32'h3b2e1a3c),
	.w3(32'h3b52d5d2),
	.w4(32'h3b441e63),
	.w5(32'hb9926c9d),
	.w6(32'h3b6ae3c1),
	.w7(32'h3b079e43),
	.w8(32'hba898b40),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba263738),
	.w1(32'hba7b396a),
	.w2(32'h3a23dbd7),
	.w3(32'hb9a25536),
	.w4(32'h3a278299),
	.w5(32'hb9b9ab43),
	.w6(32'h38fb4f30),
	.w7(32'hb94ffb53),
	.w8(32'h39173982),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0332fd),
	.w1(32'hba998287),
	.w2(32'h3a16a015),
	.w3(32'hbb7630d3),
	.w4(32'hbb3a1e99),
	.w5(32'h3a5b9022),
	.w6(32'h39b81775),
	.w7(32'hba446633),
	.w8(32'h3b05c3a2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01ae16),
	.w1(32'h3afc0800),
	.w2(32'h38e31690),
	.w3(32'hb9c719e8),
	.w4(32'hbb0c66b8),
	.w5(32'h3a11d9b6),
	.w6(32'h3a5ed275),
	.w7(32'hba81fd6b),
	.w8(32'hb9a2334d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb726ed0),
	.w1(32'h3abd9db8),
	.w2(32'h393e9502),
	.w3(32'hb722a1f8),
	.w4(32'hba35fc4a),
	.w5(32'hbb0aa42d),
	.w6(32'h3b515773),
	.w7(32'h3b493f67),
	.w8(32'h3b11a9d5),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b5d2b),
	.w1(32'hba094a84),
	.w2(32'h3a48069a),
	.w3(32'hbb3b972b),
	.w4(32'hba67fc04),
	.w5(32'hb94734f8),
	.w6(32'hbb73564f),
	.w7(32'hbb225055),
	.w8(32'h3892ce7a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e2ff4),
	.w1(32'h3adb1ec3),
	.w2(32'h3a96189b),
	.w3(32'hbaf687b4),
	.w4(32'hbb1990b0),
	.w5(32'hba1f7d67),
	.w6(32'hba64114d),
	.w7(32'hba2c09b4),
	.w8(32'h3ae5a9fa),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c26f03),
	.w1(32'h3b200490),
	.w2(32'h3b0d3d26),
	.w3(32'h3a36f94d),
	.w4(32'h3a012dca),
	.w5(32'hba48297b),
	.w6(32'h3b86f4eb),
	.w7(32'h3b60b32d),
	.w8(32'h3b0b6a0c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adce171),
	.w1(32'h3aa2d59f),
	.w2(32'h3b7e9954),
	.w3(32'h39b0ffe8),
	.w4(32'h3b336426),
	.w5(32'h3b838608),
	.w6(32'hba767bd2),
	.w7(32'h3b193615),
	.w8(32'h3b80d52d),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c8406),
	.w1(32'h3b8da21d),
	.w2(32'h3bb5aa5a),
	.w3(32'hba5b6934),
	.w4(32'h3a2a26d6),
	.w5(32'hbb0c443d),
	.w6(32'h3b047b4b),
	.w7(32'h3b38983a),
	.w8(32'h398370a7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9abe448),
	.w1(32'h3a334b2d),
	.w2(32'h3a2f97e8),
	.w3(32'hbadc5694),
	.w4(32'hba1adf82),
	.w5(32'h3ac54b36),
	.w6(32'h39bfffb8),
	.w7(32'h3a876640),
	.w8(32'h3a96578a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b392c2f),
	.w1(32'hba0228cc),
	.w2(32'h3b1d6971),
	.w3(32'hba05ca13),
	.w4(32'hbae91950),
	.w5(32'hbb05e8ff),
	.w6(32'hbaa434de),
	.w7(32'hbb98b053),
	.w8(32'hbaebf51a),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65ad79),
	.w1(32'h3b8e5fbd),
	.w2(32'h3baad9b8),
	.w3(32'h3acc4b91),
	.w4(32'h3b9a1882),
	.w5(32'h3b664e1a),
	.w6(32'h3ab9e470),
	.w7(32'h3b8d9239),
	.w8(32'h3b43646c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d4601),
	.w1(32'hba0bf91c),
	.w2(32'h3a0993e3),
	.w3(32'hba5d6008),
	.w4(32'hba56791e),
	.w5(32'hba54e03c),
	.w6(32'hba1586cd),
	.w7(32'hba9c2394),
	.w8(32'hba0df996),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7381b6),
	.w1(32'h3988d9b4),
	.w2(32'h3a0a5c76),
	.w3(32'hb9564615),
	.w4(32'hb9f7f8dc),
	.w5(32'hbaaef6f2),
	.w6(32'h3a8e8ce2),
	.w7(32'h39f22d73),
	.w8(32'hbaa40c8e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad71933),
	.w1(32'hba80c677),
	.w2(32'h39c9935e),
	.w3(32'hbb063b19),
	.w4(32'hb97c1f2f),
	.w5(32'h3aa9d203),
	.w6(32'hb9bb4224),
	.w7(32'h399e7cdb),
	.w8(32'h3ab2643e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba685c5),
	.w1(32'h3b987f6f),
	.w2(32'h3ba6eee5),
	.w3(32'h3b3756e3),
	.w4(32'h3b52648e),
	.w5(32'h3a9c84df),
	.w6(32'h39f6c7e3),
	.w7(32'h3b0c2632),
	.w8(32'hba94cd85),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb940201),
	.w1(32'hbad97311),
	.w2(32'hbaef6e77),
	.w3(32'hbb7b2cef),
	.w4(32'hbac551da),
	.w5(32'hba914fd3),
	.w6(32'hbac6f5f5),
	.w7(32'h39dde65a),
	.w8(32'h3a36945e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3ed14),
	.w1(32'h37fd9d08),
	.w2(32'hb97aa8dc),
	.w3(32'h392b210d),
	.w4(32'h3a02e353),
	.w5(32'hbad84466),
	.w6(32'hba797b01),
	.w7(32'hba792060),
	.w8(32'hba596f24),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66534b),
	.w1(32'h398b31d5),
	.w2(32'h3a1c2375),
	.w3(32'hbb7961fa),
	.w4(32'hbb12fdb0),
	.w5(32'h3b2cecc6),
	.w6(32'hbb2d8736),
	.w7(32'hba80151b),
	.w8(32'h3b09c18a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b006e3b),
	.w1(32'h3b59cd10),
	.w2(32'h3b5fb057),
	.w3(32'h3b10ea7e),
	.w4(32'h3ae49a1d),
	.w5(32'h3b37da8d),
	.w6(32'h3b0da7ae),
	.w7(32'h3b041307),
	.w8(32'h3b8c09db),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c28370),
	.w1(32'h3b051022),
	.w2(32'h3b2e4adb),
	.w3(32'hba946fcc),
	.w4(32'hbad23d7b),
	.w5(32'h3a9ab870),
	.w6(32'hb8dfd073),
	.w7(32'hb8e2e92f),
	.w8(32'h3b63601a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8475f2),
	.w1(32'h3b040bb0),
	.w2(32'hbac9fdbf),
	.w3(32'h3bcbcb44),
	.w4(32'h399e3a0c),
	.w5(32'h376e1eb4),
	.w6(32'h3b8cc687),
	.w7(32'hbbd95a90),
	.w8(32'hbb5cce27),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31101d),
	.w1(32'h3b24630f),
	.w2(32'h3b252db2),
	.w3(32'h3b41e435),
	.w4(32'h3af2857e),
	.w5(32'h3a979c36),
	.w6(32'h3abeefb4),
	.w7(32'h3a95d182),
	.w8(32'hbaaede2a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39999637),
	.w1(32'h3a0c1a63),
	.w2(32'h3a175017),
	.w3(32'h3b018d9d),
	.w4(32'h3aea6f50),
	.w5(32'hba927529),
	.w6(32'h3a53242e),
	.w7(32'h3a8263dc),
	.w8(32'hba6f72c3),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99d6b9),
	.w1(32'hba69f81e),
	.w2(32'hb8aa065e),
	.w3(32'hbbd6aba5),
	.w4(32'hbb894890),
	.w5(32'h3af70db5),
	.w6(32'hbba4780b),
	.w7(32'hbb7cc061),
	.w8(32'hba99bc5f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5a122),
	.w1(32'h3af2cc35),
	.w2(32'h3ab53db0),
	.w3(32'h3b0455ae),
	.w4(32'h3b43c0cd),
	.w5(32'h3aa51524),
	.w6(32'h39cbc1f5),
	.w7(32'h3aa56997),
	.w8(32'hbab31505),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cd3e9),
	.w1(32'hbb33b023),
	.w2(32'hb969ec53),
	.w3(32'hba1627e8),
	.w4(32'h3965f879),
	.w5(32'h3af2a7a1),
	.w6(32'hbb1204e6),
	.w7(32'hbb0e87eb),
	.w8(32'h398dda33),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a7c22),
	.w1(32'hb9cfdaef),
	.w2(32'hb99e3059),
	.w3(32'h3a562721),
	.w4(32'hb9122825),
	.w5(32'h3a45cfd6),
	.w6(32'h3b6e6cec),
	.w7(32'h3a4a204a),
	.w8(32'h3a96a052),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38668d40),
	.w1(32'h3b082726),
	.w2(32'h3ac13f03),
	.w3(32'h3b165257),
	.w4(32'h3a84533c),
	.w5(32'h3b4b1a1a),
	.w6(32'h3a66da7d),
	.w7(32'h39479621),
	.w8(32'hba8003ae),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc785c),
	.w1(32'h3a8e1995),
	.w2(32'h3b1e203f),
	.w3(32'h3b079d45),
	.w4(32'h3a5d71cd),
	.w5(32'hbb778835),
	.w6(32'h3a868148),
	.w7(32'h3aafc522),
	.w8(32'hbb524d9a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bf737),
	.w1(32'hbb1759be),
	.w2(32'hbb091779),
	.w3(32'hbace7bb8),
	.w4(32'hba62c265),
	.w5(32'h39b2f2bb),
	.w6(32'hba437a3a),
	.w7(32'hbb1d539f),
	.w8(32'h3ab92b5b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ae8d9),
	.w1(32'h3a9db671),
	.w2(32'h3b14da9f),
	.w3(32'hbae4cec1),
	.w4(32'hba220683),
	.w5(32'h39c5798a),
	.w6(32'h39aefbe5),
	.w7(32'hb957c29f),
	.w8(32'h3a8e36b8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98e3f9),
	.w1(32'h3ad80bf9),
	.w2(32'hba112799),
	.w3(32'h3a9575ca),
	.w4(32'h3ac6711c),
	.w5(32'h3b17c419),
	.w6(32'h3b4fae0d),
	.w7(32'h3a93b1e6),
	.w8(32'hbb154ea9),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9335be),
	.w1(32'h3b2b6d53),
	.w2(32'hba8dfdc1),
	.w3(32'h3b722420),
	.w4(32'h3880271e),
	.w5(32'hbb2b30e9),
	.w6(32'h3b9329fe),
	.w7(32'h3a602ba6),
	.w8(32'hb8c1fc66),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a964eae),
	.w1(32'h3a183ea9),
	.w2(32'h3b21231e),
	.w3(32'h3a972030),
	.w4(32'h3a59ad44),
	.w5(32'hb9c35d6f),
	.w6(32'h39f9aa52),
	.w7(32'h3a44ed4d),
	.w8(32'hbace2fac),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a904612),
	.w1(32'h3afadfff),
	.w2(32'h39b2d7ee),
	.w3(32'h3a91cf0b),
	.w4(32'h39a0fa3b),
	.w5(32'hbb011599),
	.w6(32'h3a1e6535),
	.w7(32'hb99887c8),
	.w8(32'h38e29f48),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384aeda4),
	.w1(32'h39885494),
	.w2(32'h39dc674f),
	.w3(32'hbb21cd62),
	.w4(32'hba84744d),
	.w5(32'h3b3eef10),
	.w6(32'hbb2a30be),
	.w7(32'hb92bf348),
	.w8(32'h3b19b886),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad1a91),
	.w1(32'h3b806085),
	.w2(32'h3b59f6b5),
	.w3(32'hbb219dbd),
	.w4(32'h3a877922),
	.w5(32'hba746444),
	.w6(32'hbabc5336),
	.w7(32'h3b9aa121),
	.w8(32'h3acf733c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82a93e),
	.w1(32'h3965c3d3),
	.w2(32'h3a775973),
	.w3(32'h3a981552),
	.w4(32'h3a596b95),
	.w5(32'h3a9b02bd),
	.w6(32'h3b0109f2),
	.w7(32'h3ad768cd),
	.w8(32'h3ab18562),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995cd36),
	.w1(32'h3b6d31ea),
	.w2(32'h3bd9f501),
	.w3(32'hbafa0ebb),
	.w4(32'h3a25a139),
	.w5(32'h3bddab91),
	.w6(32'hba0600ba),
	.w7(32'h3b20dc6a),
	.w8(32'h3b3ece45),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3738d),
	.w1(32'h3aac4feb),
	.w2(32'h39aa931f),
	.w3(32'h3ace8c3b),
	.w4(32'hb88ba28b),
	.w5(32'h3a2a99a1),
	.w6(32'h3b036487),
	.w7(32'hb9d7c563),
	.w8(32'hb8d9e978),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd78aa0),
	.w1(32'hba9782a8),
	.w2(32'hbc1849a0),
	.w3(32'hbb8df824),
	.w4(32'hbb9ca4ac),
	.w5(32'hbb7b93e7),
	.w6(32'hbab9d467),
	.w7(32'hbb616d30),
	.w8(32'h3aa756ea),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb435a93),
	.w1(32'hba92124b),
	.w2(32'h3a8ab47a),
	.w3(32'h39ec334d),
	.w4(32'hb8c1373b),
	.w5(32'h3ab8a3f4),
	.w6(32'h3af9b8ce),
	.w7(32'h3b061d97),
	.w8(32'hba3086d9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c671c),
	.w1(32'h3b1e5d38),
	.w2(32'h3b0af1c4),
	.w3(32'hbb1d5907),
	.w4(32'h3916dbd0),
	.w5(32'h3a279b7e),
	.w6(32'hba7027f3),
	.w7(32'h39a21ed5),
	.w8(32'h3b36afaa),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a891ffb),
	.w1(32'h3ac1f384),
	.w2(32'h3adb7305),
	.w3(32'hba9d8678),
	.w4(32'h3a311c3c),
	.w5(32'h3907fd8e),
	.w6(32'hbadd2b0c),
	.w7(32'h3aa04b18),
	.w8(32'h3afab43e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb222e),
	.w1(32'h3bcdcfcb),
	.w2(32'h3b3ac217),
	.w3(32'hbafd4a75),
	.w4(32'hba8dbffb),
	.w5(32'h3a033ee8),
	.w6(32'h3abf5264),
	.w7(32'h3ac73218),
	.w8(32'h3a9fc326),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c85e53),
	.w1(32'hba5fe583),
	.w2(32'hb9142a77),
	.w3(32'hbaa81e9c),
	.w4(32'hb9a5211e),
	.w5(32'hba0cf5cf),
	.w6(32'hba99b46c),
	.w7(32'hba4d6bd1),
	.w8(32'hb998c24e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c26d61),
	.w1(32'h3a99d2ff),
	.w2(32'h3a479199),
	.w3(32'h3a87d0a7),
	.w4(32'hb8f06916),
	.w5(32'hba198a30),
	.w6(32'h3a55d99b),
	.w7(32'h39d82d7f),
	.w8(32'hbb035826),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac49e24),
	.w1(32'hba86e24f),
	.w2(32'h3a81ea0b),
	.w3(32'hba9fabdd),
	.w4(32'hba8242fd),
	.w5(32'h3988304e),
	.w6(32'hb9053004),
	.w7(32'hb9b0778f),
	.w8(32'hb8ef1f9a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec4428),
	.w1(32'h3b4961e8),
	.w2(32'h3a88b45e),
	.w3(32'hbb01d5d8),
	.w4(32'hbb074ea6),
	.w5(32'h3aa6b1fd),
	.w6(32'h3b4a3a8c),
	.w7(32'h3ac59836),
	.w8(32'h3a98e2e7),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54d714),
	.w1(32'hba59eafe),
	.w2(32'hb911bd10),
	.w3(32'h398773ea),
	.w4(32'hba1c15e3),
	.w5(32'hba98c443),
	.w6(32'hba76fde7),
	.w7(32'h3abc5e20),
	.w8(32'hb9bd0b53),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b02642),
	.w1(32'h3a5e101e),
	.w2(32'h3a418e1a),
	.w3(32'hba114dab),
	.w4(32'hba00c940),
	.w5(32'h3a5956b2),
	.w6(32'h39b02b0d),
	.w7(32'h3a69e607),
	.w8(32'h3ac95f55),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa52b5a),
	.w1(32'h3b1ae580),
	.w2(32'h39bea4f1),
	.w3(32'h3a2e47cd),
	.w4(32'hb8bcb518),
	.w5(32'h395339c2),
	.w6(32'h3a36290a),
	.w7(32'hba577cb1),
	.w8(32'hba4110ae),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6a4a8),
	.w1(32'hba846e0c),
	.w2(32'hb93f24f4),
	.w3(32'h3a2171bc),
	.w4(32'hba8355d9),
	.w5(32'hba6427a5),
	.w6(32'h3a8b8284),
	.w7(32'hba9bed68),
	.w8(32'h3a3ed3d3),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba064d75),
	.w1(32'hb9dd2929),
	.w2(32'h3b07f272),
	.w3(32'h3a5cbd31),
	.w4(32'h3b82fd66),
	.w5(32'hbb2bee66),
	.w6(32'h39a573e4),
	.w7(32'h3af10fe0),
	.w8(32'hbae44cc3),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0583f),
	.w1(32'hba96580d),
	.w2(32'hba5663af),
	.w3(32'hba803e55),
	.w4(32'hb985fa26),
	.w5(32'hba06aa6a),
	.w6(32'hba041b39),
	.w7(32'h3933ccd8),
	.w8(32'h3ad0ee0b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01418a),
	.w1(32'hbb0ac704),
	.w2(32'hbba8beed),
	.w3(32'hbb92073f),
	.w4(32'hbb945dc7),
	.w5(32'hbb96d2cd),
	.w6(32'h3bb347e1),
	.w7(32'h3b5bfc48),
	.w8(32'h3b3b5479),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38afacd2),
	.w1(32'h3b6dedd7),
	.w2(32'hba0e40c3),
	.w3(32'hbb157f60),
	.w4(32'hbb69ec19),
	.w5(32'hba62f881),
	.w6(32'hbb011f3e),
	.w7(32'hbbe6eead),
	.w8(32'h39b6704c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08444c),
	.w1(32'hbb19d73f),
	.w2(32'h3a08a35e),
	.w3(32'h398ba70f),
	.w4(32'hba13bd0a),
	.w5(32'hb9b863e5),
	.w6(32'h3a49c585),
	.w7(32'h3a266e8f),
	.w8(32'h39c84799),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32e0bc),
	.w1(32'h3b08121b),
	.w2(32'h3b17aeb1),
	.w3(32'hb8e4f828),
	.w4(32'h39fe909d),
	.w5(32'h38c09ca7),
	.w6(32'h3b68cd7e),
	.w7(32'h3b801b58),
	.w8(32'hb8f5240b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba341d15),
	.w1(32'hb9e4f4a0),
	.w2(32'h3a3bb173),
	.w3(32'hba015fb7),
	.w4(32'h3a6ac90c),
	.w5(32'hb92eabb4),
	.w6(32'hba5e9442),
	.w7(32'h39e56c5e),
	.w8(32'hb99d56b5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dc9d0),
	.w1(32'h37d5dbce),
	.w2(32'h3a5d9612),
	.w3(32'hb9a23353),
	.w4(32'h39d583cd),
	.w5(32'hba8c72ba),
	.w6(32'hba833b3d),
	.w7(32'hb92e870d),
	.w8(32'h3ac143b3),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73f594),
	.w1(32'h3b954da6),
	.w2(32'h3b3fa91a),
	.w3(32'h3ae330bc),
	.w4(32'hba78471e),
	.w5(32'hbb4bab5a),
	.w6(32'h3bbbcdf7),
	.w7(32'h3b956ac9),
	.w8(32'hba0de9d9),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5de6c0),
	.w1(32'h3b6f846e),
	.w2(32'h3bd77599),
	.w3(32'h3b129284),
	.w4(32'h3b5ec7d3),
	.w5(32'h3bf83505),
	.w6(32'h3afe068e),
	.w7(32'h3b2d2a96),
	.w8(32'h3bb9d4e0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b653636),
	.w1(32'h3b482da1),
	.w2(32'h3b89dcfa),
	.w3(32'h3aacc014),
	.w4(32'h3b9b7d60),
	.w5(32'h3b825ea1),
	.w6(32'h3a1ebc97),
	.w7(32'h3b62501b),
	.w8(32'h3abddf7a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b1a04),
	.w1(32'h3a2a3333),
	.w2(32'h3af4098f),
	.w3(32'h3aece74d),
	.w4(32'h3a4b6696),
	.w5(32'h3b2bbe47),
	.w6(32'hbac1f64d),
	.w7(32'hb9a893cb),
	.w8(32'h3a98cb08),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb320a9c),
	.w1(32'hba721294),
	.w2(32'hbafbc8ca),
	.w3(32'h39b29700),
	.w4(32'hba31b6cf),
	.w5(32'hbad10372),
	.w6(32'h3b7b9129),
	.w7(32'h3b0b2d23),
	.w8(32'h3a0c1c9c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d9dcd),
	.w1(32'hbaae3463),
	.w2(32'h3ac5ce6a),
	.w3(32'hba2be21f),
	.w4(32'h3ad98a44),
	.w5(32'h3a94c834),
	.w6(32'hba3168a4),
	.w7(32'h3adefea3),
	.w8(32'h3ac88c31),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8613de),
	.w1(32'h3af7ad76),
	.w2(32'h3afae0bf),
	.w3(32'h3b8608ec),
	.w4(32'h3ac0f04a),
	.w5(32'hb9e3968b),
	.w6(32'h3b8ab698),
	.w7(32'h3690bb38),
	.w8(32'h3b29796b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb437f73),
	.w1(32'hbafe362d),
	.w2(32'hba31b60d),
	.w3(32'hb8e99820),
	.w4(32'h3b02adfb),
	.w5(32'hbb1cff04),
	.w6(32'h3bc55705),
	.w7(32'h3b3c2b11),
	.w8(32'hbab6e56f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacab3a),
	.w1(32'hbadf1489),
	.w2(32'hba92a094),
	.w3(32'hb90dded2),
	.w4(32'h393f4bb2),
	.w5(32'h3aab0911),
	.w6(32'hb89e58d4),
	.w7(32'h3aa9d9ee),
	.w8(32'h3a44c57a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1f994),
	.w1(32'h3b16cd3b),
	.w2(32'h3b6fc0c0),
	.w3(32'h3a9a801c),
	.w4(32'h3aa2d457),
	.w5(32'hbabf51d3),
	.w6(32'h3b2a15f0),
	.w7(32'h3b7513bd),
	.w8(32'h3b0ed139),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d8be8),
	.w1(32'h3b25560a),
	.w2(32'hb9f90feb),
	.w3(32'h39b2d60b),
	.w4(32'h3a4d56e8),
	.w5(32'h3b7ad6ff),
	.w6(32'hba2961f5),
	.w7(32'hba9a3ef1),
	.w8(32'h3a4cadbc),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab307dc),
	.w1(32'h3afa932d),
	.w2(32'h3b19efa1),
	.w3(32'hb907619c),
	.w4(32'h3ae854fa),
	.w5(32'h3b0b33d8),
	.w6(32'h3b06135f),
	.w7(32'h3b2ecd9b),
	.w8(32'hb9364926),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2ca7e),
	.w1(32'hbab8c4bd),
	.w2(32'hbaa53633),
	.w3(32'hb9581572),
	.w4(32'hba8d5ecf),
	.w5(32'hb988484f),
	.w6(32'h392f4fbd),
	.w7(32'hbaaaf1e6),
	.w8(32'h392519cf),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1291ad),
	.w1(32'h3b817660),
	.w2(32'h3a827083),
	.w3(32'h3a9d2745),
	.w4(32'h3a9d36c4),
	.w5(32'h3ab9fade),
	.w6(32'h3a6356f2),
	.w7(32'hb9bc3c16),
	.w8(32'h3a649ea3),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c986d),
	.w1(32'h3aa20910),
	.w2(32'h3ad40fb2),
	.w3(32'hbb364bf2),
	.w4(32'hbac140b9),
	.w5(32'hb90d84ff),
	.w6(32'h3969788c),
	.w7(32'h3a9657e3),
	.w8(32'h3ad1492c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8665e),
	.w1(32'h3a94e695),
	.w2(32'h3a32cd97),
	.w3(32'hbb96ffff),
	.w4(32'hb9bd80e3),
	.w5(32'hbb0cc8bf),
	.w6(32'hbb51a141),
	.w7(32'h3a827582),
	.w8(32'h3a9488cd),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d3b43),
	.w1(32'hb8d6c70d),
	.w2(32'hbac98ee9),
	.w3(32'hbac22417),
	.w4(32'hbad768de),
	.w5(32'h3b04d002),
	.w6(32'h3a9ea2f5),
	.w7(32'h3a0f4723),
	.w8(32'h3acdf5a5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0372c),
	.w1(32'hbb067f1f),
	.w2(32'hbb0334e5),
	.w3(32'h3b18d2c2),
	.w4(32'h38ecbfaf),
	.w5(32'h3b464da7),
	.w6(32'h38e3d566),
	.w7(32'hbb1c236c),
	.w8(32'h3aef9771),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9f1e9),
	.w1(32'h3ae135f3),
	.w2(32'h3b8e1d69),
	.w3(32'h3bdc8940),
	.w4(32'h3b88aaa2),
	.w5(32'h3b503921),
	.w6(32'h3ba56a2a),
	.w7(32'h3be3ba22),
	.w8(32'h3b4bcb56),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13cdd6),
	.w1(32'h3b010e0b),
	.w2(32'h3b08f7f8),
	.w3(32'h3a67d8f1),
	.w4(32'h3a5c98cb),
	.w5(32'h3ac33438),
	.w6(32'h3b355052),
	.w7(32'h3b520e4f),
	.w8(32'h3b4a18b3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfbf2a),
	.w1(32'h3afbae24),
	.w2(32'h3b04aa26),
	.w3(32'h39eb1174),
	.w4(32'h3acc781e),
	.w5(32'h3b6c1535),
	.w6(32'h3b0a4f0a),
	.w7(32'h3b186d9b),
	.w8(32'h3b25f745),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b245565),
	.w1(32'h3b997778),
	.w2(32'h3bc4defe),
	.w3(32'h3b9a7b0a),
	.w4(32'h39987d2b),
	.w5(32'hbaf08df2),
	.w6(32'h3b9d8f59),
	.w7(32'hbb5c7066),
	.w8(32'hba3e0dfe),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933aa1b),
	.w1(32'hb9516bb2),
	.w2(32'h3858aac2),
	.w3(32'h3950a834),
	.w4(32'hba093ac7),
	.w5(32'hba8e4d4c),
	.w6(32'h3a9ea9f5),
	.w7(32'h3a7e722b),
	.w8(32'h37cf3861),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf1a58),
	.w1(32'hba0f7fa6),
	.w2(32'h39b701ea),
	.w3(32'hba8083bb),
	.w4(32'hba3c4ae1),
	.w5(32'hba9af38b),
	.w6(32'h39f33619),
	.w7(32'h398df244),
	.w8(32'hbb1139fb),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b799cc2),
	.w1(32'hbac600fb),
	.w2(32'hba5d84e9),
	.w3(32'h3b320723),
	.w4(32'h3b8548d4),
	.w5(32'hbb9e0e8e),
	.w6(32'hb8c40330),
	.w7(32'h39e8c4e0),
	.w8(32'hb9dde027),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69ee8a),
	.w1(32'hbac82fae),
	.w2(32'hbb795604),
	.w3(32'hbafb5f47),
	.w4(32'hbb408f15),
	.w5(32'hbb518298),
	.w6(32'h3b3d805e),
	.w7(32'h3b11c2bd),
	.w8(32'hbad6a600),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb460965),
	.w1(32'hbb45f199),
	.w2(32'h3afde61c),
	.w3(32'h3a837b0c),
	.w4(32'h3b0ac73a),
	.w5(32'h387316f2),
	.w6(32'h3910f408),
	.w7(32'h3abfba24),
	.w8(32'hbad2190e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9911075),
	.w1(32'h3af6877f),
	.w2(32'h3b46bd0e),
	.w3(32'hba5afcb7),
	.w4(32'h39a46b7d),
	.w5(32'h3af53f09),
	.w6(32'hbb9f2784),
	.w7(32'hbb37416d),
	.w8(32'hba0c0e15),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02a3fe),
	.w1(32'h3b7b3963),
	.w2(32'h3b83d98a),
	.w3(32'h398d2bba),
	.w4(32'h3b1c8e65),
	.w5(32'h3b5dd432),
	.w6(32'hb96b1c2c),
	.w7(32'hba0303f5),
	.w8(32'h3ac7d40a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d8920),
	.w1(32'h3a0e413b),
	.w2(32'h3aa8a2ba),
	.w3(32'h3a2ef6d6),
	.w4(32'h39f393d3),
	.w5(32'h3b16330e),
	.w6(32'h3a2b8ff1),
	.w7(32'h39a2e449),
	.w8(32'h3b48100f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a319e),
	.w1(32'h3a62d15a),
	.w2(32'h3b5dc15f),
	.w3(32'h3ae07423),
	.w4(32'h3a9bce57),
	.w5(32'hb9f065bc),
	.w6(32'h3b5c66a8),
	.w7(32'h3b57791d),
	.w8(32'h3b08d509),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27a579),
	.w1(32'h3b999eef),
	.w2(32'h392e455d),
	.w3(32'h3b405b79),
	.w4(32'h3a96b349),
	.w5(32'h3a3db92c),
	.w6(32'h3ba937a5),
	.w7(32'h3b5b479e),
	.w8(32'h3b231532),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9ca70),
	.w1(32'hb76f1d6b),
	.w2(32'h3a7428e1),
	.w3(32'hba514bbe),
	.w4(32'hb901bf0d),
	.w5(32'hb7ca643d),
	.w6(32'h3a5c7bcd),
	.w7(32'h3b094b8b),
	.w8(32'hba3c3d24),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69aea1),
	.w1(32'hbb66a39c),
	.w2(32'hbaf802ff),
	.w3(32'hba2d428e),
	.w4(32'hbaa8e46f),
	.w5(32'hba4b4a75),
	.w6(32'hbb0b42eb),
	.w7(32'h3895704b),
	.w8(32'hbaec30a5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37abbaa6),
	.w1(32'hbafb8d80),
	.w2(32'hbafb1bcf),
	.w3(32'hbaad065d),
	.w4(32'hbb8097a9),
	.w5(32'hbb80c776),
	.w6(32'h394d96fd),
	.w7(32'hba84ee38),
	.w8(32'h3ac283b1),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81151f),
	.w1(32'h3961f7e2),
	.w2(32'hb9b4a6c0),
	.w3(32'hbabbdb78),
	.w4(32'hb9f8e8c5),
	.w5(32'hbae76e73),
	.w6(32'hbb2d861f),
	.w7(32'hbad76737),
	.w8(32'hbb4f2eb1),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e1e0),
	.w1(32'hbb9ac5b4),
	.w2(32'hbb99a77b),
	.w3(32'h3ab05572),
	.w4(32'hba0a02e9),
	.w5(32'hb9f2f366),
	.w6(32'hbaa4da3b),
	.w7(32'hbb4f4cc4),
	.w8(32'hba0bf0e6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bfec7),
	.w1(32'h38df3f3a),
	.w2(32'h3b8e9a89),
	.w3(32'hbaa3e10c),
	.w4(32'hb9d030c7),
	.w5(32'hbb920c89),
	.w6(32'h3ab01fc9),
	.w7(32'h3bc959b0),
	.w8(32'hbb2d4b82),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8298e1),
	.w1(32'hbaee12df),
	.w2(32'hbb187162),
	.w3(32'hba85d357),
	.w4(32'hbae4a55a),
	.w5(32'h3aefe38a),
	.w6(32'hbae07d85),
	.w7(32'hbaa861ec),
	.w8(32'h3a580967),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85f909),
	.w1(32'hbb4a6a0b),
	.w2(32'hb896c893),
	.w3(32'h3ba62661),
	.w4(32'h37fb534a),
	.w5(32'hb936c610),
	.w6(32'hbb66a9d8),
	.w7(32'h3baa759f),
	.w8(32'h38ae874c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4aa443),
	.w1(32'hba76fcbc),
	.w2(32'hba675154),
	.w3(32'hba432428),
	.w4(32'h3a386dfa),
	.w5(32'h3a1dcc05),
	.w6(32'h3a563ae7),
	.w7(32'h3a46411f),
	.w8(32'hba5a1751),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6d587),
	.w1(32'h39ff7d4d),
	.w2(32'h39bcacf3),
	.w3(32'h3b1410b4),
	.w4(32'h3b83ac3c),
	.w5(32'hbb6d2a97),
	.w6(32'h3ad9ada8),
	.w7(32'hba192b2b),
	.w8(32'hbad6baad),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53e29c),
	.w1(32'hba0bc1d6),
	.w2(32'hbb3dc97e),
	.w3(32'hbb40ff99),
	.w4(32'hba8c6104),
	.w5(32'h3abd4844),
	.w6(32'h3b042ff0),
	.w7(32'h3a4673fe),
	.w8(32'h3aa535fe),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d6764),
	.w1(32'hb91764ac),
	.w2(32'h3b91c5cc),
	.w3(32'hb91156fe),
	.w4(32'h3b8e4e21),
	.w5(32'hbba327e9),
	.w6(32'hbb10709d),
	.w7(32'h3b18a990),
	.w8(32'hbb42d95d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba290cf),
	.w1(32'hba8d796e),
	.w2(32'hbb86c0d2),
	.w3(32'hbb764a3b),
	.w4(32'hbbbf047d),
	.w5(32'h3ba48054),
	.w6(32'h39f3dba4),
	.w7(32'hbbadf533),
	.w8(32'h3b88c2a1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2eed6),
	.w1(32'h3ba7d69c),
	.w2(32'h3b7d494f),
	.w3(32'h3bba72df),
	.w4(32'h3ba36803),
	.w5(32'h39b0c7a3),
	.w6(32'h3b8d1011),
	.w7(32'h3b82b3be),
	.w8(32'h3a99295b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e61ac),
	.w1(32'h3b921b84),
	.w2(32'h3aa58d60),
	.w3(32'hbb280f93),
	.w4(32'hbb497b46),
	.w5(32'h3b90e925),
	.w6(32'hb8a1b32b),
	.w7(32'hbabe5be8),
	.w8(32'h3bd23e84),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921da3a),
	.w1(32'h3b0a1453),
	.w2(32'h3b0006c2),
	.w3(32'hbb134826),
	.w4(32'hbb0c2d75),
	.w5(32'h3b2640df),
	.w6(32'h3a1e9282),
	.w7(32'hbabfca0c),
	.w8(32'h3b5fda24),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59fec4),
	.w1(32'h3b4af659),
	.w2(32'h37d63782),
	.w3(32'h39b537ca),
	.w4(32'h3aace0e1),
	.w5(32'h3abf8e2a),
	.w6(32'hb9c1a442),
	.w7(32'h3aa6140d),
	.w8(32'h3aa73bf9),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb411460),
	.w1(32'h3a96f126),
	.w2(32'h3a9d85ed),
	.w3(32'h390ab954),
	.w4(32'hba334649),
	.w5(32'h3ac6e419),
	.w6(32'h3b38150d),
	.w7(32'hba659223),
	.w8(32'h3a816880),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54f86d),
	.w1(32'hba29400a),
	.w2(32'hb9401225),
	.w3(32'h3a7323a1),
	.w4(32'h39d5725d),
	.w5(32'h3af4c406),
	.w6(32'h3aa08883),
	.w7(32'h3a93d5e5),
	.w8(32'h3b3cf2ba),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98a3ef),
	.w1(32'h3baa07c1),
	.w2(32'h3b8bb752),
	.w3(32'h3b2689ec),
	.w4(32'h3b9ab3d0),
	.w5(32'hbb211651),
	.w6(32'h3ada0d44),
	.w7(32'h3b7afac0),
	.w8(32'hbbdf8ffd),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc256f),
	.w1(32'hbbc010d9),
	.w2(32'hba19b3e0),
	.w3(32'h3b44a9fe),
	.w4(32'hbb0d5d57),
	.w5(32'h39eecc8b),
	.w6(32'hbb676da3),
	.w7(32'h3ba6eaf2),
	.w8(32'hb9f456c6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cede51),
	.w1(32'h3ae1a13b),
	.w2(32'h3a9dc26e),
	.w3(32'hb96bb0f1),
	.w4(32'h3965fd7c),
	.w5(32'hbb48893a),
	.w6(32'h3b251ee8),
	.w7(32'h3b1092c7),
	.w8(32'hb9e4ea06),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba55922),
	.w1(32'hbba82d33),
	.w2(32'hba79e7d2),
	.w3(32'hbbab6dab),
	.w4(32'hba37d1b7),
	.w5(32'hbb2de228),
	.w6(32'hbbe65f39),
	.w7(32'hbb272851),
	.w8(32'hbb36a7de),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb329cb8),
	.w1(32'hbad811ec),
	.w2(32'hbaecdd7f),
	.w3(32'hbac39786),
	.w4(32'hbae73590),
	.w5(32'h3b3c637b),
	.w6(32'hba7d99cb),
	.w7(32'h39ebd265),
	.w8(32'h3b1c2baa),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a704b28),
	.w1(32'h37d5d147),
	.w2(32'hba06b584),
	.w3(32'hbaf583e5),
	.w4(32'h387aea6e),
	.w5(32'h3b7ab857),
	.w6(32'h3a97d130),
	.w7(32'h3adb0b30),
	.w8(32'hb95becb1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5944b),
	.w1(32'h3b0d0f74),
	.w2(32'hb9d72d32),
	.w3(32'h3a2a6e0e),
	.w4(32'h3a364b62),
	.w5(32'hbb0b6780),
	.w6(32'h3b4bcf9b),
	.w7(32'hbaf198ac),
	.w8(32'h3a39b762),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4fd66),
	.w1(32'hba67fc77),
	.w2(32'hbaafc4ea),
	.w3(32'hbb997665),
	.w4(32'hbb237449),
	.w5(32'h3a9dc920),
	.w6(32'hbacf3a13),
	.w7(32'hbb388334),
	.w8(32'h3a9f1889),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1886ef),
	.w1(32'h3ac2b3bd),
	.w2(32'hbb06af96),
	.w3(32'hbaa73bf4),
	.w4(32'hbae7c97b),
	.w5(32'hb9871797),
	.w6(32'h3a24f1f6),
	.w7(32'hbafebd50),
	.w8(32'h3a5ff549),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99dd07),
	.w1(32'h3c0cdde7),
	.w2(32'hbb50a985),
	.w3(32'hb8bf96c5),
	.w4(32'hbb29f8d3),
	.w5(32'h3aa6ba9e),
	.w6(32'h39771fc3),
	.w7(32'hbaa7810b),
	.w8(32'h3b457134),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba5389),
	.w1(32'h39e6d12d),
	.w2(32'h3af5e0e8),
	.w3(32'h3a392900),
	.w4(32'hba6d814b),
	.w5(32'hba41cf8f),
	.w6(32'h3ab6315c),
	.w7(32'h391480c9),
	.w8(32'h3a8b4ac1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc762bd),
	.w1(32'h3b77ffd6),
	.w2(32'hb8646f71),
	.w3(32'h3b3c839b),
	.w4(32'h3b2d9045),
	.w5(32'h3a96f8e8),
	.w6(32'h3b4600c6),
	.w7(32'h3be2dbe3),
	.w8(32'h3bae4a9c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule