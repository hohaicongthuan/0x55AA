module layer_10_featuremap_158(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb899b149),
	.w1(32'h3b2bd1fc),
	.w2(32'h3aaa001b),
	.w3(32'h3983edb1),
	.w4(32'h3b0159fd),
	.w5(32'hb9e78df5),
	.w6(32'h3aa8de2c),
	.w7(32'h3b301c0a),
	.w8(32'h3aaae3b0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06a642),
	.w1(32'h3aa0cc40),
	.w2(32'h3a098e26),
	.w3(32'h3a67a931),
	.w4(32'h3ac51b1d),
	.w5(32'h3aa86c91),
	.w6(32'h3ac90848),
	.w7(32'h3a8c0d3c),
	.w8(32'h3a6b5c66),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388cd267),
	.w1(32'hb9440a57),
	.w2(32'hba506d67),
	.w3(32'h3a5298f9),
	.w4(32'hb93da881),
	.w5(32'hba034d8c),
	.w6(32'hba038d7f),
	.w7(32'hba9820b1),
	.w8(32'hba0f1fed),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54b1f1),
	.w1(32'hba9f8f6d),
	.w2(32'hbb248381),
	.w3(32'h39596099),
	.w4(32'h3a9f1ed1),
	.w5(32'h3b64c10a),
	.w6(32'hbae0a99f),
	.w7(32'hbaeed7bd),
	.w8(32'hba4c32e4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75fb39),
	.w1(32'hba2bfb23),
	.w2(32'h3a9eb577),
	.w3(32'h39cdf743),
	.w4(32'h39db23f6),
	.w5(32'hba6e008f),
	.w6(32'hba68b25a),
	.w7(32'h3a5f731d),
	.w8(32'h3a95217b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d93bc),
	.w1(32'hba51203b),
	.w2(32'h38d85c11),
	.w3(32'h38a0585c),
	.w4(32'hba78fba4),
	.w5(32'hb9953271),
	.w6(32'hba9a3e70),
	.w7(32'hb88e0b98),
	.w8(32'hb998214f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936677d),
	.w1(32'h3a6f2748),
	.w2(32'h3954e6a3),
	.w3(32'h3a3b1c70),
	.w4(32'h3a233ca1),
	.w5(32'hb94dd915),
	.w6(32'h3a0619c5),
	.w7(32'h3a4b52a6),
	.w8(32'hb866e0f1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c52716),
	.w1(32'hbb20fc73),
	.w2(32'hbb592d79),
	.w3(32'hbb28ae51),
	.w4(32'hbafc418b),
	.w5(32'hbac65461),
	.w6(32'hbb6337ba),
	.w7(32'hbb92a148),
	.w8(32'hbb407a4f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2db9f),
	.w1(32'hbafd827b),
	.w2(32'hbaf3c59d),
	.w3(32'hbaa131dd),
	.w4(32'hbaf42aa7),
	.w5(32'hbaf4a24f),
	.w6(32'hbac342ab),
	.w7(32'hba942b4f),
	.w8(32'hba6c9ebf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb827449),
	.w1(32'hbb7ccdf0),
	.w2(32'hbbe346e1),
	.w3(32'hbaec9002),
	.w4(32'hba82f1ce),
	.w5(32'hbba0040d),
	.w6(32'hba4e2fa8),
	.w7(32'h3a725579),
	.w8(32'hbb631ea2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a661ffa),
	.w1(32'h39578299),
	.w2(32'h39ea1682),
	.w3(32'h3add0b06),
	.w4(32'h369885fa),
	.w5(32'h3a2133a1),
	.w6(32'hb9de38f4),
	.w7(32'h39539f23),
	.w8(32'h3938e331),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99802b7),
	.w1(32'hb9823f42),
	.w2(32'hb966eb50),
	.w3(32'hba3bd733),
	.w4(32'h3a8cd030),
	.w5(32'h3a50bc7d),
	.w6(32'hbb689300),
	.w7(32'hba9e8183),
	.w8(32'hbacef081),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf868e),
	.w1(32'hbb9e3cb4),
	.w2(32'hbbc6931d),
	.w3(32'hbb817942),
	.w4(32'hbb036c1e),
	.w5(32'hbb86733d),
	.w6(32'hbb7a2639),
	.w7(32'hbacd0f23),
	.w8(32'hbb53dd6b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a950ffc),
	.w1(32'hba6d0acc),
	.w2(32'hbaba3a6f),
	.w3(32'h3a99a5a9),
	.w4(32'hba37ca19),
	.w5(32'hbaf36fe3),
	.w6(32'h3963927a),
	.w7(32'hbad3131a),
	.w8(32'hbaae375d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4264d3),
	.w1(32'h3a4b41db),
	.w2(32'hbb4033e7),
	.w3(32'hbab8e34f),
	.w4(32'h3a807f5e),
	.w5(32'hbade4650),
	.w6(32'hbb02ddfc),
	.w7(32'hbb3ac3fd),
	.w8(32'hbb84dee6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fdc0e),
	.w1(32'hbaf6427e),
	.w2(32'hbb784a26),
	.w3(32'hbb2a7277),
	.w4(32'hbab74fa9),
	.w5(32'hbb5de3af),
	.w6(32'hb9f2c604),
	.w7(32'h397651c6),
	.w8(32'hbb0e071d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7d27b),
	.w1(32'hba4e728d),
	.w2(32'hbaf2a950),
	.w3(32'hba84abe3),
	.w4(32'hba8b6d79),
	.w5(32'hbac1a377),
	.w6(32'hbaa10376),
	.w7(32'hba54d5d6),
	.w8(32'h39f2dc17),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96cfd7),
	.w1(32'hbafb1d02),
	.w2(32'hbb143416),
	.w3(32'hbae4ba11),
	.w4(32'h3a1cbc94),
	.w5(32'hbaaee349),
	.w6(32'h3977882f),
	.w7(32'h3a12b361),
	.w8(32'hbabe23ad),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae90d79),
	.w1(32'hbb15e227),
	.w2(32'hbb3605f9),
	.w3(32'hb96d499d),
	.w4(32'hba9e647d),
	.w5(32'hbb25246e),
	.w6(32'hbb1951df),
	.w7(32'hbac302fe),
	.w8(32'hbb25bbff),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9adcad6),
	.w1(32'hb9348e24),
	.w2(32'hb89fd10a),
	.w3(32'h399b4111),
	.w4(32'hb90e86c9),
	.w5(32'hb993beb3),
	.w6(32'hb9440dfb),
	.w7(32'h38dce968),
	.w8(32'hb981f556),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd6a7c),
	.w1(32'hba6729b6),
	.w2(32'hba73f40f),
	.w3(32'hb9dae08c),
	.w4(32'hb88ccf8a),
	.w5(32'h38e86505),
	.w6(32'hbae8efec),
	.w7(32'hbab27f6e),
	.w8(32'hba09c6d5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54a320),
	.w1(32'hbb353a62),
	.w2(32'hbb142eff),
	.w3(32'h3956a598),
	.w4(32'h3af9bead),
	.w5(32'h3b31cf49),
	.w6(32'h3a46739e),
	.w7(32'h3a8306e7),
	.w8(32'h3ae4836f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6ee16),
	.w1(32'hba4bbd0a),
	.w2(32'hbaa7f4ef),
	.w3(32'h3ab79acd),
	.w4(32'hbb3936f0),
	.w5(32'hbb981fc6),
	.w6(32'hb9cb7e73),
	.w7(32'hbb7ceb52),
	.w8(32'hbba27ca6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d1691),
	.w1(32'hbb203a9b),
	.w2(32'hbbc12230),
	.w3(32'hb937fa3d),
	.w4(32'hbabde8ed),
	.w5(32'hbba9f3eb),
	.w6(32'hba2b92c4),
	.w7(32'h3947ea09),
	.w8(32'hbb310f3c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1b5a3),
	.w1(32'h390c5cb5),
	.w2(32'hbb1a7a06),
	.w3(32'hba93a352),
	.w4(32'h39c7a8f0),
	.w5(32'hbaaed4f8),
	.w6(32'hb8955ec9),
	.w7(32'h3a4f77d6),
	.w8(32'hbb055f8d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997ae7d),
	.w1(32'h3a46ac9d),
	.w2(32'hb9c500bc),
	.w3(32'h39669025),
	.w4(32'hba79b169),
	.w5(32'hba01d9f6),
	.w6(32'h3835ce5d),
	.w7(32'hb9ec8e3b),
	.w8(32'hba69fa93),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58faad),
	.w1(32'hb8c7bc5a),
	.w2(32'h3982d447),
	.w3(32'h39551e99),
	.w4(32'hb99e7813),
	.w5(32'hb805d18c),
	.w6(32'hb9cc422b),
	.w7(32'hb8ea6937),
	.w8(32'hb799e5fb),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d92f15),
	.w1(32'h3a0fdea6),
	.w2(32'h3933dae5),
	.w3(32'h39a28c6d),
	.w4(32'h3a5dfdf2),
	.w5(32'h39d033d7),
	.w6(32'h375442fe),
	.w7(32'h3aebce9c),
	.w8(32'h3abdc5f3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9e2eb),
	.w1(32'hb92e9bd3),
	.w2(32'h348b8c5b),
	.w3(32'h3a1f76f1),
	.w4(32'hba784153),
	.w5(32'hba86401f),
	.w6(32'hbadf7709),
	.w7(32'hba1a8e3e),
	.w8(32'hba027a50),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab71ab5),
	.w1(32'hbb4565e7),
	.w2(32'hbbc72922),
	.w3(32'hbaa366b4),
	.w4(32'hbb269e0a),
	.w5(32'hbb9ba48a),
	.w6(32'hbaae97b9),
	.w7(32'hbb1b836c),
	.w8(32'hbb89e5f8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23b448),
	.w1(32'hb9756c75),
	.w2(32'hb9a39720),
	.w3(32'hbb2cb36a),
	.w4(32'h3870b0fb),
	.w5(32'h393ca370),
	.w6(32'hba43824b),
	.w7(32'hba1376eb),
	.w8(32'h38a79c2d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cd3d63),
	.w1(32'hb9bfda35),
	.w2(32'hb99c30e7),
	.w3(32'h39931e93),
	.w4(32'hb9f57b5d),
	.w5(32'hb9e8dcbe),
	.w6(32'hba43f83e),
	.w7(32'hb9d7c07e),
	.w8(32'hba129319),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf493a),
	.w1(32'hb9c9e5dc),
	.w2(32'hba4be349),
	.w3(32'hba62d786),
	.w4(32'h3acda938),
	.w5(32'hba896081),
	.w6(32'h3aad12d3),
	.w7(32'h3ae8fbdc),
	.w8(32'hba637079),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925e5b7),
	.w1(32'hb9f70e00),
	.w2(32'h38ea5310),
	.w3(32'hb9a78cad),
	.w4(32'hba04768c),
	.w5(32'hbac43f28),
	.w6(32'h393d3c96),
	.w7(32'h3a8a5bbf),
	.w8(32'hbb06a6a6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadba7de),
	.w1(32'h39a62971),
	.w2(32'hb9b3d108),
	.w3(32'hbafe1ac4),
	.w4(32'h39f98baf),
	.w5(32'h39a74086),
	.w6(32'hba429006),
	.w7(32'h39be820a),
	.w8(32'hb9bc39df),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8c2ba),
	.w1(32'hba593a1e),
	.w2(32'hba8726c0),
	.w3(32'h3a04cdcc),
	.w4(32'h37c34f65),
	.w5(32'hba39a7f8),
	.w6(32'hba49a65b),
	.w7(32'hb9f13070),
	.w8(32'hba81dfd4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a360a7),
	.w1(32'h3a001522),
	.w2(32'hbad1693d),
	.w3(32'hb97bb60a),
	.w4(32'h3a2ab800),
	.w5(32'hbac7c2b0),
	.w6(32'h3a4767ca),
	.w7(32'h3ac00aa6),
	.w8(32'hbaee5552),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc1b5b),
	.w1(32'h3b8b9d2b),
	.w2(32'h3b7d5fb1),
	.w3(32'h3aae58de),
	.w4(32'h3b8fa53c),
	.w5(32'h3b70d653),
	.w6(32'h39982e37),
	.w7(32'h3b9b2275),
	.w8(32'h3b944e7f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa42128),
	.w1(32'h3b1ef5e3),
	.w2(32'h3ba53136),
	.w3(32'hba8b6f49),
	.w4(32'hb99badce),
	.w5(32'h3ac38ca6),
	.w6(32'hbb0564cc),
	.w7(32'hbaaf8df1),
	.w8(32'h3a720bd7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d71da6),
	.w1(32'h3a95460c),
	.w2(32'h3a3e2d85),
	.w3(32'h3a7cf553),
	.w4(32'h3b01845a),
	.w5(32'h3aaa7885),
	.w6(32'h3a944838),
	.w7(32'h3ac7c539),
	.w8(32'h39b908d0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6ce31),
	.w1(32'hbb24aae4),
	.w2(32'hbb6b4eb8),
	.w3(32'h39fd7ec5),
	.w4(32'hbb3356c1),
	.w5(32'hbb5887e8),
	.w6(32'hbb07d9fa),
	.w7(32'hbb80f4d7),
	.w8(32'hbb5d17a7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd7fd8),
	.w1(32'h381a07fe),
	.w2(32'h38a1a9ef),
	.w3(32'hbb061e1b),
	.w4(32'h3907a3fe),
	.w5(32'h38e5a2bd),
	.w6(32'h38d1cc6a),
	.w7(32'hb830755b),
	.w8(32'hba328ab8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a400c11),
	.w1(32'h396a32b7),
	.w2(32'hb964419c),
	.w3(32'hba1468b7),
	.w4(32'hb8da515c),
	.w5(32'hba278dcc),
	.w6(32'hba08f1b9),
	.w7(32'h39a3df0d),
	.w8(32'hb8c9f6ec),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8686e5),
	.w1(32'hba8af50d),
	.w2(32'hbba6419c),
	.w3(32'hba3d4d49),
	.w4(32'h3b0f100a),
	.w5(32'hbb19ff5a),
	.w6(32'h3ac46592),
	.w7(32'h3a8941b3),
	.w8(32'hbb87026d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e40b39),
	.w1(32'hba2e9183),
	.w2(32'hbb8c8aa4),
	.w3(32'h3af82da5),
	.w4(32'h3a4e67f6),
	.w5(32'hbb874c2e),
	.w6(32'h3adf9a07),
	.w7(32'h3b5168a8),
	.w8(32'h38f5c17b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39b2e9),
	.w1(32'hbae1413c),
	.w2(32'hbbd5d0e9),
	.w3(32'hbae9da1b),
	.w4(32'hb8d2583e),
	.w5(32'hbba8a459),
	.w6(32'h3a0dc6e8),
	.w7(32'h3ab7e86c),
	.w8(32'hbb70115c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab402bb),
	.w1(32'hbb023219),
	.w2(32'hbbc37028),
	.w3(32'hbb1db57c),
	.w4(32'h3a5554d5),
	.w5(32'hbaefca5a),
	.w6(32'hbb22ec53),
	.w7(32'hbb2f3e5b),
	.w8(32'hbb94d4ec),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1b64a),
	.w1(32'hbbb33a78),
	.w2(32'hbbc89cc5),
	.w3(32'hbb9d4bd1),
	.w4(32'hbb1d6a4c),
	.w5(32'hbb95b5de),
	.w6(32'hbbe8d472),
	.w7(32'hbbbd69a6),
	.w8(32'hbbc6c93d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38562d33),
	.w1(32'hb9264e02),
	.w2(32'hba43d0d9),
	.w3(32'hb99d78d6),
	.w4(32'hb996e283),
	.w5(32'hbab0de6d),
	.w6(32'h39ea57a5),
	.w7(32'h398cf5aa),
	.w8(32'hba818192),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90cdd33),
	.w1(32'h396d5cfe),
	.w2(32'hba17f1c3),
	.w3(32'hb9df7e4f),
	.w4(32'hb9a4659e),
	.w5(32'hba22c2e6),
	.w6(32'hba77d423),
	.w7(32'hbb029682),
	.w8(32'hbad5323b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67baaa),
	.w1(32'h3aaea299),
	.w2(32'h3978cb63),
	.w3(32'h3a7de3d2),
	.w4(32'h3a036cc6),
	.w5(32'hba041c75),
	.w6(32'h3a88f129),
	.w7(32'hb9ddd9cb),
	.w8(32'hbb0f5c06),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6dca37),
	.w1(32'hbadef3ad),
	.w2(32'hbb89fa5a),
	.w3(32'hba0829d4),
	.w4(32'h3a88a5e1),
	.w5(32'hbaed4ad1),
	.w6(32'h3ad81819),
	.w7(32'h3995cdb7),
	.w8(32'hbae5b345),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b515139),
	.w1(32'hb9f9efea),
	.w2(32'hb94a2352),
	.w3(32'h39bf7ec3),
	.w4(32'hb98d4c4a),
	.w5(32'h39049325),
	.w6(32'hba3e7370),
	.w7(32'h3a4a083e),
	.w8(32'hba0bf4af),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba788366),
	.w1(32'hbb5588f4),
	.w2(32'hbb5ab947),
	.w3(32'h3a9e640d),
	.w4(32'hb9d2ff6b),
	.w5(32'hbb973a6f),
	.w6(32'hb92f1e15),
	.w7(32'h3a9fc74a),
	.w8(32'hbae593fe),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06016f),
	.w1(32'hb9aa1c83),
	.w2(32'hb9ba0ec3),
	.w3(32'h3b035019),
	.w4(32'hb9f3212f),
	.w5(32'hba51de1a),
	.w6(32'hba0565ba),
	.w7(32'hb976eea5),
	.w8(32'h39baccec),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a4e77),
	.w1(32'hbadfe742),
	.w2(32'hb9c82906),
	.w3(32'hb9f2cda8),
	.w4(32'hba8a6966),
	.w5(32'hb90fd081),
	.w6(32'hbb1addc3),
	.w7(32'hbb2eb2cf),
	.w8(32'hbad1e24b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebaa06),
	.w1(32'hbaf4a401),
	.w2(32'hbb186cdf),
	.w3(32'hba152e79),
	.w4(32'hbaaeecbd),
	.w5(32'hbac2191f),
	.w6(32'hba8b2f30),
	.w7(32'hbb135b72),
	.w8(32'hbadf85f5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee8ca0),
	.w1(32'h3a49688e),
	.w2(32'hb9cc416d),
	.w3(32'hbacbdf65),
	.w4(32'hb99ac4c6),
	.w5(32'hb985a35c),
	.w6(32'hba0abd2d),
	.w7(32'hbad4449f),
	.w8(32'hb9855723),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8527cb),
	.w1(32'h3a8d6af1),
	.w2(32'h3a6185b0),
	.w3(32'hbab35ded),
	.w4(32'h3a72745c),
	.w5(32'h3a8bdc00),
	.w6(32'hb96f863b),
	.w7(32'h3995ef1f),
	.w8(32'h399ebc24),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8b704),
	.w1(32'hba37ff4e),
	.w2(32'hba743dcd),
	.w3(32'h39ab5920),
	.w4(32'hba73fa44),
	.w5(32'hba8ea3ea),
	.w6(32'hba9ec9b8),
	.w7(32'hba83c73e),
	.w8(32'hba2458b2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb139971),
	.w1(32'hbad07a8e),
	.w2(32'hbb2aaade),
	.w3(32'hba65b3b4),
	.w4(32'hba769891),
	.w5(32'hbaf5b08b),
	.w6(32'hb63f5b4c),
	.w7(32'hb9133c82),
	.w8(32'hba81012e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39f59d),
	.w1(32'hba320a87),
	.w2(32'hba0f8d70),
	.w3(32'h39bf08a4),
	.w4(32'hba358f08),
	.w5(32'hb9dfe0bc),
	.w6(32'hba1ae76b),
	.w7(32'hb9825b81),
	.w8(32'hba1b1c15),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391fc820),
	.w1(32'hb98b0513),
	.w2(32'h3a9e5367),
	.w3(32'hb92b6492),
	.w4(32'hb95c9ea5),
	.w5(32'hba6bd26c),
	.w6(32'h3ad01e5a),
	.w7(32'h3aa3ef28),
	.w8(32'h38da90e3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8de310),
	.w1(32'h3a561ba8),
	.w2(32'h3a2e2459),
	.w3(32'hbafe3985),
	.w4(32'h3a878f8d),
	.w5(32'h3a83f37b),
	.w6(32'h3a22c1da),
	.w7(32'h3a6b95c4),
	.w8(32'h3a2556b4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86dd0b),
	.w1(32'hb8608940),
	.w2(32'h3a081497),
	.w3(32'h3ad0949a),
	.w4(32'hb9496179),
	.w5(32'h3a2f703a),
	.w6(32'hb98ef9e0),
	.w7(32'h39ae3b05),
	.w8(32'h3a011b1e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985cd48),
	.w1(32'hba49ec03),
	.w2(32'hbadacbf5),
	.w3(32'h396a9e57),
	.w4(32'hb9e578f7),
	.w5(32'hb9d4a1c3),
	.w6(32'h3a8318d5),
	.w7(32'hba932302),
	.w8(32'hb98c1f1b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6315cf),
	.w1(32'hbb849ca4),
	.w2(32'hbb813170),
	.w3(32'h3abb2146),
	.w4(32'hbb167339),
	.w5(32'hbb3edeb2),
	.w6(32'hbb539e23),
	.w7(32'hbb84ff14),
	.w8(32'hbb871106),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb155083),
	.w1(32'hbad28299),
	.w2(32'hbbb4f9ec),
	.w3(32'hbb16e9c4),
	.w4(32'hbb16d4e7),
	.w5(32'hbbee7aa8),
	.w6(32'hb9370d08),
	.w7(32'h3a5237a8),
	.w8(32'hbb252e79),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06c07b),
	.w1(32'h39e2d664),
	.w2(32'hba493f02),
	.w3(32'hba9dc6cf),
	.w4(32'h3a83c787),
	.w5(32'hb8b65ce4),
	.w6(32'h392a7a1a),
	.w7(32'h3b21db19),
	.w8(32'h3a98783b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3ab79),
	.w1(32'h3b529dd5),
	.w2(32'hbbac30f6),
	.w3(32'h3b1774e5),
	.w4(32'h3b38f4b2),
	.w5(32'hbac27aa4),
	.w6(32'h3bc03945),
	.w7(32'h3bb34e92),
	.w8(32'hba162b19),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d39b9),
	.w1(32'h3a4a2412),
	.w2(32'hb8626660),
	.w3(32'h3a79cd75),
	.w4(32'h3a172df9),
	.w5(32'hb9040a9c),
	.w6(32'h3a48e073),
	.w7(32'h3a25259e),
	.w8(32'h394a7db0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38273d1f),
	.w1(32'hb9e370b3),
	.w2(32'hb97e86e6),
	.w3(32'h39b52899),
	.w4(32'hb9d61108),
	.w5(32'hb95dfcc2),
	.w6(32'hba640f72),
	.w7(32'hba7527b4),
	.w8(32'hba0cdb69),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fd3ff0),
	.w1(32'hba31048e),
	.w2(32'hba16a0b7),
	.w3(32'hb7f06fc6),
	.w4(32'hba3e43fc),
	.w5(32'hba04677b),
	.w6(32'hba676c90),
	.w7(32'hba8b77fd),
	.w8(32'hba097f12),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2db563),
	.w1(32'hba4f90ac),
	.w2(32'hba43c50b),
	.w3(32'h3893b8fa),
	.w4(32'hb9813ce6),
	.w5(32'hba140cac),
	.w6(32'hbab2878b),
	.w7(32'hbab11864),
	.w8(32'hba63d3b9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37ff39),
	.w1(32'h3a1b8071),
	.w2(32'hb9046afd),
	.w3(32'hb91a13cb),
	.w4(32'h3a4bb40d),
	.w5(32'h39b1ebeb),
	.w6(32'h3a2d852b),
	.w7(32'h3a908f8d),
	.w8(32'h39e04f49),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e33de),
	.w1(32'hbad59144),
	.w2(32'hb9c91d37),
	.w3(32'h3a030f04),
	.w4(32'h3a91311a),
	.w5(32'h3a97e5ec),
	.w6(32'hbb4ec9f0),
	.w7(32'hbb90a79e),
	.w8(32'hbb47b80d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f2574),
	.w1(32'hbb300d03),
	.w2(32'hbb82c71a),
	.w3(32'hbaa92ac1),
	.w4(32'hbb096b42),
	.w5(32'hbb242e64),
	.w6(32'hbade150f),
	.w7(32'hbad44580),
	.w8(32'hbb635891),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d912f),
	.w1(32'hbb93bdf7),
	.w2(32'hbb859e79),
	.w3(32'hbb8b2f52),
	.w4(32'hbb0e64b6),
	.w5(32'hbb41e2f2),
	.w6(32'hbb7cc2eb),
	.w7(32'hbab8443f),
	.w8(32'hbb27de54),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29176e),
	.w1(32'hbabaf67b),
	.w2(32'hbb905ab9),
	.w3(32'h3a4f036a),
	.w4(32'hbacace27),
	.w5(32'hbb68861a),
	.w6(32'h3a53994b),
	.w7(32'h3a01c2f0),
	.w8(32'hbac5a358),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb057c3d),
	.w1(32'hba5dd512),
	.w2(32'hbb38d49f),
	.w3(32'hb9b3475e),
	.w4(32'hba5a2e9b),
	.w5(32'hbb256340),
	.w6(32'hbad316c9),
	.w7(32'hba7d8e9a),
	.w8(32'hba521eb2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c7023),
	.w1(32'hbb2cece1),
	.w2(32'hbb81a015),
	.w3(32'hb7eae711),
	.w4(32'hbb0cf502),
	.w5(32'hbb86913a),
	.w6(32'hbaf070d9),
	.w7(32'hbad77d70),
	.w8(32'hbae068f2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb540a52),
	.w1(32'hbb299cc4),
	.w2(32'hbac455c4),
	.w3(32'hbb155b06),
	.w4(32'hba66657b),
	.w5(32'hba3c74cd),
	.w6(32'hbb08e8e9),
	.w7(32'hba585bc1),
	.w8(32'hba87f0e2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5426d2),
	.w1(32'hb94b4ffe),
	.w2(32'h3988f1f6),
	.w3(32'h3a592fc2),
	.w4(32'hb93d3d43),
	.w5(32'h396e7dfa),
	.w6(32'hb99af996),
	.w7(32'h37d94196),
	.w8(32'hb9a4ee11),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39047d19),
	.w1(32'h3a104ec9),
	.w2(32'h3a5c8bb4),
	.w3(32'hb9a67916),
	.w4(32'h3a0c3b58),
	.w5(32'h3a4116f5),
	.w6(32'h3952abd5),
	.w7(32'h3a476c56),
	.w8(32'h3a303224),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da4da6),
	.w1(32'hba16b7cb),
	.w2(32'hbb3cd904),
	.w3(32'h3a021922),
	.w4(32'h393a15ce),
	.w5(32'hbb49fc30),
	.w6(32'hba2cb4ff),
	.w7(32'hb70cb39f),
	.w8(32'h3a05811e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a0ad5),
	.w1(32'hb93acdad),
	.w2(32'h39c53296),
	.w3(32'hba84a3c3),
	.w4(32'h3a852526),
	.w5(32'h3aa62453),
	.w6(32'h392e9d69),
	.w7(32'hb9ef6130),
	.w8(32'h3906544d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a357b12),
	.w1(32'h3a357225),
	.w2(32'h3a267f72),
	.w3(32'h3a146c25),
	.w4(32'h3a998a11),
	.w5(32'hb94e94b8),
	.w6(32'h3a2f9196),
	.w7(32'h3a552532),
	.w8(32'hb9c0cfa3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c69a9),
	.w1(32'h37a93791),
	.w2(32'hb95b4257),
	.w3(32'hba835653),
	.w4(32'hb9f8f420),
	.w5(32'hb85b1960),
	.w6(32'hbaaf6e9e),
	.w7(32'hba337b43),
	.w8(32'h370f9ffa),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a9cea),
	.w1(32'h3a510f28),
	.w2(32'hbaf0e4b7),
	.w3(32'h3b18b3c6),
	.w4(32'h39b01b48),
	.w5(32'hbb253b46),
	.w6(32'h3a9d064b),
	.w7(32'h3aa10cc4),
	.w8(32'hb9dcb2c3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e641c),
	.w1(32'hbb12fb99),
	.w2(32'hbb01a74f),
	.w3(32'hbb791a6c),
	.w4(32'hba743c8a),
	.w5(32'hbafcfc61),
	.w6(32'hbba0c50c),
	.w7(32'hbb27c35a),
	.w8(32'hbac899f2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa64f0),
	.w1(32'hb993dcf9),
	.w2(32'hb96b6bb7),
	.w3(32'hba3f2413),
	.w4(32'h390603dd),
	.w5(32'h38f1f631),
	.w6(32'hbad19f51),
	.w7(32'hb7d7b9ac),
	.w8(32'hb916c427),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96e7cc),
	.w1(32'h39be2b62),
	.w2(32'hba943a0c),
	.w3(32'hb95ee863),
	.w4(32'hba282db4),
	.w5(32'hbb0982da),
	.w6(32'h3ab965ae),
	.w7(32'h39d51863),
	.w8(32'hba8b99a0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e3e2d),
	.w1(32'h3b167e7a),
	.w2(32'h3a8b2e5c),
	.w3(32'h3b29e6ec),
	.w4(32'h3b30fc40),
	.w5(32'h3ace9271),
	.w6(32'h3b424270),
	.w7(32'h3b5c25b8),
	.w8(32'h3b3c637b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ab58a),
	.w1(32'h39d4f724),
	.w2(32'hbb80c73b),
	.w3(32'h3b987d4a),
	.w4(32'h3a96be5b),
	.w5(32'hbb4ef0ba),
	.w6(32'h3b22703e),
	.w7(32'h3ae3aeb0),
	.w8(32'hba89f17a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaca254),
	.w1(32'h3af6a550),
	.w2(32'hb9ee3488),
	.w3(32'h3ad26dba),
	.w4(32'h3ad00170),
	.w5(32'hb9abdf10),
	.w6(32'h3b08fafe),
	.w7(32'h3ac773ec),
	.w8(32'hba102493),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1edf9),
	.w1(32'hb91d75f5),
	.w2(32'h3a8bd76f),
	.w3(32'h3a923ee3),
	.w4(32'h3ac4c9ae),
	.w5(32'h3a59a140),
	.w6(32'hb98feb21),
	.w7(32'h3a99a957),
	.w8(32'hba0c1c4d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e8ceb),
	.w1(32'hbb02a71b),
	.w2(32'hba935178),
	.w3(32'h3b2866a4),
	.w4(32'hbaa970c9),
	.w5(32'h39902cf8),
	.w6(32'hbae50364),
	.w7(32'hbab55cca),
	.w8(32'h38caea11),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a984db4),
	.w1(32'h3aafdc7d),
	.w2(32'hbb41a7f6),
	.w3(32'h3b64bd62),
	.w4(32'h3b032182),
	.w5(32'hbb5231f5),
	.w6(32'h3b36376e),
	.w7(32'h3b239183),
	.w8(32'hbb41980d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b476a9d),
	.w1(32'h3ae0f4e5),
	.w2(32'h3a7147b3),
	.w3(32'h3adb765c),
	.w4(32'h3b553eb1),
	.w5(32'h3b115003),
	.w6(32'hba1a9138),
	.w7(32'h3abf6a23),
	.w8(32'h399e671e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a015402),
	.w1(32'h3a04b022),
	.w2(32'hbae4176d),
	.w3(32'hba2e6a53),
	.w4(32'hba2748d5),
	.w5(32'hbb122cf1),
	.w6(32'hbb2ad9d9),
	.w7(32'hbaa2233a),
	.w8(32'hbb6ed249),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a792e49),
	.w1(32'h3bf98f8c),
	.w2(32'h3b8b4856),
	.w3(32'h3984d484),
	.w4(32'h3bd2adf6),
	.w5(32'h3b31377a),
	.w6(32'h3b3eec68),
	.w7(32'h3b7295e2),
	.w8(32'hb87b55ed),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37725d),
	.w1(32'hba88976f),
	.w2(32'hbbc32611),
	.w3(32'h3b2f7592),
	.w4(32'h3a3c0538),
	.w5(32'hbb4371d5),
	.w6(32'h3b294dd0),
	.w7(32'hb9a685f1),
	.w8(32'hbb32f205),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b338909),
	.w1(32'h399afc77),
	.w2(32'hbb40143c),
	.w3(32'h3b422056),
	.w4(32'h3aa4386b),
	.w5(32'hbafa46f1),
	.w6(32'h3a9649a6),
	.w7(32'h3a5ddbe4),
	.w8(32'hba6e9519),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8d90a),
	.w1(32'h3aa442b3),
	.w2(32'hba489869),
	.w3(32'h3a995be8),
	.w4(32'h3a82a148),
	.w5(32'h392d7193),
	.w6(32'hba36a65b),
	.w7(32'hbaa69482),
	.w8(32'hbb2137d9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb199b7a),
	.w1(32'hbb82862b),
	.w2(32'hbbaf21f6),
	.w3(32'hbaafc7ec),
	.w4(32'hbb0a09c0),
	.w5(32'hbb9d47a2),
	.w6(32'hbac28787),
	.w7(32'hbafda719),
	.w8(32'hbacdc952),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb099466),
	.w1(32'hba83b015),
	.w2(32'hbb02b7aa),
	.w3(32'hbaecb255),
	.w4(32'hba52beae),
	.w5(32'hba7177e1),
	.w6(32'hba2941b4),
	.w7(32'h3a14716c),
	.w8(32'hb94358e0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bb6e9),
	.w1(32'h391bd529),
	.w2(32'hb9e9b34a),
	.w3(32'hb9d72752),
	.w4(32'hb70cc29f),
	.w5(32'h389e2ef9),
	.w6(32'hba5cd1ea),
	.w7(32'hba0a96ea),
	.w8(32'h39b80291),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba933dd6),
	.w1(32'hb9d03872),
	.w2(32'hb9b6a8c2),
	.w3(32'h388c68e0),
	.w4(32'h394c94d3),
	.w5(32'h3a2d4d4e),
	.w6(32'hbadc2283),
	.w7(32'hbabaa7f1),
	.w8(32'hba38b668),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac58f67),
	.w1(32'hbaad801f),
	.w2(32'hbb532e53),
	.w3(32'h3a2397c3),
	.w4(32'hba3b4100),
	.w5(32'hbb17d2de),
	.w6(32'hbb5e8424),
	.w7(32'hbb4299bc),
	.w8(32'hbb745e1b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e5741),
	.w1(32'hb9934138),
	.w2(32'hbae2f1c6),
	.w3(32'h3a9e797c),
	.w4(32'h3adb51a6),
	.w5(32'hbb1e391b),
	.w6(32'h3ab36589),
	.w7(32'h3ac0d9fa),
	.w8(32'hbaf73c00),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42de25),
	.w1(32'h393f599a),
	.w2(32'hba08ba9d),
	.w3(32'h39e1280b),
	.w4(32'h39a9f900),
	.w5(32'hb9d33145),
	.w6(32'hbac78dc9),
	.w7(32'hba1d88b7),
	.w8(32'hbb1e0db2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947879d),
	.w1(32'h3a241f25),
	.w2(32'h39b32cd1),
	.w3(32'hbabb1751),
	.w4(32'hb931434f),
	.w5(32'hbb3aa2fb),
	.w6(32'h3a6f97ec),
	.w7(32'h3a50b46e),
	.w8(32'hb8c6fe52),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed0674),
	.w1(32'hba345f1f),
	.w2(32'hba8408b2),
	.w3(32'hbb26e817),
	.w4(32'hba1db1d5),
	.w5(32'hb9bdabc6),
	.w6(32'hba91f43b),
	.w7(32'h39865d00),
	.w8(32'h39a719d0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf75b2),
	.w1(32'hbafac3cd),
	.w2(32'hbb8c0486),
	.w3(32'hbae37406),
	.w4(32'hbae3b692),
	.w5(32'hbb74ab20),
	.w6(32'hba6d99d0),
	.w7(32'hbb165882),
	.w8(32'hbb8622a4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac24642),
	.w1(32'hba9ebac5),
	.w2(32'hbb18a5c2),
	.w3(32'hb9e6d2f0),
	.w4(32'hba4a6a8c),
	.w5(32'hbb56e7a9),
	.w6(32'hba963cd9),
	.w7(32'hba1f3ce1),
	.w8(32'hbb180285),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab240a),
	.w1(32'hba822c4b),
	.w2(32'hba91ab1d),
	.w3(32'hbae8d571),
	.w4(32'hba836199),
	.w5(32'hba7aac05),
	.w6(32'hbaa142e8),
	.w7(32'hbac39c53),
	.w8(32'hba14bd5b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f59b63),
	.w1(32'hb981c7de),
	.w2(32'hb930a1f9),
	.w3(32'hb999eb57),
	.w4(32'hb98c49af),
	.w5(32'hb9ba81cf),
	.w6(32'hba23e751),
	.w7(32'hba29c4d0),
	.w8(32'hb8edafbd),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9d9a2),
	.w1(32'hb876d247),
	.w2(32'hb8f768c4),
	.w3(32'h3809f5e0),
	.w4(32'hb72ba9b1),
	.w5(32'hb96eb9cf),
	.w6(32'hba3fddbd),
	.w7(32'hba0da707),
	.w8(32'h3774f7f2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39831709),
	.w1(32'h38941aa9),
	.w2(32'hba94c9ce),
	.w3(32'h38e07371),
	.w4(32'hba0362c8),
	.w5(32'hb95401fd),
	.w6(32'h382df112),
	.w7(32'hba33b26d),
	.w8(32'hb9f7a09d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b082b),
	.w1(32'hba22e497),
	.w2(32'hbb9058b1),
	.w3(32'hba136cb0),
	.w4(32'hb9aef1d6),
	.w5(32'hbb62a4ec),
	.w6(32'h3aec8a03),
	.w7(32'h3a3b4357),
	.w8(32'hbad4316c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ca0fa),
	.w1(32'hb9947e9e),
	.w2(32'hb8e57b81),
	.w3(32'h3ac24b69),
	.w4(32'h3a24b156),
	.w5(32'h3a1c5f81),
	.w6(32'hb9d355bc),
	.w7(32'h3984f099),
	.w8(32'h398f36ec),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cec2b),
	.w1(32'hba83455f),
	.w2(32'hbaba4287),
	.w3(32'hb9933871),
	.w4(32'h39bf47ea),
	.w5(32'hba809fd9),
	.w6(32'hba4d48bb),
	.w7(32'h3a0579cd),
	.w8(32'hba78d24f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08ee70),
	.w1(32'hba00349f),
	.w2(32'h3a429022),
	.w3(32'hbaf5edcf),
	.w4(32'hba92c8c5),
	.w5(32'h3a1060fd),
	.w6(32'hbb634ab4),
	.w7(32'hbb33ba5f),
	.w8(32'hbad86ab5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85e5c81),
	.w1(32'hb9e539df),
	.w2(32'hb48fb0db),
	.w3(32'hb974d6aa),
	.w4(32'h3a2e16c2),
	.w5(32'h3a042ca8),
	.w6(32'h3ae0ab36),
	.w7(32'h3a1b24a0),
	.w8(32'h3a9c41eb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad05c29),
	.w1(32'hba65828c),
	.w2(32'h3aeaba0e),
	.w3(32'hb8f82e20),
	.w4(32'hb96ad04c),
	.w5(32'h3aad2497),
	.w6(32'hbaa159cc),
	.w7(32'h3a84586f),
	.w8(32'h39a9fe0f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a978c3d),
	.w1(32'hba1fc7e3),
	.w2(32'hba0b137e),
	.w3(32'h3b0750b5),
	.w4(32'hb8d3334a),
	.w5(32'h38386511),
	.w6(32'hbace2358),
	.w7(32'hba91d076),
	.w8(32'hb93f1ef7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94938bf),
	.w1(32'hba1f7183),
	.w2(32'hb9c16353),
	.w3(32'h3a0a343b),
	.w4(32'h391dc6ca),
	.w5(32'h3946e794),
	.w6(32'hba0f0a0d),
	.w7(32'hb9925857),
	.w8(32'hb9be61ac),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab562bf),
	.w1(32'hba973622),
	.w2(32'hbb1f163b),
	.w3(32'hba407d3d),
	.w4(32'hbaad9cb1),
	.w5(32'hbb49b455),
	.w6(32'hb92bb742),
	.w7(32'hb9b1e176),
	.w8(32'hbad7ba82),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba901e66),
	.w1(32'hbb0d7fd2),
	.w2(32'hbb66113f),
	.w3(32'h3998cd01),
	.w4(32'hba20512d),
	.w5(32'hbb378936),
	.w6(32'h3a867b25),
	.w7(32'h3a8772f4),
	.w8(32'hbaa4f8e1),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3783ed93),
	.w1(32'h36b861dc),
	.w2(32'h36854a77),
	.w3(32'h379baf4c),
	.w4(32'hb6f475c2),
	.w5(32'hb680c25f),
	.w6(32'h37c3f447),
	.w7(32'hb709ded1),
	.w8(32'h3712e4c6),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68d033),
	.w1(32'hba3813f7),
	.w2(32'hba8a86c7),
	.w3(32'hbaa511bc),
	.w4(32'hba2bd302),
	.w5(32'hb9e5234c),
	.w6(32'hba471973),
	.w7(32'hba2a71ee),
	.w8(32'hba070b14),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bc3922),
	.w1(32'h3a4d79e5),
	.w2(32'h395118b3),
	.w3(32'hb9c972ff),
	.w4(32'hb892a4ee),
	.w5(32'hba501c46),
	.w6(32'hba283903),
	.w7(32'hb92d8480),
	.w8(32'hba638e47),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ad46c),
	.w1(32'hba484ef4),
	.w2(32'hbabc3482),
	.w3(32'h3933086a),
	.w4(32'hb698d59a),
	.w5(32'hba964c00),
	.w6(32'h37089aa6),
	.w7(32'h3867943c),
	.w8(32'hbaa4be67),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8c2ec),
	.w1(32'h39c17c18),
	.w2(32'hba65db0b),
	.w3(32'h37f20cd8),
	.w4(32'h3a04934d),
	.w5(32'hb9f3d2b6),
	.w6(32'h394afac2),
	.w7(32'h3a7cb58a),
	.w8(32'h3a12e760),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d1a92),
	.w1(32'hbb066775),
	.w2(32'hbb5a821a),
	.w3(32'hba9bdae6),
	.w4(32'hba79cd48),
	.w5(32'hbb57fb8b),
	.w6(32'hb9d4a760),
	.w7(32'h38524b93),
	.w8(32'hbb284284),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e964d),
	.w1(32'h3a39f4f1),
	.w2(32'hb9d21d00),
	.w3(32'h3a272bb5),
	.w4(32'h3a4a29bd),
	.w5(32'hb8bd4ee5),
	.w6(32'h3a2a5edc),
	.w7(32'h3a779137),
	.w8(32'hb842ef4b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fd3ac),
	.w1(32'hba436d70),
	.w2(32'hbac22848),
	.w3(32'h3804923f),
	.w4(32'h3a232cfb),
	.w5(32'hb99084f4),
	.w6(32'h3aa2b9a1),
	.w7(32'h3b03db65),
	.w8(32'h3948c6d3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ccd9c5),
	.w1(32'hb908544e),
	.w2(32'hbaf01cee),
	.w3(32'h389cda99),
	.w4(32'h39ff8200),
	.w5(32'hbb0b11ef),
	.w6(32'hb9b6dffc),
	.w7(32'h39f55c16),
	.w8(32'hbaba549f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ea8c66),
	.w1(32'h398e7f02),
	.w2(32'hba1e26d2),
	.w3(32'hb9949f26),
	.w4(32'h390b43a6),
	.w5(32'hb996f22c),
	.w6(32'hb90499e5),
	.w7(32'h39e31cdd),
	.w8(32'hb95b00ad),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89ee5a),
	.w1(32'h39b2b451),
	.w2(32'hbaf1fc80),
	.w3(32'h3a7f2d57),
	.w4(32'h3a002c43),
	.w5(32'hbabc9e23),
	.w6(32'h3a97a4cc),
	.w7(32'h3a07b77f),
	.w8(32'hba926247),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30549e),
	.w1(32'hba031df0),
	.w2(32'hba70d972),
	.w3(32'hb93382f3),
	.w4(32'hb7eb76be),
	.w5(32'hba430f85),
	.w6(32'hb9a38f09),
	.w7(32'hb919ce9b),
	.w8(32'hba44a2fa),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14b95b),
	.w1(32'h3a406769),
	.w2(32'h387d220a),
	.w3(32'hba4b0b9c),
	.w4(32'h3a4d74cb),
	.w5(32'h3a57c7ba),
	.w6(32'h39fde7b8),
	.w7(32'hb91b02a2),
	.w8(32'hba783f29),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17218d),
	.w1(32'h3affb56f),
	.w2(32'h3ab64da5),
	.w3(32'h3b1a779e),
	.w4(32'h3b02c72c),
	.w5(32'h3a86f261),
	.w6(32'h3b0500a2),
	.w7(32'h3acf9180),
	.w8(32'h396fa7d5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3795ea33),
	.w1(32'h3791c597),
	.w2(32'h378a76b8),
	.w3(32'h3701a1cc),
	.w4(32'h373593cb),
	.w5(32'h37fd36b4),
	.w6(32'h36aaae40),
	.w7(32'h379e04a7),
	.w8(32'h37ad4244),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bb4f8f),
	.w1(32'h3719ac42),
	.w2(32'h376bd5ff),
	.w3(32'h380e3b81),
	.w4(32'h379c3c93),
	.w5(32'h374ddd9c),
	.w6(32'h37e9bd96),
	.w7(32'h37933a22),
	.w8(32'h36a7d714),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f431a7),
	.w1(32'hb9d01723),
	.w2(32'hba775f5d),
	.w3(32'hba16eed9),
	.w4(32'hb8dac8a7),
	.w5(32'hb923e393),
	.w6(32'hb9b4c4bf),
	.w7(32'hb9db14ea),
	.w8(32'hb9f17adf),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18aefd),
	.w1(32'h3b00d676),
	.w2(32'hb8f5e204),
	.w3(32'h3b1e7634),
	.w4(32'h3b573595),
	.w5(32'h3a548eb8),
	.w6(32'h3b52908b),
	.w7(32'h3b7abcde),
	.w8(32'h3a979d17),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88379b),
	.w1(32'hbb796cf3),
	.w2(32'hbb531c8c),
	.w3(32'hbb86ced0),
	.w4(32'hbb1bf5b5),
	.w5(32'hbb0b4848),
	.w6(32'hbb9f799c),
	.w7(32'hbb532ec9),
	.w8(32'hbb451ee5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37937a6d),
	.w1(32'hb666e0cf),
	.w2(32'h364bab46),
	.w3(32'h37a4479d),
	.w4(32'hb5bda7d6),
	.w5(32'h341a3db3),
	.w6(32'h37ee2b89),
	.w7(32'h36f4f183),
	.w8(32'hb683f025),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba913ad2),
	.w1(32'hbadeee4b),
	.w2(32'hbb6dd7bb),
	.w3(32'h3951d567),
	.w4(32'hba0e28d6),
	.w5(32'hbb4d24e7),
	.w6(32'hba1899d1),
	.w7(32'hb886a965),
	.w8(32'hbaf776d1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c52c8),
	.w1(32'hb9ce756d),
	.w2(32'hba9ebb39),
	.w3(32'h3a334922),
	.w4(32'hb9816357),
	.w5(32'hbaa9ee95),
	.w6(32'h38b84edc),
	.w7(32'hb952404a),
	.w8(32'hba7c513c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60af0b),
	.w1(32'hbb70d7e1),
	.w2(32'hbba5614f),
	.w3(32'hbb2d0fe3),
	.w4(32'hbaebbda4),
	.w5(32'hbb6c4213),
	.w6(32'hbb17a5b8),
	.w7(32'hba48b570),
	.w8(32'hbb0362ea),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac78f05),
	.w1(32'h3a7fa85f),
	.w2(32'hbb093500),
	.w3(32'h3a64e90f),
	.w4(32'h3a37ac58),
	.w5(32'hbb023df0),
	.w6(32'h3adf7a65),
	.w7(32'h3af92760),
	.w8(32'hb985317f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b333ad5),
	.w1(32'h3b6cc5e5),
	.w2(32'h3b2c55ff),
	.w3(32'h3ae8c4c0),
	.w4(32'h3b0c69cf),
	.w5(32'h3ad7293c),
	.w6(32'h3a7d4206),
	.w7(32'h3a71e3a7),
	.w8(32'h382fa009),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3829f1),
	.w1(32'h3af617c0),
	.w2(32'h3ab992be),
	.w3(32'h3b5e1a86),
	.w4(32'h3b16690c),
	.w5(32'h3ae6a6aa),
	.w6(32'h3b3c7fb8),
	.w7(32'h3aa755b9),
	.w8(32'h3a20d5e7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb5fb7),
	.w1(32'hba4fc8fe),
	.w2(32'hbb45c51a),
	.w3(32'hb739ec58),
	.w4(32'h39c8b772),
	.w5(32'hbb1e8ed2),
	.w6(32'h3a2b7511),
	.w7(32'h3ac7a710),
	.w8(32'hba251d96),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b334472),
	.w1(32'h3b814b90),
	.w2(32'h3b271193),
	.w3(32'h3b74abc4),
	.w4(32'h3b8d4275),
	.w5(32'h3b45316c),
	.w6(32'h3b72edae),
	.w7(32'h3b91577b),
	.w8(32'h3b31decb),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37acb565),
	.w1(32'h3a210327),
	.w2(32'h3a97118f),
	.w3(32'hb9f05101),
	.w4(32'h394def4c),
	.w5(32'h3a4c5a2a),
	.w6(32'hb9c5ee18),
	.w7(32'h3a14a5af),
	.w8(32'h3a8946ca),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9403de6),
	.w1(32'hb9871614),
	.w2(32'hb98f281f),
	.w3(32'hb9235c74),
	.w4(32'hb9eaeea2),
	.w5(32'hb9fed585),
	.w6(32'hb98fce39),
	.w7(32'hb921d59a),
	.w8(32'hb9aeb558),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ed1892),
	.w1(32'h37b0ae06),
	.w2(32'hb81971fd),
	.w3(32'h38c0b335),
	.w4(32'hb873a070),
	.w5(32'hb8c0936e),
	.w6(32'hb8c438bd),
	.w7(32'hb97c9ebe),
	.w8(32'hb995e825),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380e1bbf),
	.w1(32'hb86a0d06),
	.w2(32'hbab1fc3f),
	.w3(32'h3982ef87),
	.w4(32'h394528b6),
	.w5(32'hbaa3fa99),
	.w6(32'h3809da40),
	.w7(32'h3a18c61f),
	.w8(32'hba3ab4a8),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d20d6d),
	.w1(32'hb882b657),
	.w2(32'hb623d5a1),
	.w3(32'hb793274b),
	.w4(32'hb83610e8),
	.w5(32'hb639c76d),
	.w6(32'h37a66f93),
	.w7(32'hb750e1bf),
	.w8(32'hb6ea57ad),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b7546),
	.w1(32'h39fceeb7),
	.w2(32'hba568f3a),
	.w3(32'h3a4c98ad),
	.w4(32'h39f0a61b),
	.w5(32'hba526763),
	.w6(32'h3a8e4c74),
	.w7(32'h3aaa68bf),
	.w8(32'h396a63ed),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391bda04),
	.w1(32'h3959c35b),
	.w2(32'hb93be948),
	.w3(32'h371c4571),
	.w4(32'h399462f7),
	.w5(32'hb88eea3c),
	.w6(32'h391bc101),
	.w7(32'h39c173a5),
	.w8(32'h39960d7d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3adff8),
	.w1(32'hbacb6e70),
	.w2(32'hb9d998de),
	.w3(32'hbb7f3625),
	.w4(32'hbaf9dd43),
	.w5(32'hbab915d2),
	.w6(32'hbac80798),
	.w7(32'hba10e185),
	.w8(32'hba91ea94),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390eef6f),
	.w1(32'h396784f7),
	.w2(32'h38ea49e4),
	.w3(32'h377809d7),
	.w4(32'h3985bf33),
	.w5(32'h3949d3e8),
	.w6(32'h38ec00dc),
	.w7(32'h397bb773),
	.w8(32'h397d588e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39676538),
	.w1(32'h3947c2fb),
	.w2(32'h38eab624),
	.w3(32'h396b92da),
	.w4(32'h3997be6f),
	.w5(32'h39e763dc),
	.w6(32'h36d15389),
	.w7(32'hb76c7df1),
	.w8(32'h399f631f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e2778),
	.w1(32'h3b05c844),
	.w2(32'hba72aff9),
	.w3(32'h3b4685bd),
	.w4(32'h3b49786c),
	.w5(32'h394c79ec),
	.w6(32'h3b4d37c7),
	.w7(32'h3b256c50),
	.w8(32'hb9b7bbe1),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0309d3),
	.w1(32'hbaaceaa0),
	.w2(32'hbb94f8e2),
	.w3(32'hba34fc1a),
	.w4(32'hbb1e5c92),
	.w5(32'hbbe1536b),
	.w6(32'h3a4561d4),
	.w7(32'h3a5369a6),
	.w8(32'hbb4a79b4),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a0f5bb),
	.w1(32'h3a0353df),
	.w2(32'h3a20324b),
	.w3(32'hba63e8c6),
	.w4(32'hb9bb1862),
	.w5(32'hb916a526),
	.w6(32'hba76b197),
	.w7(32'hb920032a),
	.w8(32'h3a29bcb6),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba712fdd),
	.w1(32'h38e53880),
	.w2(32'hbace0b5d),
	.w3(32'hba66852c),
	.w4(32'h3a32dc27),
	.w5(32'hba3f2501),
	.w6(32'hba4f1c7f),
	.w7(32'h3a045385),
	.w8(32'hba9164ec),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ed8421),
	.w1(32'h38ecdf9b),
	.w2(32'h38589289),
	.w3(32'hb8f5a170),
	.w4(32'h39a0e1e2),
	.w5(32'h3981a61a),
	.w6(32'hb994d623),
	.w7(32'h3819caaa),
	.w8(32'hb88aa161),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57a100),
	.w1(32'hbb4b121c),
	.w2(32'hbb9c8a03),
	.w3(32'hb9e28e1a),
	.w4(32'hba35cc80),
	.w5(32'hbb42d167),
	.w6(32'h3a2efc73),
	.w7(32'h3ae704a1),
	.w8(32'hbb00d08d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba182fa7),
	.w1(32'hb9a405a5),
	.w2(32'hbaacf75f),
	.w3(32'hb9aab5f8),
	.w4(32'hb9029890),
	.w5(32'hbab30698),
	.w6(32'hb9bf5a9c),
	.w7(32'h3a097f02),
	.w8(32'hba1f0b74),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1628a3),
	.w1(32'hbb1e6aee),
	.w2(32'hbb8f3b03),
	.w3(32'hba6bd136),
	.w4(32'hba924bcc),
	.w5(32'hbb8fe6bb),
	.w6(32'hba03542c),
	.w7(32'hb9bd773c),
	.w8(32'hbb56967c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9cac7),
	.w1(32'h3a178f3e),
	.w2(32'hb8a8b41a),
	.w3(32'h39b7fd10),
	.w4(32'h3a486915),
	.w5(32'h3941ae23),
	.w6(32'h3a36e820),
	.w7(32'h3a6a0607),
	.w8(32'h3a092d94),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0da8e),
	.w1(32'h3a1a7442),
	.w2(32'hbae4f016),
	.w3(32'h3b034d97),
	.w4(32'h3a4ada3e),
	.w5(32'hbaf15fe7),
	.w6(32'h3b0d86f2),
	.w7(32'h3ab851b4),
	.w8(32'hba33b5eb),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382cabb7),
	.w1(32'h37292215),
	.w2(32'h379c94f1),
	.w3(32'h37accdf6),
	.w4(32'h3555e3b3),
	.w5(32'h378fbea7),
	.w6(32'h36ead8e6),
	.w7(32'hb7aa3dd8),
	.w8(32'h36c74108),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88d0c08),
	.w1(32'hb9dddd82),
	.w2(32'hba58be58),
	.w3(32'hb9223928),
	.w4(32'hb9c1daa8),
	.w5(32'hba304468),
	.w6(32'hb8b143e3),
	.w7(32'hba0f9a40),
	.w8(32'hba615040),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac667f),
	.w1(32'h39cee208),
	.w2(32'hb8d34054),
	.w3(32'h397ea00c),
	.w4(32'h39a248dc),
	.w5(32'hb81e22cd),
	.w6(32'h3916eb6d),
	.w7(32'hb7550e02),
	.w8(32'hb944b301),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07cad3),
	.w1(32'hbaff134d),
	.w2(32'hbb263533),
	.w3(32'hba8ec66d),
	.w4(32'hbab83f25),
	.w5(32'hbaecf705),
	.w6(32'hbb13f065),
	.w7(32'hbad37744),
	.w8(32'hbb0dc790),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379301f0),
	.w1(32'h3608a39d),
	.w2(32'h360ff400),
	.w3(32'h378ff4c8),
	.w4(32'h362cb5a4),
	.w5(32'hb4e91ce1),
	.w6(32'h3761758e),
	.w7(32'h36cd2d9c),
	.w8(32'h365b53c7),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39411434),
	.w1(32'h39cf81b6),
	.w2(32'h393c82ea),
	.w3(32'h392e63e9),
	.w4(32'h39ab1043),
	.w5(32'h39412825),
	.w6(32'h38d1e8c2),
	.w7(32'h39444e4b),
	.w8(32'hb8193297),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c4dba),
	.w1(32'h38076f18),
	.w2(32'h38270070),
	.w3(32'hba65c060),
	.w4(32'hb8b5c60e),
	.w5(32'hb8bb6855),
	.w6(32'hba13dea5),
	.w7(32'h38d068e2),
	.w8(32'h376302df),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952cf9d),
	.w1(32'h3a3a4f62),
	.w2(32'hba699512),
	.w3(32'hba01c12b),
	.w4(32'h3a233ae9),
	.w5(32'hba32762a),
	.w6(32'hb8f9fab3),
	.w7(32'h3a2e172a),
	.w8(32'hb99e9ea0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a88442),
	.w1(32'h35abe264),
	.w2(32'h37e57108),
	.w3(32'h393d2721),
	.w4(32'h38b0ab3a),
	.w5(32'h368b7b4a),
	.w6(32'h39869a84),
	.w7(32'h392c186c),
	.w8(32'h387e0f74),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a17a58),
	.w1(32'hb9aa57fc),
	.w2(32'hba055237),
	.w3(32'hb9c4a8a0),
	.w4(32'hb9e90640),
	.w5(32'hb9fe0d02),
	.w6(32'hb89528f9),
	.w7(32'hb8fe5a8c),
	.w8(32'hb9ba766a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6b798),
	.w1(32'hbb9dabbe),
	.w2(32'hbc23087e),
	.w3(32'hbb4e1cba),
	.w4(32'hbabd7a7f),
	.w5(32'hbbb79634),
	.w6(32'h3b21356f),
	.w7(32'h3b750ddc),
	.w8(32'hbb65559c),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2fccf),
	.w1(32'h3b24d653),
	.w2(32'h3a0e039b),
	.w3(32'h3b2e2f5a),
	.w4(32'h3b7c7dc7),
	.w5(32'h3a6ad12a),
	.w6(32'h3b5668a8),
	.w7(32'h3b8628cf),
	.w8(32'h3a1e662f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de992e),
	.w1(32'h399ae62e),
	.w2(32'hb85db82d),
	.w3(32'h39a2d317),
	.w4(32'h39497e29),
	.w5(32'h38944d7d),
	.w6(32'h3967d3f4),
	.w7(32'h39271934),
	.w8(32'h37d2cbc2),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f77d41),
	.w1(32'hb826a29b),
	.w2(32'hb7e099db),
	.w3(32'hb826a614),
	.w4(32'hb87f93c7),
	.w5(32'hb7cb8e64),
	.w6(32'hb8befd2c),
	.w7(32'hb89fc579),
	.w8(32'hb84dfe82),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923cdef),
	.w1(32'h3862e60e),
	.w2(32'h3965d587),
	.w3(32'h390e905b),
	.w4(32'h38ce5b63),
	.w5(32'h39558ae8),
	.w6(32'hb81f451a),
	.w7(32'hb90d1305),
	.w8(32'hb9306f5e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388439e9),
	.w1(32'h37c9a098),
	.w2(32'h3807c1e1),
	.w3(32'h3865327e),
	.w4(32'h3776b386),
	.w5(32'h38017b0c),
	.w6(32'h3648233f),
	.w7(32'hb85f382c),
	.w8(32'hb74d000f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a961080),
	.w1(32'h3a801e77),
	.w2(32'hb89eac70),
	.w3(32'h3a30efab),
	.w4(32'h3a3aec22),
	.w5(32'hb91359a6),
	.w6(32'h39da81c3),
	.w7(32'h39439d5e),
	.w8(32'hb9a0d2b7),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fd984),
	.w1(32'h3b2ede1a),
	.w2(32'h3928e12f),
	.w3(32'h3a6d9f82),
	.w4(32'h3aa62503),
	.w5(32'hba88d451),
	.w6(32'h3a878cda),
	.w7(32'h3b1bc0a6),
	.w8(32'h39c4be0a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fcf82),
	.w1(32'hbb483529),
	.w2(32'hbb38cbdb),
	.w3(32'hba806331),
	.w4(32'hba4c55ea),
	.w5(32'hbafb7eb0),
	.w6(32'hbac3c007),
	.w7(32'hb8ebe980),
	.w8(32'hbb0ff2ce),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383e634d),
	.w1(32'hb85101fc),
	.w2(32'hb9063c74),
	.w3(32'hba706801),
	.w4(32'hba0ecbda),
	.w5(32'hb9d2a04d),
	.w6(32'hb9af7c8b),
	.w7(32'hb9f4d13a),
	.w8(32'hb9b8e2b3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb688899),
	.w1(32'hbb4a1c46),
	.w2(32'hbb9a8649),
	.w3(32'hbb38f433),
	.w4(32'hbabf1da9),
	.w5(32'hbb3f558e),
	.w6(32'hbb419001),
	.w7(32'hba768c47),
	.w8(32'hbb2e0dc0),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f11e8a),
	.w1(32'hba80be6c),
	.w2(32'hbab1dde2),
	.w3(32'hb9dfed6d),
	.w4(32'hba47dcbb),
	.w5(32'hba8d8d40),
	.w6(32'hba371f97),
	.w7(32'hba4d567c),
	.w8(32'hba0e89e8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f62384),
	.w1(32'h37c4aad9),
	.w2(32'h37c9df3a),
	.w3(32'h37a65596),
	.w4(32'h3778a5e1),
	.w5(32'h37a86157),
	.w6(32'h37d2342a),
	.w7(32'h37841b6c),
	.w8(32'h37d630fe),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7840a85),
	.w1(32'hb8788e03),
	.w2(32'hb869a99f),
	.w3(32'h38148e88),
	.w4(32'hb88c50a6),
	.w5(32'hb816066b),
	.w6(32'h38212531),
	.w7(32'hb7959fae),
	.w8(32'hb781328e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385a1250),
	.w1(32'h36b4fc5f),
	.w2(32'h382367e5),
	.w3(32'h3829a2ce),
	.w4(32'hb7751943),
	.w5(32'h37e6abf0),
	.w6(32'h382be87a),
	.w7(32'hb79b4aca),
	.w8(32'h3817bde5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacac704),
	.w1(32'hb9a7d820),
	.w2(32'hb9a2f103),
	.w3(32'hba0802bc),
	.w4(32'h3a00f85f),
	.w5(32'hba1ab712),
	.w6(32'hb901fe3e),
	.w7(32'hb983f57a),
	.w8(32'hba7c255b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ee7d6),
	.w1(32'h3b0d559e),
	.w2(32'h3b0a02f9),
	.w3(32'h3a4a26de),
	.w4(32'h3b155c1d),
	.w5(32'h3b040796),
	.w6(32'h3a84258f),
	.w7(32'h3b12a6d9),
	.w8(32'h3af901c6),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4e9b4),
	.w1(32'h39c6ad50),
	.w2(32'hba6fe439),
	.w3(32'h39bb596d),
	.w4(32'h3a3d8316),
	.w5(32'hba04db5f),
	.w6(32'h3a01f57c),
	.w7(32'h3a9b2041),
	.w8(32'h398bc7fd),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1f65d),
	.w1(32'hb889af22),
	.w2(32'hb8d85247),
	.w3(32'hba00bae7),
	.w4(32'hb9e2dedf),
	.w5(32'hb9131353),
	.w6(32'hb9fb8c0c),
	.w7(32'hb9fbec10),
	.w8(32'hb8fcd665),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39976d51),
	.w1(32'h39ffdd84),
	.w2(32'hba3c6ffa),
	.w3(32'hb70beb3c),
	.w4(32'h3a3c5745),
	.w5(32'hb948337e),
	.w6(32'hb99548be),
	.w7(32'h39a272ae),
	.w8(32'hba101fb6),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5fdd1),
	.w1(32'hb99807a3),
	.w2(32'hbad100af),
	.w3(32'h39ab4abf),
	.w4(32'h3a0a7d5e),
	.w5(32'hbac30c4e),
	.w6(32'h395e7e60),
	.w7(32'h3a005abd),
	.w8(32'hbaa3aa6d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa3797),
	.w1(32'hbbceeb39),
	.w2(32'hbbeca2fb),
	.w3(32'hbbb4936a),
	.w4(32'hbb8c6c39),
	.w5(32'hbbb0da3b),
	.w6(32'hbbb0562a),
	.w7(32'hbb42d27a),
	.w8(32'hbbd225c2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b090c8),
	.w1(32'hb7a7870e),
	.w2(32'hb77a9b18),
	.w3(32'h376a2e45),
	.w4(32'hb75d8d5f),
	.w5(32'hb7848c6b),
	.w6(32'h37b73656),
	.w7(32'hb724b264),
	.w8(32'hb6e8c4d1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d9a2bd),
	.w1(32'hb7402221),
	.w2(32'h37b4748f),
	.w3(32'h37814dc9),
	.w4(32'hb7aff606),
	.w5(32'h36fd8ce0),
	.w6(32'h383943d2),
	.w7(32'h3827bce4),
	.w8(32'h3674169c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5defbe),
	.w1(32'h378b8a2a),
	.w2(32'hbac37b9b),
	.w3(32'hba2f5d10),
	.w4(32'h39039f77),
	.w5(32'hbab4c5a3),
	.w6(32'h38ef8499),
	.w7(32'h3a978dfc),
	.w8(32'hba0cf296),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f8910),
	.w1(32'h3a720fa2),
	.w2(32'hbb38f14f),
	.w3(32'h3a5352e7),
	.w4(32'hb8f0f307),
	.w5(32'hbb9acf38),
	.w6(32'h3ab7a02a),
	.w7(32'h3b139ed2),
	.w8(32'hba0700ca),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4a995),
	.w1(32'hbb0234f0),
	.w2(32'hbb720839),
	.w3(32'hb92d01f8),
	.w4(32'hba7faabd),
	.w5(32'hbb5f5508),
	.w6(32'h3a61ecd5),
	.w7(32'h39d60b8d),
	.w8(32'hbb0c139d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8579b13),
	.w1(32'hb765d6d9),
	.w2(32'hb7829c6e),
	.w3(32'hb8af434f),
	.w4(32'hb8c6696c),
	.w5(32'hb88b0713),
	.w6(32'hb89ed8cb),
	.w7(32'hb8f04de2),
	.w8(32'hb8974ae2),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38376a73),
	.w1(32'h37d48ff1),
	.w2(32'h37f0807c),
	.w3(32'h386cc4dc),
	.w4(32'hb6c38716),
	.w5(32'h3741e2f9),
	.w6(32'h37b90e14),
	.w7(32'hb7f6852b),
	.w8(32'hb7288b16),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391fb877),
	.w1(32'h39b0e4fa),
	.w2(32'h39025e99),
	.w3(32'h38bcf2cc),
	.w4(32'h3926fe7a),
	.w5(32'h371f144a),
	.w6(32'hb83afc71),
	.w7(32'hb81ce01e),
	.w8(32'hb77d7c8a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d62ee0),
	.w1(32'hb955228f),
	.w2(32'hba18734e),
	.w3(32'hba6d2cd6),
	.w4(32'hba1657de),
	.w5(32'hba9ba61e),
	.w6(32'hb9ae0ae3),
	.w7(32'hb95e6113),
	.w8(32'hb9fede05),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc631ef),
	.w1(32'hbba3cf7d),
	.w2(32'hbbb9dac8),
	.w3(32'hbb8c0dbd),
	.w4(32'hbb5d679f),
	.w5(32'hbb9d3b75),
	.w6(32'hbb7c7a78),
	.w7(32'hba01c4d8),
	.w8(32'hbb2e54e1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a917c02),
	.w1(32'hb9ae0b8c),
	.w2(32'hbacfd531),
	.w3(32'h3a4bc712),
	.w4(32'h3a3c3c95),
	.w5(32'hb984cc86),
	.w6(32'hb931f3b4),
	.w7(32'hba2e656b),
	.w8(32'hba333629),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5552ef),
	.w1(32'h3af56687),
	.w2(32'h3a8ef981),
	.w3(32'h39890409),
	.w4(32'h3a9f1860),
	.w5(32'h3a283d85),
	.w6(32'h398d098d),
	.w7(32'h3a93c9f0),
	.w8(32'h3a079c40),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb056cb6),
	.w1(32'hba8e4d7a),
	.w2(32'hbb1f33b3),
	.w3(32'hba86fb1b),
	.w4(32'h394a77a1),
	.w5(32'hbac56451),
	.w6(32'h3916dbb9),
	.w7(32'h3abe4dcb),
	.w8(32'h390e4e9b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ac9a11),
	.w1(32'h376ce34d),
	.w2(32'h37a7f123),
	.w3(32'h378e6fec),
	.w4(32'h373bed64),
	.w5(32'h3798f1a9),
	.w6(32'h379fe058),
	.w7(32'h379401fe),
	.w8(32'h37df1145),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f140e9),
	.w1(32'hb71c992d),
	.w2(32'hb6728a24),
	.w3(32'hb6f498b8),
	.w4(32'hb765b0cb),
	.w5(32'hb6563b74),
	.w6(32'h34537b46),
	.w7(32'hb6d9caf9),
	.w8(32'h36733d7a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c871a4),
	.w1(32'h380b20aa),
	.w2(32'h378a8e0e),
	.w3(32'hb6e05234),
	.w4(32'h36f67eaf),
	.w5(32'hb59c1752),
	.w6(32'h3752f453),
	.w7(32'h371e808d),
	.w8(32'h36814533),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380070d6),
	.w1(32'h37125c3e),
	.w2(32'hb56ffbf9),
	.w3(32'h37d2b57b),
	.w4(32'h37852c03),
	.w5(32'h36be88b0),
	.w6(32'h371c7ddd),
	.w7(32'h36de33cf),
	.w8(32'h368073e2),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9060113),
	.w1(32'h391a70b1),
	.w2(32'h387fa0c0),
	.w3(32'hb98e7422),
	.w4(32'h368d94d6),
	.w5(32'hb8abb76f),
	.w6(32'hb9a93dee),
	.w7(32'hb7e5481f),
	.w8(32'hb70f8c7a),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c2063),
	.w1(32'h36df96ec),
	.w2(32'hbb27cf95),
	.w3(32'h3a674408),
	.w4(32'hb9df2e08),
	.w5(32'hbb723b3d),
	.w6(32'h3abe2ddb),
	.w7(32'h39eb5e5d),
	.w8(32'hbad67b79),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fb937),
	.w1(32'hb8b4020d),
	.w2(32'hbaa49c84),
	.w3(32'hba3bb095),
	.w4(32'hba4d6246),
	.w5(32'hba80fb31),
	.w6(32'hb8226c18),
	.w7(32'hb9804a2b),
	.w8(32'hba7ab2d9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74f9467),
	.w1(32'hb464fbcc),
	.w2(32'h37656ce8),
	.w3(32'hb7be8bf4),
	.w4(32'hb638a2c7),
	.w5(32'h3791c677),
	.w6(32'hb7c8547a),
	.w7(32'h36dcf622),
	.w8(32'h3699fb9e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb305071),
	.w1(32'hbb341613),
	.w2(32'hbb842a7d),
	.w3(32'hbb1f8107),
	.w4(32'hbadaca7c),
	.w5(32'hbb5d808d),
	.w6(32'hbb62e1fb),
	.w7(32'hbb15f971),
	.w8(32'hbb45b3d9),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0eda1c),
	.w1(32'hba2210b7),
	.w2(32'hbaa8f2fc),
	.w3(32'hb990dbf7),
	.w4(32'hba1b2c1d),
	.w5(32'hbaad773b),
	.w6(32'hb9f3e159),
	.w7(32'hba5046fc),
	.w8(32'hbaa79769),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8405f31),
	.w1(32'hb88df5dc),
	.w2(32'h3680eced),
	.w3(32'hb89929f0),
	.w4(32'hb8737d4f),
	.w5(32'hb7bb12d3),
	.w6(32'hb88b902a),
	.w7(32'hb868405a),
	.w8(32'h37dd1345),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba700e06),
	.w1(32'hba0034ba),
	.w2(32'hba927ca3),
	.w3(32'hba095690),
	.w4(32'hb93a2adf),
	.w5(32'hba4766f1),
	.w6(32'hba6a1f79),
	.w7(32'h38398ef0),
	.w8(32'hba31e892),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399151a6),
	.w1(32'h39a9c921),
	.w2(32'h39a36bde),
	.w3(32'h399ee22c),
	.w4(32'h39b9f7b5),
	.w5(32'h39a5920d),
	.w6(32'h39534fe0),
	.w7(32'h397856a9),
	.w8(32'h39596a9a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987419c),
	.w1(32'hb94254a9),
	.w2(32'hb9dee9ba),
	.w3(32'hb9ad195a),
	.w4(32'hb9240ea2),
	.w5(32'hb9d908ee),
	.w6(32'hb98f2bd3),
	.w7(32'hb8551241),
	.w8(32'hb9563220),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e82374),
	.w1(32'h379b1cc0),
	.w2(32'h35d80f54),
	.w3(32'h37c56223),
	.w4(32'h37062bf8),
	.w5(32'h34383fea),
	.w6(32'h3743dcca),
	.w7(32'h36a1c530),
	.w8(32'h3700b293),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3752511d),
	.w1(32'h36884d20),
	.w2(32'h38010e41),
	.w3(32'h37b661f6),
	.w4(32'h3790320a),
	.w5(32'h38200d41),
	.w6(32'h3806b596),
	.w7(32'h37f60efa),
	.w8(32'h383b9222),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94508d0),
	.w1(32'h39cc578a),
	.w2(32'h398784c1),
	.w3(32'hb98c8a94),
	.w4(32'h39afdeac),
	.w5(32'h38d83fac),
	.w6(32'hb8a401bf),
	.w7(32'h39e9519d),
	.w8(32'h39397d2e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba979d66),
	.w1(32'hbadc6454),
	.w2(32'hbb9ea0d0),
	.w3(32'h3861d0e2),
	.w4(32'hbac56594),
	.w5(32'hbba51b62),
	.w6(32'h3a0444aa),
	.w7(32'h39f1a827),
	.w8(32'hbb3646b2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39061da4),
	.w1(32'hb9865a04),
	.w2(32'hbb2bf183),
	.w3(32'h3a81aa79),
	.w4(32'h39a640c9),
	.w5(32'hbb15a355),
	.w6(32'h3aa54b5d),
	.w7(32'h3ab4dbf9),
	.w8(32'hba328f11),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb410941),
	.w1(32'hbb242a60),
	.w2(32'hbb668537),
	.w3(32'hbaa4176a),
	.w4(32'hba83671a),
	.w5(32'hbb5bbed7),
	.w6(32'hba489261),
	.w7(32'hb5b67de5),
	.w8(32'hbb232027),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3828d298),
	.w1(32'h389389f0),
	.w2(32'h38d3a9f6),
	.w3(32'hb76aa7c3),
	.w4(32'h3853338c),
	.w5(32'h38dd11f0),
	.w6(32'hb5f78474),
	.w7(32'h38a687cb),
	.w8(32'h38fff457),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3777a58d),
	.w1(32'h371dd41f),
	.w2(32'h374dbf40),
	.w3(32'hb64f7268),
	.w4(32'h3646443f),
	.w5(32'h37346684),
	.w6(32'h367e96d8),
	.w7(32'h34c090a2),
	.w8(32'h36ff80e8),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d37f18),
	.w1(32'hb803dfe0),
	.w2(32'hb811ea1b),
	.w3(32'h37f8c6a8),
	.w4(32'hb86cef9a),
	.w5(32'hb88a1640),
	.w6(32'h3840fee3),
	.w7(32'hb7ff89b6),
	.w8(32'hb894cee7),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e48dd6),
	.w1(32'h35161424),
	.w2(32'h37321e64),
	.w3(32'hb632e96f),
	.w4(32'h3608214c),
	.w5(32'h37950857),
	.w6(32'hb6ea0855),
	.w7(32'hb614c0d1),
	.w8(32'h37078a4a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae07f7d),
	.w1(32'h3a35de4a),
	.w2(32'hbac5db2c),
	.w3(32'h3b01e095),
	.w4(32'h3a767038),
	.w5(32'hba9646d0),
	.w6(32'h3adc5609),
	.w7(32'h3a83e9cc),
	.w8(32'hba2c383f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1663eb),
	.w1(32'hb9f7d454),
	.w2(32'hb9c2ce97),
	.w3(32'hba0aa8f8),
	.w4(32'hba1042f9),
	.w5(32'hba10fd1d),
	.w6(32'hba0b2a94),
	.w7(32'hba2ba849),
	.w8(32'hba68d593),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b19bde),
	.w1(32'h3924095b),
	.w2(32'h39f1e0f0),
	.w3(32'h39146b4d),
	.w4(32'hb90903c0),
	.w5(32'h39875797),
	.w6(32'h38de99a5),
	.w7(32'hb854a5d6),
	.w8(32'h3850ebb6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f773b2),
	.w1(32'h391ec32b),
	.w2(32'h399aafa5),
	.w3(32'hb9212cc7),
	.w4(32'h37ffb52f),
	.w5(32'h399000eb),
	.w6(32'hb95101bf),
	.w7(32'h390a7b5c),
	.w8(32'h39adb082),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d12c80),
	.w1(32'hb8146298),
	.w2(32'hb5ade5d4),
	.w3(32'h374967b4),
	.w4(32'hb614696d),
	.w5(32'hb720919b),
	.w6(32'h374944f8),
	.w7(32'h381e66d0),
	.w8(32'h382625bc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9741c1),
	.w1(32'hba916a1c),
	.w2(32'hb9de8d6e),
	.w3(32'hba3f03e3),
	.w4(32'hb9a0f3d7),
	.w5(32'hb936a19e),
	.w6(32'hba803d7a),
	.w7(32'hb9a5203c),
	.w8(32'hba4e88bb),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3737b03f),
	.w1(32'h3782b119),
	.w2(32'hb6de06e1),
	.w3(32'hb81447bd),
	.w4(32'hb7e57277),
	.w5(32'hb7a5c845),
	.w6(32'hb83cd7c6),
	.w7(32'hb7f61511),
	.w8(32'hb712e92d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f6992c),
	.w1(32'hba49a64a),
	.w2(32'hbb07fa94),
	.w3(32'h3a04a776),
	.w4(32'hb9d90eab),
	.w5(32'hba9b6ac9),
	.w6(32'h3a147413),
	.w7(32'h3a8967c6),
	.w8(32'h38ae6c1a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8942dc2),
	.w1(32'h3a2830b6),
	.w2(32'hbb6a7bb3),
	.w3(32'hb802ee54),
	.w4(32'h3b25e361),
	.w5(32'h39b7da59),
	.w6(32'h3bb4a149),
	.w7(32'h3b810a5f),
	.w8(32'h3b05955a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06a806),
	.w1(32'h3a448227),
	.w2(32'hb956904a),
	.w3(32'h3b585eb2),
	.w4(32'h3ad4353d),
	.w5(32'h3a293f01),
	.w6(32'h3b015be0),
	.w7(32'h3ba84350),
	.w8(32'h3b2b2a0a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule