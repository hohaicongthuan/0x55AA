module layer_10_featuremap_328(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1c337),
	.w1(32'h3ae66983),
	.w2(32'h3b9d04bf),
	.w3(32'h3b4636d0),
	.w4(32'h3b87bc44),
	.w5(32'h3856e90b),
	.w6(32'h3bb770e2),
	.w7(32'h3c027536),
	.w8(32'hba8f29f9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3763f),
	.w1(32'hbb92b886),
	.w2(32'h3acabf1b),
	.w3(32'h39ee4657),
	.w4(32'h3b9cd35c),
	.w5(32'h3bda3d4b),
	.w6(32'hb936455f),
	.w7(32'hba6b0745),
	.w8(32'h3b944f05),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3fa7e),
	.w1(32'h3afbdda2),
	.w2(32'h3b0dc064),
	.w3(32'hbb9a7b9d),
	.w4(32'hbb713863),
	.w5(32'hbb29883c),
	.w6(32'hbb1c9491),
	.w7(32'hbb502201),
	.w8(32'hbb370f48),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10f36c),
	.w1(32'hbac088ce),
	.w2(32'hba0304bf),
	.w3(32'hbafa32e5),
	.w4(32'hbabb522c),
	.w5(32'hbb12c130),
	.w6(32'hbb3fe3cc),
	.w7(32'hbad6cc58),
	.w8(32'hbbaf88ab),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b4b24),
	.w1(32'hbb29e957),
	.w2(32'h3a3f323d),
	.w3(32'hbaa319a9),
	.w4(32'h38ae2cc4),
	.w5(32'hbb305e60),
	.w6(32'hbb570e87),
	.w7(32'hbb33b597),
	.w8(32'hbb17f739),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e2d27),
	.w1(32'hba636080),
	.w2(32'h38fb6186),
	.w3(32'hba817525),
	.w4(32'hb9e30d78),
	.w5(32'hba7e1af0),
	.w6(32'h3a1add43),
	.w7(32'hba04946c),
	.w8(32'hb9912340),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e2a5e),
	.w1(32'hbbd6912e),
	.w2(32'hbbe2c7a2),
	.w3(32'h3ad44b25),
	.w4(32'hbac5cc30),
	.w5(32'hbbf64f23),
	.w6(32'hbb167e96),
	.w7(32'hbb9da2a1),
	.w8(32'hbbdb35dd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96ab80),
	.w1(32'hb95d3781),
	.w2(32'hbbc9a18e),
	.w3(32'hbb92cee1),
	.w4(32'hbb966a67),
	.w5(32'hbacc5d47),
	.w6(32'hbb02b683),
	.w7(32'hbbc2fd5e),
	.w8(32'hbb568ba5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc1c71),
	.w1(32'h3af105af),
	.w2(32'h3b038c74),
	.w3(32'h3adb08b8),
	.w4(32'h3b286379),
	.w5(32'hbb82a6be),
	.w6(32'h3b413cf9),
	.w7(32'h3b25af69),
	.w8(32'hbb55342e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb75193),
	.w1(32'hba008633),
	.w2(32'hbbad410c),
	.w3(32'hbb20d807),
	.w4(32'h3ab0e16a),
	.w5(32'hbb389bd0),
	.w6(32'hbbafe1c9),
	.w7(32'hbb124681),
	.w8(32'hbbad50fb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9a622),
	.w1(32'h3b2be62b),
	.w2(32'h3ad551d5),
	.w3(32'hba6ddd09),
	.w4(32'hb9dcda29),
	.w5(32'h3a528028),
	.w6(32'h3b44f051),
	.w7(32'hb8e0fbec),
	.w8(32'h3a4fc2f5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9008e1),
	.w1(32'h3bdbc25f),
	.w2(32'hbb45df09),
	.w3(32'hbba7bc7a),
	.w4(32'hbb5706af),
	.w5(32'hbb459cc8),
	.w6(32'hbc027a61),
	.w7(32'hbb0fc11f),
	.w8(32'hbbb0c1c8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a1492),
	.w1(32'hb9cabe7e),
	.w2(32'hbbf7a5ed),
	.w3(32'h3abe83a5),
	.w4(32'h3b489cf8),
	.w5(32'hbb672b30),
	.w6(32'h3a6058d4),
	.w7(32'h3aacbc1e),
	.w8(32'hbc07c76f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5badb),
	.w1(32'hbbb902f7),
	.w2(32'hba7315ea),
	.w3(32'h3b4097dc),
	.w4(32'h3b85bf19),
	.w5(32'h36fe57b8),
	.w6(32'h3b6aff5c),
	.w7(32'h3b906862),
	.w8(32'h3add15da),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11c73e),
	.w1(32'h3b5191e4),
	.w2(32'h3b2a11cd),
	.w3(32'hbad28530),
	.w4(32'h3b90a155),
	.w5(32'h3b5843f4),
	.w6(32'hbb06937c),
	.w7(32'h3a848b30),
	.w8(32'h3a17af05),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dcf87),
	.w1(32'hbc15ddbd),
	.w2(32'hbb1d1acf),
	.w3(32'hbb4e821f),
	.w4(32'h3be14432),
	.w5(32'h3a199789),
	.w6(32'hbb9f1c92),
	.w7(32'h3b40dcd9),
	.w8(32'hbbe2dd28),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92705ef),
	.w1(32'h39960edc),
	.w2(32'h3b968377),
	.w3(32'h3af1b1cb),
	.w4(32'h3ba2608a),
	.w5(32'hb990b5a1),
	.w6(32'h3b27366b),
	.w7(32'h3b9e9fd2),
	.w8(32'h3a326d51),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae5415),
	.w1(32'hb8ff76c7),
	.w2(32'hbbd072b4),
	.w3(32'hb902b6fd),
	.w4(32'hbb19da09),
	.w5(32'hbc234a88),
	.w6(32'hbba83cde),
	.w7(32'hbbec47fa),
	.w8(32'hbc00ed7f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fd2ea),
	.w1(32'h3a995990),
	.w2(32'hbb3af2d0),
	.w3(32'hba4cf6d9),
	.w4(32'hba1c5bc5),
	.w5(32'hbb2a588d),
	.w6(32'hbaccc5be),
	.w7(32'hba9310f9),
	.w8(32'hbb96096f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d8010),
	.w1(32'h3a126b72),
	.w2(32'hb9f72f9c),
	.w3(32'h3ac197e3),
	.w4(32'hb9c49a33),
	.w5(32'hb9880393),
	.w6(32'h3a04b671),
	.w7(32'hba2a6ab9),
	.w8(32'hba9597a3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913710b),
	.w1(32'hbc2024fc),
	.w2(32'hba81b68a),
	.w3(32'hbbbfaa77),
	.w4(32'h3ae3d77b),
	.w5(32'hbb76638f),
	.w6(32'hbbc42405),
	.w7(32'h3ad405a0),
	.w8(32'hbba8a027),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba85e61),
	.w1(32'hbab0ca13),
	.w2(32'hba236b77),
	.w3(32'hbb1bc0d6),
	.w4(32'h3a24d0f4),
	.w5(32'h3ab89bfa),
	.w6(32'hbb9621e4),
	.w7(32'hbb2a87bc),
	.w8(32'h3ab8de8a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ab24e),
	.w1(32'h3bd1a2dc),
	.w2(32'hbb1628d1),
	.w3(32'hbb8da6cc),
	.w4(32'h3b671994),
	.w5(32'hbc0a60a4),
	.w6(32'hbc5a8ca6),
	.w7(32'hbc116ffc),
	.w8(32'hbca5beec),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6776e),
	.w1(32'h3b6549e3),
	.w2(32'h39185d52),
	.w3(32'hbb1c99c1),
	.w4(32'h3c56f829),
	.w5(32'h3a8a4796),
	.w6(32'hbb503149),
	.w7(32'h3b91b42f),
	.w8(32'hbb866a9f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28012b),
	.w1(32'h3afb267c),
	.w2(32'h3b9f531d),
	.w3(32'hbc1c37e5),
	.w4(32'hbaa54df6),
	.w5(32'h3bedbe0c),
	.w6(32'hbc3ed778),
	.w7(32'hbafc4938),
	.w8(32'hb9524431),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7fa372),
	.w1(32'h382a6146),
	.w2(32'h3a9e30f0),
	.w3(32'hb9dacd13),
	.w4(32'h3aafa11b),
	.w5(32'hbad3b61d),
	.w6(32'hbb4ca31f),
	.w7(32'h36d71cc9),
	.w8(32'hbb178c23),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12706c),
	.w1(32'hbae6bd8c),
	.w2(32'hbaf10acd),
	.w3(32'hbb1701d2),
	.w4(32'hbad75471),
	.w5(32'hbacc7a1d),
	.w6(32'hbb0e30bd),
	.w7(32'hbadbe946),
	.w8(32'h38336cc1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27ccf9),
	.w1(32'hbab51e19),
	.w2(32'h3b939a9d),
	.w3(32'hbb81838f),
	.w4(32'h3b9ade78),
	.w5(32'hbb685f32),
	.w6(32'h39f2d2a0),
	.w7(32'h3bc10968),
	.w8(32'hbb50ce13),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b6487),
	.w1(32'hb7ee0da3),
	.w2(32'h3ba7eb2f),
	.w3(32'h3a88dc06),
	.w4(32'h3ba70add),
	.w5(32'h3aead75e),
	.w6(32'hb9f40c27),
	.w7(32'h3bbe9cf8),
	.w8(32'h395c1dfe),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93032d),
	.w1(32'h3be0b3b5),
	.w2(32'h3b9060a7),
	.w3(32'hb98c8a36),
	.w4(32'hbaf5161a),
	.w5(32'h3aecb094),
	.w6(32'h3a94ffa1),
	.w7(32'hbb8758ee),
	.w8(32'h39b15885),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0809ad),
	.w1(32'hbaaea227),
	.w2(32'hbbd8596f),
	.w3(32'h3a04671f),
	.w4(32'hba834704),
	.w5(32'h391f45ba),
	.w6(32'hbb4d1c27),
	.w7(32'hbba29397),
	.w8(32'h3a228a0e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb947638c),
	.w1(32'h3be48e74),
	.w2(32'h3b9370b9),
	.w3(32'hb7b4a369),
	.w4(32'hbb41250c),
	.w5(32'h3a38f0eb),
	.w6(32'h3ae0f25a),
	.w7(32'hba906401),
	.w8(32'h3b2966de),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cded35),
	.w1(32'h3b082ac9),
	.w2(32'hbace6671),
	.w3(32'h3b4016e8),
	.w4(32'h3b4018c0),
	.w5(32'h3a7043db),
	.w6(32'hb9907fdc),
	.w7(32'hba3e45cc),
	.w8(32'hba59aac9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4ca2c),
	.w1(32'h3abc1c8a),
	.w2(32'h3b8ef0d2),
	.w3(32'h3aa4b25d),
	.w4(32'h3ba735a4),
	.w5(32'hba5d7dc8),
	.w6(32'hba37397e),
	.w7(32'h3b49a6c4),
	.w8(32'hbaa7bd32),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381ce214),
	.w1(32'h3b0635a0),
	.w2(32'h3a458edb),
	.w3(32'h3b70133c),
	.w4(32'h3b147753),
	.w5(32'h3b58ea56),
	.w6(32'h3b853cee),
	.w7(32'h3b5a77ac),
	.w8(32'h3b87706f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16eefa),
	.w1(32'h3b464cca),
	.w2(32'h3b0ae376),
	.w3(32'h3b5f00fc),
	.w4(32'h3bdd1e20),
	.w5(32'h3b0acd2c),
	.w6(32'h3b2fb335),
	.w7(32'h3b7f6ed2),
	.w8(32'h3a7fa46b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a5ba6),
	.w1(32'h3bb41c82),
	.w2(32'hbc32cfc4),
	.w3(32'hbba5dedc),
	.w4(32'h3c38137f),
	.w5(32'hbbb1853b),
	.w6(32'hbc96027b),
	.w7(32'h3a67f344),
	.w8(32'hbc308d0d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ccfd8),
	.w1(32'h3b66f7a4),
	.w2(32'h3c2b5043),
	.w3(32'hbc320b2f),
	.w4(32'hbae4c9e9),
	.w5(32'h3c356e94),
	.w6(32'hbc583127),
	.w7(32'hbbc5fce3),
	.w8(32'h3c09a32d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7acd0),
	.w1(32'h3b197d89),
	.w2(32'h3c5bda0d),
	.w3(32'hbc05f762),
	.w4(32'h3abd0392),
	.w5(32'h3b67991b),
	.w6(32'hbc041aee),
	.w7(32'hba1b4f9a),
	.w8(32'hbb27780e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb970185),
	.w1(32'hba9437d4),
	.w2(32'h3ac34dd3),
	.w3(32'hbb90c4e1),
	.w4(32'h3ac5fe62),
	.w5(32'h3a28c30d),
	.w6(32'hbbc50161),
	.w7(32'h3a331c8f),
	.w8(32'hba6f3c32),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba931c55),
	.w1(32'hbaa2bfcf),
	.w2(32'h3a6affe0),
	.w3(32'hbba660d1),
	.w4(32'hba156e0b),
	.w5(32'h3a1569ee),
	.w6(32'hbb144db5),
	.w7(32'h3b08ee6f),
	.w8(32'hbb063a10),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d16096),
	.w1(32'hb708b06a),
	.w2(32'h3af45605),
	.w3(32'hb9ab676d),
	.w4(32'h3a8a1af9),
	.w5(32'hbb9281a3),
	.w6(32'hbb328c39),
	.w7(32'hb9d90826),
	.w8(32'hbb5cfdc7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88de2f),
	.w1(32'hbb454de4),
	.w2(32'hbb11c8cc),
	.w3(32'hbbde5cd8),
	.w4(32'hbb900cd9),
	.w5(32'hbb2a0870),
	.w6(32'hbbc7250f),
	.w7(32'hbb55d766),
	.w8(32'hbb945d73),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc70e5),
	.w1(32'hb9845371),
	.w2(32'hbb509936),
	.w3(32'hbb72d8be),
	.w4(32'h3babc39a),
	.w5(32'hbba2e0f0),
	.w6(32'hbbc9c343),
	.w7(32'hbbcc977f),
	.w8(32'hbc2b6761),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba82cd),
	.w1(32'h3a672528),
	.w2(32'hb9f52013),
	.w3(32'hbbb99743),
	.w4(32'h3a55ddd9),
	.w5(32'h3ba45346),
	.w6(32'hbc23a97e),
	.w7(32'hbb736483),
	.w8(32'hbb8a34e9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b594a),
	.w1(32'h3bb1e420),
	.w2(32'h3a852723),
	.w3(32'hb9d63fa2),
	.w4(32'h3badf1ff),
	.w5(32'h3b051a28),
	.w6(32'hbc600d61),
	.w7(32'hbb1f80c5),
	.w8(32'hbbc00f48),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82ed43),
	.w1(32'h3b0faab6),
	.w2(32'hba78aa40),
	.w3(32'hbaf89377),
	.w4(32'hba5fbe43),
	.w5(32'h3a0aa280),
	.w6(32'hbbd5eb21),
	.w7(32'hbb8e1547),
	.w8(32'hbb128e52),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7aaf3),
	.w1(32'h3b906f9f),
	.w2(32'hbbd4b8c2),
	.w3(32'h3bd17ed2),
	.w4(32'h3b736af8),
	.w5(32'hbb99e7b3),
	.w6(32'hbb2fc410),
	.w7(32'hbb91a3fc),
	.w8(32'hbb90a22e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7b813),
	.w1(32'h3bb960b4),
	.w2(32'h3b78e993),
	.w3(32'h3b2de01f),
	.w4(32'h3b434217),
	.w5(32'hbb2a0dbc),
	.w6(32'h3c054cb1),
	.w7(32'h3b9c7d8f),
	.w8(32'hbb8bcbdd),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7543c5),
	.w1(32'hbb0db102),
	.w2(32'hbaabcf15),
	.w3(32'hbb20c11c),
	.w4(32'hbaffe6a6),
	.w5(32'hba1a232f),
	.w6(32'hbbadfde6),
	.w7(32'hbbad7211),
	.w8(32'hbb18649c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d567f),
	.w1(32'h3942348a),
	.w2(32'hb8ca4d59),
	.w3(32'hbb2d02b1),
	.w4(32'hba9988d8),
	.w5(32'hba0c7d7c),
	.w6(32'hba0e174e),
	.w7(32'hbaedb054),
	.w8(32'hb9a1eb89),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83b6a9),
	.w1(32'hbb07fa53),
	.w2(32'hbb040f20),
	.w3(32'hbb88b419),
	.w4(32'hbb09165f),
	.w5(32'h3ad2327d),
	.w6(32'hbbb03c2f),
	.w7(32'hbb8c2e0f),
	.w8(32'hbb630f6b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fb332c),
	.w1(32'h3aa2d708),
	.w2(32'h3b709255),
	.w3(32'hbb41972f),
	.w4(32'h3b6795a8),
	.w5(32'h37c23de2),
	.w6(32'hba7008d5),
	.w7(32'h3b8e20d0),
	.w8(32'hbaf770d4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a8c65),
	.w1(32'h3b55db79),
	.w2(32'hbc1ba71c),
	.w3(32'h3b8d4b4e),
	.w4(32'h3a2458f0),
	.w5(32'hbc01afdd),
	.w6(32'hbbcb3e20),
	.w7(32'hbbb24ebd),
	.w8(32'hbc101cbb),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe1d17),
	.w1(32'hba9601db),
	.w2(32'hbad08e50),
	.w3(32'hbb17dce2),
	.w4(32'hbb40925a),
	.w5(32'hbb3803b7),
	.w6(32'hbb62df11),
	.w7(32'hbb67984e),
	.w8(32'hbb5de7e4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90b9ee),
	.w1(32'h3a1222ad),
	.w2(32'h3b40c7d8),
	.w3(32'h3b8a5b7d),
	.w4(32'h3b42e8d1),
	.w5(32'hbad947ab),
	.w6(32'h3b3ba84f),
	.w7(32'h3a574e1f),
	.w8(32'hbb369689),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf18f7),
	.w1(32'hb98fe98c),
	.w2(32'h3a6bd84d),
	.w3(32'h38b3bc6f),
	.w4(32'h3b28ec9a),
	.w5(32'h3afcc589),
	.w6(32'hbaa89bda),
	.w7(32'h3b051eba),
	.w8(32'h3ab5d216),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe129c),
	.w1(32'hb9b8f709),
	.w2(32'h3af117f4),
	.w3(32'hbadd144a),
	.w4(32'h3b2f333b),
	.w5(32'hbb002bf8),
	.w6(32'hba87c79f),
	.w7(32'h3b50a8a7),
	.w8(32'hbb2e6be3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2aae1a),
	.w1(32'hb91bff11),
	.w2(32'hb9018ae0),
	.w3(32'hbad7d675),
	.w4(32'hbae5b004),
	.w5(32'hba947ace),
	.w6(32'hbb8bf0cf),
	.w7(32'hbba16817),
	.w8(32'hbb31c184),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18c8eb),
	.w1(32'hb94d90ae),
	.w2(32'hbb035350),
	.w3(32'h3ab426e9),
	.w4(32'hbba8edee),
	.w5(32'hbaf16dc4),
	.w6(32'hba188a91),
	.w7(32'hbb662a7d),
	.w8(32'h3b07991d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad959fa),
	.w1(32'h3b2a10d9),
	.w2(32'h3a075daf),
	.w3(32'hb982805f),
	.w4(32'h3a8afb30),
	.w5(32'hbb65f0bc),
	.w6(32'h3a9487f4),
	.w7(32'hba8a7718),
	.w8(32'hbbd84d72),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd047e),
	.w1(32'hbb2b4d5d),
	.w2(32'h3ad4938c),
	.w3(32'hba757087),
	.w4(32'h3a852790),
	.w5(32'hbb3d4574),
	.w6(32'hbb2c0cd4),
	.w7(32'hbb5ea3bc),
	.w8(32'hbba23a63),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a048912),
	.w1(32'hbabcb2ac),
	.w2(32'hbada297b),
	.w3(32'h38b6e5a9),
	.w4(32'hb9ca73a8),
	.w5(32'hbad5f1ce),
	.w6(32'hba432548),
	.w7(32'hbb0efbfd),
	.w8(32'hbb012eaf),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94f930),
	.w1(32'h3aef755c),
	.w2(32'h3b2bf77b),
	.w3(32'h3b462b38),
	.w4(32'h3b81f2a0),
	.w5(32'hbb7fa6a1),
	.w6(32'h3b343afc),
	.w7(32'h3b614891),
	.w8(32'hbb045c3d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab52906),
	.w1(32'hba9d3b63),
	.w2(32'h3927b199),
	.w3(32'h3ad35434),
	.w4(32'h3ae60779),
	.w5(32'hb907e45b),
	.w6(32'h3a222d4c),
	.w7(32'hb8fd1a78),
	.w8(32'h387729d0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86b281),
	.w1(32'h3b2961c2),
	.w2(32'h3aecb620),
	.w3(32'hb75a9999),
	.w4(32'hb9fb2f5a),
	.w5(32'h3ba91a93),
	.w6(32'hb90818c3),
	.w7(32'h3adb956c),
	.w8(32'h3b89c35f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e636d),
	.w1(32'hbbadf044),
	.w2(32'hbc1f374c),
	.w3(32'h3b855de0),
	.w4(32'h3a8dfb86),
	.w5(32'hbbf87f69),
	.w6(32'h3b3b6bec),
	.w7(32'hb95f069f),
	.w8(32'hbc1becc5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1fd72),
	.w1(32'hbb410309),
	.w2(32'hbc11871e),
	.w3(32'hbc2f7e41),
	.w4(32'hbb8e26ab),
	.w5(32'hbbd71dd7),
	.w6(32'hbc9dfd1e),
	.w7(32'hbc83c2b5),
	.w8(32'hbc5dd3f2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41d8a2),
	.w1(32'hbb334075),
	.w2(32'hbbbf9c17),
	.w3(32'hbb0d475e),
	.w4(32'hbb17bccf),
	.w5(32'hbb9a9987),
	.w6(32'hbc2ec960),
	.w7(32'hbc3d6c37),
	.w8(32'hbc2d57ec),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b437c),
	.w1(32'h3bb27548),
	.w2(32'h3c26782e),
	.w3(32'hbc54f4aa),
	.w4(32'h3b530aaa),
	.w5(32'h3c2a85c3),
	.w6(32'hbc81136a),
	.w7(32'hbb48abd4),
	.w8(32'h3a3c3004),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5321c),
	.w1(32'hba0ab497),
	.w2(32'hb8c1c9a5),
	.w3(32'hbac4117c),
	.w4(32'hbabbd320),
	.w5(32'h3b9b7b1e),
	.w6(32'hba46701a),
	.w7(32'hb9a3eef6),
	.w8(32'h3b50e766),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b902dbf),
	.w1(32'hbbae347d),
	.w2(32'h3b90ca45),
	.w3(32'hbb193184),
	.w4(32'h3aed24ce),
	.w5(32'hb9d1ba33),
	.w6(32'hbb0342e1),
	.w7(32'h3bb84b7a),
	.w8(32'h3a72cca8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0a08a),
	.w1(32'h38f9249d),
	.w2(32'hb9ee8a24),
	.w3(32'hba253a53),
	.w4(32'h3afe507f),
	.w5(32'h3b23fa99),
	.w6(32'hb9adf724),
	.w7(32'h3b67989d),
	.w8(32'h3ade45fa),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d6dc7),
	.w1(32'hba373168),
	.w2(32'hbb34c001),
	.w3(32'h3b1dd024),
	.w4(32'h3a86e694),
	.w5(32'hba844a25),
	.w6(32'hbb1c58fe),
	.w7(32'hba901cd1),
	.w8(32'hb9e770b3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fc781),
	.w1(32'hba60c4b9),
	.w2(32'h3bc2800c),
	.w3(32'hbb6de416),
	.w4(32'h3aab9208),
	.w5(32'h3b3b2107),
	.w6(32'hba056dc4),
	.w7(32'h3bd9aee8),
	.w8(32'h3b396779),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad8bf1),
	.w1(32'h3aa13757),
	.w2(32'hbb9b59aa),
	.w3(32'h3a2ab6d7),
	.w4(32'hba43e9bd),
	.w5(32'hbb9b7240),
	.w6(32'hba899c8b),
	.w7(32'hbb2aff72),
	.w8(32'hbbd5feb6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8c5d5),
	.w1(32'h3b96d332),
	.w2(32'hbb0c39e2),
	.w3(32'hbaf48cd4),
	.w4(32'h3b2b486a),
	.w5(32'hbb4c863c),
	.w6(32'hbb457ee6),
	.w7(32'hbb085ccb),
	.w8(32'hbc0dabe9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6f66f),
	.w1(32'h39bb7148),
	.w2(32'h3a172c8a),
	.w3(32'hbb9b23ae),
	.w4(32'h3b08ab32),
	.w5(32'h3b84e5ea),
	.w6(32'hbbb6e901),
	.w7(32'hba52f6c7),
	.w8(32'h3b387d3f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3896a09b),
	.w1(32'h3a83889c),
	.w2(32'hbb3f898e),
	.w3(32'hba8ca0bd),
	.w4(32'hbb6711c5),
	.w5(32'h384160d5),
	.w6(32'hb9e036a5),
	.w7(32'hbb19597a),
	.w8(32'hbb028dfe),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c6c8e),
	.w1(32'h39898ad2),
	.w2(32'h3898988e),
	.w3(32'h3b0abf6b),
	.w4(32'h3bf08419),
	.w5(32'hbbb758e7),
	.w6(32'h3b62735e),
	.w7(32'h3bcfb609),
	.w8(32'hbbf4c995),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8a5b),
	.w1(32'h39ffdda7),
	.w2(32'hbab73fc1),
	.w3(32'hbb7de2d2),
	.w4(32'hbb0ea0e0),
	.w5(32'h3a267ed1),
	.w6(32'hbb3b0662),
	.w7(32'hbb550beb),
	.w8(32'h3a5b8765),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8845f1),
	.w1(32'h3a1e56bc),
	.w2(32'hbb91358a),
	.w3(32'hba95de83),
	.w4(32'hbaf4f05e),
	.w5(32'hbbfcd1c2),
	.w6(32'hbb4d6ee0),
	.w7(32'hbb59435d),
	.w8(32'hbc0a7e73),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51d80f),
	.w1(32'hb92b96a7),
	.w2(32'hb93ccdb2),
	.w3(32'hbb793a4b),
	.w4(32'hbb0ac5f4),
	.w5(32'hbbc4874c),
	.w6(32'h3a53012c),
	.w7(32'hbac2ca64),
	.w8(32'hbbbc397f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd537f2),
	.w1(32'hbbcdc314),
	.w2(32'hbb98a69a),
	.w3(32'hbbb7dcc7),
	.w4(32'hbb5cd396),
	.w5(32'hba94cbef),
	.w6(32'hbbaa3876),
	.w7(32'hbb55cdf9),
	.w8(32'hbaf31af7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb548615),
	.w1(32'hbaacdf08),
	.w2(32'h3a276195),
	.w3(32'hbaff8540),
	.w4(32'hbb22566b),
	.w5(32'hba16b360),
	.w6(32'hbadf64fb),
	.w7(32'hbae8bb3c),
	.w8(32'h39a57c59),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac94d8a),
	.w1(32'h3a922767),
	.w2(32'h3bcf87ef),
	.w3(32'hbb00f03c),
	.w4(32'h3a8047bb),
	.w5(32'h3a2e2d71),
	.w6(32'hba561b26),
	.w7(32'h3ad39332),
	.w8(32'h39eff530),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc348b),
	.w1(32'h3b154575),
	.w2(32'h3bb10382),
	.w3(32'hbc041640),
	.w4(32'h3b428752),
	.w5(32'h3aeba015),
	.w6(32'hbc23b3a5),
	.w7(32'hba5fa138),
	.w8(32'hba79e30b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0385f9),
	.w1(32'h3a05bc13),
	.w2(32'hba915e52),
	.w3(32'hba5178e3),
	.w4(32'hba9c6547),
	.w5(32'hb94dcfc3),
	.w6(32'h3a0434a2),
	.w7(32'hb989e8d0),
	.w8(32'hbab30e92),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9db4b2),
	.w1(32'hbaeac3a8),
	.w2(32'hbacfc855),
	.w3(32'hbb89c39e),
	.w4(32'h3a3e116f),
	.w5(32'hba9350d3),
	.w6(32'hbbb78428),
	.w7(32'hbb4e28bc),
	.w8(32'hbb1b1b5f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61fa60),
	.w1(32'h3c0d542b),
	.w2(32'hbb0c99bd),
	.w3(32'h3b5a4040),
	.w4(32'hbabfd394),
	.w5(32'hbc2db482),
	.w6(32'hbac3f713),
	.w7(32'hbc1bbbf8),
	.w8(32'hbc87317a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfae261),
	.w1(32'h3b7298d7),
	.w2(32'h3c0f66eb),
	.w3(32'h3b1bfee6),
	.w4(32'h3bcc7001),
	.w5(32'h3aec6e4c),
	.w6(32'h3b11ab44),
	.w7(32'h3b6b2a6b),
	.w8(32'hba1aaa40),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98df86),
	.w1(32'h3badf1f9),
	.w2(32'hbc112c6e),
	.w3(32'h3c046af5),
	.w4(32'h3afcd6f7),
	.w5(32'hbbb72be1),
	.w6(32'h3ae4491e),
	.w7(32'hbb97b0f1),
	.w8(32'hbc3e6e48),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc048852),
	.w1(32'h3b8b24a2),
	.w2(32'h3ba89deb),
	.w3(32'hbae88a63),
	.w4(32'h3b04ef9f),
	.w5(32'h3b82cf17),
	.w6(32'hbb66c3ac),
	.w7(32'hbb365e30),
	.w8(32'h39da6537),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d02a2),
	.w1(32'hbc06aa50),
	.w2(32'hbc4d7a03),
	.w3(32'hbb5633cd),
	.w4(32'hbbb6238f),
	.w5(32'hbbe7a786),
	.w6(32'hbc133e32),
	.w7(32'hbc2c56c9),
	.w8(32'hbc275af2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacecf4),
	.w1(32'hbbb13444),
	.w2(32'hbbd8c721),
	.w3(32'hbbabf3f0),
	.w4(32'hbb9ffc16),
	.w5(32'hbafab738),
	.w6(32'hbb99a4f5),
	.w7(32'hbb8632c7),
	.w8(32'hb92fa525),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c1ee5),
	.w1(32'h3b574f3f),
	.w2(32'h3c16a279),
	.w3(32'hbbf516b8),
	.w4(32'hbb3605a8),
	.w5(32'h3b47fe01),
	.w6(32'hbb09aa24),
	.w7(32'h3b1aec5b),
	.w8(32'h3b41c9ea),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09c401),
	.w1(32'hbad9a053),
	.w2(32'hbb35edeb),
	.w3(32'hba72ef34),
	.w4(32'hbb5a9abf),
	.w5(32'hbb1627d2),
	.w6(32'hba9d3d06),
	.w7(32'hbb407282),
	.w8(32'hbb9b18ad),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ededc),
	.w1(32'h3bad8a23),
	.w2(32'hbba15fc7),
	.w3(32'h3b92b57e),
	.w4(32'h3b977c04),
	.w5(32'hbb0f3b8e),
	.w6(32'h3a9aec09),
	.w7(32'hbb2d4f3c),
	.w8(32'hbbd1302d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998008e),
	.w1(32'h3840f9b3),
	.w2(32'hbbc0431f),
	.w3(32'hbb0fafe7),
	.w4(32'h39151a49),
	.w5(32'hbbb4d343),
	.w6(32'hbc05afe3),
	.w7(32'hbb88143f),
	.w8(32'hbc3bc150),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1ed1b),
	.w1(32'h3b7abb65),
	.w2(32'hbc1a3dea),
	.w3(32'hbbcfed77),
	.w4(32'h3c0af65a),
	.w5(32'hbb3110c3),
	.w6(32'hbc9bde23),
	.w7(32'hbaa61c02),
	.w8(32'hbc7be68d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37d47d),
	.w1(32'h3b307d7d),
	.w2(32'h3c37c614),
	.w3(32'hbc01c77b),
	.w4(32'h3bbea73e),
	.w5(32'h3c5612b2),
	.w6(32'hbc21791b),
	.w7(32'h3ab2e2e0),
	.w8(32'h3c19211d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ca636),
	.w1(32'h3be3ea97),
	.w2(32'h3b9857aa),
	.w3(32'hbb5a1609),
	.w4(32'h3b6dbb8e),
	.w5(32'h3b72e558),
	.w6(32'hbb35a456),
	.w7(32'h3adcc8ee),
	.w8(32'h38f8572a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8c4ae),
	.w1(32'hb7def9e4),
	.w2(32'hbc061eed),
	.w3(32'h38e15ec8),
	.w4(32'h3b65205a),
	.w5(32'hbaa7ba3c),
	.w6(32'hbbe91172),
	.w7(32'hbac33cfc),
	.w8(32'hbc13c5de),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f7108),
	.w1(32'hba1c4eb2),
	.w2(32'hbaa1c999),
	.w3(32'hba6405ef),
	.w4(32'h3ab68cab),
	.w5(32'h396adc00),
	.w6(32'hba3627c0),
	.w7(32'hb9bd5e9e),
	.w8(32'h3abb9484),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc445985),
	.w1(32'hbb8fde21),
	.w2(32'hbc7a58a6),
	.w3(32'hbc431f57),
	.w4(32'hbb00bd8c),
	.w5(32'hbabd5140),
	.w6(32'hbc1a1c66),
	.w7(32'h3a012c62),
	.w8(32'hbc17734f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850d4e),
	.w1(32'hbb1d1be5),
	.w2(32'hbb2a3213),
	.w3(32'h3ac8a741),
	.w4(32'h3a5045ea),
	.w5(32'hbb6da0d3),
	.w6(32'hbba64ad2),
	.w7(32'h3a52755f),
	.w8(32'hbb28b122),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd67ae),
	.w1(32'hb8c20663),
	.w2(32'hba85dfce),
	.w3(32'hbae046b3),
	.w4(32'h39b7dff8),
	.w5(32'hb99bb095),
	.w6(32'hbac1e96a),
	.w7(32'h37cc64a3),
	.w8(32'h39e66abc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa0e21),
	.w1(32'hba70c55d),
	.w2(32'hbb097a32),
	.w3(32'hb9d2a73c),
	.w4(32'h393dcda8),
	.w5(32'h3a8fde94),
	.w6(32'hbaa84178),
	.w7(32'hbab1954e),
	.w8(32'hbb6e11c9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2dcc6),
	.w1(32'h3b1840a9),
	.w2(32'h39c99382),
	.w3(32'h3aecb051),
	.w4(32'h3ba05b39),
	.w5(32'h3b101215),
	.w6(32'hbbb9626c),
	.w7(32'hbab6ef4a),
	.w8(32'hbba08a54),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fa910),
	.w1(32'hba4300ab),
	.w2(32'h3a314cd2),
	.w3(32'hbabdeebe),
	.w4(32'h3b3f3a95),
	.w5(32'h3a851258),
	.w6(32'hbbb14635),
	.w7(32'h39a1e6bd),
	.w8(32'hba6fd972),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ab75),
	.w1(32'hbaab011d),
	.w2(32'h3b6476d4),
	.w3(32'hbb053399),
	.w4(32'hba3ec782),
	.w5(32'h3acd9a4c),
	.w6(32'hbba0cb2d),
	.w7(32'hbad10787),
	.w8(32'hbae23761),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9355bb),
	.w1(32'hb92e0c90),
	.w2(32'h397638cb),
	.w3(32'hba577889),
	.w4(32'h39f71525),
	.w5(32'h3ac3f7c9),
	.w6(32'hbaf3ac01),
	.w7(32'hbab12222),
	.w8(32'hbad8849e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6833f8),
	.w1(32'h3b99a62a),
	.w2(32'h3b3b4ed8),
	.w3(32'hbb94cd94),
	.w4(32'h3b060380),
	.w5(32'h3a24a79e),
	.w6(32'hbc198a2e),
	.w7(32'hbba1ebcd),
	.w8(32'hbbbb0608),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8febe),
	.w1(32'hbbf88b3a),
	.w2(32'hbc409a6b),
	.w3(32'h3ae87d77),
	.w4(32'h39acb13e),
	.w5(32'hbbd1f8cf),
	.w6(32'hba202892),
	.w7(32'hbb407cdd),
	.w8(32'hbbc8a4ed),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07fc9a),
	.w1(32'h3ac343fd),
	.w2(32'hbaed53ca),
	.w3(32'hba8773fd),
	.w4(32'hba58a5e3),
	.w5(32'h39983e9e),
	.w6(32'hbb5e5314),
	.w7(32'hbb2aad24),
	.w8(32'hbb5f4e9f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04ef6e),
	.w1(32'hbb2a6a6c),
	.w2(32'hb9a86c60),
	.w3(32'h3aa02f26),
	.w4(32'h38a3c50d),
	.w5(32'h3adf9cdf),
	.w6(32'hb8b74a2d),
	.w7(32'hb9ed154f),
	.w8(32'h3b1916b7),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ee652),
	.w1(32'h3aa755a4),
	.w2(32'hb833bb5c),
	.w3(32'h3b02dc84),
	.w4(32'h3a8cd576),
	.w5(32'h386ab343),
	.w6(32'h3b043f28),
	.w7(32'h3aa58c1b),
	.w8(32'h3a73d373),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3856f),
	.w1(32'h390ef2c7),
	.w2(32'h3ad68805),
	.w3(32'hbac709a5),
	.w4(32'h3924de62),
	.w5(32'h3aef7c3f),
	.w6(32'h3a3167dc),
	.w7(32'h398f5660),
	.w8(32'hba9c930f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bace8),
	.w1(32'hba80e054),
	.w2(32'hbaa27bf7),
	.w3(32'h3b46f499),
	.w4(32'h3b298eb9),
	.w5(32'h3ae33481),
	.w6(32'hbaab262e),
	.w7(32'hba2d56fa),
	.w8(32'h3a2a1b89),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae43c45),
	.w1(32'h3b887b16),
	.w2(32'h3b47893d),
	.w3(32'hbadf98ea),
	.w4(32'h3b828cea),
	.w5(32'h3ad3eeef),
	.w6(32'hbb1cb799),
	.w7(32'h396d599f),
	.w8(32'hbb2e47e6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68f96c),
	.w1(32'hba0dacf7),
	.w2(32'hb8b909af),
	.w3(32'hba5a6426),
	.w4(32'hb900fa88),
	.w5(32'hb8ba9704),
	.w6(32'hba7a7d3e),
	.w7(32'h38466621),
	.w8(32'hba89bdae),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81dbde0),
	.w1(32'h3a322371),
	.w2(32'hbb021e08),
	.w3(32'h3b12b2c2),
	.w4(32'h3a9457bb),
	.w5(32'hba434292),
	.w6(32'hbad7bd30),
	.w7(32'h39c992e7),
	.w8(32'hbbdbbb09),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb950e45),
	.w1(32'h3bb64fcd),
	.w2(32'h3c055623),
	.w3(32'h39c09f55),
	.w4(32'h3b301bbb),
	.w5(32'h3b92ec54),
	.w6(32'hbbe0f121),
	.w7(32'hbc038854),
	.w8(32'h3a1ad43f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b828c),
	.w1(32'hbb778019),
	.w2(32'hba9eaea2),
	.w3(32'hba604520),
	.w4(32'hbb7ac81a),
	.w5(32'h3b853c47),
	.w6(32'h3b8eeccc),
	.w7(32'h3a6d57d6),
	.w8(32'hbb92b44d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926c9ae),
	.w1(32'h3a033c59),
	.w2(32'hb835b34e),
	.w3(32'h3c1533be),
	.w4(32'h3be7107c),
	.w5(32'hb9949687),
	.w6(32'hbb50d755),
	.w7(32'hbb17f782),
	.w8(32'hb9e9c050),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa706dd),
	.w1(32'h3a5857e0),
	.w2(32'hba02a590),
	.w3(32'h3a688817),
	.w4(32'h3a9527ef),
	.w5(32'hb9588caf),
	.w6(32'h3aab5576),
	.w7(32'hba86aaff),
	.w8(32'hba86ee58),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba798ea1),
	.w1(32'hbb013ab0),
	.w2(32'hba0d2bdd),
	.w3(32'h39cba821),
	.w4(32'h3a9aad95),
	.w5(32'h3a8d4991),
	.w6(32'hba5fe418),
	.w7(32'h3a4573e3),
	.w8(32'hba9dc18c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21748f),
	.w1(32'h3b975faa),
	.w2(32'hbbc27a62),
	.w3(32'h3b38e16d),
	.w4(32'h3ab9417d),
	.w5(32'hbb2bea58),
	.w6(32'hbbc5f963),
	.w7(32'hbbfe0f96),
	.w8(32'hbc10287c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cca680),
	.w1(32'hbb82b23c),
	.w2(32'hbbf0281f),
	.w3(32'h3b9de2fe),
	.w4(32'h3b2e62a0),
	.w5(32'hbbc50848),
	.w6(32'hbb83f109),
	.w7(32'hbb71a7b4),
	.w8(32'hbb8e5c30),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad52f59),
	.w1(32'hb9e01886),
	.w2(32'hba46b6a9),
	.w3(32'h3a1d3a40),
	.w4(32'hb958d08b),
	.w5(32'hba822579),
	.w6(32'h3997f997),
	.w7(32'h3a210fc1),
	.w8(32'hbb61e5b5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d7f15),
	.w1(32'hba03f346),
	.w2(32'hbaf2e046),
	.w3(32'hba735856),
	.w4(32'hb9c5dcff),
	.w5(32'hb953e28a),
	.w6(32'hbb3ea5a6),
	.w7(32'hbb7d0cb8),
	.w8(32'hbad2c234),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2484b1),
	.w1(32'hb8c328c4),
	.w2(32'h3a13d185),
	.w3(32'hba7ffcbc),
	.w4(32'h3a6fb258),
	.w5(32'hbafc93de),
	.w6(32'hba84d8dc),
	.w7(32'h3aa28e7a),
	.w8(32'hbb977d9f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc70385),
	.w1(32'hbbcb75d4),
	.w2(32'hbb76f90e),
	.w3(32'hbae879f7),
	.w4(32'hba72cd37),
	.w5(32'h3a618bce),
	.w6(32'hbb97244f),
	.w7(32'hbb689c3a),
	.w8(32'hbb64e037),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbf47f),
	.w1(32'hbb9435ac),
	.w2(32'hbb5abf00),
	.w3(32'h3b122aeb),
	.w4(32'h3b48e1dc),
	.w5(32'h3a86cfc3),
	.w6(32'hbab7ac0a),
	.w7(32'hba7a8cbe),
	.w8(32'hba8a5d5b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f99b1),
	.w1(32'hb9f04dd2),
	.w2(32'hbbdd613c),
	.w3(32'h3bb3b559),
	.w4(32'h3b6ea116),
	.w5(32'hbb4a6efb),
	.w6(32'hbb378b24),
	.w7(32'hbb81e322),
	.w8(32'hbb8f7ca5),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb816e3c),
	.w1(32'h3ad6cae7),
	.w2(32'h3b6db393),
	.w3(32'hba5f60e7),
	.w4(32'h3a8a81c0),
	.w5(32'h3ba44c91),
	.w6(32'hbadd64fb),
	.w7(32'h3a02943c),
	.w8(32'h3acf8d5a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1bd78),
	.w1(32'hbae0acb1),
	.w2(32'hbb62ed0e),
	.w3(32'h3a8346cd),
	.w4(32'h3b01eacb),
	.w5(32'hb953d24c),
	.w6(32'hbb657459),
	.w7(32'hbb3f0251),
	.w8(32'hbbd42114),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16a149),
	.w1(32'hbac677da),
	.w2(32'hbbd56f2e),
	.w3(32'h3b2ab4a6),
	.w4(32'h3b556047),
	.w5(32'hbb37bd46),
	.w6(32'hbb876649),
	.w7(32'hbaddd84d),
	.w8(32'hbbfc8dee),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13c936),
	.w1(32'h3aaf4be5),
	.w2(32'h3a5a9aea),
	.w3(32'h3a0af381),
	.w4(32'h3b31fac6),
	.w5(32'h39ef2408),
	.w6(32'hbbdec45b),
	.w7(32'hbb08a3e3),
	.w8(32'hbb7694dc),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a858d4b),
	.w1(32'hbaa9c899),
	.w2(32'hbb67917e),
	.w3(32'h3ab4b25c),
	.w4(32'h3ac8e037),
	.w5(32'hbb74f015),
	.w6(32'hbb4c3bf6),
	.w7(32'hbb4a02d8),
	.w8(32'hbbc3a351),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05cbe2),
	.w1(32'hbad3feee),
	.w2(32'hbb1bc092),
	.w3(32'hbb02e69f),
	.w4(32'hbaa8ec65),
	.w5(32'hba8b399e),
	.w6(32'hbb675fe1),
	.w7(32'hbb575ca9),
	.w8(32'hba093327),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d7b8f),
	.w1(32'h3b0b4397),
	.w2(32'h3c1d5679),
	.w3(32'hbbe59f49),
	.w4(32'h3a22ac49),
	.w5(32'h3be65109),
	.w6(32'hba4b05d0),
	.w7(32'h3b2f4ad5),
	.w8(32'h3b38696b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fdc8d),
	.w1(32'hbb234f77),
	.w2(32'hb982cf61),
	.w3(32'hbada3d7f),
	.w4(32'hbaeda462),
	.w5(32'hbb5c514d),
	.w6(32'hbba0a963),
	.w7(32'hbb496584),
	.w8(32'hbb25b851),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f3f57),
	.w1(32'hbb41cb51),
	.w2(32'hbb4b007c),
	.w3(32'hbb154916),
	.w4(32'h3ac63bac),
	.w5(32'hb9054f6b),
	.w6(32'hbb4f89b7),
	.w7(32'hba99d112),
	.w8(32'hbabb0b65),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d992f0),
	.w1(32'hbaef3994),
	.w2(32'hb9db4fed),
	.w3(32'h398f303b),
	.w4(32'hb839b394),
	.w5(32'hba09d5b5),
	.w6(32'hba57c401),
	.w7(32'h3a11bad1),
	.w8(32'hba8bd1e6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba133d3e),
	.w1(32'hba2a51c5),
	.w2(32'hba903719),
	.w3(32'h3a691ca7),
	.w4(32'h3b05d5bb),
	.w5(32'h3adf9f2a),
	.w6(32'hbb586972),
	.w7(32'hb9af8e83),
	.w8(32'hba3b0380),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb745028),
	.w1(32'h3aa5ab86),
	.w2(32'h3b4023bc),
	.w3(32'hbb3e3ad3),
	.w4(32'h3af7a21a),
	.w5(32'h3b6c4df1),
	.w6(32'hbc096a5a),
	.w7(32'hbac05246),
	.w8(32'hb9feebb7),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2de680),
	.w1(32'hb890a531),
	.w2(32'hbb967eee),
	.w3(32'h3ac5fc75),
	.w4(32'h3b228a34),
	.w5(32'hbb014e3a),
	.w6(32'hbb768b83),
	.w7(32'hba152a54),
	.w8(32'hbb2ae3dd),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3daf6),
	.w1(32'hbb5d11ab),
	.w2(32'hbad647b1),
	.w3(32'hbb6a3e18),
	.w4(32'hba6001b0),
	.w5(32'h3b195b7d),
	.w6(32'hbb34f650),
	.w7(32'hba4f8cf5),
	.w8(32'h3b1afbe1),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f1be5),
	.w1(32'h3b50fb8c),
	.w2(32'hbab728c7),
	.w3(32'h3b487e2d),
	.w4(32'h3b57f926),
	.w5(32'h39e9e213),
	.w6(32'hba74b2e7),
	.w7(32'h3a0a255b),
	.w8(32'hbb6444a9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64629a),
	.w1(32'h3b1c337f),
	.w2(32'h3a4d80c1),
	.w3(32'h3a4468ef),
	.w4(32'h3af51fed),
	.w5(32'hbb5f435e),
	.w6(32'hba89e9ac),
	.w7(32'h3a319421),
	.w8(32'hbae4e933),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ad179),
	.w1(32'hbb23436d),
	.w2(32'hbc1c04a9),
	.w3(32'h3a65dfad),
	.w4(32'h3a8544ce),
	.w5(32'hba0f3eae),
	.w6(32'hbb886d1f),
	.w7(32'hbb5d9f35),
	.w8(32'hbbb997cb),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29a282),
	.w1(32'h3a1335f8),
	.w2(32'h3b18b1fd),
	.w3(32'h3b8acfb3),
	.w4(32'h3bc565f7),
	.w5(32'h3ac29270),
	.w6(32'hbb5f63a2),
	.w7(32'hbb0150a7),
	.w8(32'hbb8afc6e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c1b99),
	.w1(32'hbb5b7508),
	.w2(32'hbb27e97e),
	.w3(32'hbb58a56e),
	.w4(32'hbb4d208c),
	.w5(32'h39326ac5),
	.w6(32'hbb13a05f),
	.w7(32'hbb02ccea),
	.w8(32'hb9e82c86),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93a353),
	.w1(32'h3a9c2d29),
	.w2(32'h3a620392),
	.w3(32'hbaa829e5),
	.w4(32'h3a28f679),
	.w5(32'h3afaca9b),
	.w6(32'h3ace564a),
	.w7(32'h3aaaae12),
	.w8(32'hba668d89),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b584c),
	.w1(32'hb80658d9),
	.w2(32'h3a925e7b),
	.w3(32'hba683e53),
	.w4(32'h3affd270),
	.w5(32'h3b3a1dad),
	.w6(32'hbbc922a2),
	.w7(32'hbb3e512c),
	.w8(32'h3ace6d59),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b42fa),
	.w1(32'h3a3b21fe),
	.w2(32'h3a488bb2),
	.w3(32'h3a4f6336),
	.w4(32'h3b982871),
	.w5(32'h399a8a85),
	.w6(32'hba83eb89),
	.w7(32'h3a48ccaf),
	.w8(32'hbb5f0758),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb296d0d),
	.w1(32'h3b68ce1c),
	.w2(32'h3b0aecfb),
	.w3(32'h391c369d),
	.w4(32'h3aa28060),
	.w5(32'h3b9b2a74),
	.w6(32'hbac75a44),
	.w7(32'h3ad37b74),
	.w8(32'h3b1d5d4d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4208aa),
	.w1(32'hb933829e),
	.w2(32'hbab6c55d),
	.w3(32'h3ac05a42),
	.w4(32'hbb34ccad),
	.w5(32'hb7bfacd6),
	.w6(32'h39c75294),
	.w7(32'hbad27d89),
	.w8(32'hbb2b7a5d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89817c),
	.w1(32'h3a8b2551),
	.w2(32'h3abb85bb),
	.w3(32'h3aabccda),
	.w4(32'h3a80302f),
	.w5(32'hb997f945),
	.w6(32'h3b34d50d),
	.w7(32'hbad7b467),
	.w8(32'hbaa51f0f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ed150),
	.w1(32'h38e35143),
	.w2(32'hbb5b9463),
	.w3(32'h3a72a17a),
	.w4(32'h3a9ce0c8),
	.w5(32'hbb483544),
	.w6(32'hbae987f5),
	.w7(32'hba0aaa9a),
	.w8(32'hbbac0e10),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77ad0f),
	.w1(32'hbb3511dc),
	.w2(32'hbbb212e0),
	.w3(32'h3a085fb5),
	.w4(32'hba47c1ff),
	.w5(32'h3a9f2010),
	.w6(32'hbb80e66a),
	.w7(32'hba476ba7),
	.w8(32'hb8623e07),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb426059),
	.w1(32'hba886c8d),
	.w2(32'hb97f3f0d),
	.w3(32'hba6437e2),
	.w4(32'h3aa136ed),
	.w5(32'h3b063b18),
	.w6(32'hbb6c7c1d),
	.w7(32'hbabc1895),
	.w8(32'hba87e4de),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb812830),
	.w1(32'hbbd3e458),
	.w2(32'hbb2266ec),
	.w3(32'h3a9a9edf),
	.w4(32'hba9428f3),
	.w5(32'h3ae44d63),
	.w6(32'hba6348ee),
	.w7(32'h3b0eee13),
	.w8(32'h3ac9c7ec),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2394dc),
	.w1(32'h3b1e90aa),
	.w2(32'hba0c4be1),
	.w3(32'h3aa815b1),
	.w4(32'h3b3661f0),
	.w5(32'h3ae69f65),
	.w6(32'hb95b6b99),
	.w7(32'h3b42ccc8),
	.w8(32'hbb11445a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe80d1),
	.w1(32'hbb1c6d2b),
	.w2(32'hbab38d85),
	.w3(32'h3ae6b503),
	.w4(32'h3b3af8a5),
	.w5(32'h39fea7d0),
	.w6(32'hba996b17),
	.w7(32'hb91a9e40),
	.w8(32'h3a33a59c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d2df4),
	.w1(32'hbbe06395),
	.w2(32'hbb8999f6),
	.w3(32'hbac84c10),
	.w4(32'hbaddff29),
	.w5(32'h3a4df44e),
	.w6(32'h3b2edaee),
	.w7(32'h3b81c009),
	.w8(32'h3b1ec5b1),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d6748),
	.w1(32'hb99a995d),
	.w2(32'h3ad1c26c),
	.w3(32'hbb455913),
	.w4(32'h3b812b2e),
	.w5(32'h3aa0ba39),
	.w6(32'hbb37058d),
	.w7(32'h3a72aa82),
	.w8(32'hba3ebd6c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e5227),
	.w1(32'h3bce846b),
	.w2(32'hba865a1e),
	.w3(32'hbb17bd39),
	.w4(32'h3aef4a08),
	.w5(32'hbbb54424),
	.w6(32'hbc3164b2),
	.w7(32'hbbb8c757),
	.w8(32'hbc23b137),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaca582),
	.w1(32'hbac06891),
	.w2(32'hba9f1e26),
	.w3(32'hba9400f7),
	.w4(32'hb94348b6),
	.w5(32'hba2b6b58),
	.w6(32'hbaba0507),
	.w7(32'h3a556fef),
	.w8(32'hb9d17630),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f2113),
	.w1(32'h3ae7716c),
	.w2(32'h3b2a3b78),
	.w3(32'hbb720e76),
	.w4(32'h3ad24249),
	.w5(32'hba86ebce),
	.w6(32'hbb86ca31),
	.w7(32'hb80ccc2e),
	.w8(32'hbae63e80),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d8d31),
	.w1(32'hba017eb0),
	.w2(32'hb9c8b776),
	.w3(32'hb971f407),
	.w4(32'h37a4f3d3),
	.w5(32'hbb0425ab),
	.w6(32'h3a405111),
	.w7(32'h3a8711a2),
	.w8(32'h37b0a216),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7cee1),
	.w1(32'hbb32eb19),
	.w2(32'hbbbf562b),
	.w3(32'hbb46b7bc),
	.w4(32'h3b1730e4),
	.w5(32'hbb8975c2),
	.w6(32'hbbd1d81f),
	.w7(32'hbba81125),
	.w8(32'hbc0eed58),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31b0ae),
	.w1(32'hbaec0c4a),
	.w2(32'hbb61a28d),
	.w3(32'hbadf07ec),
	.w4(32'h3970f721),
	.w5(32'hbaea2264),
	.w6(32'hbb71b601),
	.w7(32'hbb029076),
	.w8(32'hbad0030a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1889aa),
	.w1(32'h392f9045),
	.w2(32'hbbc02d05),
	.w3(32'hbab3fc70),
	.w4(32'hb9a2e9a4),
	.w5(32'hbb1bfcec),
	.w6(32'hbae1921b),
	.w7(32'hbb51b492),
	.w8(32'hbb93cbd6),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d4f50),
	.w1(32'h3a17499f),
	.w2(32'h3af9df1f),
	.w3(32'h3a91b7dd),
	.w4(32'h3a43f80a),
	.w5(32'hba1c2044),
	.w6(32'h3a6d836f),
	.w7(32'h3a8dd96a),
	.w8(32'hbaa7a46f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf50f7b),
	.w1(32'hbb4de47a),
	.w2(32'hbb83f999),
	.w3(32'h3a30c638),
	.w4(32'hbb043405),
	.w5(32'hb9a6c360),
	.w6(32'hbaddb63c),
	.w7(32'hbb85d6ab),
	.w8(32'hba95c7d3),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20c058),
	.w1(32'hb9b3952c),
	.w2(32'h390bd8b9),
	.w3(32'h3a5b0a5c),
	.w4(32'h3ad0bd85),
	.w5(32'hbb5af360),
	.w6(32'h3a162a95),
	.w7(32'h3ad1d89e),
	.w8(32'hbb15a14e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cfdba),
	.w1(32'hbbaa9beb),
	.w2(32'hbb33b504),
	.w3(32'hbb1ec6a9),
	.w4(32'hb9d79494),
	.w5(32'h3a85f181),
	.w6(32'hbbbfa49f),
	.w7(32'hbac4ee2b),
	.w8(32'h3a8d0909),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9194f70),
	.w1(32'h3a85cc69),
	.w2(32'h3b1b61ef),
	.w3(32'h3a333aa9),
	.w4(32'h3a7e4be2),
	.w5(32'h39eb140a),
	.w6(32'hba0c4a37),
	.w7(32'h3a6e9078),
	.w8(32'hbb67fe00),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4049d4),
	.w1(32'hbafd93e0),
	.w2(32'hbbb0c8c8),
	.w3(32'hbaeb4c49),
	.w4(32'hbb354447),
	.w5(32'hb9b91960),
	.w6(32'hbb971459),
	.w7(32'hbbb72761),
	.w8(32'hbb3887af),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e8ae0),
	.w1(32'h3a5ac6ee),
	.w2(32'hbad5f302),
	.w3(32'h3aeee79c),
	.w4(32'h3a4aabfc),
	.w5(32'hb9ae47aa),
	.w6(32'h3b2dcada),
	.w7(32'h3a645899),
	.w8(32'hbb000efe),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391ae862),
	.w1(32'hb9921487),
	.w2(32'h394e73d5),
	.w3(32'h3a8aa819),
	.w4(32'h397c1b6f),
	.w5(32'hb9ae714d),
	.w6(32'hbafc3783),
	.w7(32'hbb13a066),
	.w8(32'hbabdf046),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacad76f),
	.w1(32'hbaab5f7a),
	.w2(32'hbac9f7c5),
	.w3(32'hba9689d1),
	.w4(32'h3ac6a327),
	.w5(32'h385ff5a8),
	.w6(32'hbb9f2182),
	.w7(32'hbb713439),
	.w8(32'hb8200e4b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f10718),
	.w1(32'h3ac36b0b),
	.w2(32'hbb020092),
	.w3(32'hba928c81),
	.w4(32'h3b4249df),
	.w5(32'hbb1010bf),
	.w6(32'hbb453eb5),
	.w7(32'h37ad3f04),
	.w8(32'hbb761f16),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fc9d4),
	.w1(32'h3b769b3c),
	.w2(32'hbae1894c),
	.w3(32'hbbb10ae9),
	.w4(32'h3b5e0543),
	.w5(32'h3ad5a0fd),
	.w6(32'hbba58d74),
	.w7(32'h3b174f8b),
	.w8(32'h3865dc74),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h359c1386),
	.w1(32'hba736fea),
	.w2(32'hba09efe9),
	.w3(32'hb89082f4),
	.w4(32'h39353eba),
	.w5(32'h3b61f829),
	.w6(32'hbaabaf5e),
	.w7(32'h3a2697d1),
	.w8(32'hba87269d),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd592f),
	.w1(32'h3b21b0a8),
	.w2(32'hbb807921),
	.w3(32'h3b33e604),
	.w4(32'h3b91b165),
	.w5(32'hbc0a90e3),
	.w6(32'hbb697549),
	.w7(32'hbaf6c271),
	.w8(32'hbc218dd7),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc020555),
	.w1(32'hbb0690a0),
	.w2(32'hbaf3a7a2),
	.w3(32'hbb205bea),
	.w4(32'h3a228489),
	.w5(32'h3a12eecf),
	.w6(32'hbb6c6cf1),
	.w7(32'hbb1ff46f),
	.w8(32'hbba43b51),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998b533),
	.w1(32'hba717bd5),
	.w2(32'hbae50a7d),
	.w3(32'hbb2d9110),
	.w4(32'hbb0aaeb1),
	.w5(32'h3a6de83d),
	.w6(32'hbb118567),
	.w7(32'hbac2c0e4),
	.w8(32'hbb290960),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade7ecd),
	.w1(32'hba89a663),
	.w2(32'hba2ce57b),
	.w3(32'h39e4e5fc),
	.w4(32'h3acd30bb),
	.w5(32'h3ac70aba),
	.w6(32'hbae550e1),
	.w7(32'hbb1ed8a3),
	.w8(32'h3ac7d1d5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a392d),
	.w1(32'hba296450),
	.w2(32'hba4578d3),
	.w3(32'h3ac0b1e7),
	.w4(32'h3ae7c9b0),
	.w5(32'h3a430408),
	.w6(32'h39a1695a),
	.w7(32'h3a8c5d0b),
	.w8(32'h3a8e6f05),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba492ef8),
	.w1(32'h3af8759a),
	.w2(32'h39ba163c),
	.w3(32'h3ad89002),
	.w4(32'h3b0a6dbe),
	.w5(32'hbad60600),
	.w6(32'hba0f0045),
	.w7(32'h39f042a7),
	.w8(32'hbb8f1c9b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fe526),
	.w1(32'h3b48f442),
	.w2(32'hba8c5c2b),
	.w3(32'h3ad189de),
	.w4(32'h3a20140e),
	.w5(32'h3a5f7d71),
	.w6(32'hbb7bb5a9),
	.w7(32'hbb8f0905),
	.w8(32'hb8c7bac8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e0cab),
	.w1(32'h3a0f1b2a),
	.w2(32'hba13debb),
	.w3(32'h3a221a98),
	.w4(32'h3a27d647),
	.w5(32'hbb2dc246),
	.w6(32'hbb722318),
	.w7(32'hbb30266e),
	.w8(32'hbb8debf0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae9b93),
	.w1(32'h3a21bfd5),
	.w2(32'h3a267c22),
	.w3(32'hbbdc2b2b),
	.w4(32'h3a82ea8d),
	.w5(32'h39bb048d),
	.w6(32'hbba39045),
	.w7(32'h39b737d0),
	.w8(32'h3a9a3481),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a5d3f),
	.w1(32'hbb345526),
	.w2(32'h39848d4e),
	.w3(32'hba9ca483),
	.w4(32'h3a777af1),
	.w5(32'h385e6a6c),
	.w6(32'hbb02aa72),
	.w7(32'h398a1c11),
	.w8(32'hbaf9e6ec),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9998460),
	.w1(32'h3af4d01e),
	.w2(32'hbafcfb70),
	.w3(32'h3b8213c5),
	.w4(32'h3b8e3a85),
	.w5(32'hb9745b07),
	.w6(32'hbbcf10ca),
	.w7(32'h3817e67c),
	.w8(32'hbb183d3f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6989c6),
	.w1(32'h3b22acb9),
	.w2(32'h3ab98671),
	.w3(32'hbadab5da),
	.w4(32'hb9abd8e7),
	.w5(32'hbb2fa2e6),
	.w6(32'hbb1b3ec8),
	.w7(32'h3a1e3485),
	.w8(32'hbb865205),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac12ac6),
	.w1(32'hba3d42d2),
	.w2(32'hba3128b6),
	.w3(32'hbb821465),
	.w4(32'hbb203081),
	.w5(32'hbbceba76),
	.w6(32'h39a32204),
	.w7(32'h3b07022a),
	.w8(32'h3b58f59e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f46fcc),
	.w1(32'hbb6ce735),
	.w2(32'hbb6df08b),
	.w3(32'hbc484bfa),
	.w4(32'hbc0891aa),
	.w5(32'hbb596581),
	.w6(32'h3b2f2a51),
	.w7(32'h3b1b2459),
	.w8(32'hb9d65374),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3916f99d),
	.w1(32'hba13cecb),
	.w2(32'hba94c8ec),
	.w3(32'h3ae6a58c),
	.w4(32'h39b99dcb),
	.w5(32'h3a3e12c3),
	.w6(32'hba434356),
	.w7(32'h39be1300),
	.w8(32'hba9e90bf),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb241311),
	.w1(32'hbac35d70),
	.w2(32'hba8d2d1e),
	.w3(32'h39dcafda),
	.w4(32'h3b544cc4),
	.w5(32'h3a03aba6),
	.w6(32'hbbd59f1b),
	.w7(32'hbb20f903),
	.w8(32'hbb86d073),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa09d0),
	.w1(32'hbac4fa51),
	.w2(32'hb9a47f16),
	.w3(32'hbb53fcc5),
	.w4(32'h39fb0639),
	.w5(32'h3b76dd93),
	.w6(32'hbc1827c1),
	.w7(32'hbbd568ac),
	.w8(32'hbb029013),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3d1d4),
	.w1(32'h3b11f19e),
	.w2(32'h3a8dbbb1),
	.w3(32'hb9968ad2),
	.w4(32'h3aff6bfb),
	.w5(32'hb7cbe09a),
	.w6(32'hbb4b1ada),
	.w7(32'hba4e5938),
	.w8(32'hbb29d3fa),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cd766),
	.w1(32'hbb3fd62f),
	.w2(32'hbb1e2efb),
	.w3(32'hbac4adde),
	.w4(32'hbae877c5),
	.w5(32'h3aa85c44),
	.w6(32'hbb4d6cb8),
	.w7(32'hba9f3d8b),
	.w8(32'h3a272126),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbb76f),
	.w1(32'hbabcbe85),
	.w2(32'h3ac91452),
	.w3(32'hbb32a512),
	.w4(32'h3b0dc070),
	.w5(32'h3b310b55),
	.w6(32'hbb211759),
	.w7(32'hbaaea96e),
	.w8(32'hbaef1b0b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadacd30),
	.w1(32'hba9f2b55),
	.w2(32'hbb1aa577),
	.w3(32'h3b162bf0),
	.w4(32'h3a519930),
	.w5(32'hba0c1a80),
	.w6(32'hbaca3d63),
	.w7(32'hba8d7b64),
	.w8(32'hbb025d36),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb861f1d),
	.w1(32'h3b0d5dcd),
	.w2(32'hba9acd8f),
	.w3(32'hbaa56414),
	.w4(32'h3b571b8e),
	.w5(32'h3a1ec2b7),
	.w6(32'hbb5142ba),
	.w7(32'hba36b823),
	.w8(32'hbb43e432),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba093109),
	.w1(32'hbac15cf3),
	.w2(32'hbae6d611),
	.w3(32'h3a595126),
	.w4(32'h38fbf96c),
	.w5(32'h3b179994),
	.w6(32'hbb3a1b27),
	.w7(32'hba6b0fd5),
	.w8(32'h3b5210d5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af65361),
	.w1(32'h3b1a1054),
	.w2(32'h3a7de9b3),
	.w3(32'h3a70dd27),
	.w4(32'h39bd691e),
	.w5(32'h3a79640b),
	.w6(32'h3b1da7b9),
	.w7(32'h3b116087),
	.w8(32'hba5a2d69),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cad7e),
	.w1(32'h3b77965e),
	.w2(32'hb9d8ec7d),
	.w3(32'hba3da95a),
	.w4(32'h3b9144fd),
	.w5(32'h39d0a9e0),
	.w6(32'hbc1e6ff3),
	.w7(32'hbb9d5b42),
	.w8(32'hbbe4012c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d3525),
	.w1(32'h3baf47b9),
	.w2(32'hba610e51),
	.w3(32'hbac9d878),
	.w4(32'hba551ea9),
	.w5(32'hbbba11c7),
	.w6(32'hbbe28d38),
	.w7(32'hbb8faf33),
	.w8(32'hbc19425e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0a4bf),
	.w1(32'h3a5528a0),
	.w2(32'hb95204db),
	.w3(32'hba583bd5),
	.w4(32'h3ae425c2),
	.w5(32'hba8aa152),
	.w6(32'hbbabd9bc),
	.w7(32'hbb5e290d),
	.w8(32'hbb7385e7),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12609a),
	.w1(32'hbb6b1ff2),
	.w2(32'hbc2cb58f),
	.w3(32'h391705ba),
	.w4(32'hba19b1ec),
	.w5(32'hbb1522b6),
	.w6(32'h3b2bd527),
	.w7(32'hbb25cedb),
	.w8(32'hbadc349c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f28dc),
	.w1(32'h3ae71d72),
	.w2(32'h3a41702c),
	.w3(32'h3b059735),
	.w4(32'h3a10a9ac),
	.w5(32'h3a1bf098),
	.w6(32'h3b62b13f),
	.w7(32'h3aded807),
	.w8(32'h3a0cb830),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f59324),
	.w1(32'hbad946f4),
	.w2(32'hbab9817c),
	.w3(32'h3ac950eb),
	.w4(32'h3aab1249),
	.w5(32'hba838451),
	.w6(32'h3a43ee22),
	.w7(32'h3a9e4342),
	.w8(32'hbb15740c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b392457),
	.w1(32'h3c446c2b),
	.w2(32'hbaf3c4a3),
	.w3(32'h3b88729c),
	.w4(32'h3bd7aa30),
	.w5(32'hbb6827d1),
	.w6(32'hbc043229),
	.w7(32'hb92986df),
	.w8(32'hbbb852e8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927c81e),
	.w1(32'hbb11241e),
	.w2(32'hbbbc3c06),
	.w3(32'h3b1453e7),
	.w4(32'h3b38fbde),
	.w5(32'hbbf46921),
	.w6(32'hbb8cdbf2),
	.w7(32'hba4e622f),
	.w8(32'hbbd6666e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d86f7),
	.w1(32'h3b904953),
	.w2(32'hbb960c72),
	.w3(32'h3a872f39),
	.w4(32'h3b8f03aa),
	.w5(32'hbb8f5142),
	.w6(32'hbb9a98e3),
	.w7(32'hbafcbb41),
	.w8(32'hbbf878d9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafb0c3),
	.w1(32'hbb629372),
	.w2(32'hba7b9912),
	.w3(32'hbb91e8bb),
	.w4(32'hb95a146f),
	.w5(32'h3b75ee7d),
	.w6(32'hbbba6d77),
	.w7(32'hbb012294),
	.w8(32'hba45bde5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb82125),
	.w1(32'hbaa99892),
	.w2(32'h3aa2245d),
	.w3(32'hbab4ad7c),
	.w4(32'h3b339f06),
	.w5(32'h3b8de4cc),
	.w6(32'hbba5dc77),
	.w7(32'hbb4d9937),
	.w8(32'hbb3d3372),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fff0e),
	.w1(32'hbb00e753),
	.w2(32'hbb00016c),
	.w3(32'h39dce30a),
	.w4(32'h39a98136),
	.w5(32'h3a8ff18f),
	.w6(32'hb980079d),
	.w7(32'h3a8ee659),
	.w8(32'hbb3f0bb9),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53a405),
	.w1(32'hba5c44dd),
	.w2(32'hba1c3301),
	.w3(32'h3a449513),
	.w4(32'h3b1d4898),
	.w5(32'h3aeff189),
	.w6(32'hb9c500f0),
	.w7(32'hbb00313d),
	.w8(32'hb93f6896),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99af56b),
	.w1(32'hba9fb2c6),
	.w2(32'hb678997e),
	.w3(32'hba07ab48),
	.w4(32'h3a949888),
	.w5(32'hbb071bc7),
	.w6(32'hba478921),
	.w7(32'hb9cce12b),
	.w8(32'h3993644b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90bb8a),
	.w1(32'h3a8d4a5d),
	.w2(32'hba9b89a5),
	.w3(32'h3a925dba),
	.w4(32'hbb559b20),
	.w5(32'hb7dcf99c),
	.w6(32'h3aa63128),
	.w7(32'hba841a7f),
	.w8(32'hb99b16e2),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba363bf0),
	.w1(32'hbb00f60e),
	.w2(32'hbb79cb68),
	.w3(32'h39eec964),
	.w4(32'hba2d6c53),
	.w5(32'hbb6df91e),
	.w6(32'hb90b938a),
	.w7(32'hbb3b8f23),
	.w8(32'hbba3a35e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c111c),
	.w1(32'h3a982955),
	.w2(32'hbba74c89),
	.w3(32'hbb78cc18),
	.w4(32'hbb38e4e4),
	.w5(32'hbb22996a),
	.w6(32'hbc2d0c5a),
	.w7(32'hbbe07588),
	.w8(32'hbbd6e912),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7252b),
	.w1(32'h3aa16fb4),
	.w2(32'h39fb6fd2),
	.w3(32'hbb601942),
	.w4(32'h3a862cab),
	.w5(32'hbaf39f0b),
	.w6(32'hbaf98970),
	.w7(32'hbb19284e),
	.w8(32'hb9d2cc02),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90ed14),
	.w1(32'hbb140e7b),
	.w2(32'hbb69f5f3),
	.w3(32'h3aef682c),
	.w4(32'h3ba23356),
	.w5(32'h3a87becd),
	.w6(32'h3bb5fc35),
	.w7(32'h3b71dedf),
	.w8(32'h368cabbb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a102ef8),
	.w1(32'h3af1a7b0),
	.w2(32'hbbdcab68),
	.w3(32'h3a9a5769),
	.w4(32'h3bc7e0e7),
	.w5(32'hbb824aff),
	.w6(32'hbbce258f),
	.w7(32'hbb3994d6),
	.w8(32'hbbe363da),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb5319),
	.w1(32'hba1bb683),
	.w2(32'hbba3d86d),
	.w3(32'h3abad4a7),
	.w4(32'h3a9dbb00),
	.w5(32'hba53301f),
	.w6(32'hbb34b183),
	.w7(32'hbb122b3b),
	.w8(32'hbc0f4a45),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7e497),
	.w1(32'hbb1f10e4),
	.w2(32'hbb1e71ac),
	.w3(32'hbb3e78a8),
	.w4(32'hbbfcd2ff),
	.w5(32'h39d66eae),
	.w6(32'hbc03ebfe),
	.w7(32'hbbc89706),
	.w8(32'h3b1821e5),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88a251),
	.w1(32'h3b084aef),
	.w2(32'hbaf70de2),
	.w3(32'h3917f6ba),
	.w4(32'h39c11c5a),
	.w5(32'hbb6abc30),
	.w6(32'h37d90237),
	.w7(32'hba9a2c9a),
	.w8(32'hbc0e4cfe),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39ce86),
	.w1(32'h3add4418),
	.w2(32'hbb9b1c2a),
	.w3(32'hbbb20984),
	.w4(32'hbba2b900),
	.w5(32'h3b24fcd2),
	.w6(32'hba4bd3f7),
	.w7(32'h3a088acb),
	.w8(32'hba2da668),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40fa96),
	.w1(32'hbadb8a6c),
	.w2(32'h394a3ba8),
	.w3(32'hb9996716),
	.w4(32'hbaedb423),
	.w5(32'h3a7a9bd0),
	.w6(32'h3ac165da),
	.w7(32'hbb107355),
	.w8(32'hba2e0a01),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e95e62),
	.w1(32'hbafc3c90),
	.w2(32'hbb3e6887),
	.w3(32'h39d9a6eb),
	.w4(32'hb98fd5c6),
	.w5(32'hba00eb9e),
	.w6(32'h39b35187),
	.w7(32'hbb286720),
	.w8(32'h3b7d59ed),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ced36),
	.w1(32'hbae31d2f),
	.w2(32'hbc0a4204),
	.w3(32'h38ac6e11),
	.w4(32'h3ad0d8c2),
	.w5(32'hbbbf3beb),
	.w6(32'h3bbb960d),
	.w7(32'hbb66dcd1),
	.w8(32'hbb6a2e2a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8ab69),
	.w1(32'h3836d547),
	.w2(32'hbb8e2e58),
	.w3(32'hbbb4d5db),
	.w4(32'h3b28e15f),
	.w5(32'h3b387f07),
	.w6(32'h39503392),
	.w7(32'hbaeb34b3),
	.w8(32'h3b1896fc),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980722c),
	.w1(32'hb9fc4168),
	.w2(32'hbb8ee050),
	.w3(32'hbae0c03e),
	.w4(32'h39c9570f),
	.w5(32'hbb9f448d),
	.w6(32'hba466062),
	.w7(32'h3aa423c7),
	.w8(32'hbc1cb21d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba35117),
	.w1(32'h3b92d5d0),
	.w2(32'hbba0f419),
	.w3(32'hbacef2b2),
	.w4(32'hb9b39e1d),
	.w5(32'hbb4df13f),
	.w6(32'h385387b8),
	.w7(32'hbabfd5eb),
	.w8(32'hbb8bd9f6),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88dc60),
	.w1(32'h3a0ca852),
	.w2(32'hbaff4fc2),
	.w3(32'h3af0d1f0),
	.w4(32'hbac58578),
	.w5(32'h3ae321de),
	.w6(32'hbb46a13d),
	.w7(32'hbb55214a),
	.w8(32'hbb34bbd7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67eedb),
	.w1(32'h3a85d347),
	.w2(32'h3bd3ab24),
	.w3(32'h3aef690b),
	.w4(32'h3b8b6e27),
	.w5(32'hbb8006e5),
	.w6(32'hb9c659df),
	.w7(32'h3aa7bfb2),
	.w8(32'hb99711f0),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3abefc),
	.w1(32'hbb420ec8),
	.w2(32'hba4971b7),
	.w3(32'hbb893207),
	.w4(32'hbb0745b0),
	.w5(32'h3bd1ab29),
	.w6(32'h3b14a653),
	.w7(32'h3b1d033b),
	.w8(32'h3bab964f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c6c69),
	.w1(32'hb9a89882),
	.w2(32'h3a61ea20),
	.w3(32'h3bed4c73),
	.w4(32'h3b79c1e8),
	.w5(32'h3b6300f0),
	.w6(32'hba9b13f2),
	.w7(32'hbac0a054),
	.w8(32'h3b790211),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2d3d2),
	.w1(32'h3aa575f1),
	.w2(32'h3aaaa9d3),
	.w3(32'h3abff473),
	.w4(32'h3a79b873),
	.w5(32'h3b46fc11),
	.w6(32'h3b455caa),
	.w7(32'h3af4e33f),
	.w8(32'h3ac0b20b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a327679),
	.w1(32'hbaf094a2),
	.w2(32'hbbccb0c6),
	.w3(32'h3b454f44),
	.w4(32'hba552163),
	.w5(32'hbbaa80f4),
	.w6(32'hbb267268),
	.w7(32'hbbaa39c6),
	.w8(32'hbbcb8b5c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef7bbd),
	.w1(32'hbb56f346),
	.w2(32'hbb83d792),
	.w3(32'hbb2d9004),
	.w4(32'h37baf710),
	.w5(32'h3a0c7e7a),
	.w6(32'h3a4671c0),
	.w7(32'hbb4ee7c2),
	.w8(32'h3a906f4d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80fad0),
	.w1(32'h3bace55d),
	.w2(32'h3bb28a36),
	.w3(32'hbb5c053a),
	.w4(32'hbaa71d79),
	.w5(32'h3afa6a33),
	.w6(32'h3b2e39c4),
	.w7(32'h3bcfcf49),
	.w8(32'hba02fa54),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eefe7),
	.w1(32'hbbb02681),
	.w2(32'hba96dcbb),
	.w3(32'h3ae04f5b),
	.w4(32'hbba8142a),
	.w5(32'hbbf0cbc9),
	.w6(32'hba3b0e62),
	.w7(32'hbba1d340),
	.w8(32'hb9360cb2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d2fb4),
	.w1(32'hbb19285e),
	.w2(32'hbb7b8cfc),
	.w3(32'hbc094305),
	.w4(32'h3ba857fb),
	.w5(32'h3ba391c7),
	.w6(32'h3c17cff7),
	.w7(32'h3b67b945),
	.w8(32'h3a092e79),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2872ba),
	.w1(32'h3b584604),
	.w2(32'h3a33a309),
	.w3(32'h3b54b084),
	.w4(32'h3ac29800),
	.w5(32'hbc00b2aa),
	.w6(32'h3a4f0fe7),
	.w7(32'hbb78011f),
	.w8(32'hbb99c0cc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad56986),
	.w1(32'hb9084064),
	.w2(32'hbb296a19),
	.w3(32'hbbd9a962),
	.w4(32'h3a6b6b4b),
	.w5(32'h3b8af347),
	.w6(32'h3b9c809c),
	.w7(32'h3bce95f9),
	.w8(32'h3b03cc50),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68f327),
	.w1(32'hbbf39fb4),
	.w2(32'hbc25ff60),
	.w3(32'h3bfdc397),
	.w4(32'h3a880450),
	.w5(32'hb89d1af5),
	.w6(32'hbab9a1be),
	.w7(32'hbc0c4902),
	.w8(32'hbc31cbca),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ada0d),
	.w1(32'hbaa50ad1),
	.w2(32'h3b2733db),
	.w3(32'hbb08c668),
	.w4(32'hbb89eaa2),
	.w5(32'h3b0fe3f0),
	.w6(32'hbb519502),
	.w7(32'hbb657af2),
	.w8(32'hb9eef16c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba878e6f),
	.w1(32'h3b84fad2),
	.w2(32'h3bcd0794),
	.w3(32'hbb040213),
	.w4(32'h3aaae788),
	.w5(32'hba1fa3ab),
	.w6(32'hbc17fd43),
	.w7(32'hbafb9101),
	.w8(32'hbb46f099),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule