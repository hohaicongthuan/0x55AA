module layer_10_featuremap_504(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d40c9),
	.w1(32'h3a9835dd),
	.w2(32'hba49f6df),
	.w3(32'hba7ea284),
	.w4(32'h3a871ccd),
	.w5(32'h3a0fbb57),
	.w6(32'hba9d7e83),
	.w7(32'h3a691d68),
	.w8(32'h3aac544d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00c3ec),
	.w1(32'hba9270ed),
	.w2(32'hbb2f546e),
	.w3(32'h3ac9d895),
	.w4(32'hba92f8d1),
	.w5(32'hbb229872),
	.w6(32'h3aa8d0ab),
	.w7(32'hbaac5809),
	.w8(32'hbb56a459),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d3fd9),
	.w1(32'hb9cfb1c3),
	.w2(32'h3a44aebe),
	.w3(32'hbaa6a23c),
	.w4(32'hbad68df2),
	.w5(32'hbab73318),
	.w6(32'hbada9554),
	.w7(32'h39ae22f9),
	.w8(32'hb815bbf2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b245613),
	.w1(32'hb8c81af5),
	.w2(32'h39db1916),
	.w3(32'h39c0d95e),
	.w4(32'hbb0167b6),
	.w5(32'h3b03b3b0),
	.w6(32'h3a2db291),
	.w7(32'hba2ea092),
	.w8(32'h3a835298),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba626d4a),
	.w1(32'h3a63be3d),
	.w2(32'h3a98ae1b),
	.w3(32'hb998e77a),
	.w4(32'h3ab9ba03),
	.w5(32'h3a31359a),
	.w6(32'hb8993ff0),
	.w7(32'h3a612aa7),
	.w8(32'hb6b205c6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b86d26),
	.w1(32'hb878fb15),
	.w2(32'hb95e9a72),
	.w3(32'h3b241776),
	.w4(32'hba89db12),
	.w5(32'h39b4f461),
	.w6(32'h3a86d85e),
	.w7(32'hbac0689a),
	.w8(32'hba88fed6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2241ca),
	.w1(32'h3b962b69),
	.w2(32'h3ba768ec),
	.w3(32'h3aed22d3),
	.w4(32'h3b2c898d),
	.w5(32'h3b51aed5),
	.w6(32'h399bc85b),
	.w7(32'h3af449fa),
	.w8(32'h3b22860c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23e657),
	.w1(32'hbae9c312),
	.w2(32'h3aa99ee6),
	.w3(32'h3a16be28),
	.w4(32'hba16a6bf),
	.w5(32'hb9381dbd),
	.w6(32'hbba0f435),
	.w7(32'h3ab11495),
	.w8(32'h3bc841a0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e472d),
	.w1(32'h38af9bc2),
	.w2(32'h3b323411),
	.w3(32'hba431c4f),
	.w4(32'hb98e5910),
	.w5(32'h3a7cbda4),
	.w6(32'hbab63a56),
	.w7(32'h3aa219a3),
	.w8(32'h3a62d366),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0fb2e),
	.w1(32'hb7b927a9),
	.w2(32'h3b53a7ec),
	.w3(32'h3b82c9c1),
	.w4(32'h3b29a9db),
	.w5(32'h3ba8e7cd),
	.w6(32'h3b37900e),
	.w7(32'h3b78891e),
	.w8(32'h3b22d88e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38859940),
	.w1(32'hba84f82e),
	.w2(32'hb9cdb363),
	.w3(32'h3a1ba7b6),
	.w4(32'h38bec7ef),
	.w5(32'hba267933),
	.w6(32'hb9a79382),
	.w7(32'h3914de4a),
	.w8(32'hb7854ad7),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2de670),
	.w1(32'h3b6ef405),
	.w2(32'h3bc66150),
	.w3(32'hba0f4896),
	.w4(32'h3b36cec9),
	.w5(32'h3bc15b89),
	.w6(32'hbb85dadd),
	.w7(32'h3ac1b56a),
	.w8(32'h3b95eb5b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39850199),
	.w1(32'h3a99742e),
	.w2(32'h3a8176c0),
	.w3(32'h3b0a1355),
	.w4(32'h3b6c3af4),
	.w5(32'h3b6f7e47),
	.w6(32'h3b46e151),
	.w7(32'h3b1d9848),
	.w8(32'h3aaf0700),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcc08e),
	.w1(32'h3a57ffe3),
	.w2(32'h3ac42368),
	.w3(32'hba626da8),
	.w4(32'h3a85543a),
	.w5(32'hbacf2717),
	.w6(32'h39897d0f),
	.w7(32'h3a8c0ddb),
	.w8(32'hba35c8f8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e1a98),
	.w1(32'hbb3b8d35),
	.w2(32'hbb78ec87),
	.w3(32'h3b84fb6b),
	.w4(32'hbaf81a1b),
	.w5(32'hbb9723c8),
	.w6(32'h3a64f582),
	.w7(32'hbb33c088),
	.w8(32'hbb5cab2e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb2b3c),
	.w1(32'h3aefd03e),
	.w2(32'h3b6b017f),
	.w3(32'h39eab3a7),
	.w4(32'h3aec4dcd),
	.w5(32'h3ba06403),
	.w6(32'hba3a8bef),
	.w7(32'h3b23a200),
	.w8(32'h3ba88572),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cb24a),
	.w1(32'hba8fb9ee),
	.w2(32'hba5ed1ef),
	.w3(32'h37e94513),
	.w4(32'hbaf661c8),
	.w5(32'hbabb1997),
	.w6(32'hba3729c8),
	.w7(32'hbadf5183),
	.w8(32'hba85078c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76b4ef),
	.w1(32'hb83f66bd),
	.w2(32'h3b20e050),
	.w3(32'hbb1e8f56),
	.w4(32'h3b87b7fa),
	.w5(32'h3b74d8e5),
	.w6(32'hbb587366),
	.w7(32'h3bde87ee),
	.w8(32'h3c1d676b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02ae2f),
	.w1(32'hb8fd1f73),
	.w2(32'h3b2df39f),
	.w3(32'hba96513f),
	.w4(32'h3b014b2f),
	.w5(32'h3b0a268a),
	.w6(32'h3aeb4477),
	.w7(32'h3b981b34),
	.w8(32'h3b840c5f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38e77d),
	.w1(32'hba241fb9),
	.w2(32'hba572a9d),
	.w3(32'h3a9cdc77),
	.w4(32'hbaded9be),
	.w5(32'h3a8567f2),
	.w6(32'hba120f97),
	.w7(32'hb9c7a3d6),
	.w8(32'h398eaa95),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38041075),
	.w1(32'hba13eed0),
	.w2(32'h39b6388e),
	.w3(32'hba510540),
	.w4(32'h3aa41b3a),
	.w5(32'h3b03bd87),
	.w6(32'hbafb8746),
	.w7(32'h3a4d28ed),
	.w8(32'h3a6d304f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8af79),
	.w1(32'hb9b4381d),
	.w2(32'hbaa6b261),
	.w3(32'h38fd80ba),
	.w4(32'hbaee1287),
	.w5(32'h384b2b3b),
	.w6(32'h396df8b0),
	.w7(32'hb9bb9cee),
	.w8(32'hbabd9730),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c7e4e),
	.w1(32'hbc040578),
	.w2(32'h3b34ffc2),
	.w3(32'hbb7b8801),
	.w4(32'hbb85dc39),
	.w5(32'h3a599da8),
	.w6(32'h3b0f4402),
	.w7(32'h3b201f40),
	.w8(32'h3b5412d7),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59013a),
	.w1(32'h393b4f85),
	.w2(32'h3979e55a),
	.w3(32'hb9188ea9),
	.w4(32'h3a920811),
	.w5(32'h3ac13456),
	.w6(32'h39a57a15),
	.w7(32'h3a9e802d),
	.w8(32'h3a7f6a19),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f2816),
	.w1(32'h395502bd),
	.w2(32'hbb760b66),
	.w3(32'h3ba2520c),
	.w4(32'h3a74ba3a),
	.w5(32'hbba0a789),
	.w6(32'h3bb13013),
	.w7(32'hbace0f12),
	.w8(32'hbb8d32a3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e511f),
	.w1(32'hb9c9e61c),
	.w2(32'hbaf75885),
	.w3(32'hba9cf8d7),
	.w4(32'hba37bae8),
	.w5(32'h3a84e214),
	.w6(32'hbb0d20eb),
	.w7(32'hba2aa4e7),
	.w8(32'hb982d630),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad48921),
	.w1(32'h3a8448cc),
	.w2(32'h3a127ff4),
	.w3(32'h3a4446b6),
	.w4(32'h3a9f4223),
	.w5(32'hb931bf4d),
	.w6(32'h3b30a70b),
	.w7(32'hba5ede29),
	.w8(32'h3a1d645e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb100823),
	.w1(32'h3b34a2e9),
	.w2(32'h3b639098),
	.w3(32'h3adbebe9),
	.w4(32'h39ec7bf0),
	.w5(32'hbb237278),
	.w6(32'hbb628f40),
	.w7(32'hbb785ec1),
	.w8(32'hbbb0938f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8744e1d),
	.w1(32'hba8ca941),
	.w2(32'hb9b1f538),
	.w3(32'hba7a6ecf),
	.w4(32'hba526447),
	.w5(32'hba3bd406),
	.w6(32'hba1e84fe),
	.w7(32'hbaaeb030),
	.w8(32'hba0d108d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2327aa),
	.w1(32'h3b8ab54a),
	.w2(32'h3b01a39b),
	.w3(32'h3b996cc6),
	.w4(32'h3b8411b9),
	.w5(32'hba93341d),
	.w6(32'h3ae7dd16),
	.w7(32'hb9ee2afb),
	.w8(32'hbbd5ef45),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af06684),
	.w1(32'h39715daf),
	.w2(32'hb8e604ad),
	.w3(32'h3b0760ec),
	.w4(32'h3921a613),
	.w5(32'h3aa740ad),
	.w6(32'h3acd96f1),
	.w7(32'h38ffac8c),
	.w8(32'hb8599353),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a22b74),
	.w1(32'h39e87829),
	.w2(32'h39f8da8a),
	.w3(32'hbaaedf9a),
	.w4(32'hb9db4032),
	.w5(32'hbb1c8a94),
	.w6(32'hb83f6096),
	.w7(32'h394e8ac0),
	.w8(32'hb8b1223f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad37de2),
	.w1(32'hba8fbe6a),
	.w2(32'hba9173b2),
	.w3(32'h3a672b85),
	.w4(32'hbacfc565),
	.w5(32'hbb03d0a1),
	.w6(32'h3a025eb5),
	.w7(32'h3a270ad0),
	.w8(32'hba3fd0cd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba513516),
	.w1(32'h3a174842),
	.w2(32'h3a86ae5f),
	.w3(32'h39a95c77),
	.w4(32'h3a45d031),
	.w5(32'h3a8b6c94),
	.w6(32'hba1cfeb5),
	.w7(32'hbace7e5c),
	.w8(32'hbaad17f2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f39ac),
	.w1(32'hba43e409),
	.w2(32'hb85f4908),
	.w3(32'h3a172e2c),
	.w4(32'hbac8a4bd),
	.w5(32'h38a9669f),
	.w6(32'h3847d096),
	.w7(32'hba20c8b5),
	.w8(32'h39fea988),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f87f2),
	.w1(32'h3a44a6af),
	.w2(32'h3a82beee),
	.w3(32'hba348112),
	.w4(32'h3a6eae52),
	.w5(32'h3b46af29),
	.w6(32'hbb1bba35),
	.w7(32'h3ad33f3f),
	.w8(32'h3b068022),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c2437),
	.w1(32'hbba83757),
	.w2(32'h3bbce121),
	.w3(32'h3b8a18ed),
	.w4(32'hbab907a5),
	.w5(32'h3bc53ae4),
	.w6(32'hba038f2a),
	.w7(32'hbacf4930),
	.w8(32'h3bfa00a9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b133b6f),
	.w1(32'h3acb4028),
	.w2(32'hbbe45fac),
	.w3(32'h3bc2a037),
	.w4(32'h381260dd),
	.w5(32'hbbfdface),
	.w6(32'h3b42c8d7),
	.w7(32'hbb106873),
	.w8(32'hbc1ebb83),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9076a3),
	.w1(32'h3ae6a805),
	.w2(32'hbbf9a6a5),
	.w3(32'h3b95ad31),
	.w4(32'h38e56a1c),
	.w5(32'hbc397bdd),
	.w6(32'h3b21d2db),
	.w7(32'hbb74895d),
	.w8(32'hbc4493c5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af14eb2),
	.w1(32'h39a2ac94),
	.w2(32'hbb07f061),
	.w3(32'h3afc9dbc),
	.w4(32'hb8e7f26a),
	.w5(32'hba98282b),
	.w6(32'h3b081eb2),
	.w7(32'hbae5fb00),
	.w8(32'hbae9b2fe),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9057429),
	.w1(32'hbacd1763),
	.w2(32'hbaf4189a),
	.w3(32'hba60da72),
	.w4(32'h3a2cd518),
	.w5(32'hb9796fb1),
	.w6(32'h3a491e6f),
	.w7(32'hb9f752cd),
	.w8(32'hbb443dc1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83a571),
	.w1(32'h391d33da),
	.w2(32'h3abb73b0),
	.w3(32'hbaa0ddbb),
	.w4(32'h3a7fa62e),
	.w5(32'h3ac86eb8),
	.w6(32'hb96a0a90),
	.w7(32'hba0b7b9c),
	.w8(32'h3a841992),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2e1b5),
	.w1(32'hba5edb2e),
	.w2(32'hba0163ce),
	.w3(32'hba7c6240),
	.w4(32'hba31b61a),
	.w5(32'h3ac395fa),
	.w6(32'hbb1eb94c),
	.w7(32'hba2aae7b),
	.w8(32'hba9e4584),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88389c),
	.w1(32'h3b3daaf1),
	.w2(32'h3b93151a),
	.w3(32'hba549ce9),
	.w4(32'h3b7c3a57),
	.w5(32'h3baea911),
	.w6(32'h3b151de4),
	.w7(32'h3b9d4dea),
	.w8(32'h3bca53a3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18cbf9),
	.w1(32'h377bb7b4),
	.w2(32'hba8fb297),
	.w3(32'h3b2cc283),
	.w4(32'h3b016e62),
	.w5(32'hb99fed2c),
	.w6(32'h3b10952c),
	.w7(32'hbaab3324),
	.w8(32'hbb36493f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba294729),
	.w1(32'hba7a2344),
	.w2(32'hbae472ad),
	.w3(32'h3a318b16),
	.w4(32'h3b07430e),
	.w5(32'h3aeb1b8d),
	.w6(32'h3afde1be),
	.w7(32'h3af442a6),
	.w8(32'h37fadde3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a6adb),
	.w1(32'hba071f62),
	.w2(32'h39bb474b),
	.w3(32'h3a88c10d),
	.w4(32'h3ac615a5),
	.w5(32'h3a510795),
	.w6(32'hba07ddf9),
	.w7(32'hb99e1ad8),
	.w8(32'hba130f27),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6da0c),
	.w1(32'hbad53b60),
	.w2(32'h3b75bfa1),
	.w3(32'hbb2c83d9),
	.w4(32'h3b92dbc4),
	.w5(32'h3bd2f399),
	.w6(32'hbb0eafad),
	.w7(32'h3c0a4463),
	.w8(32'h3c08ce0e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e21022),
	.w1(32'h3a064b7e),
	.w2(32'h3a069ef4),
	.w3(32'hba512bd1),
	.w4(32'h3ab5baae),
	.w5(32'hb9a7d723),
	.w6(32'h3a069078),
	.w7(32'h3b03a0ed),
	.w8(32'hba0bed6c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e688ec),
	.w1(32'hba96ad99),
	.w2(32'h3ab0aec1),
	.w3(32'h3a9592d1),
	.w4(32'h3a8f1af2),
	.w5(32'h3afd17f3),
	.w6(32'hba1d8c8a),
	.w7(32'hb99e87fe),
	.w8(32'h3a95468e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af71517),
	.w1(32'hbaa49b97),
	.w2(32'hb8eca16c),
	.w3(32'h3acaac7a),
	.w4(32'hbad6c815),
	.w5(32'h3aed53e0),
	.w6(32'h3af84a39),
	.w7(32'hbb23fa7b),
	.w8(32'hba911f9e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7cd08),
	.w1(32'hb9a92e11),
	.w2(32'h3a90b005),
	.w3(32'hbaa18217),
	.w4(32'hba35374b),
	.w5(32'h3ac7358d),
	.w6(32'hb9a50048),
	.w7(32'h3aaa9186),
	.w8(32'h3a10b000),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6f830),
	.w1(32'h3a7225a6),
	.w2(32'h3a9103b9),
	.w3(32'hba640eae),
	.w4(32'h3ae351a7),
	.w5(32'h3abf6d46),
	.w6(32'hbb2131cd),
	.w7(32'h3b044d46),
	.w8(32'h3a921cb2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbce86),
	.w1(32'h3a348ffd),
	.w2(32'h3b905b79),
	.w3(32'h3944f57f),
	.w4(32'h3b847feb),
	.w5(32'h3b5f982e),
	.w6(32'h3935b556),
	.w7(32'h3bd38ed7),
	.w8(32'h3bd7834b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7efde4),
	.w1(32'h3aa2f61a),
	.w2(32'h3abc9142),
	.w3(32'hb88b2cb8),
	.w4(32'hb7074748),
	.w5(32'h3aaeb284),
	.w6(32'h39efa515),
	.w7(32'hba90c513),
	.w8(32'h3b14e858),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1dee90),
	.w1(32'h3a986806),
	.w2(32'hb7c9561a),
	.w3(32'h3abcc857),
	.w4(32'h3a8aae8c),
	.w5(32'hbb57b701),
	.w6(32'h3a9fbf1f),
	.w7(32'h3aa30397),
	.w8(32'hba563510),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39710555),
	.w1(32'h3a9824cf),
	.w2(32'h38c68836),
	.w3(32'h393e14ab),
	.w4(32'h3a8d2f1b),
	.w5(32'hb98fb969),
	.w6(32'hba08e570),
	.w7(32'h39ccdd35),
	.w8(32'hb9d54c47),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe4323),
	.w1(32'hb9fe928f),
	.w2(32'hb97538ea),
	.w3(32'h3b01255e),
	.w4(32'hba628d26),
	.w5(32'h3ac339e8),
	.w6(32'h3a6dd8e2),
	.w7(32'hb9d15737),
	.w8(32'hbadca573),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9e1dc),
	.w1(32'hb8813f5d),
	.w2(32'h3a481a5d),
	.w3(32'hb966f222),
	.w4(32'h39844c4a),
	.w5(32'h3b0f1460),
	.w6(32'hb9ac239d),
	.w7(32'hb9947a88),
	.w8(32'h3a9147c8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88844a),
	.w1(32'hbac002c6),
	.w2(32'hba4b8c06),
	.w3(32'h3a120ac1),
	.w4(32'hba1f56d0),
	.w5(32'hba51f4d3),
	.w6(32'h3a056deb),
	.w7(32'hba784b16),
	.w8(32'hba973227),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae78a3d),
	.w1(32'h3b1c20fb),
	.w2(32'h3b4ad3b3),
	.w3(32'hbb02469f),
	.w4(32'h3af9907d),
	.w5(32'h3b81255c),
	.w6(32'hb9fedfb9),
	.w7(32'h3ae49f3d),
	.w8(32'h3baeca1b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4737eb),
	.w1(32'hb9092a17),
	.w2(32'h3af2920a),
	.w3(32'hbafa7c41),
	.w4(32'h3a648410),
	.w5(32'h3a8bed5c),
	.w6(32'h3ae357de),
	.w7(32'h3ad7061c),
	.w8(32'h3b81df6e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b220394),
	.w1(32'hbb5c29fd),
	.w2(32'hbab1e85c),
	.w3(32'h3a69fc48),
	.w4(32'hbb55a033),
	.w5(32'hb8ba692c),
	.w6(32'h3a2d9194),
	.w7(32'hbb28fe29),
	.w8(32'hb62262ff),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7e4be),
	.w1(32'h3a0a9bda),
	.w2(32'h3a914929),
	.w3(32'hba951d18),
	.w4(32'hb8d63279),
	.w5(32'h3860271b),
	.w6(32'hba03f778),
	.w7(32'hb8002931),
	.w8(32'hba4ae454),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25719a),
	.w1(32'h3b8856d7),
	.w2(32'h3b04d06c),
	.w3(32'h38552372),
	.w4(32'h3b46b02a),
	.w5(32'hb9ea860d),
	.w6(32'h39095a00),
	.w7(32'h3b33d9f8),
	.w8(32'h3aa7292c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20be74),
	.w1(32'h3a8377e1),
	.w2(32'h3a4bbb81),
	.w3(32'h3aeb8c56),
	.w4(32'h3b062a2f),
	.w5(32'h39587cd6),
	.w6(32'h3b6f4696),
	.w7(32'h3b088945),
	.w8(32'h3b08d39a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcb537),
	.w1(32'h3b7deace),
	.w2(32'h3bc5e39b),
	.w3(32'h3b5a4ee4),
	.w4(32'h3a9edd44),
	.w5(32'h3b636d5f),
	.w6(32'hb9833451),
	.w7(32'h3b94e6ee),
	.w8(32'h3b4ef6ac),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeaefca),
	.w1(32'h3aeb41fc),
	.w2(32'h3a6e0687),
	.w3(32'hbb4df679),
	.w4(32'hb90d7463),
	.w5(32'h3b0532e3),
	.w6(32'hba6dd3a8),
	.w7(32'h3b8d9fd1),
	.w8(32'h3bd60a43),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc1822),
	.w1(32'h3a3fe1f7),
	.w2(32'h3b456d98),
	.w3(32'hba285771),
	.w4(32'h3b0cc4cb),
	.w5(32'h3b9abad3),
	.w6(32'h3ad42637),
	.w7(32'h3b7049bf),
	.w8(32'h3be8d214),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8890e5),
	.w1(32'h3c5b11f1),
	.w2(32'h3c54597f),
	.w3(32'h3ba872ed),
	.w4(32'h3b94f06e),
	.w5(32'h3bfbd830),
	.w6(32'h3bf76051),
	.w7(32'h3b355aa1),
	.w8(32'hbbd195d3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc83cd4),
	.w1(32'h3a8662fe),
	.w2(32'hbb957ba1),
	.w3(32'h3b57add9),
	.w4(32'h3af9d0f7),
	.w5(32'hbb0a4606),
	.w6(32'h3c5d87da),
	.w7(32'hba41b76d),
	.w8(32'hba9ff8f5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b4ef0),
	.w1(32'h3b4544c1),
	.w2(32'hb9af5c03),
	.w3(32'hb9f678f1),
	.w4(32'hbc033bd9),
	.w5(32'hbae8669f),
	.w6(32'hb83be3de),
	.w7(32'hbb14f28c),
	.w8(32'hbb44363b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20e6e3),
	.w1(32'h3965b714),
	.w2(32'h3a80f08f),
	.w3(32'hbaa8938f),
	.w4(32'hbb8c3df8),
	.w5(32'h3b714706),
	.w6(32'h39ebf259),
	.w7(32'hbb0a5cab),
	.w8(32'h3b1bc5e2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d8f18),
	.w1(32'hba551d31),
	.w2(32'h3aa7794e),
	.w3(32'h3b815145),
	.w4(32'h3b722347),
	.w5(32'h3b140aa4),
	.w6(32'h3a3ae975),
	.w7(32'hba42b98a),
	.w8(32'h3b28aab7),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35f80f),
	.w1(32'h38b199c6),
	.w2(32'hb98a4977),
	.w3(32'hba9839a4),
	.w4(32'h3b84e901),
	.w5(32'h3c3a7f05),
	.w6(32'hb911b6db),
	.w7(32'hbbbc0505),
	.w8(32'h3c11a7a0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e32b5),
	.w1(32'h3b631d42),
	.w2(32'h3b217979),
	.w3(32'hb9cb80c5),
	.w4(32'hbb1eba2a),
	.w5(32'h3c0a8454),
	.w6(32'h3b67adc1),
	.w7(32'hba998764),
	.w8(32'h3a54172c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c80d6),
	.w1(32'h3b623773),
	.w2(32'h3b90c2a3),
	.w3(32'hba8b97a8),
	.w4(32'h3b9e267e),
	.w5(32'h3b758186),
	.w6(32'hbab6b665),
	.w7(32'h3bf42ce6),
	.w8(32'h3c20d792),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e527fc),
	.w1(32'hbb943e61),
	.w2(32'hbb875588),
	.w3(32'h3ace934c),
	.w4(32'hbbbcca2a),
	.w5(32'hbbe3fc24),
	.w6(32'h3b4442ce),
	.w7(32'hb928ba25),
	.w8(32'hbc12eb1c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbda2a3),
	.w1(32'hbab31420),
	.w2(32'h3b1e798f),
	.w3(32'hbaf0f1f1),
	.w4(32'h3b263d5e),
	.w5(32'hbb34e2f2),
	.w6(32'hbbd03527),
	.w7(32'hb9e92068),
	.w8(32'h3b1cf7d1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07fd04),
	.w1(32'h3bba5a3c),
	.w2(32'h3a06ad16),
	.w3(32'h3b647f52),
	.w4(32'h3b9d9015),
	.w5(32'h3c115c58),
	.w6(32'h3a9416d0),
	.w7(32'h3aa9305e),
	.w8(32'h3c307fd2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a0143),
	.w1(32'h3bff22b0),
	.w2(32'h3c2ab918),
	.w3(32'h3b369c1d),
	.w4(32'h3b9f5c49),
	.w5(32'h3b745a6f),
	.w6(32'h3c212e2b),
	.w7(32'h3be2ec38),
	.w8(32'h3a7bebd9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54063c),
	.w1(32'h3a8bb932),
	.w2(32'hbaf10440),
	.w3(32'h3ba149c5),
	.w4(32'hbb137811),
	.w5(32'hbb22a885),
	.w6(32'h3ab70e3c),
	.w7(32'hb7a73236),
	.w8(32'hb9ce4e1c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac66d79),
	.w1(32'h3b53626b),
	.w2(32'h399e1cc4),
	.w3(32'hba4c75eb),
	.w4(32'h3a92b3da),
	.w5(32'hb92cb739),
	.w6(32'hbbc37b1c),
	.w7(32'hbb0b8168),
	.w8(32'hba7acf8e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49cd75),
	.w1(32'h3b844654),
	.w2(32'h39a4ed01),
	.w3(32'h3b3b3f77),
	.w4(32'h3c67ef38),
	.w5(32'h3c3432da),
	.w6(32'h3b133b3f),
	.w7(32'h3bf42d5d),
	.w8(32'h3b88d340),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b1cad),
	.w1(32'h39b87811),
	.w2(32'hb90c485e),
	.w3(32'h3c9678c8),
	.w4(32'hbaef11a0),
	.w5(32'h3b959ebc),
	.w6(32'hba3a3b56),
	.w7(32'hbaa4f6af),
	.w8(32'hba9ffda5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89ac918),
	.w1(32'h3b8237a4),
	.w2(32'h3b1ebd61),
	.w3(32'h3b6bfd6e),
	.w4(32'h39bf300f),
	.w5(32'h3c0afe61),
	.w6(32'hbb6b79c2),
	.w7(32'h3bbf6199),
	.w8(32'h3c01aca0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aead284),
	.w1(32'hbb92d910),
	.w2(32'hbc2f2a77),
	.w3(32'h3c055dfa),
	.w4(32'h3bc01544),
	.w5(32'h3c6bb3cb),
	.w6(32'h3b8e8272),
	.w7(32'hbbdca784),
	.w8(32'h3c0e76e7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7dfde),
	.w1(32'hbb83b6f9),
	.w2(32'hbc01cc12),
	.w3(32'h39147f72),
	.w4(32'h3b972a0f),
	.w5(32'h3bde4c35),
	.w6(32'h3b5ce19c),
	.w7(32'hbb8d573a),
	.w8(32'h3bec58e1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc126b28),
	.w1(32'h3aa2fa82),
	.w2(32'h3b0ce33c),
	.w3(32'hbb847f6d),
	.w4(32'h3b87518c),
	.w5(32'h3bda812e),
	.w6(32'h3b1aa290),
	.w7(32'h3ba2fbc8),
	.w8(32'h3beeb464),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3e132),
	.w1(32'hbba0e2ea),
	.w2(32'h3c00e139),
	.w3(32'h3ae73f91),
	.w4(32'hbb348840),
	.w5(32'h38e0d551),
	.w6(32'h3b9202ef),
	.w7(32'h3b511341),
	.w8(32'h3b95ae90),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bc8bb),
	.w1(32'hba28a32d),
	.w2(32'hbb589e7f),
	.w3(32'h3b7e8ac8),
	.w4(32'hbada1bf5),
	.w5(32'hb9c49f80),
	.w6(32'hbb85244a),
	.w7(32'h3b9a6955),
	.w8(32'hbc06f36f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb483db),
	.w1(32'h3b432704),
	.w2(32'h3c0ea207),
	.w3(32'hbb977c47),
	.w4(32'h3b918e51),
	.w5(32'h3bef0249),
	.w6(32'hbbe57bed),
	.w7(32'hbb03f306),
	.w8(32'h3af8936e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dda9e),
	.w1(32'h3b48153b),
	.w2(32'hbb6fa76b),
	.w3(32'h3c15d822),
	.w4(32'hbb5979ad),
	.w5(32'hbbb6aafb),
	.w6(32'h3bb89fd5),
	.w7(32'hbbbd7319),
	.w8(32'hbba305ad),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54b466),
	.w1(32'h3bc4984b),
	.w2(32'h3bd02dc4),
	.w3(32'h3b599085),
	.w4(32'h3bb04906),
	.w5(32'h3b1e7d50),
	.w6(32'hba777030),
	.w7(32'h3b1082e2),
	.w8(32'h3bca4c0d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8723a1),
	.w1(32'h3b61bbc9),
	.w2(32'hb9ca6640),
	.w3(32'h3b886c00),
	.w4(32'h3c3bd261),
	.w5(32'h3bacbe6c),
	.w6(32'h3bac437e),
	.w7(32'h3b369ac3),
	.w8(32'h3c260bdd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d23bb0),
	.w1(32'hbb819b4d),
	.w2(32'hbb86b640),
	.w3(32'h3bfcdb65),
	.w4(32'hbaa4098a),
	.w5(32'hbbfd1b33),
	.w6(32'h3bcaf445),
	.w7(32'hbb104183),
	.w8(32'hbc06a3d2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab15dd5),
	.w1(32'hbb11b381),
	.w2(32'hbbad4fbe),
	.w3(32'hbade0a21),
	.w4(32'h3b4aac70),
	.w5(32'hbb0e7762),
	.w6(32'hbac1f300),
	.w7(32'hbb167d6a),
	.w8(32'h3bbf1cac),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb049bcb),
	.w1(32'hbb45267e),
	.w2(32'h3b79869f),
	.w3(32'h3b4512bd),
	.w4(32'h3bb8ba2e),
	.w5(32'h3bda070a),
	.w6(32'h3bb62cdf),
	.w7(32'h3bc959b2),
	.w8(32'h3c05f6c1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a5b1c),
	.w1(32'h3b274629),
	.w2(32'h3c5efbae),
	.w3(32'h3b277942),
	.w4(32'hbb7a7cf9),
	.w5(32'h397c46e1),
	.w6(32'hbbb13496),
	.w7(32'h3b07d4b5),
	.w8(32'hbb2c545f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdeced),
	.w1(32'hbc12f739),
	.w2(32'hbaf645fb),
	.w3(32'h3b80d805),
	.w4(32'hbb155628),
	.w5(32'h3b7d3882),
	.w6(32'hbbe14036),
	.w7(32'hb90641b7),
	.w8(32'h3b1a57eb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b819592),
	.w1(32'hbb5be728),
	.w2(32'hbc2ca826),
	.w3(32'h39da8299),
	.w4(32'h3b882290),
	.w5(32'hbb0d0879),
	.w6(32'h3ad276fb),
	.w7(32'hbc3abcaf),
	.w8(32'hbc02afd9),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c7205),
	.w1(32'h3b2b01a0),
	.w2(32'h392507d1),
	.w3(32'h3b0f1c31),
	.w4(32'h3bebdcb3),
	.w5(32'h3b84832c),
	.w6(32'h3bf89301),
	.w7(32'hbb233233),
	.w8(32'hba7a39d6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb37fb),
	.w1(32'hba45c793),
	.w2(32'h3bd37868),
	.w3(32'h3a8eaa56),
	.w4(32'h3b228888),
	.w5(32'h3b74f30b),
	.w6(32'hbb1ec5ac),
	.w7(32'h3b967faa),
	.w8(32'h3bb8d967),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc44dc),
	.w1(32'hbc15ffba),
	.w2(32'hbb92eea8),
	.w3(32'hbb9329fb),
	.w4(32'hbb40c08b),
	.w5(32'hbba88399),
	.w6(32'hbb412cff),
	.w7(32'h39670982),
	.w8(32'hbb3d40b7),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2544f),
	.w1(32'hbbe9f708),
	.w2(32'hbbaf0c6f),
	.w3(32'hbb3c5a24),
	.w4(32'hbc0b0dc8),
	.w5(32'h3b1326b0),
	.w6(32'hbbfe99ba),
	.w7(32'hbbf94f4b),
	.w8(32'hbb4c6ace),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe91270),
	.w1(32'h391f2c9e),
	.w2(32'h3b07c635),
	.w3(32'hbbd9b473),
	.w4(32'hba85472d),
	.w5(32'h3adccb37),
	.w6(32'hbba93840),
	.w7(32'h3b974fab),
	.w8(32'h3bc8f7e6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba3024),
	.w1(32'h3a647a91),
	.w2(32'hbb19e7e7),
	.w3(32'h3a45f384),
	.w4(32'hba5007ba),
	.w5(32'hbba43f5b),
	.w6(32'h3b636bbf),
	.w7(32'hbae28f24),
	.w8(32'hb7c827e0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba981380),
	.w1(32'h3c0b2e33),
	.w2(32'h3c93bbd2),
	.w3(32'hbac0fe5d),
	.w4(32'h3a31963b),
	.w5(32'h3be3d6ed),
	.w6(32'hbb295a7c),
	.w7(32'hba1ef0fc),
	.w8(32'hbbcf48fd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdefb99),
	.w1(32'h3b5ecbd0),
	.w2(32'h3bc54e62),
	.w3(32'h3cbc2939),
	.w4(32'h3b97d40d),
	.w5(32'h3c2303bb),
	.w6(32'h3bcd0319),
	.w7(32'h3ba790ec),
	.w8(32'h33ee0280),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01f4f8),
	.w1(32'h3bf3c3e9),
	.w2(32'hbbf06919),
	.w3(32'h3ba38cb7),
	.w4(32'hb9846708),
	.w5(32'h3c916616),
	.w6(32'h3b376e36),
	.w7(32'hbc2e6259),
	.w8(32'hbb813f53),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12be83),
	.w1(32'h3bc236e6),
	.w2(32'h3b09e768),
	.w3(32'h3bcb97dc),
	.w4(32'hbb7d31a8),
	.w5(32'hb794a530),
	.w6(32'h3c028998),
	.w7(32'hbb8e5e79),
	.w8(32'hbbfbfff2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3be5e3),
	.w1(32'hba0b94e8),
	.w2(32'h3b6b789e),
	.w3(32'h3c96155b),
	.w4(32'hbb60910b),
	.w5(32'hbb28d4cc),
	.w6(32'h39cf66d8),
	.w7(32'h3b76c47b),
	.w8(32'hbb406412),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7341db),
	.w1(32'h381d6cbc),
	.w2(32'h3b5202da),
	.w3(32'h3bbeb37e),
	.w4(32'h3baa6804),
	.w5(32'h3b909c06),
	.w6(32'h3b63437c),
	.w7(32'h3a8f74d5),
	.w8(32'h3b9a08d9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c0ee4),
	.w1(32'h382e56c7),
	.w2(32'hba88d7d0),
	.w3(32'h3aa57bc5),
	.w4(32'h3b7c7822),
	.w5(32'h3bd0a612),
	.w6(32'hbb360bfc),
	.w7(32'hba569ca0),
	.w8(32'h3ab3873f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48a337),
	.w1(32'h3b488bce),
	.w2(32'h3b7dfcd9),
	.w3(32'hbbe33902),
	.w4(32'h3b459961),
	.w5(32'hbb819e95),
	.w6(32'h3ab0c4af),
	.w7(32'hbb8a2100),
	.w8(32'hbb16093e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4faa7e),
	.w1(32'h3a4c5a65),
	.w2(32'h3ac661d6),
	.w3(32'h3b08839d),
	.w4(32'h3948f3d7),
	.w5(32'hba5bbe34),
	.w6(32'h3bec73a6),
	.w7(32'hb936205c),
	.w8(32'h3aa66927),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bf076),
	.w1(32'h3bba0b87),
	.w2(32'hbae430d2),
	.w3(32'h3ad4426f),
	.w4(32'h398589e7),
	.w5(32'h3b48e383),
	.w6(32'h3bb2ef1d),
	.w7(32'h3aaa205e),
	.w8(32'h3aaa806b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6cbc02),
	.w1(32'hba8267ad),
	.w2(32'hba548641),
	.w3(32'h3b84264c),
	.w4(32'hbb137ec4),
	.w5(32'hbbc271f7),
	.w6(32'h3bc8e520),
	.w7(32'h3b0f7ff4),
	.w8(32'h3a91ee0e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad258b4),
	.w1(32'hbb2e6def),
	.w2(32'h3a255f67),
	.w3(32'hbb32c070),
	.w4(32'hbb17ac04),
	.w5(32'hbaa73638),
	.w6(32'h3a8a3444),
	.w7(32'hbb7059ea),
	.w8(32'h3acf9801),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74f209),
	.w1(32'hbb4f4d96),
	.w2(32'h3a1c6d3f),
	.w3(32'hbac2bf54),
	.w4(32'hbb3efc09),
	.w5(32'h3b869336),
	.w6(32'hba97f9eb),
	.w7(32'hbb21c3a4),
	.w8(32'hbbaf74ed),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad071c),
	.w1(32'hbad8b1c6),
	.w2(32'hba33f46b),
	.w3(32'hbaeffda7),
	.w4(32'h3aee38a3),
	.w5(32'hb9b22da1),
	.w6(32'hbb658da6),
	.w7(32'hb9dc95e4),
	.w8(32'h3a81dcda),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe450f),
	.w1(32'h3b663b0a),
	.w2(32'h3c3dfc29),
	.w3(32'hbb8af0ff),
	.w4(32'h3b8d0bf6),
	.w5(32'h3b1595c7),
	.w6(32'h3a069dfb),
	.w7(32'h3b639754),
	.w8(32'h3a2b77e4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf79235),
	.w1(32'hba50a6ce),
	.w2(32'hbbfc45e0),
	.w3(32'h3ba4d447),
	.w4(32'h3bbc5ffa),
	.w5(32'hbb6ebd4c),
	.w6(32'h3ba20aab),
	.w7(32'hbb7e7d9c),
	.w8(32'hbb870e95),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae8228),
	.w1(32'hbb13ec46),
	.w2(32'h3ad1d792),
	.w3(32'hbb09ac83),
	.w4(32'hbc06ff8c),
	.w5(32'hbbea4dbe),
	.w6(32'hbaee836f),
	.w7(32'hbbccbbe8),
	.w8(32'hbba9f5c5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5bdf4),
	.w1(32'h3b0f69c5),
	.w2(32'hbb0a5037),
	.w3(32'hb9e4cd6b),
	.w4(32'hbc040c6d),
	.w5(32'h3b15b208),
	.w6(32'hbc203485),
	.w7(32'hb94e912f),
	.w8(32'hbb9d8eee),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826f0f),
	.w1(32'h3ae50016),
	.w2(32'hbb84c15a),
	.w3(32'hbaed4f4c),
	.w4(32'h3b233bdf),
	.w5(32'h395c4718),
	.w6(32'hbab1a0f2),
	.w7(32'hbb235554),
	.w8(32'hbaab79f7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb363e8b),
	.w1(32'hbb269b9b),
	.w2(32'hbb325e7a),
	.w3(32'hbb1fa7fe),
	.w4(32'hbc09ac75),
	.w5(32'hbbae62a9),
	.w6(32'h3b245eeb),
	.w7(32'hbb18ddfa),
	.w8(32'hbc317678),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa670c),
	.w1(32'h3c304d1f),
	.w2(32'h3b5e2506),
	.w3(32'hbb3d942f),
	.w4(32'h3c487879),
	.w5(32'h3af210dc),
	.w6(32'hbbf022dc),
	.w7(32'h3bec5229),
	.w8(32'h3aa561d5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f1bb8),
	.w1(32'hb9f42ee5),
	.w2(32'h3af260aa),
	.w3(32'h3b969fa5),
	.w4(32'h3b9273bd),
	.w5(32'h3c02685b),
	.w6(32'h3a67713d),
	.w7(32'h3bb82fd5),
	.w8(32'h3c1e8857),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ba5d4),
	.w1(32'hbb79834d),
	.w2(32'hb9fd90c0),
	.w3(32'hbafe9642),
	.w4(32'h3b1cb995),
	.w5(32'hbb2953a7),
	.w6(32'h3a8c83b0),
	.w7(32'hbacbc980),
	.w8(32'h3a1c0f77),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44331b),
	.w1(32'h3c1d9823),
	.w2(32'hbb8c10f6),
	.w3(32'hbaad89f1),
	.w4(32'h3b3ab181),
	.w5(32'h3c29f588),
	.w6(32'hbb1a388e),
	.w7(32'hbae1ff98),
	.w8(32'hbb3f7df6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc72fd),
	.w1(32'hbad158cb),
	.w2(32'h3991055c),
	.w3(32'h3ad06e05),
	.w4(32'hbbc228db),
	.w5(32'hbb7e9c75),
	.w6(32'h3be772db),
	.w7(32'hbb86dca5),
	.w8(32'hbb6f7547),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb460634),
	.w1(32'hbadfe7d5),
	.w2(32'h3b7a56fa),
	.w3(32'hbb961145),
	.w4(32'h3b74ac1e),
	.w5(32'h3b4caf48),
	.w6(32'h3b5b0c20),
	.w7(32'h3b180605),
	.w8(32'h3aa49d9d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd578ec),
	.w1(32'h3ad2fb52),
	.w2(32'hbaabfdd0),
	.w3(32'h3ba6f974),
	.w4(32'h3b945b9f),
	.w5(32'hbb954d14),
	.w6(32'hba82589b),
	.w7(32'hbb04f737),
	.w8(32'h395e13ae),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8132dd),
	.w1(32'hbb6e5f2b),
	.w2(32'h3aac3729),
	.w3(32'hbb6d0678),
	.w4(32'hba7d8988),
	.w5(32'h3a938dc1),
	.w6(32'hba1674e1),
	.w7(32'h3a603a1b),
	.w8(32'h3b492865),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb30cab),
	.w1(32'h3b010633),
	.w2(32'hbaccb79b),
	.w3(32'hbb17ef5f),
	.w4(32'hbb9c9ba6),
	.w5(32'hbc5b87b2),
	.w6(32'hbaddce4b),
	.w7(32'hbb2e23f4),
	.w8(32'hbc1aa8e1),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ffae2),
	.w1(32'hbb26795e),
	.w2(32'h3bb5ded2),
	.w3(32'hbac85199),
	.w4(32'h39c91918),
	.w5(32'h3bdac775),
	.w6(32'hbbcdb15c),
	.w7(32'hbab83af6),
	.w8(32'h3bb81e6f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d099f),
	.w1(32'hb9f10c15),
	.w2(32'h3b0b356c),
	.w3(32'hbbbb1c0b),
	.w4(32'h3bee7bf2),
	.w5(32'h3adf723e),
	.w6(32'h3b37f4bd),
	.w7(32'h3b825aad),
	.w8(32'h3bb8ec43),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cb949),
	.w1(32'h3b00c4b6),
	.w2(32'h3b113648),
	.w3(32'hbba22743),
	.w4(32'hbbda350c),
	.w5(32'h3b7194e0),
	.w6(32'h3adbe371),
	.w7(32'hbbe0081f),
	.w8(32'hbbf50ef1),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c2903),
	.w1(32'h3b3b4ec1),
	.w2(32'h3bc4f341),
	.w3(32'h3c0135d1),
	.w4(32'hba44f8ca),
	.w5(32'hb99a3290),
	.w6(32'hbb5c0d67),
	.w7(32'hbb38c090),
	.w8(32'h3b01d4df),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f0d19),
	.w1(32'hbb93552f),
	.w2(32'hbb4fa2b3),
	.w3(32'hbab2e3c9),
	.w4(32'hbb862686),
	.w5(32'hbc04b33b),
	.w6(32'hbb217d88),
	.w7(32'hbb1042ef),
	.w8(32'hbb027c9d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a3887),
	.w1(32'hba554922),
	.w2(32'hbb93bfe9),
	.w3(32'h3b752804),
	.w4(32'h3b3efa44),
	.w5(32'hbb80d441),
	.w6(32'h3b8dc9b9),
	.w7(32'hbb5d99aa),
	.w8(32'hbc10a898),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bff032),
	.w1(32'h3b0d52ed),
	.w2(32'hbb27227f),
	.w3(32'h399ca195),
	.w4(32'h39c05d45),
	.w5(32'h3b0dd767),
	.w6(32'hbb289e19),
	.w7(32'h3b4c1d29),
	.w8(32'h3a0bf425),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32697c),
	.w1(32'h3b17a476),
	.w2(32'h3b7c16cb),
	.w3(32'h3b4f4391),
	.w4(32'hbb416d89),
	.w5(32'hb93aed7e),
	.w6(32'hbab2bf0c),
	.w7(32'h3a24ad1a),
	.w8(32'hbb45bb63),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b454d7b),
	.w1(32'hbb11d938),
	.w2(32'hbacdde58),
	.w3(32'h3aeaec5c),
	.w4(32'hbbd0116e),
	.w5(32'hb9b4d6ee),
	.w6(32'h38b23b16),
	.w7(32'hbbb3b675),
	.w8(32'hbbb76c91),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00697a),
	.w1(32'hba09da3c),
	.w2(32'h39955cd1),
	.w3(32'h3a3a1e9e),
	.w4(32'h3a458280),
	.w5(32'h39da9cfa),
	.w6(32'hbba6f57c),
	.w7(32'h3bb015b7),
	.w8(32'h3b95def0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa871fc),
	.w1(32'hbb501b8c),
	.w2(32'hbb8b3539),
	.w3(32'hbb278165),
	.w4(32'hbb0d92d4),
	.w5(32'hbba2d77b),
	.w6(32'hbb29fa29),
	.w7(32'hbb6bcad0),
	.w8(32'hbb84d072),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7e2f7),
	.w1(32'hbb0e42cb),
	.w2(32'hbb91a52e),
	.w3(32'hb901e1c1),
	.w4(32'h3b085e47),
	.w5(32'h3c7c7edd),
	.w6(32'hba523130),
	.w7(32'h3b81d0e7),
	.w8(32'h3bead22e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7570c4),
	.w1(32'h3ac1b9c2),
	.w2(32'h3a4eee6d),
	.w3(32'h3b4b5fd2),
	.w4(32'h3b5e38f7),
	.w5(32'hbacfdb95),
	.w6(32'h3b9b935b),
	.w7(32'hbb81fb6f),
	.w8(32'h3abc556b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c7290),
	.w1(32'h3ab2484c),
	.w2(32'h3ac1c4e9),
	.w3(32'hb981d17d),
	.w4(32'h3b7cbbaf),
	.w5(32'h3bc9efb5),
	.w6(32'hbb2bbbb8),
	.w7(32'h3bd28891),
	.w8(32'h3bb2385f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c6a05),
	.w1(32'h3b38ea95),
	.w2(32'h3abb82aa),
	.w3(32'h3a800735),
	.w4(32'hba2d34a3),
	.w5(32'h38446a5f),
	.w6(32'h3ad5a934),
	.w7(32'hbb1d7be0),
	.w8(32'hbb6a66e8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ad93d),
	.w1(32'h39f89f52),
	.w2(32'h3aa9d4f4),
	.w3(32'h3bc12857),
	.w4(32'h3bc477c8),
	.w5(32'h3b6347b8),
	.w6(32'h3b00c06f),
	.w7(32'h3b48bec6),
	.w8(32'h3b8b8b13),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1962f),
	.w1(32'hbaf0f587),
	.w2(32'hbb168692),
	.w3(32'h3ba1ec12),
	.w4(32'hbbd27519),
	.w5(32'hbb68fb39),
	.w6(32'h3ba5bad3),
	.w7(32'h3ba146bb),
	.w8(32'hbbf45cbd),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba315584),
	.w1(32'hba05ef1e),
	.w2(32'h3bad55e5),
	.w3(32'hb95b78d2),
	.w4(32'hbaec3f84),
	.w5(32'h3bb6d168),
	.w6(32'hbb4416c6),
	.w7(32'hbaaffe92),
	.w8(32'hbb5b0a24),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8679c0),
	.w1(32'hbb965634),
	.w2(32'hbba09d2a),
	.w3(32'h3c31c319),
	.w4(32'hbbe07fa3),
	.w5(32'hbbb2a7a4),
	.w6(32'h3b771192),
	.w7(32'hbba8bbd5),
	.w8(32'hbb925e9f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea2568),
	.w1(32'h3af04bc6),
	.w2(32'h3bb28ce8),
	.w3(32'hbb9a78ed),
	.w4(32'h3a1aab25),
	.w5(32'h3a20098f),
	.w6(32'h39cb04b6),
	.w7(32'h3b717452),
	.w8(32'hbb511362),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90dd1f),
	.w1(32'hbb1b56f7),
	.w2(32'hbb424b5b),
	.w3(32'hbaa21304),
	.w4(32'hbb62a20f),
	.w5(32'hbabf66ba),
	.w6(32'hbada2fdf),
	.w7(32'h3b414cac),
	.w8(32'h3ba42462),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a8955),
	.w1(32'h39ee565a),
	.w2(32'hba88b7d5),
	.w3(32'h3b39e10e),
	.w4(32'hbb521fd9),
	.w5(32'hbba81959),
	.w6(32'hbacc545c),
	.w7(32'hbb822cb7),
	.w8(32'hbabf5bca),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5ddfc),
	.w1(32'h3a28141c),
	.w2(32'h39858897),
	.w3(32'h3a3f0d5e),
	.w4(32'hbb26dde1),
	.w5(32'h3bb639b9),
	.w6(32'hbba91fef),
	.w7(32'h3aaab07b),
	.w8(32'h3aa3f909),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb977811),
	.w1(32'hba722d15),
	.w2(32'h38916633),
	.w3(32'h3aa96ba0),
	.w4(32'hbb093cec),
	.w5(32'h3b87b0f6),
	.w6(32'h3a2ebb63),
	.w7(32'hb8ee4cfe),
	.w8(32'hb9bf7fe2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7b14c),
	.w1(32'hbb7104e3),
	.w2(32'hba494ad9),
	.w3(32'h3a189645),
	.w4(32'h3b85aa62),
	.w5(32'h3b8312e0),
	.w6(32'h381b8cfa),
	.w7(32'h3a732897),
	.w8(32'h3bf5c8d2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf21948),
	.w1(32'hba8b5abf),
	.w2(32'h3bc6300c),
	.w3(32'hb9d0983e),
	.w4(32'hbb4db10f),
	.w5(32'hbbc8772c),
	.w6(32'h3a94b47d),
	.w7(32'h3b041fbd),
	.w8(32'h3a575167),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f39e4),
	.w1(32'hbb6d8f20),
	.w2(32'hbb26d187),
	.w3(32'h3b21749c),
	.w4(32'hbbadc1f8),
	.w5(32'hbc2419eb),
	.w6(32'h3bcaf7ee),
	.w7(32'hba9a9f41),
	.w8(32'hbb6ba430),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b023d88),
	.w1(32'h3b15ea11),
	.w2(32'h3b18e434),
	.w3(32'hbb6af425),
	.w4(32'hbafe4fb0),
	.w5(32'hbb30f5c0),
	.w6(32'hbbc97fc9),
	.w7(32'hbb4b9f27),
	.w8(32'hba9fb951),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b439c64),
	.w1(32'h3b34c376),
	.w2(32'h3b97c10c),
	.w3(32'h3a3fe7da),
	.w4(32'h3a6697fe),
	.w5(32'h3c274879),
	.w6(32'h3aac5df4),
	.w7(32'h3a89bc16),
	.w8(32'h3bad5e1f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c89cd),
	.w1(32'hbb729a37),
	.w2(32'h3a1e6c24),
	.w3(32'h3c23c856),
	.w4(32'hbae39365),
	.w5(32'hbacb79b7),
	.w6(32'h3bee7dcb),
	.w7(32'hbb977c08),
	.w8(32'hba94f5c1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e39b3),
	.w1(32'h3ae9d552),
	.w2(32'hba82eabe),
	.w3(32'hbb452e83),
	.w4(32'h3a028e3b),
	.w5(32'h3c089e92),
	.w6(32'hbb878bbb),
	.w7(32'hbb8908b1),
	.w8(32'hbb42881b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a15687),
	.w1(32'h3aa5bd7b),
	.w2(32'h3a635180),
	.w3(32'h3aa65557),
	.w4(32'h3adca243),
	.w5(32'h3bb7f066),
	.w6(32'h3b04f147),
	.w7(32'hbbcd1328),
	.w8(32'hbb89cc7f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5160c),
	.w1(32'hbc4d624b),
	.w2(32'h3b4cef56),
	.w3(32'hbb2b3668),
	.w4(32'hba0cfd70),
	.w5(32'hbae2078f),
	.w6(32'hba9aaf5e),
	.w7(32'hbac302d6),
	.w8(32'h3bea2939),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae8576),
	.w1(32'h3b15e71a),
	.w2(32'hb8fd9dc3),
	.w3(32'hbbd4c033),
	.w4(32'h3a7be5d7),
	.w5(32'hb93a129e),
	.w6(32'hbb826bc7),
	.w7(32'hbbb65a79),
	.w8(32'hb7809c19),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65d783),
	.w1(32'hbbb9d2be),
	.w2(32'hbabf122e),
	.w3(32'h3b17bba7),
	.w4(32'hbb55d68b),
	.w5(32'hbb877b61),
	.w6(32'hbb21d3cc),
	.w7(32'hbb8f0319),
	.w8(32'hbaf3e4e5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe9276),
	.w1(32'hba34179a),
	.w2(32'hba079459),
	.w3(32'hbabf75f6),
	.w4(32'hba9ccde1),
	.w5(32'h3981971c),
	.w6(32'h3a498ba9),
	.w7(32'hbb122a1d),
	.w8(32'h399b5f65),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05a3a9),
	.w1(32'hbb28f63b),
	.w2(32'hbae36277),
	.w3(32'hbbb99710),
	.w4(32'h3b96a074),
	.w5(32'hbb87e9f6),
	.w6(32'hbadabcb6),
	.w7(32'h39e32894),
	.w8(32'hbb090b01),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bc675),
	.w1(32'h396e2c8b),
	.w2(32'hbb0a93e0),
	.w3(32'hbb758f7a),
	.w4(32'hbb723fd5),
	.w5(32'hb9af27de),
	.w6(32'hbbcda334),
	.w7(32'h3b47fa17),
	.w8(32'hb8727489),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ccabe),
	.w1(32'h3c846f8a),
	.w2(32'h3b48ae2a),
	.w3(32'hbaa8c6a0),
	.w4(32'h3c231b48),
	.w5(32'h3c974190),
	.w6(32'hbb2ad244),
	.w7(32'h3bf7b0fd),
	.w8(32'h3c4e9fcd),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca518),
	.w1(32'h3b06cac6),
	.w2(32'h3b0d37a8),
	.w3(32'h3c627eb2),
	.w4(32'hbb060788),
	.w5(32'h3b55f8c0),
	.w6(32'h3c335cfa),
	.w7(32'hbad84edb),
	.w8(32'hba449bfa),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d0e9d),
	.w1(32'hbba020ab),
	.w2(32'h3bb1657b),
	.w3(32'h3a6e4933),
	.w4(32'hbb810636),
	.w5(32'hbac3356e),
	.w6(32'h3b9d2d5e),
	.w7(32'hba4fd181),
	.w8(32'hba15a226),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0cac0),
	.w1(32'h3b864c65),
	.w2(32'h3bf0bc5c),
	.w3(32'h3aa15121),
	.w4(32'hbb09b802),
	.w5(32'h39e084ff),
	.w6(32'h3a1641f8),
	.w7(32'h3ae38921),
	.w8(32'hbb13d6bc),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fd922),
	.w1(32'h3bb7cc27),
	.w2(32'h3b1fc260),
	.w3(32'h3bcfa739),
	.w4(32'h3bc1ee10),
	.w5(32'hbbedcf43),
	.w6(32'hb9c346ed),
	.w7(32'h3b72055d),
	.w8(32'h3987d2c4),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b780d28),
	.w1(32'hbb0b7464),
	.w2(32'hbbb51fe3),
	.w3(32'hbb2ea011),
	.w4(32'hb93a6519),
	.w5(32'h3b252642),
	.w6(32'hba1247ab),
	.w7(32'hbb31659d),
	.w8(32'h3ba5bf0b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98527e),
	.w1(32'hb96f6f4d),
	.w2(32'h3b8865b4),
	.w3(32'hba1bcc96),
	.w4(32'hb8e0bc0b),
	.w5(32'hbb5f32fa),
	.w6(32'h3b92a4a7),
	.w7(32'h3992541c),
	.w8(32'hbae7a610),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08269a),
	.w1(32'hbb2495fb),
	.w2(32'hbb2a414b),
	.w3(32'hbaf4c03a),
	.w4(32'hba1313dd),
	.w5(32'hbbe30b85),
	.w6(32'hbb699820),
	.w7(32'h3b0c5002),
	.w8(32'hb81f37d9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac632ce),
	.w1(32'hbbbd276d),
	.w2(32'hbb536307),
	.w3(32'hbb751a61),
	.w4(32'hbbc2a3a0),
	.w5(32'h3b2c7885),
	.w6(32'hbb8f9ccf),
	.w7(32'hbaec149a),
	.w8(32'hbb56cab4),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb658f5),
	.w1(32'h3a138708),
	.w2(32'h3ac97f99),
	.w3(32'hbb69b35e),
	.w4(32'h3c0e56d7),
	.w5(32'h3bf371b8),
	.w6(32'hbb42c550),
	.w7(32'h3ba0186f),
	.w8(32'h3c49187b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56c9b9),
	.w1(32'h3b44fa79),
	.w2(32'h3b7a3519),
	.w3(32'hba7e2c73),
	.w4(32'h3b50a1fd),
	.w5(32'hbbd9d78e),
	.w6(32'h3b58705b),
	.w7(32'h3be5ef5f),
	.w8(32'h3a90857b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3889a),
	.w1(32'hbb20694a),
	.w2(32'h3b9c00b2),
	.w3(32'hba1c5611),
	.w4(32'hba0db77f),
	.w5(32'h3ade9471),
	.w6(32'hbaee7960),
	.w7(32'h3aaa625d),
	.w8(32'h3bbd1ab7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37b2d6),
	.w1(32'hb9d3b92c),
	.w2(32'hbb3a056c),
	.w3(32'hbaa8ac13),
	.w4(32'h3ba5f44a),
	.w5(32'h3a6f00b5),
	.w6(32'hbb8c39e9),
	.w7(32'h392cdff0),
	.w8(32'hbaab21b5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75b0af),
	.w1(32'h3b610e08),
	.w2(32'h3af7fa0e),
	.w3(32'hbb9d49c0),
	.w4(32'h3b73070c),
	.w5(32'h3cb8c8f5),
	.w6(32'h3a148199),
	.w7(32'h3b3b1a21),
	.w8(32'h3ad9aefb),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb371b39),
	.w1(32'h3c46a647),
	.w2(32'h3c027cdf),
	.w3(32'h3c11335f),
	.w4(32'h3b8c5723),
	.w5(32'h3c835345),
	.w6(32'h3c2b97bc),
	.w7(32'hbbc88ad5),
	.w8(32'hbc48334f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b718e96),
	.w1(32'h3b982025),
	.w2(32'h3bf5b7e6),
	.w3(32'h3cd2e725),
	.w4(32'h3abf4ee6),
	.w5(32'h3c06ec5b),
	.w6(32'h3babbd45),
	.w7(32'hb9bd5304),
	.w8(32'h3ab5a9f2),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f86dc),
	.w1(32'h3af1e25b),
	.w2(32'h3aa46750),
	.w3(32'h3be15b3f),
	.w4(32'h3b6e2807),
	.w5(32'h3b385b48),
	.w6(32'hbab4b297),
	.w7(32'h3a8f732e),
	.w8(32'h3ac85b37),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7001ad),
	.w1(32'hb9baf2e7),
	.w2(32'hbaad4905),
	.w3(32'hbaf50593),
	.w4(32'hba0a90be),
	.w5(32'hbb6d2adb),
	.w6(32'hbb8213ee),
	.w7(32'hbabb2995),
	.w8(32'h3accf2be),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d3e1d),
	.w1(32'h3b84b736),
	.w2(32'h3b8f8271),
	.w3(32'hbb339063),
	.w4(32'h3b8fe519),
	.w5(32'h3b0cdb81),
	.w6(32'h3a4cf19c),
	.w7(32'h3b9a98f3),
	.w8(32'h3b2d0716),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a0415),
	.w1(32'h3a28a245),
	.w2(32'h3b6bdbc3),
	.w3(32'h3b34174e),
	.w4(32'h3ac74fea),
	.w5(32'h3b8d0412),
	.w6(32'h3b419ebb),
	.w7(32'hbba64871),
	.w8(32'hba5acfcb),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54adbf),
	.w1(32'hbc0ab9dd),
	.w2(32'hbc0843e5),
	.w3(32'h3a83e8c8),
	.w4(32'hbb6d4214),
	.w5(32'hbbb15ee4),
	.w6(32'hbb14475e),
	.w7(32'hba9c7d79),
	.w8(32'h3b29b9f3),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc282b32),
	.w1(32'h3bd05995),
	.w2(32'h3c1b2a0a),
	.w3(32'hbbcccf98),
	.w4(32'h3a718728),
	.w5(32'h3b9031bb),
	.w6(32'hb9844eb0),
	.w7(32'h3bd32ef7),
	.w8(32'h3b0f4233),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b448801),
	.w1(32'hbb8b0a29),
	.w2(32'hbb918e88),
	.w3(32'h3bdbf24a),
	.w4(32'hba86fc90),
	.w5(32'hbb9f4dad),
	.w6(32'h3b15ee74),
	.w7(32'hbb74ec5e),
	.w8(32'hb78d0c23),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31ed72),
	.w1(32'hba683361),
	.w2(32'h3abfaba6),
	.w3(32'hba250872),
	.w4(32'h39b01dc5),
	.w5(32'h3b0389d4),
	.w6(32'h3b150d23),
	.w7(32'h3b1cd4d5),
	.w8(32'h3b3958dd),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58fb5d),
	.w1(32'hb9c8fbfd),
	.w2(32'h3a21f416),
	.w3(32'hbab46db7),
	.w4(32'h3a894b06),
	.w5(32'h3a97b7d2),
	.w6(32'hba46946b),
	.w7(32'h3a084473),
	.w8(32'h3acc494c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9578c59),
	.w1(32'h39deeac4),
	.w2(32'h38262614),
	.w3(32'hba14875c),
	.w4(32'hba1bd5e0),
	.w5(32'hbb03f901),
	.w6(32'hb99c3702),
	.w7(32'hb998c57e),
	.w8(32'h390c2ac2),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925b9a5),
	.w1(32'hba47951c),
	.w2(32'h3a434b7d),
	.w3(32'h387a876d),
	.w4(32'hb7f806ae),
	.w5(32'h3a027bd2),
	.w6(32'h3a7f9482),
	.w7(32'hb8049def),
	.w8(32'h391b03bb),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39d8d8),
	.w1(32'h3a077ce7),
	.w2(32'h3a163948),
	.w3(32'hba33cf20),
	.w4(32'h391f48b9),
	.w5(32'hb9f13f5a),
	.w6(32'hba3fc0da),
	.w7(32'hb937a681),
	.w8(32'hb91c974b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94cfbf4),
	.w1(32'h3a67f2e0),
	.w2(32'h3ab8dfae),
	.w3(32'h39919a64),
	.w4(32'h3a190613),
	.w5(32'h39363793),
	.w6(32'h39ddd948),
	.w7(32'h3a9f2f45),
	.w8(32'h3ab1ce9c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa22ae5),
	.w1(32'h39afaf83),
	.w2(32'hba392247),
	.w3(32'h39efdc94),
	.w4(32'h3a53c120),
	.w5(32'hb80cb6a5),
	.w6(32'h3a474ebf),
	.w7(32'h37ea977a),
	.w8(32'hba25aa37),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968d38c),
	.w1(32'h39d01cca),
	.w2(32'h3853898a),
	.w3(32'h3af16793),
	.w4(32'h3a601399),
	.w5(32'h39ddf4de),
	.w6(32'h3ab6155b),
	.w7(32'hb8a05864),
	.w8(32'hba76d07a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb0c2c),
	.w1(32'hba0b9be4),
	.w2(32'h38a8b543),
	.w3(32'h39ca7b6c),
	.w4(32'hb9952001),
	.w5(32'h3a8d07d5),
	.w6(32'hb99a2435),
	.w7(32'hb970f5a4),
	.w8(32'h3a06453d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39caac53),
	.w1(32'h3a945838),
	.w2(32'hb98070da),
	.w3(32'h3b6b13d4),
	.w4(32'h3aab3657),
	.w5(32'hba02aabb),
	.w6(32'h3b350337),
	.w7(32'hb92bf1c2),
	.w8(32'hbac634aa),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d8a17),
	.w1(32'hba0c8ff9),
	.w2(32'h3a2213ab),
	.w3(32'h3a06c515),
	.w4(32'h39482e77),
	.w5(32'h3a1143e5),
	.w6(32'h3a443f90),
	.w7(32'h3a1ef583),
	.w8(32'h3a4049a2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba423b51),
	.w1(32'h3b440bce),
	.w2(32'h3af4bfee),
	.w3(32'h3b1e3b86),
	.w4(32'h3ba7f583),
	.w5(32'h3b20820c),
	.w6(32'h3b2d8f4e),
	.w7(32'h3b8990bd),
	.w8(32'h3b4a0724),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19ccc4),
	.w1(32'h39c92b99),
	.w2(32'hb84398be),
	.w3(32'h391386a4),
	.w4(32'hb8df8728),
	.w5(32'hb96a06b9),
	.w6(32'h3a55a29b),
	.w7(32'h3926877d),
	.w8(32'h38b915e4),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933c961),
	.w1(32'h38f141d0),
	.w2(32'h39d3313a),
	.w3(32'h37b60c3b),
	.w4(32'h394af706),
	.w5(32'hb869c9ed),
	.w6(32'h38e1b568),
	.w7(32'h39b9d28d),
	.w8(32'h3a13710f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b193e97),
	.w1(32'h3a871275),
	.w2(32'h3acac717),
	.w3(32'h39231328),
	.w4(32'h3a8a1015),
	.w5(32'h3b15ca8b),
	.w6(32'h3b0aa618),
	.w7(32'h3b026ca4),
	.w8(32'h3b6c484a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373c41ba),
	.w1(32'hbaacff37),
	.w2(32'h39c9ca67),
	.w3(32'hba9911cb),
	.w4(32'hba130d4b),
	.w5(32'h3a93b3ac),
	.w6(32'h3abd7012),
	.w7(32'h3a0378f4),
	.w8(32'h3b3ee1ed),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac00f43),
	.w1(32'hba881d41),
	.w2(32'hba2f4088),
	.w3(32'h3aaba573),
	.w4(32'h3a28f4ab),
	.w5(32'h39a5a5df),
	.w6(32'h3b0c7f14),
	.w7(32'h3a44a9a2),
	.w8(32'hba4789e2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b605de1),
	.w1(32'h3b516447),
	.w2(32'h3c01ae26),
	.w3(32'h3b11f15b),
	.w4(32'h3b269d81),
	.w5(32'h3b9625d8),
	.w6(32'h3ae79249),
	.w7(32'h3b758418),
	.w8(32'h3b558de9),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cf3cc1),
	.w1(32'hba028e77),
	.w2(32'hba051171),
	.w3(32'hb98d851c),
	.w4(32'hb9709262),
	.w5(32'hbaaed76d),
	.w6(32'hb9c49f78),
	.w7(32'h38dd5b09),
	.w8(32'hba30383a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb889a5fe),
	.w1(32'h38ae5086),
	.w2(32'h3a089b3b),
	.w3(32'h3889269e),
	.w4(32'h3a7cde4b),
	.w5(32'h3a0013a2),
	.w6(32'h39bc96cd),
	.w7(32'h3a96b628),
	.w8(32'h3a338067),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c0896),
	.w1(32'h396f9fff),
	.w2(32'h3b9e9bdf),
	.w3(32'hbb9c8641),
	.w4(32'hba78fbc2),
	.w5(32'h3ba5b5ad),
	.w6(32'hbb91ae06),
	.w7(32'hb9d94fa1),
	.w8(32'h3b37f5ef),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e427ab),
	.w1(32'h3a626069),
	.w2(32'h3b949568),
	.w3(32'hbb4526cd),
	.w4(32'h3b848ad5),
	.w5(32'h3bba0934),
	.w6(32'hbab81f90),
	.w7(32'h3bbd9412),
	.w8(32'h3c06edf4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69effa),
	.w1(32'hba9a865b),
	.w2(32'h3b64060f),
	.w3(32'hbb45ace1),
	.w4(32'hba839ab3),
	.w5(32'h3b7db366),
	.w6(32'hbb4d9123),
	.w7(32'h3a889b0e),
	.w8(32'h3ba92b56),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a772e14),
	.w1(32'h39a0cd06),
	.w2(32'hbaa5c709),
	.w3(32'h3ac35fb9),
	.w4(32'h38a056df),
	.w5(32'hbac21a52),
	.w6(32'h3a9152a7),
	.w7(32'hbadc6336),
	.w8(32'hbb4dea37),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19b95c),
	.w1(32'hb8f3f51e),
	.w2(32'hbb0c38c0),
	.w3(32'h3b838162),
	.w4(32'h38443fdc),
	.w5(32'hbb016e51),
	.w6(32'h3b1200b1),
	.w7(32'hbb1887f6),
	.w8(32'hbb96b124),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4af1f),
	.w1(32'h39b6247f),
	.w2(32'h3a326ce8),
	.w3(32'h3a2cc492),
	.w4(32'hb9ebe658),
	.w5(32'hba251a67),
	.w6(32'h3a2a3c00),
	.w7(32'hba156b08),
	.w8(32'h396dc757),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998411f),
	.w1(32'hb9a74bdd),
	.w2(32'hb822cb33),
	.w3(32'h396183bd),
	.w4(32'hb870de49),
	.w5(32'hba99b4e9),
	.w6(32'h3932ae61),
	.w7(32'h39ce9564),
	.w8(32'h3893f85d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d233b9),
	.w1(32'h3ab282f8),
	.w2(32'h3abf07af),
	.w3(32'hb9f944ad),
	.w4(32'hba035e01),
	.w5(32'hbaa93b3e),
	.w6(32'h3a28c490),
	.w7(32'h39d98846),
	.w8(32'h3a064b42),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d4c72),
	.w1(32'hb8908472),
	.w2(32'hb9ceebbc),
	.w3(32'hba1b3589),
	.w4(32'h39ed54d5),
	.w5(32'hba076db7),
	.w6(32'hb9ad0776),
	.w7(32'h39d89f6e),
	.w8(32'hb93e318f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ae3e1),
	.w1(32'h39b0335e),
	.w2(32'hba812c73),
	.w3(32'hb98a0187),
	.w4(32'hba3c425c),
	.w5(32'hba71a653),
	.w6(32'hba9324e4),
	.w7(32'hb96e5a02),
	.w8(32'hba4507fd),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2da4a6),
	.w1(32'hba25500e),
	.w2(32'h39abd795),
	.w3(32'hbb18b15b),
	.w4(32'h391d388c),
	.w5(32'h3997ad7e),
	.w6(32'h39946f3b),
	.w7(32'h3a9e0343),
	.w8(32'h3af29d39),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902e633),
	.w1(32'hba2f43fd),
	.w2(32'h3915f5f9),
	.w3(32'h39bd481d),
	.w4(32'hb8964a42),
	.w5(32'hb9d5c0c2),
	.w6(32'h3a19ff67),
	.w7(32'hb8976f01),
	.w8(32'hb98225f7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39299080),
	.w1(32'h389cb279),
	.w2(32'hb7bc0074),
	.w3(32'h386b4868),
	.w4(32'h398284a5),
	.w5(32'h3a445020),
	.w6(32'hb96660be),
	.w7(32'hb9b1d578),
	.w8(32'h39dbea97),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf9f24),
	.w1(32'hbb34bc5f),
	.w2(32'h3ba7a724),
	.w3(32'hbb0c1f8e),
	.w4(32'h3a4272d2),
	.w5(32'h3b8a8f6f),
	.w6(32'hbb91a4d2),
	.w7(32'h3b688eaa),
	.w8(32'h3bdbac01),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a363e62),
	.w1(32'h3a3ed0ba),
	.w2(32'h392fd925),
	.w3(32'h3a86456a),
	.w4(32'h3999ff20),
	.w5(32'h399357ac),
	.w6(32'h3a93c329),
	.w7(32'h3a167d8a),
	.w8(32'h3b06655c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fb130),
	.w1(32'h399af673),
	.w2(32'h3a01356b),
	.w3(32'hba5be4fe),
	.w4(32'h3a4a424b),
	.w5(32'h3895b3f1),
	.w6(32'hb830fa8b),
	.w7(32'h3a5348dc),
	.w8(32'h3a7179c4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953ac64),
	.w1(32'hb9897947),
	.w2(32'h3b07b1cd),
	.w3(32'h39523f92),
	.w4(32'h39d14aa0),
	.w5(32'h3ae2aecc),
	.w6(32'h38d30a21),
	.w7(32'h3ad6beca),
	.w8(32'h3af67a7b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c5ace3),
	.w1(32'h39c0d53e),
	.w2(32'h39bf7549),
	.w3(32'h38d1853f),
	.w4(32'h391e5db2),
	.w5(32'h391d2006),
	.w6(32'h38e08269),
	.w7(32'h3967a054),
	.w8(32'h399df689),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a189856),
	.w1(32'h37ca5ebd),
	.w2(32'h39bb8c10),
	.w3(32'h3930b341),
	.w4(32'h37499bd4),
	.w5(32'hb72c3b8e),
	.w6(32'h3a254e47),
	.w7(32'h39a1b386),
	.w8(32'h38f4d3af),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbd629),
	.w1(32'hb8154f0b),
	.w2(32'hb98844c2),
	.w3(32'h39c1c6ca),
	.w4(32'h38d7f4fe),
	.w5(32'h384f5415),
	.w6(32'hb8954810),
	.w7(32'h3a3f17af),
	.w8(32'h3a35ee4a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f19412),
	.w1(32'h37d6760e),
	.w2(32'hb9fef50c),
	.w3(32'h399d2e00),
	.w4(32'h3a1e0d42),
	.w5(32'h3a89493b),
	.w6(32'h3806d6e7),
	.w7(32'h39078733),
	.w8(32'h3943f8c1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a836a87),
	.w1(32'h3ab4c4e0),
	.w2(32'h3a53bee2),
	.w3(32'h3ae01aa5),
	.w4(32'h3a865cfa),
	.w5(32'hb9b83d26),
	.w6(32'h3afff091),
	.w7(32'h3a467c36),
	.w8(32'hba169657),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4efdd),
	.w1(32'h3a8740b1),
	.w2(32'h3b15dea0),
	.w3(32'h3b56dd30),
	.w4(32'h3b1d145b),
	.w5(32'h3b18440a),
	.w6(32'h3ab5da4c),
	.w7(32'h3af13193),
	.w8(32'h3a6342d9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba637337),
	.w1(32'h39a986c1),
	.w2(32'h3b31693c),
	.w3(32'hba4b44ee),
	.w4(32'h3ace2f80),
	.w5(32'h3a84cb48),
	.w6(32'hba39cba9),
	.w7(32'h3a821b8e),
	.w8(32'h3b089181),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5d743),
	.w1(32'h3a063dbb),
	.w2(32'h3b4c03b9),
	.w3(32'hba8b302b),
	.w4(32'h3af64a3f),
	.w5(32'h3b02254c),
	.w6(32'hba262dbc),
	.w7(32'h3b38afbc),
	.w8(32'h3b2a9b7e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cc5484),
	.w1(32'h39cda5da),
	.w2(32'h387f4672),
	.w3(32'hba243bf0),
	.w4(32'h39bb0fd7),
	.w5(32'h39822fd5),
	.w6(32'hba927498),
	.w7(32'h39c33a53),
	.w8(32'h3a1aa9a8),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3865110e),
	.w1(32'hb8956af8),
	.w2(32'hb97139da),
	.w3(32'h3866a8a0),
	.w4(32'hba19f404),
	.w5(32'hb9d1da9b),
	.w6(32'h3904d404),
	.w7(32'hb9816b70),
	.w8(32'hb9f02f89),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6199e),
	.w1(32'h3a083606),
	.w2(32'h3a86930a),
	.w3(32'hb9046e18),
	.w4(32'h398a6e1a),
	.w5(32'h3ac5a82d),
	.w6(32'hba25f837),
	.w7(32'h39b794f4),
	.w8(32'h3a4b4a34),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39326972),
	.w1(32'h39b584f7),
	.w2(32'hb9504101),
	.w3(32'h3a92365a),
	.w4(32'hb9a36c73),
	.w5(32'hb95f4d3e),
	.w6(32'h3a046cf7),
	.w7(32'hb9af1e93),
	.w8(32'hb8feadcf),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9469332),
	.w1(32'h39154395),
	.w2(32'h3afaec5b),
	.w3(32'hba06c338),
	.w4(32'h3a6bfa30),
	.w5(32'h3a6c5ea6),
	.w6(32'h3aa6a96e),
	.w7(32'h3b56a694),
	.w8(32'h3b597ab7),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0501ff),
	.w1(32'hb8dca217),
	.w2(32'hb98390e3),
	.w3(32'h39fe2cb8),
	.w4(32'hba0b8505),
	.w5(32'hba487182),
	.w6(32'h39bf2ee7),
	.w7(32'hba0f793a),
	.w8(32'hb932c747),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba386c),
	.w1(32'h38c55284),
	.w2(32'h382cca44),
	.w3(32'hba230acc),
	.w4(32'hb8c3aaff),
	.w5(32'h3747115a),
	.w6(32'hb9ff3b20),
	.w7(32'hb86b6156),
	.w8(32'hb99159dc),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d4b944),
	.w1(32'hba0308b6),
	.w2(32'h3a30effa),
	.w3(32'h394ef120),
	.w4(32'h380a1968),
	.w5(32'hb8ab625d),
	.w6(32'hb919a2fa),
	.w7(32'h3a0379e0),
	.w8(32'h3a91a5f9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ef5c60),
	.w1(32'hba0e72e9),
	.w2(32'hba050ad1),
	.w3(32'h3a2bdc02),
	.w4(32'hb9f43057),
	.w5(32'hbad5ce26),
	.w6(32'h38e1b481),
	.w7(32'hb8d955f5),
	.w8(32'hb9f3378f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a59e62),
	.w1(32'h394c4ff2),
	.w2(32'h3994aa25),
	.w3(32'hb9ac85a3),
	.w4(32'h391f79dd),
	.w5(32'h3a13f186),
	.w6(32'h39a20707),
	.w7(32'h3a5d936b),
	.w8(32'h3a65f061),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb975f93f),
	.w1(32'h394b6cf9),
	.w2(32'hb8f348a8),
	.w3(32'hba151ff7),
	.w4(32'hb8a34843),
	.w5(32'h39c9034e),
	.w6(32'hb9d507bd),
	.w7(32'hb853858a),
	.w8(32'h39931cf4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb331895),
	.w1(32'h3a93872a),
	.w2(32'h3ad8c011),
	.w3(32'h3b143698),
	.w4(32'h39a34385),
	.w5(32'h3a41bc84),
	.w6(32'h3b276017),
	.w7(32'h3aecdf2e),
	.w8(32'h3b45c0bf),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ad44c),
	.w1(32'hb958218f),
	.w2(32'h382d6967),
	.w3(32'hba1344b0),
	.w4(32'hb9bd6c54),
	.w5(32'h3a5431fc),
	.w6(32'hb9ba5ebf),
	.w7(32'hba8335d4),
	.w8(32'hb9fd2923),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7770bd),
	.w1(32'h3b2b4409),
	.w2(32'h3b6cef7e),
	.w3(32'hb79820d8),
	.w4(32'h3adc3a8f),
	.w5(32'h3b0697cd),
	.w6(32'h3b1ca4d4),
	.w7(32'h3ac98373),
	.w8(32'h3b2505c3),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule