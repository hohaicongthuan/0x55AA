module layer_10_featuremap_410(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb842aa2a),
	.w1(32'h3a04f964),
	.w2(32'h39a0169d),
	.w3(32'h3a7b98a2),
	.w4(32'h3a25aaef),
	.w5(32'h3a031de7),
	.w6(32'h3aae57ca),
	.w7(32'h3893017b),
	.w8(32'h3a50ded3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c533b),
	.w1(32'hbb1b761e),
	.w2(32'hbb4a7059),
	.w3(32'hba9ac8de),
	.w4(32'hbaf6806d),
	.w5(32'hba6fcf8c),
	.w6(32'hbb1482e3),
	.w7(32'hbb25fdf2),
	.w8(32'hbad90ae4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b23174),
	.w1(32'hba300402),
	.w2(32'hb9ea3d13),
	.w3(32'hb9359338),
	.w4(32'hba1b33ba),
	.w5(32'hba583bee),
	.w6(32'hba025a05),
	.w7(32'hba2a6cc0),
	.w8(32'h38241670),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945daae),
	.w1(32'h393ff4a9),
	.w2(32'h3a20f308),
	.w3(32'h3949789f),
	.w4(32'h3828f7a0),
	.w5(32'hb5b48f1d),
	.w6(32'h39b81355),
	.w7(32'hb98903d8),
	.w8(32'hba298030),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993be89),
	.w1(32'hba574905),
	.w2(32'hba17affa),
	.w3(32'hba348587),
	.w4(32'hba44993c),
	.w5(32'hba1bdc5b),
	.w6(32'hba54de8c),
	.w7(32'hbabd664e),
	.w8(32'hb9eded9f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b29fdc),
	.w1(32'h38ff49b1),
	.w2(32'hb9c553dc),
	.w3(32'hba24f4d7),
	.w4(32'hb808e12c),
	.w5(32'hb9194170),
	.w6(32'hb9f7c577),
	.w7(32'hb9b26e5b),
	.w8(32'hba12228b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81fa8d),
	.w1(32'h39d58886),
	.w2(32'h3ab62819),
	.w3(32'hbadc3126),
	.w4(32'h3a05d873),
	.w5(32'h3ab89687),
	.w6(32'hba870143),
	.w7(32'h3a64ba2f),
	.w8(32'h3aea64c7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d2581),
	.w1(32'h3bcc2570),
	.w2(32'h3bab9b11),
	.w3(32'h3b99cd32),
	.w4(32'h3ba24e6d),
	.w5(32'h3a11cc5b),
	.w6(32'h3bc80cda),
	.w7(32'h3bd0c435),
	.w8(32'h3ba6508d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b8a51),
	.w1(32'hb97a1d38),
	.w2(32'h39e75036),
	.w3(32'hba526610),
	.w4(32'hb9a81304),
	.w5(32'h3a0e9af8),
	.w6(32'hba4c9328),
	.w7(32'hba8328a0),
	.w8(32'h3a27f457),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f018a),
	.w1(32'hb971fef4),
	.w2(32'hbad478c6),
	.w3(32'h39e259de),
	.w4(32'hbada73ee),
	.w5(32'hbaa55764),
	.w6(32'h3b0e4009),
	.w7(32'hb90d2891),
	.w8(32'hb9ca66de),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d484d4),
	.w1(32'hb977f85e),
	.w2(32'h391cba66),
	.w3(32'hba891679),
	.w4(32'hb9bf38ca),
	.w5(32'h3a882396),
	.w6(32'hba32a297),
	.w7(32'hb7c03a92),
	.w8(32'h3a210d32),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9828c29),
	.w1(32'h3a8a94eb),
	.w2(32'h3b333103),
	.w3(32'hba523ece),
	.w4(32'h3a2ebdde),
	.w5(32'h3b3ba656),
	.w6(32'hb9fb56d3),
	.w7(32'h3a77a44a),
	.w8(32'h3b36a06f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c52bc),
	.w1(32'hba85cb61),
	.w2(32'h39807c58),
	.w3(32'hb7dd0b0c),
	.w4(32'hba8201e0),
	.w5(32'h3a413bc8),
	.w6(32'hbad580ca),
	.w7(32'hba3c9c5f),
	.w8(32'h3a264203),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c407c),
	.w1(32'h395e9ffb),
	.w2(32'h3a29d642),
	.w3(32'h39d02453),
	.w4(32'h3a42dfd1),
	.w5(32'h3a064f6e),
	.w6(32'h3a679860),
	.w7(32'h3a719981),
	.w8(32'h3aa3109f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba616b84),
	.w1(32'hbab70aba),
	.w2(32'hb9fd603f),
	.w3(32'hbac37c15),
	.w4(32'hbafb099a),
	.w5(32'hb74abc59),
	.w6(32'hb7cae7fa),
	.w7(32'hba465b2a),
	.w8(32'h38bc9774),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c58602),
	.w1(32'hbaeb3fc2),
	.w2(32'hba98c049),
	.w3(32'h3932d92c),
	.w4(32'hbac3490e),
	.w5(32'hb9992525),
	.w6(32'h3b4b0a73),
	.w7(32'h3b0a2e6a),
	.w8(32'h3adac1b6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08184c),
	.w1(32'hb9f29129),
	.w2(32'hb63b0e36),
	.w3(32'hb86349ae),
	.w4(32'h3846d5e1),
	.w5(32'hb901dad6),
	.w6(32'h3a0fa8af),
	.w7(32'h3a1de391),
	.w8(32'h37b5a405),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baecd28),
	.w1(32'h3c372e18),
	.w2(32'h3c3657c0),
	.w3(32'h3bc9ca92),
	.w4(32'h3c253110),
	.w5(32'h3bf3b3ac),
	.w6(32'h3c3cb0ce),
	.w7(32'h3c3fd5b2),
	.w8(32'h3c5857c8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7f0af),
	.w1(32'h3b496aba),
	.w2(32'h3b34a1cc),
	.w3(32'h3b074560),
	.w4(32'h3b66ce50),
	.w5(32'h3b299c98),
	.w6(32'h3b7a62a4),
	.w7(32'h3b80b720),
	.w8(32'h3b385bcc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb963bc9f),
	.w1(32'hb886e795),
	.w2(32'h39c1df47),
	.w3(32'h3965134c),
	.w4(32'hba227ade),
	.w5(32'h3a32d9a1),
	.w6(32'hb8f43642),
	.w7(32'h38a1041f),
	.w8(32'hb9dd26bd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0e61d),
	.w1(32'h3a1d201b),
	.w2(32'h3896d1e6),
	.w3(32'hb854fed3),
	.w4(32'h39396d0d),
	.w5(32'h38f10aea),
	.w6(32'h3851bac3),
	.w7(32'hb9d80187),
	.w8(32'hb91208bd),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa7e2f),
	.w1(32'hba379d7a),
	.w2(32'hba18b6a1),
	.w3(32'hbab48da8),
	.w4(32'hba1978a0),
	.w5(32'hb9d5159f),
	.w6(32'hbaffcbc1),
	.w7(32'hba6a7f6b),
	.w8(32'hba910eb2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ecdbb),
	.w1(32'h3c2a8b9b),
	.w2(32'h3c4a346d),
	.w3(32'h3c0158fd),
	.w4(32'h3c1253ed),
	.w5(32'h3c02ff72),
	.w6(32'h3c8629b2),
	.w7(32'h3c7b5f44),
	.w8(32'h3c32b845),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a996545),
	.w1(32'hbaa7f0c1),
	.w2(32'hbb410890),
	.w3(32'h39dda9a6),
	.w4(32'hbb1de26e),
	.w5(32'hbb5f47ee),
	.w6(32'h3a841c47),
	.w7(32'hba35b727),
	.w8(32'hbaede33a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91be870),
	.w1(32'hbb35e724),
	.w2(32'hbb72397d),
	.w3(32'hba996b85),
	.w4(32'hbb4f1583),
	.w5(32'hbb19e741),
	.w6(32'hbb1e068d),
	.w7(32'hbb5904d3),
	.w8(32'hbafe0754),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7534d1),
	.w1(32'h39dc8c2b),
	.w2(32'h379e6ece),
	.w3(32'hba506669),
	.w4(32'h39cb23fd),
	.w5(32'hb94c7b78),
	.w6(32'h397e0e72),
	.w7(32'h3a0d93f2),
	.w8(32'h3983ab8d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2649f3),
	.w1(32'h39b8fe30),
	.w2(32'hb8fcc9dc),
	.w3(32'h3a07b4ff),
	.w4(32'hb9edd5b9),
	.w5(32'hb98e0cb7),
	.w6(32'h39e74321),
	.w7(32'hb84f77de),
	.w8(32'h39d4b316),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaddacf),
	.w1(32'hbb04d56f),
	.w2(32'hba6fc6e7),
	.w3(32'hbb2c22ce),
	.w4(32'hbb3425a2),
	.w5(32'hba0c9eff),
	.w6(32'hbb89a9fd),
	.w7(32'hbb6c543e),
	.w8(32'hbae3af61),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3885512a),
	.w1(32'hba1c4c49),
	.w2(32'hb9710f89),
	.w3(32'hba11cc57),
	.w4(32'hb99e1d1a),
	.w5(32'hb9c5644e),
	.w6(32'hba24db7e),
	.w7(32'hb9037fdb),
	.w8(32'hba3facb4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99780c5),
	.w1(32'hbb18ee62),
	.w2(32'hbb15f8d1),
	.w3(32'hbaa80c47),
	.w4(32'hbb63f9bb),
	.w5(32'hbae18450),
	.w6(32'hbb299665),
	.w7(32'hbb7e99c8),
	.w8(32'hbb3547e7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc8afb),
	.w1(32'h38535996),
	.w2(32'h399bc794),
	.w3(32'h3a08f873),
	.w4(32'hba0a71f2),
	.w5(32'hb9b6bfc0),
	.w6(32'h393f9c15),
	.w7(32'hb9a39cb5),
	.w8(32'hba041b8f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3860c920),
	.w1(32'hba027e85),
	.w2(32'hb9ed40d1),
	.w3(32'hb885900a),
	.w4(32'hb96030f2),
	.w5(32'h38a7b919),
	.w6(32'h399ad1d8),
	.w7(32'hb91710b0),
	.w8(32'h37c7ac26),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe7350),
	.w1(32'h39e51464),
	.w2(32'h39addef9),
	.w3(32'h3a3c64e8),
	.w4(32'h39d8e99c),
	.w5(32'hba2035f4),
	.w6(32'h3ab1bb3a),
	.w7(32'h39d4b146),
	.w8(32'h3a2c7ec6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89d9ff),
	.w1(32'hb9c17d08),
	.w2(32'hba98219c),
	.w3(32'h38d366c5),
	.w4(32'hba0731dd),
	.w5(32'hba3f48a1),
	.w6(32'hb892587c),
	.w7(32'hb8b6e4e1),
	.w8(32'hb9c47690),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39472026),
	.w1(32'h3a26745a),
	.w2(32'h3a1259cf),
	.w3(32'hb984578f),
	.w4(32'h3a2a429f),
	.w5(32'h38d715ca),
	.w6(32'hb9141991),
	.w7(32'h3a21f563),
	.w8(32'h3a683f38),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c718bf),
	.w1(32'h39ac3bc1),
	.w2(32'h3938a677),
	.w3(32'h3a3d13a6),
	.w4(32'h39d9ba5f),
	.w5(32'h38dc589f),
	.w6(32'h3b315b5e),
	.w7(32'h39423f0f),
	.w8(32'h3a0af894),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a25cd),
	.w1(32'hba0553b0),
	.w2(32'h3a8d9f66),
	.w3(32'hba4c226c),
	.w4(32'h39c0ba4b),
	.w5(32'h3afba78b),
	.w6(32'h3b593425),
	.w7(32'h3b4f650b),
	.w8(32'h3b5dcf9e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f949a),
	.w1(32'hbbd596e1),
	.w2(32'hbbe11239),
	.w3(32'hbb921000),
	.w4(32'hbc051410),
	.w5(32'hbb79e4ab),
	.w6(32'hbc091aa6),
	.w7(32'hbbedfb63),
	.w8(32'hbbc19fa1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4750e4),
	.w1(32'hbbb49570),
	.w2(32'hbb88e8c2),
	.w3(32'hbbeb8ada),
	.w4(32'hbbe1d1b1),
	.w5(32'hbacad8e8),
	.w6(32'hbc4b1c31),
	.w7(32'hbbe71019),
	.w8(32'hbb6edd81),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2c158),
	.w1(32'hba92e363),
	.w2(32'hba6d8733),
	.w3(32'hba62138d),
	.w4(32'hba7a3856),
	.w5(32'hba493fce),
	.w6(32'hbaaadd6e),
	.w7(32'hba4f2270),
	.w8(32'hba559b0e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376f6cc3),
	.w1(32'h39d76e1b),
	.w2(32'h3a068baa),
	.w3(32'hb953e242),
	.w4(32'hb78b3f83),
	.w5(32'h3a9153ed),
	.w6(32'hb9b50362),
	.w7(32'h3a39ce1e),
	.w8(32'h3a5aaed6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c71c70),
	.w1(32'hb933421b),
	.w2(32'hba1e457a),
	.w3(32'h3977219d),
	.w4(32'hb9bc8d99),
	.w5(32'h393c8868),
	.w6(32'h39124970),
	.w7(32'hb9a96a0f),
	.w8(32'hb9fd61e8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a424c58),
	.w1(32'h3a360457),
	.w2(32'hb953114a),
	.w3(32'h3a927c73),
	.w4(32'h3a2e5e4c),
	.w5(32'hb8532c5e),
	.w6(32'h3a20bfac),
	.w7(32'h374e65ea),
	.w8(32'hb92c1952),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83b08c),
	.w1(32'h3adaf569),
	.w2(32'h3a8093cb),
	.w3(32'h3b39fa01),
	.w4(32'h3b06a61e),
	.w5(32'h39d26b20),
	.w6(32'h3bafe6ff),
	.w7(32'h3b917025),
	.w8(32'h3ad6546b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac4f81),
	.w1(32'hba457c03),
	.w2(32'hbab48964),
	.w3(32'h399a5391),
	.w4(32'hbb1a32c1),
	.w5(32'hbac141ee),
	.w6(32'h386b8a80),
	.w7(32'hbb2067b5),
	.w8(32'hbac5a4ca),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28a386),
	.w1(32'hbaeb0117),
	.w2(32'hbb152a39),
	.w3(32'hb8c17ab6),
	.w4(32'hbb36af87),
	.w5(32'hbb07d0ab),
	.w6(32'h3a0e7307),
	.w7(32'hbaf2bd9f),
	.w8(32'hbabb89f4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982dc84),
	.w1(32'hb997a59a),
	.w2(32'h3a56fe05),
	.w3(32'h39d78eee),
	.w4(32'hb9cb2595),
	.w5(32'hb99bb1f6),
	.w6(32'h3b7adc93),
	.w7(32'h3ab86cd5),
	.w8(32'h3a55efd2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a7013),
	.w1(32'h3c153f5d),
	.w2(32'h3c52ad46),
	.w3(32'h3b77b099),
	.w4(32'h3c09f794),
	.w5(32'h3c0481f0),
	.w6(32'h3c293981),
	.w7(32'h3c218601),
	.w8(32'h3c371100),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a6486),
	.w1(32'hb975cca8),
	.w2(32'h38c2dd68),
	.w3(32'hba331d77),
	.w4(32'hb9b72915),
	.w5(32'hb97a0b29),
	.w6(32'hb911dc1e),
	.w7(32'hb9b032da),
	.w8(32'h390a39f4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e6d65),
	.w1(32'h3903c355),
	.w2(32'h3a5ed585),
	.w3(32'h3a3b537c),
	.w4(32'h3a20a11d),
	.w5(32'h3a565a86),
	.w6(32'h3ac301d4),
	.w7(32'h3a854a9a),
	.w8(32'h3ac7c2de),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f72e4),
	.w1(32'h38ba4b03),
	.w2(32'h397aecb2),
	.w3(32'h39fbb00a),
	.w4(32'h38cfc313),
	.w5(32'h38d0f8bf),
	.w6(32'hb8a5e4ba),
	.w7(32'hb9bab000),
	.w8(32'h39b00e2f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375d6bb6),
	.w1(32'h39495604),
	.w2(32'h3a5610d3),
	.w3(32'hb9341251),
	.w4(32'hb71b4dc3),
	.w5(32'h3a7190cd),
	.w6(32'h3715c407),
	.w7(32'hb7e69d76),
	.w8(32'h3a59e396),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19e6dd),
	.w1(32'h3ad879e0),
	.w2(32'h3af4b3df),
	.w3(32'h3a541bdc),
	.w4(32'h3a92e449),
	.w5(32'h39efd409),
	.w6(32'h3a8e1c5d),
	.w7(32'h3acdd0b1),
	.w8(32'h3ad9604a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6efc6e),
	.w1(32'h3bddf0db),
	.w2(32'h3bb8967d),
	.w3(32'h3bd14015),
	.w4(32'h3be8104e),
	.w5(32'h3b35127a),
	.w6(32'h3c08ce02),
	.w7(32'h3c042e9c),
	.w8(32'h3bbfac96),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381bc2fb),
	.w1(32'h3935df7f),
	.w2(32'h39d03b42),
	.w3(32'h39cd5d2b),
	.w4(32'h39aafa89),
	.w5(32'hb9e06528),
	.w6(32'h3a954e49),
	.w7(32'h3a82fdaa),
	.w8(32'h3a70e14d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0464ed),
	.w1(32'hba14c0b4),
	.w2(32'hba21f127),
	.w3(32'hba70f661),
	.w4(32'hb9c1b5c5),
	.w5(32'hb9baaf1a),
	.w6(32'hba1f589b),
	.w7(32'hb9949b46),
	.w8(32'h39d9ad6c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea577a),
	.w1(32'h39a9f491),
	.w2(32'h38a5553b),
	.w3(32'hb80f5cb0),
	.w4(32'h39c000b1),
	.w5(32'h3989ffeb),
	.w6(32'hb85cd3a5),
	.w7(32'h39716df2),
	.w8(32'h381bab9f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3896ff8c),
	.w1(32'h3820be45),
	.w2(32'hba7c0acb),
	.w3(32'hb9a2ab1e),
	.w4(32'h3953f1a8),
	.w5(32'hb9f8f66b),
	.w6(32'hb956c2cc),
	.w7(32'hba26ef8d),
	.w8(32'hba726460),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994a49c),
	.w1(32'hb9a3ffca),
	.w2(32'hba016307),
	.w3(32'hba665d8e),
	.w4(32'hba12780b),
	.w5(32'hba731e4a),
	.w6(32'hbabf2bbc),
	.w7(32'hba14cc7e),
	.w8(32'hba80cdc9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00d214),
	.w1(32'hb98171ef),
	.w2(32'h399103f9),
	.w3(32'hba863ab2),
	.w4(32'hb9c47512),
	.w5(32'h39c342c6),
	.w6(32'hba55c4e4),
	.w7(32'h39f426e7),
	.w8(32'h398b479a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e00fa),
	.w1(32'h3b1ff53d),
	.w2(32'h3b2af98c),
	.w3(32'h3b2fb9ee),
	.w4(32'h3b06d6bb),
	.w5(32'h3af94e3e),
	.w6(32'h3b71b373),
	.w7(32'h3b5bbe70),
	.w8(32'h3b7f37b2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e5087),
	.w1(32'h3b529ea9),
	.w2(32'h3b126c6d),
	.w3(32'h3b47fd2c),
	.w4(32'h3b587b45),
	.w5(32'h3b61b4d4),
	.w6(32'h3b9d1fb9),
	.w7(32'h3b6cb382),
	.w8(32'h3b3ab7ae),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c9b51e),
	.w1(32'hb9c4472f),
	.w2(32'hb9bd6b60),
	.w3(32'h38305e6d),
	.w4(32'hb9aa1144),
	.w5(32'hb8d5258e),
	.w6(32'h37e7e4f5),
	.w7(32'hb9b34d79),
	.w8(32'hb9c076b8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df06cf),
	.w1(32'h39c01975),
	.w2(32'h39bd659f),
	.w3(32'h39b6b179),
	.w4(32'h3a0a2d3d),
	.w5(32'h39f1753a),
	.w6(32'h39ec8bc5),
	.w7(32'h3985f250),
	.w8(32'h39e33950),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80aedfc),
	.w1(32'h3a55b330),
	.w2(32'h3a42da37),
	.w3(32'h390d0275),
	.w4(32'h39fdc4d3),
	.w5(32'h378561d6),
	.w6(32'h3970069a),
	.w7(32'h3a22e1bb),
	.w8(32'h3a19705c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cb35b),
	.w1(32'hb9945f74),
	.w2(32'hb956c212),
	.w3(32'h3a3c40bb),
	.w4(32'h37cfeefe),
	.w5(32'h3a1fc203),
	.w6(32'h3a3f43d0),
	.w7(32'hb92b28e7),
	.w8(32'h38a67478),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6037f),
	.w1(32'h3a92cee3),
	.w2(32'h3a834aae),
	.w3(32'hb9c583e2),
	.w4(32'h3a31636d),
	.w5(32'hb6cbde4b),
	.w6(32'h3aba5cea),
	.w7(32'h3b04dbe5),
	.w8(32'h398f6f7c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cb287),
	.w1(32'hbab2af6d),
	.w2(32'hbabb23d9),
	.w3(32'hba8b289f),
	.w4(32'hbac515a4),
	.w5(32'hb9f0e1aa),
	.w6(32'hb93a4823),
	.w7(32'hb9bde44e),
	.w8(32'h3af788bc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b666763),
	.w1(32'h3baadc66),
	.w2(32'h3b8e9c1d),
	.w3(32'h3b5d7ab5),
	.w4(32'h3b9376f5),
	.w5(32'h3b8cb9ec),
	.w6(32'h3c057fd3),
	.w7(32'h3bef40b2),
	.w8(32'h3bdcd885),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5ac08),
	.w1(32'hbc0b3b8e),
	.w2(32'hbb8c6eb2),
	.w3(32'hbb2d7a0d),
	.w4(32'hbbb5ec32),
	.w5(32'hba90a8a4),
	.w6(32'hbb811118),
	.w7(32'hbbef30fa),
	.w8(32'hbbccd17e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91fc2a),
	.w1(32'h3c3d1736),
	.w2(32'h3ba1f46b),
	.w3(32'h3b41a35a),
	.w4(32'h3bb67b2c),
	.w5(32'hbaac562b),
	.w6(32'h3aaeef13),
	.w7(32'h3b532f26),
	.w8(32'hb9a23a8e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b948495),
	.w1(32'h3b53a362),
	.w2(32'h3afe560d),
	.w3(32'hba314d77),
	.w4(32'hbb1b2507),
	.w5(32'h3b07ce7e),
	.w6(32'hbb0bc591),
	.w7(32'hbacb92f2),
	.w8(32'h397ce44e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90d512),
	.w1(32'h3b7eee07),
	.w2(32'h3a040053),
	.w3(32'h3ba62967),
	.w4(32'h3c1ee741),
	.w5(32'h3b1782ae),
	.w6(32'hbaccef3f),
	.w7(32'h3c17e519),
	.w8(32'h3b7dc0d2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f7fe2),
	.w1(32'h3a900e32),
	.w2(32'h3b937abf),
	.w3(32'h3a1229a6),
	.w4(32'h3b9482d4),
	.w5(32'h3bba2a9a),
	.w6(32'h3ae87ebe),
	.w7(32'h3b836fea),
	.w8(32'h3b800b25),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8a46f),
	.w1(32'h39ca8780),
	.w2(32'hbb006b8b),
	.w3(32'h39f9c0b8),
	.w4(32'hbad8627d),
	.w5(32'hbb822292),
	.w6(32'h3814d7c5),
	.w7(32'hba482797),
	.w8(32'hbb387096),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaafe8e),
	.w1(32'h3ba0602f),
	.w2(32'h3c5ca642),
	.w3(32'hbaa767b2),
	.w4(32'h3c4b4438),
	.w5(32'h3c6aa2c2),
	.w6(32'h3b17c5fa),
	.w7(32'h3c2b3450),
	.w8(32'h3bf45f91),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0303ca),
	.w1(32'h3bae0f47),
	.w2(32'h3c3e2c48),
	.w3(32'h3c888eab),
	.w4(32'h3c1a1519),
	.w5(32'h3c65af94),
	.w6(32'h3c329534),
	.w7(32'h3c2696ac),
	.w8(32'h3c8faf09),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c9c2d),
	.w1(32'h3b262aca),
	.w2(32'hba875f79),
	.w3(32'hbb95e45b),
	.w4(32'h3b351462),
	.w5(32'hbafe981e),
	.w6(32'hbbd98120),
	.w7(32'h3b352aa3),
	.w8(32'h3b97b8c4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9195b7),
	.w1(32'hbabc3e3d),
	.w2(32'h3a7c4b33),
	.w3(32'h3b7772c9),
	.w4(32'h39fa0606),
	.w5(32'h3b6f270e),
	.w6(32'h3b5fa8ab),
	.w7(32'h399ace12),
	.w8(32'h3bcacd03),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0024de),
	.w1(32'hbb09eca1),
	.w2(32'h38e9e459),
	.w3(32'h3b69bb47),
	.w4(32'hbb31a5f8),
	.w5(32'hb9cf1e0d),
	.w6(32'h3b2b61d9),
	.w7(32'hbafcd10f),
	.w8(32'h3a1d2ea0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80345d),
	.w1(32'hba986baa),
	.w2(32'h394d7f3d),
	.w3(32'hbb68b8f7),
	.w4(32'h3a4009ca),
	.w5(32'h3a5bccfb),
	.w6(32'hba24f1ba),
	.w7(32'h3a984d46),
	.w8(32'h3b14325b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26b7da),
	.w1(32'h3beabaa4),
	.w2(32'h3b6d4a8a),
	.w3(32'h3baeb48c),
	.w4(32'h3c0539fa),
	.w5(32'hbb3473d2),
	.w6(32'h3c095495),
	.w7(32'h3c3b72bb),
	.w8(32'h3aa43c26),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba865dc5),
	.w1(32'h3b1ba230),
	.w2(32'hb8c1f0b3),
	.w3(32'hbb395c29),
	.w4(32'h3a9fd9c1),
	.w5(32'h3979a51c),
	.w6(32'hbb1557b7),
	.w7(32'h3ab56474),
	.w8(32'h3a95a9e2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53abc7),
	.w1(32'h3bc2140d),
	.w2(32'hba7ccf38),
	.w3(32'hb73fdc7f),
	.w4(32'h3be4215d),
	.w5(32'h3bad2bb6),
	.w6(32'hba368f39),
	.w7(32'h3bde5943),
	.w8(32'h3b5c57cd),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c13a1),
	.w1(32'h3aee92d9),
	.w2(32'hbabebf61),
	.w3(32'h3a9b4ea9),
	.w4(32'h3ba8b221),
	.w5(32'hbb56dcfe),
	.w6(32'h3a2b369c),
	.w7(32'h3c2526c8),
	.w8(32'hbad99c8b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b540194),
	.w1(32'h3b3ac112),
	.w2(32'h39239936),
	.w3(32'h3a60d9bc),
	.w4(32'hbb25645e),
	.w5(32'h3b5eb7d1),
	.w6(32'hbaa52bd1),
	.w7(32'hbb6fb991),
	.w8(32'h3944dc15),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff3123),
	.w1(32'hbb514d16),
	.w2(32'hbbea9bda),
	.w3(32'hbbb29ff8),
	.w4(32'hbb13ac43),
	.w5(32'hbaf50c79),
	.w6(32'hbc0646a6),
	.w7(32'hbb747e2f),
	.w8(32'h3b5dea5c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3910833c),
	.w1(32'hbbcc2c42),
	.w2(32'hbbdb2ffc),
	.w3(32'hbad3c081),
	.w4(32'hbbfde45b),
	.w5(32'hbb901e27),
	.w6(32'h3c211fb1),
	.w7(32'hbba13284),
	.w8(32'h3b879968),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39b7bc),
	.w1(32'h3bf7fd46),
	.w2(32'h3bfb2914),
	.w3(32'h3a94a84c),
	.w4(32'h3b6eb968),
	.w5(32'h3a8109a6),
	.w6(32'h3c765973),
	.w7(32'h39f8cd88),
	.w8(32'hba6dbad5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25d6df),
	.w1(32'h3c1bef54),
	.w2(32'h3b8c9cc6),
	.w3(32'h3c0a494e),
	.w4(32'h3c0068ed),
	.w5(32'hba1b30e9),
	.w6(32'h3c6ae0a6),
	.w7(32'h3c031dfe),
	.w8(32'h3b5c07b7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc427e),
	.w1(32'h3b7e250b),
	.w2(32'h3b0a99de),
	.w3(32'hbc1b5bf4),
	.w4(32'h3c06e19f),
	.w5(32'hbae0ac2c),
	.w6(32'hbbf33c91),
	.w7(32'h3b5c4466),
	.w8(32'hbb887eaf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a45e8),
	.w1(32'hb9d747c5),
	.w2(32'h3bb57365),
	.w3(32'hbb8ccd25),
	.w4(32'hbb9ec252),
	.w5(32'h3b536abf),
	.w6(32'hba464c84),
	.w7(32'hbbbb3038),
	.w8(32'hbb09d5c8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42f2b1),
	.w1(32'hbbc898cd),
	.w2(32'hbbb7f199),
	.w3(32'hbb171ac7),
	.w4(32'hbc14da64),
	.w5(32'hbbbe9723),
	.w6(32'hba817a97),
	.w7(32'hbbe9f749),
	.w8(32'hbc104289),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc54f8),
	.w1(32'h3b430705),
	.w2(32'h3b6c4f3c),
	.w3(32'h3bcefae8),
	.w4(32'h3b2ece0a),
	.w5(32'h3b62e8ca),
	.w6(32'h3baed044),
	.w7(32'h3ae566ab),
	.w8(32'h3b0946d2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4b121),
	.w1(32'h3c7074b0),
	.w2(32'h3c10638d),
	.w3(32'h3b01c175),
	.w4(32'hbbada9c1),
	.w5(32'hbbd20091),
	.w6(32'h3a734add),
	.w7(32'hbb2634bf),
	.w8(32'hbb381a92),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bd81e),
	.w1(32'hbbf259ea),
	.w2(32'hb9f4a184),
	.w3(32'hbc25d272),
	.w4(32'hbbea990c),
	.w5(32'h3b47e3a5),
	.w6(32'hbb2f9dcf),
	.w7(32'hbc08bf29),
	.w8(32'hbb77a8a4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a199130),
	.w1(32'h3bf8b228),
	.w2(32'h3b47b9c1),
	.w3(32'hbb301735),
	.w4(32'h3ae109b7),
	.w5(32'hbb54ee5e),
	.w6(32'h3ac0044e),
	.w7(32'h3b8560a2),
	.w8(32'hbaafc3e5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba68f07),
	.w1(32'hbb8741ce),
	.w2(32'h3b7f5dbe),
	.w3(32'h3b06fd5c),
	.w4(32'hbb404d5a),
	.w5(32'h3ba22a0d),
	.w6(32'h3bc90811),
	.w7(32'hbb87d48f),
	.w8(32'h3b677677),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e27f26),
	.w1(32'h3a7d918d),
	.w2(32'h3b8a7bea),
	.w3(32'hbb142d85),
	.w4(32'h3b3474c9),
	.w5(32'h3b492d5d),
	.w6(32'hbb5c8f7f),
	.w7(32'h3a17fbe6),
	.w8(32'h3a38e120),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ae864),
	.w1(32'h3b301b75),
	.w2(32'h3bab77d2),
	.w3(32'h398a0e85),
	.w4(32'h3b89abf1),
	.w5(32'h3bd4f281),
	.w6(32'h3b9e3847),
	.w7(32'h3c4cf361),
	.w8(32'h3c02f64d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba802ff3),
	.w1(32'h3b385de9),
	.w2(32'h3bde29d7),
	.w3(32'h3b6f25d4),
	.w4(32'hbbb2830c),
	.w5(32'hbb99565b),
	.w6(32'hbbe33483),
	.w7(32'hbbff598e),
	.w8(32'hbad0e7b5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc699e6),
	.w1(32'hbba0c42b),
	.w2(32'hbbd00fbf),
	.w3(32'hbb8fe908),
	.w4(32'hbc1625f5),
	.w5(32'hbb8d3652),
	.w6(32'hbb21b16b),
	.w7(32'hbb8a4964),
	.w8(32'hbbac749f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab958a3),
	.w1(32'h3b6a209c),
	.w2(32'h3b2126d0),
	.w3(32'h3b4c2dac),
	.w4(32'hb98eb9fe),
	.w5(32'hbac7d46c),
	.w6(32'h3b96fcfc),
	.w7(32'h3b843b23),
	.w8(32'h3ab713c4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3a759),
	.w1(32'h3c205601),
	.w2(32'h3ace7e98),
	.w3(32'hbb9b7917),
	.w4(32'h3c31e7b7),
	.w5(32'hba572956),
	.w6(32'h3bb3cfd8),
	.w7(32'h3c31eb86),
	.w8(32'h3aba362b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6436ab),
	.w1(32'h3bfcd068),
	.w2(32'h3c904336),
	.w3(32'h3b02d84a),
	.w4(32'h3c21a865),
	.w5(32'h3c637358),
	.w6(32'h3bdb022b),
	.w7(32'h3c4a54bf),
	.w8(32'h3c775247),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac80e85),
	.w1(32'hbb7e139b),
	.w2(32'h3875ad6f),
	.w3(32'h3ab51e22),
	.w4(32'hbbc4f81c),
	.w5(32'hbb5cbe2c),
	.w6(32'hb9fa1a20),
	.w7(32'hbbfce35c),
	.w8(32'hbb7b6d42),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86da88),
	.w1(32'hbb1ed694),
	.w2(32'hba89e575),
	.w3(32'hbbb793ff),
	.w4(32'hbb86b180),
	.w5(32'hbbac5f54),
	.w6(32'hbbd0c865),
	.w7(32'h397f48d7),
	.w8(32'hbad836aa),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912dc5b),
	.w1(32'hbaa5add2),
	.w2(32'h3b7a6698),
	.w3(32'h3b849452),
	.w4(32'hbb4fce5d),
	.w5(32'h3b0fcd10),
	.w6(32'h3b8997cb),
	.w7(32'hbbd5b10f),
	.w8(32'hbb776ae7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b2248),
	.w1(32'hbb9b23fe),
	.w2(32'hbb25503d),
	.w3(32'h3a4198c9),
	.w4(32'hbb543618),
	.w5(32'hbaeddc28),
	.w6(32'h3a948c44),
	.w7(32'hbb01ba8d),
	.w8(32'h3a257f90),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba303787),
	.w1(32'hbac40d1a),
	.w2(32'h3a63b05e),
	.w3(32'h3b6c951c),
	.w4(32'hbb447f62),
	.w5(32'hba163bdb),
	.w6(32'h3ae720bf),
	.w7(32'hbb98d989),
	.w8(32'hbba46dda),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af66cc7),
	.w1(32'h3719fc41),
	.w2(32'h3bcfeb9d),
	.w3(32'h3af31f10),
	.w4(32'h3b62db9b),
	.w5(32'h3b84ce03),
	.w6(32'hbb79f880),
	.w7(32'hba89b8e6),
	.w8(32'hb9f5e503),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e3cd5),
	.w1(32'h37738552),
	.w2(32'hbb1c3550),
	.w3(32'hb9c7e1a8),
	.w4(32'hbb84e50a),
	.w5(32'hbbaa2995),
	.w6(32'hbbb63150),
	.w7(32'hbb1276ea),
	.w8(32'hbb43e1b4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5790a),
	.w1(32'hbb367218),
	.w2(32'hbb12d006),
	.w3(32'hbc01ce32),
	.w4(32'hbb54ee0b),
	.w5(32'hbac6787c),
	.w6(32'hbbbbcc7c),
	.w7(32'h3b49a52f),
	.w8(32'h3b058576),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968d065),
	.w1(32'h3b9be86e),
	.w2(32'h3c05064d),
	.w3(32'h38fa423e),
	.w4(32'h3c1ee591),
	.w5(32'h3c8b2c29),
	.w6(32'h3bba144c),
	.w7(32'h3b597c79),
	.w8(32'h3bf023e4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394fa778),
	.w1(32'h3b299c9a),
	.w2(32'h3b2b5b56),
	.w3(32'h3c030f34),
	.w4(32'hba5ce29a),
	.w5(32'h3bad3bb8),
	.w6(32'hbaeb789e),
	.w7(32'hbb65f0a8),
	.w8(32'h3bfbc3f9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3464af),
	.w1(32'h3ac3ee98),
	.w2(32'hb94ef3f9),
	.w3(32'h3989938d),
	.w4(32'h3a9a4adc),
	.w5(32'hbb76ffd4),
	.w6(32'h3b5664f2),
	.w7(32'h3a08a0ab),
	.w8(32'h3a988a10),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b7e53),
	.w1(32'h371f5c56),
	.w2(32'hb9b083bd),
	.w3(32'hba9fa99d),
	.w4(32'hbaa3c6c2),
	.w5(32'hbbb9f95d),
	.w6(32'hb9ffbe9d),
	.w7(32'h3a7968a9),
	.w8(32'hbb4b6945),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd255b),
	.w1(32'hbac1492e),
	.w2(32'h39b87d4e),
	.w3(32'h3a8697f4),
	.w4(32'h3b58e45e),
	.w5(32'hba214b19),
	.w6(32'hbbc024d5),
	.w7(32'h3a0770d2),
	.w8(32'hbbd7288f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c675a),
	.w1(32'hbb9acefa),
	.w2(32'hbad1e49a),
	.w3(32'h3ad049c4),
	.w4(32'hbb719a45),
	.w5(32'hbb4f4778),
	.w6(32'hbbb431c4),
	.w7(32'hbb6ae6d6),
	.w8(32'h3ac7c548),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af25ea4),
	.w1(32'hb98aafbf),
	.w2(32'h38f2ba04),
	.w3(32'hbb06ef78),
	.w4(32'hbb955819),
	.w5(32'hba982dd0),
	.w6(32'h3b81bba9),
	.w7(32'hbbe1ba27),
	.w8(32'hbb24e25a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36e257),
	.w1(32'hba67d282),
	.w2(32'h3a342e09),
	.w3(32'hb949ef06),
	.w4(32'h393b7fa0),
	.w5(32'h3b4e1c79),
	.w6(32'h3b1713ef),
	.w7(32'hbaca449c),
	.w8(32'h3a2d07a7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81bbf9),
	.w1(32'hbbd8942e),
	.w2(32'h3a638a29),
	.w3(32'h3acf9d2e),
	.w4(32'h3b403475),
	.w5(32'h3b77e868),
	.w6(32'h3b7749cb),
	.w7(32'h3b2de168),
	.w8(32'h3b7b1a12),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0511ac),
	.w1(32'h3aee7b7a),
	.w2(32'hbba32ef0),
	.w3(32'hba6c73ba),
	.w4(32'hbbc1c9a0),
	.w5(32'hbbc1e167),
	.w6(32'hbb54996e),
	.w7(32'hb8c93f9e),
	.w8(32'hba85ec58),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6513f9),
	.w1(32'hba6eab99),
	.w2(32'h39841a65),
	.w3(32'hbb537292),
	.w4(32'hbbe711e0),
	.w5(32'hbb3ed2aa),
	.w6(32'h3bbb86eb),
	.w7(32'hbb200766),
	.w8(32'hbb8a7c74),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90d6c1),
	.w1(32'hb9bbf988),
	.w2(32'h3aa0055e),
	.w3(32'h3a044c61),
	.w4(32'hbae9e3b9),
	.w5(32'h378131e0),
	.w6(32'h3a4627df),
	.w7(32'hbb22bb0a),
	.w8(32'hbb834b69),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a81e63),
	.w1(32'h37a325f4),
	.w2(32'h3b3e1e54),
	.w3(32'h3c03321b),
	.w4(32'h3b8b4619),
	.w5(32'h3bd39cc1),
	.w6(32'h3857ffbd),
	.w7(32'hba268a98),
	.w8(32'hbb3bb069),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0f0c7),
	.w1(32'h3c519eff),
	.w2(32'h3bab5522),
	.w3(32'h3ba5f3b4),
	.w4(32'h3a88faac),
	.w5(32'hbbbbf073),
	.w6(32'hbae9bc76),
	.w7(32'h3b286f21),
	.w8(32'hba41b9d4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0aa69),
	.w1(32'h3c54abd4),
	.w2(32'h3bd097ed),
	.w3(32'h3aa0e932),
	.w4(32'h3bbccf60),
	.w5(32'h39e6237d),
	.w6(32'h3b35dbbe),
	.w7(32'h3b6a51b2),
	.w8(32'hba1d059a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c7a84),
	.w1(32'hba670e8c),
	.w2(32'h3b0e6cd3),
	.w3(32'h3a24dc99),
	.w4(32'hbaf56d25),
	.w5(32'hbae22f77),
	.w6(32'h3a0fe345),
	.w7(32'hbb1912a9),
	.w8(32'hbb2e6cc6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395bd5d4),
	.w1(32'h3b1b53a0),
	.w2(32'h3b9a4d6c),
	.w3(32'hbbc68fb4),
	.w4(32'h39f7a9d9),
	.w5(32'h3c0744fa),
	.w6(32'hbb029369),
	.w7(32'hbb6a4688),
	.w8(32'h3c47d20b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82ec1d),
	.w1(32'h38bcb77d),
	.w2(32'h3bcfde43),
	.w3(32'h3bb89e78),
	.w4(32'h3ba48da9),
	.w5(32'h3b86e1d7),
	.w6(32'h3c1710e3),
	.w7(32'h3b906beb),
	.w8(32'h3b05436a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baecbe4),
	.w1(32'hbb17be52),
	.w2(32'h3a752786),
	.w3(32'h3b97aa5d),
	.w4(32'h3b4c3a26),
	.w5(32'h3c278782),
	.w6(32'hbb6f7ee5),
	.w7(32'hbb86686c),
	.w8(32'h3aa66489),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb770d7c),
	.w1(32'hba8fc0f8),
	.w2(32'hba474007),
	.w3(32'h3bf9161b),
	.w4(32'hb8713a44),
	.w5(32'h39d66e19),
	.w6(32'h3b24bfef),
	.w7(32'h3a22eeda),
	.w8(32'h3a19e2b3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cf9016),
	.w1(32'h3ba95569),
	.w2(32'hbb4a6ca4),
	.w3(32'h3b35d21b),
	.w4(32'hbb8069d0),
	.w5(32'hbbd91002),
	.w6(32'h3abed407),
	.w7(32'hb99a2a48),
	.w8(32'hbb8e6aa0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadad00),
	.w1(32'h3b1329d8),
	.w2(32'h3bfe0e63),
	.w3(32'h3b106826),
	.w4(32'h3ba3405b),
	.w5(32'h3c070494),
	.w6(32'h3bba781e),
	.w7(32'h3c2a751d),
	.w8(32'h3c550819),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fe7bb),
	.w1(32'h3abb6f24),
	.w2(32'hb6ab76f3),
	.w3(32'h3af8631c),
	.w4(32'h3a98d7d3),
	.w5(32'h39e02524),
	.w6(32'h3b52df81),
	.w7(32'hbbc1c16c),
	.w8(32'hbb53b927),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399dd22a),
	.w1(32'h3c1da542),
	.w2(32'h3c1e8a70),
	.w3(32'h3ac9e707),
	.w4(32'h3c382b9e),
	.w5(32'h3c3a39ed),
	.w6(32'hb9dae7d8),
	.w7(32'h3bcf0195),
	.w8(32'h3c22d591),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b680593),
	.w1(32'h3ba3ad65),
	.w2(32'h3bd0b94f),
	.w3(32'h3b3ce56c),
	.w4(32'h3b6e8ada),
	.w5(32'h3b2b2a0c),
	.w6(32'h3abe9439),
	.w7(32'h3b1b81eb),
	.w8(32'h3adc1650),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cf6bd),
	.w1(32'hbbeab9c5),
	.w2(32'hbc2dcb9b),
	.w3(32'h3b9aa55e),
	.w4(32'h3aadf44c),
	.w5(32'hbaef3e45),
	.w6(32'h3b731cf0),
	.w7(32'h3c062fa4),
	.w8(32'h3c14b164),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc091616),
	.w1(32'hbba7650a),
	.w2(32'hb93d2d5c),
	.w3(32'hbaccebc5),
	.w4(32'hbbb22717),
	.w5(32'hbbd250c4),
	.w6(32'h3c1d68bd),
	.w7(32'hbb38fc6a),
	.w8(32'hbb44eed3),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44ba08),
	.w1(32'h3b1e1903),
	.w2(32'h3998ea4c),
	.w3(32'hbba65e78),
	.w4(32'h3adc66af),
	.w5(32'hba7811fb),
	.w6(32'hbb33342e),
	.w7(32'hb9b7b963),
	.w8(32'hb8ddf89d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12fb26),
	.w1(32'h39cb0495),
	.w2(32'hbb0785b5),
	.w3(32'hbb948b81),
	.w4(32'hb7b1cd4b),
	.w5(32'hb7ec8911),
	.w6(32'hbbcdd9d5),
	.w7(32'h3a6f376c),
	.w8(32'hb66eeaa4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba98307),
	.w1(32'h3bf52a22),
	.w2(32'h3b150c0e),
	.w3(32'h3bbfd641),
	.w4(32'h3bb1b2ed),
	.w5(32'h3a80ada1),
	.w6(32'h3b83c41f),
	.w7(32'h3c532942),
	.w8(32'h3ad9337f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06bbc4),
	.w1(32'h3a3861e0),
	.w2(32'h3b75464f),
	.w3(32'h3ba7e6f3),
	.w4(32'h3b059a64),
	.w5(32'h3adbb80b),
	.w6(32'h3aab8bfd),
	.w7(32'h3b97b034),
	.w8(32'h3abff4ef),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89ae73),
	.w1(32'hbbaff771),
	.w2(32'hbb36837d),
	.w3(32'h3b272e55),
	.w4(32'hba2c3cbc),
	.w5(32'hbb4172c4),
	.w6(32'h3b1e80e7),
	.w7(32'h3b744f16),
	.w8(32'h3a1736fc),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1d2e4),
	.w1(32'hbbab82d3),
	.w2(32'hb9a42d49),
	.w3(32'hbb613b79),
	.w4(32'hbba37a24),
	.w5(32'h3b4b6cc9),
	.w6(32'hbb9b11c2),
	.w7(32'hbba9cb15),
	.w8(32'h3b5b528f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb60add),
	.w1(32'h3ab3bad4),
	.w2(32'hba0e9184),
	.w3(32'h3a11d0d7),
	.w4(32'hbb0ef26e),
	.w5(32'hbb985291),
	.w6(32'h3b4c2edc),
	.w7(32'h3b092042),
	.w8(32'hbb32baec),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea579b),
	.w1(32'h3b9f7cbd),
	.w2(32'hbb63cdfb),
	.w3(32'hbad2cc3f),
	.w4(32'h3c49088e),
	.w5(32'hbb378e6c),
	.w6(32'hbae456bc),
	.w7(32'h3c92c668),
	.w8(32'hbaddee37),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7c303),
	.w1(32'h39f64c1e),
	.w2(32'hbb85b666),
	.w3(32'hba0d2d50),
	.w4(32'hbbb19d74),
	.w5(32'hbc0c1980),
	.w6(32'hbb890aee),
	.w7(32'hbae4eb03),
	.w8(32'hbb8b5ab5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad493af),
	.w1(32'h3b31d713),
	.w2(32'hbb9c98dc),
	.w3(32'hba4e6a73),
	.w4(32'h3b63dbce),
	.w5(32'hbb44b992),
	.w6(32'h3b00420a),
	.w7(32'h3ba7555b),
	.w8(32'hbaf6cfc3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf397c7),
	.w1(32'hba066361),
	.w2(32'hbb2d6e0d),
	.w3(32'h3936e3b8),
	.w4(32'hb9f5c6a1),
	.w5(32'hb855c754),
	.w6(32'hbb00ba3a),
	.w7(32'h3afb5189),
	.w8(32'h3acc7396),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b613757),
	.w1(32'h3c1569b6),
	.w2(32'h3aee20f7),
	.w3(32'h3c01f3fe),
	.w4(32'h3c025ce0),
	.w5(32'h3a128e06),
	.w6(32'h3bd4ea27),
	.w7(32'h3c21378b),
	.w8(32'h3af2dbed),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad02857),
	.w1(32'hbafbc6d3),
	.w2(32'hbb061c50),
	.w3(32'hbb66dab1),
	.w4(32'hbb89111c),
	.w5(32'hbbae4994),
	.w6(32'hbb24d23c),
	.w7(32'hbc0c8406),
	.w8(32'hbbb4972c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c128f77),
	.w1(32'hbc1a3556),
	.w2(32'hbbd4f83d),
	.w3(32'h3ba934ac),
	.w4(32'hbbeca299),
	.w5(32'hbb5b1ef6),
	.w6(32'h3afe4a61),
	.w7(32'hbb83e542),
	.w8(32'hba966abb),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8d853),
	.w1(32'hba98404f),
	.w2(32'h3a6d0cf7),
	.w3(32'hbae14f77),
	.w4(32'hbb888357),
	.w5(32'hba8fa2f8),
	.w6(32'hbad4213a),
	.w7(32'hbb566152),
	.w8(32'hbafe37d0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a4ec8),
	.w1(32'hbb586af1),
	.w2(32'hba01d14c),
	.w3(32'h3a8cfd18),
	.w4(32'hbb0e66ed),
	.w5(32'h38c7fc7d),
	.w6(32'h3accd703),
	.w7(32'hba438551),
	.w8(32'hba9de928),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b539af8),
	.w1(32'hbc022887),
	.w2(32'hbc0a3a93),
	.w3(32'h3b0b86c2),
	.w4(32'hbbc1a3bf),
	.w5(32'hbb415e38),
	.w6(32'h3bab4efc),
	.w7(32'hbb0e6363),
	.w8(32'h3b59967a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7212a),
	.w1(32'hbac97a77),
	.w2(32'hbad7e5a7),
	.w3(32'h3a126b98),
	.w4(32'hbbbb9efe),
	.w5(32'hbbecb5cd),
	.w6(32'hba821082),
	.w7(32'hbaa3a539),
	.w8(32'hbbd20c30),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a06f5),
	.w1(32'h38e5d3fd),
	.w2(32'h3b9526f4),
	.w3(32'hbb6cdfca),
	.w4(32'hbaeded5a),
	.w5(32'hb9e31d6a),
	.w6(32'hbb2279eb),
	.w7(32'h3b275e0d),
	.w8(32'h3b1d542d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add97a7),
	.w1(32'hbab49294),
	.w2(32'h3b43c069),
	.w3(32'hbb927810),
	.w4(32'hbb1cb90b),
	.w5(32'h3b77eee7),
	.w6(32'hbbab129b),
	.w7(32'hbaefd4e5),
	.w8(32'h3bacf1b8),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b1193),
	.w1(32'h391595c9),
	.w2(32'hbb33c050),
	.w3(32'h3b9d95a6),
	.w4(32'h3ab2c599),
	.w5(32'hbadc74b1),
	.w6(32'h3c0f14ce),
	.w7(32'h3b3c9357),
	.w8(32'h3b21c4c5),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52a7b4),
	.w1(32'hbacc4690),
	.w2(32'hbb2fa245),
	.w3(32'hbb880fef),
	.w4(32'h3960903a),
	.w5(32'h39aff0e7),
	.w6(32'h3aac68e9),
	.w7(32'h3b8b116f),
	.w8(32'h3ac8aab8),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b1da4),
	.w1(32'hbb6c913e),
	.w2(32'hbc09aa17),
	.w3(32'hbb5f3c42),
	.w4(32'hb9aaef9e),
	.w5(32'hbb4bd552),
	.w6(32'hb94a4c85),
	.w7(32'h3b744f31),
	.w8(32'hbaf072df),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb770a41),
	.w1(32'hbaebfe31),
	.w2(32'h3a91eca8),
	.w3(32'hbadb5974),
	.w4(32'hb8d10e91),
	.w5(32'h3bbccde6),
	.w6(32'hbb12d6fd),
	.w7(32'hbb5a4a47),
	.w8(32'h3b69bbe3),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03bd66),
	.w1(32'h39f9a295),
	.w2(32'h3aa72d3f),
	.w3(32'hbb060bed),
	.w4(32'h3bf68a74),
	.w5(32'h3ba42ee2),
	.w6(32'hbb10296b),
	.w7(32'h3a79feaa),
	.w8(32'h3b9363a1),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9ce12),
	.w1(32'hbac2c09a),
	.w2(32'h3ae8d03a),
	.w3(32'hbbdc7aeb),
	.w4(32'hba6e6040),
	.w5(32'h3ba60598),
	.w6(32'hbba729c0),
	.w7(32'hbb8c4d0c),
	.w8(32'h3c20a675),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d418a),
	.w1(32'hb9ecc6a7),
	.w2(32'h3b1cd38d),
	.w3(32'h3bbf9f18),
	.w4(32'hbb7ad6c5),
	.w5(32'h3b1dfe06),
	.w6(32'h3be90df0),
	.w7(32'hbbd5d190),
	.w8(32'hbaae8614),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3d4aa),
	.w1(32'hbb21cbc0),
	.w2(32'hba8fc8b9),
	.w3(32'hbb16d41e),
	.w4(32'hbaeed508),
	.w5(32'h3b4d56d9),
	.w6(32'hbb60d2eb),
	.w7(32'hbb54f2e7),
	.w8(32'h3b66e640),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3e7fe),
	.w1(32'h3c38f511),
	.w2(32'h3b925c44),
	.w3(32'h3c1388c8),
	.w4(32'h3b626a9d),
	.w5(32'h39becd6c),
	.w6(32'h3c8254a4),
	.w7(32'h3c237e25),
	.w8(32'h3b4cd63c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a9ea0),
	.w1(32'hbba95902),
	.w2(32'hbb73be27),
	.w3(32'hbb1b7191),
	.w4(32'hbc10be31),
	.w5(32'hbb825007),
	.w6(32'hba76dfa8),
	.w7(32'hbbae1f8a),
	.w8(32'hbb97e153),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0b555),
	.w1(32'hbb2b6590),
	.w2(32'hbb297649),
	.w3(32'h3a8a9bbf),
	.w4(32'hba6b92a2),
	.w5(32'h39d4a178),
	.w6(32'hba69b5d6),
	.w7(32'hbb95aa51),
	.w8(32'hbaf31c4a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11a7d9),
	.w1(32'hbb73b3ac),
	.w2(32'hbb23effa),
	.w3(32'hba09bedb),
	.w4(32'hbb266531),
	.w5(32'h3b751d69),
	.w6(32'h389fd329),
	.w7(32'hbb99cbe1),
	.w8(32'hbadc4caa),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae82f50),
	.w1(32'h3a40fe19),
	.w2(32'h3ae7bbeb),
	.w3(32'h3b0d3ca3),
	.w4(32'h3ad242fb),
	.w5(32'h3b05fc46),
	.w6(32'h3a10b83e),
	.w7(32'h39c74c1f),
	.w8(32'hba1971ff),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31d1c9),
	.w1(32'hba121495),
	.w2(32'h3b98ec8f),
	.w3(32'hba5a0aec),
	.w4(32'hb9ac849d),
	.w5(32'h3b608824),
	.w6(32'h39406390),
	.w7(32'h3afd4524),
	.w8(32'h3aad1773),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba51599),
	.w1(32'h3be529b6),
	.w2(32'h3bccbfdc),
	.w3(32'h3b199e1e),
	.w4(32'h3b4de356),
	.w5(32'h3b2ce81b),
	.w6(32'h3bd7f023),
	.w7(32'h3b441b98),
	.w8(32'h3b6b94ac),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39256114),
	.w1(32'hbbb94ef1),
	.w2(32'hbba04c84),
	.w3(32'h37de5c5e),
	.w4(32'hbbcfd0d4),
	.w5(32'hbb8189c7),
	.w6(32'hba703a70),
	.w7(32'hbbb4cd26),
	.w8(32'hbb82ad69),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03c5ab),
	.w1(32'h3b9f1165),
	.w2(32'h3ba4776b),
	.w3(32'h3b4e991f),
	.w4(32'h3b730fef),
	.w5(32'h3ba40747),
	.w6(32'h3b58d32f),
	.w7(32'h3b2b1680),
	.w8(32'h3b6b3670),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badc942),
	.w1(32'hbb448545),
	.w2(32'h3b4ae527),
	.w3(32'h3b84c229),
	.w4(32'hbbc62bdf),
	.w5(32'h39e3180a),
	.w6(32'hb9a408c6),
	.w7(32'hbbc6cebd),
	.w8(32'hba0daec6),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9df6a8),
	.w1(32'hbad67286),
	.w2(32'hbb226d45),
	.w3(32'h3ae63a89),
	.w4(32'hbb49fc27),
	.w5(32'hbb95d692),
	.w6(32'h3b0b208b),
	.w7(32'hbb6ebe30),
	.w8(32'hbb616428),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2558e9),
	.w1(32'h3b16c0c7),
	.w2(32'hbb87d735),
	.w3(32'hbbc54591),
	.w4(32'h3b05e58c),
	.w5(32'hbb4922c3),
	.w6(32'hbb8735bf),
	.w7(32'hba0ed51d),
	.w8(32'hbb85eae3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd7a0d),
	.w1(32'hbb6ace04),
	.w2(32'hbab6020e),
	.w3(32'h3a7d3c59),
	.w4(32'hbb7891d2),
	.w5(32'hbae8352e),
	.w6(32'hba9f5135),
	.w7(32'hb9f42e40),
	.w8(32'h3b0be231),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c2818),
	.w1(32'hba20ac00),
	.w2(32'hbbc80e87),
	.w3(32'hb782ad3d),
	.w4(32'h3a8c686a),
	.w5(32'hbb88e5c2),
	.w6(32'h3bb16427),
	.w7(32'h38b74c5b),
	.w8(32'h3bb3481b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27b821),
	.w1(32'hba5f4611),
	.w2(32'hbb8c7873),
	.w3(32'h398071c7),
	.w4(32'h3b2c92cf),
	.w5(32'hba3c370b),
	.w6(32'h3bed3fb6),
	.w7(32'hbb089786),
	.w8(32'h3ba5e31c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad36aec),
	.w1(32'h3aa82ceb),
	.w2(32'hbb652950),
	.w3(32'h3bda6b1e),
	.w4(32'h3bc6e07d),
	.w5(32'h3a953337),
	.w6(32'h3c13ef8a),
	.w7(32'h3aa84150),
	.w8(32'h3c24b6d1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1baef),
	.w1(32'h3b45c9c9),
	.w2(32'h3adbe9dc),
	.w3(32'hba770b8d),
	.w4(32'hba3f5b8f),
	.w5(32'hbb8a1e28),
	.w6(32'h3bc95b31),
	.w7(32'h3b20b793),
	.w8(32'hba87df8e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb966b3c9),
	.w1(32'hbb57ca00),
	.w2(32'hbaf5cb1a),
	.w3(32'hba905589),
	.w4(32'hbaf5f6e1),
	.w5(32'hb7ea84bd),
	.w6(32'h3a3db09f),
	.w7(32'hbaf54d41),
	.w8(32'hba86987b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88c155),
	.w1(32'h3bf172e9),
	.w2(32'h3a856368),
	.w3(32'hbb8d53ef),
	.w4(32'h3c2ce4b5),
	.w5(32'h3a872727),
	.w6(32'hbb807b58),
	.w7(32'h3c154b59),
	.w8(32'h3acb1d01),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b320dbb),
	.w1(32'h3b21c5a7),
	.w2(32'h3b9974ba),
	.w3(32'h3bb46014),
	.w4(32'h3a88607f),
	.w5(32'h3b4c625c),
	.w6(32'h3bfb2e95),
	.w7(32'hbb234cfa),
	.w8(32'h3a2cc258),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf19c78),
	.w1(32'hbc042486),
	.w2(32'hbbe61258),
	.w3(32'hbb2b9f1e),
	.w4(32'hbbe6c531),
	.w5(32'hbb3d3268),
	.w6(32'hbb940447),
	.w7(32'hbc1d9ede),
	.w8(32'hbc017aee),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7a69c),
	.w1(32'h3ab188c0),
	.w2(32'h3a108136),
	.w3(32'hbb745a77),
	.w4(32'hba7f63c5),
	.w5(32'hbb27513a),
	.w6(32'hbb398200),
	.w7(32'h3accd41c),
	.w8(32'hbb0bf36a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2220f0),
	.w1(32'h3b629474),
	.w2(32'hbb6bf8bb),
	.w3(32'hba96881b),
	.w4(32'h3beab621),
	.w5(32'h3ba760a8),
	.w6(32'hba858054),
	.w7(32'h3ad4875d),
	.w8(32'h3ad2b2d4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac67636),
	.w1(32'h3aa2f9d2),
	.w2(32'h3a68fa64),
	.w3(32'h3ba49b92),
	.w4(32'hbb2ee2ed),
	.w5(32'hbbd459cb),
	.w6(32'h3bc46293),
	.w7(32'hbab1caff),
	.w8(32'hb992166f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f42cf),
	.w1(32'h3ac54721),
	.w2(32'h3b013e48),
	.w3(32'hbb5ee8b2),
	.w4(32'h3a8409ee),
	.w5(32'h3a207a3d),
	.w6(32'h3994d63b),
	.w7(32'h3ac95382),
	.w8(32'h3a8b65f5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f1d2b),
	.w1(32'hbb5b0248),
	.w2(32'h3ab5ce8a),
	.w3(32'h3b51f0bb),
	.w4(32'hbbb6ce89),
	.w5(32'h3b9a2ad6),
	.w6(32'h3b46c338),
	.w7(32'hbb2a655e),
	.w8(32'h3b584d21),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b129c42),
	.w1(32'hbb1e1779),
	.w2(32'hbb84d60c),
	.w3(32'h3b7a6402),
	.w4(32'hbb84d6e5),
	.w5(32'hbb940a4a),
	.w6(32'h3b9da76f),
	.w7(32'hbb2c7806),
	.w8(32'h3abd08f3),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a713c4d),
	.w1(32'h3aea8575),
	.w2(32'h3bd31781),
	.w3(32'h3ab777bb),
	.w4(32'h3b3f6191),
	.w5(32'h3b0472a2),
	.w6(32'h39ca36c5),
	.w7(32'hbb6f9d56),
	.w8(32'hbab2e203),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6a796),
	.w1(32'hbb8ca148),
	.w2(32'hbbd1745d),
	.w3(32'hbac29155),
	.w4(32'hbb6df4f1),
	.w5(32'hbb16aa41),
	.w6(32'h3ab4afc4),
	.w7(32'hbbab6e9d),
	.w8(32'h3a7c99b7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1691bc),
	.w1(32'h3b8238ab),
	.w2(32'hbb7736ba),
	.w3(32'hbb8c68e8),
	.w4(32'hba867999),
	.w5(32'hbb09ec59),
	.w6(32'hbb2ab1e3),
	.w7(32'hbb2233bf),
	.w8(32'h3bd2a983),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36b1ae),
	.w1(32'h3ba1bd99),
	.w2(32'h3badbda5),
	.w3(32'h3ba88a96),
	.w4(32'h3b407623),
	.w5(32'h3c2009b7),
	.w6(32'h3bf63332),
	.w7(32'h3b60e61e),
	.w8(32'h3ba8d088),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bb18d),
	.w1(32'hb99707ec),
	.w2(32'hbc1f7832),
	.w3(32'h3b8700ec),
	.w4(32'hbbc231f3),
	.w5(32'hbbe4cdc4),
	.w6(32'hbb123afd),
	.w7(32'hbb353baa),
	.w8(32'hbbe42d56),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1da111),
	.w1(32'h3c0376ad),
	.w2(32'h3b23fbc7),
	.w3(32'hbc60fcea),
	.w4(32'h3a985ed0),
	.w5(32'hba91dd30),
	.w6(32'hbafd15dc),
	.w7(32'hbab8c713),
	.w8(32'h3bb2f3c3),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd8bce),
	.w1(32'hbbdd20c4),
	.w2(32'h3baa57d4),
	.w3(32'h3b90034b),
	.w4(32'h3bd26304),
	.w5(32'h3d1ee487),
	.w6(32'h3b92d798),
	.w7(32'h3bd4d68f),
	.w8(32'h3c5b6c3b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5022a),
	.w1(32'h3b9406d3),
	.w2(32'h3bc5e511),
	.w3(32'h3c530ef1),
	.w4(32'hbb5c3150),
	.w5(32'hbc9aa12e),
	.w6(32'h3aff0d7b),
	.w7(32'hbc10560d),
	.w8(32'hbb933933),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1042d6),
	.w1(32'hbb6d2e2c),
	.w2(32'hbb40afa7),
	.w3(32'hbc455508),
	.w4(32'hbc4a0ee0),
	.w5(32'h3b03e617),
	.w6(32'h3b355eb3),
	.w7(32'hbc0e3aec),
	.w8(32'hbb39e19b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba714b2a),
	.w1(32'hbb4e0ad2),
	.w2(32'hb9047922),
	.w3(32'h3b6510bb),
	.w4(32'hbbc4b5cf),
	.w5(32'hbb9968b0),
	.w6(32'hbb18bba2),
	.w7(32'hbad866bc),
	.w8(32'h3b78079c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af64ec7),
	.w1(32'hbb9929d6),
	.w2(32'hbc5148c7),
	.w3(32'h3bfc16b6),
	.w4(32'h3c0a0022),
	.w5(32'hbbb3b985),
	.w6(32'h3bf51bb8),
	.w7(32'h3b41a5ca),
	.w8(32'h3ad8e15a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc115367),
	.w1(32'hbbfb526a),
	.w2(32'hbc8c1109),
	.w3(32'h3a86ff43),
	.w4(32'hbcb99f3d),
	.w5(32'hbcb37ab0),
	.w6(32'hba951ace),
	.w7(32'hbc371d10),
	.w8(32'hbc63380d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf17bae),
	.w1(32'h3b230498),
	.w2(32'h3c174041),
	.w3(32'hbc884ba0),
	.w4(32'h3b71689f),
	.w5(32'h3b6ee0e0),
	.w6(32'h3a7a6842),
	.w7(32'h3c055ab3),
	.w8(32'h3aa02b3a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b787b48),
	.w1(32'h3bf7e57a),
	.w2(32'h3c24cd9f),
	.w3(32'h3b3116f0),
	.w4(32'h3bbd74f1),
	.w5(32'h3a8ca17d),
	.w6(32'hbbcf3b7f),
	.w7(32'h3c17d076),
	.w8(32'hbb3681d1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b9997),
	.w1(32'hbb4a3519),
	.w2(32'h3bc93852),
	.w3(32'hbb497eb3),
	.w4(32'hba2ea2b9),
	.w5(32'h3c02ad05),
	.w6(32'h3ac443ef),
	.w7(32'h3b3c1073),
	.w8(32'h3b0e5324),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3612ba),
	.w1(32'h3b4b0fb1),
	.w2(32'hbba6f326),
	.w3(32'h39e0a6c0),
	.w4(32'hbb120ab1),
	.w5(32'hbb68127e),
	.w6(32'hbb1dbd0d),
	.w7(32'hbaffbf1c),
	.w8(32'hbbcd07be),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc108988),
	.w1(32'hbb034f58),
	.w2(32'h3b01ad15),
	.w3(32'hbc490d2a),
	.w4(32'hba4bf28e),
	.w5(32'h3bfdde61),
	.w6(32'hbc0e99fd),
	.w7(32'hbb5354a6),
	.w8(32'h3bd17463),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a297a2f),
	.w1(32'hbabd0cf2),
	.w2(32'h3c3ce99a),
	.w3(32'h3bb70b83),
	.w4(32'hbbf3995a),
	.w5(32'h3a5e2211),
	.w6(32'h3c6cb56b),
	.w7(32'h3c61f6d5),
	.w8(32'h3c902a28),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d132bc),
	.w1(32'hbbfcebf6),
	.w2(32'hbba9a9af),
	.w3(32'hbbdf551a),
	.w4(32'hbb21b37e),
	.w5(32'hba307d5c),
	.w6(32'hbbe76f79),
	.w7(32'hbbe44da3),
	.w8(32'hbbc7ccc5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d9244),
	.w1(32'hbbb9c05e),
	.w2(32'hbc35fbda),
	.w3(32'hbae4e78f),
	.w4(32'h3b956677),
	.w5(32'hbc1c44ee),
	.w6(32'hba960848),
	.w7(32'h39b74de8),
	.w8(32'hbbfd8aa4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f41d8),
	.w1(32'hbbf54891),
	.w2(32'hbc1e0bc9),
	.w3(32'h3ba04ec3),
	.w4(32'h3c050da8),
	.w5(32'h3d0135ac),
	.w6(32'hba021461),
	.w7(32'h3ae6896e),
	.w8(32'h3c1563cc),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacad841),
	.w1(32'h3af715bf),
	.w2(32'hbaddd264),
	.w3(32'h3cd22214),
	.w4(32'hba49b772),
	.w5(32'h3b7a43a7),
	.w6(32'hbad0a546),
	.w7(32'h3a4b5914),
	.w8(32'h3c87b14f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb65a0d),
	.w1(32'hbbfe23fd),
	.w2(32'hbc023473),
	.w3(32'h3b8546b0),
	.w4(32'hba75f59c),
	.w5(32'hbbc80c62),
	.w6(32'h392b342e),
	.w7(32'hba82a995),
	.w8(32'hbb1316f4),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6d524),
	.w1(32'h3c02bf95),
	.w2(32'h3c1e1aef),
	.w3(32'h3b8e8278),
	.w4(32'h3bf777f1),
	.w5(32'h3bb3b674),
	.w6(32'h3bcef806),
	.w7(32'h3aff7592),
	.w8(32'h3af41b0d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11a7a6),
	.w1(32'h38741161),
	.w2(32'h3ba00198),
	.w3(32'h3b7bf618),
	.w4(32'h3a814afb),
	.w5(32'h3b07d515),
	.w6(32'h3bc0d1b6),
	.w7(32'h3be30c44),
	.w8(32'h3b1927c0),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd6b60),
	.w1(32'hbb4a8c31),
	.w2(32'hbc9786ba),
	.w3(32'h3ac520e0),
	.w4(32'hbca65f61),
	.w5(32'hbca33bbb),
	.w6(32'h39f3da8b),
	.w7(32'hbbe439c2),
	.w8(32'hbc5bef88),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28ddc4),
	.w1(32'h3b17131e),
	.w2(32'hbb4e035b),
	.w3(32'hbc22971f),
	.w4(32'hbb678ebd),
	.w5(32'h38e85960),
	.w6(32'h3af2bca4),
	.w7(32'hbb3bc2b7),
	.w8(32'h387ab227),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b658c),
	.w1(32'hbc0a4b9f),
	.w2(32'h3a209045),
	.w3(32'hbb23d80f),
	.w4(32'hbaf9d3fb),
	.w5(32'hba6b9400),
	.w6(32'h3b1aceaa),
	.w7(32'h3b14186e),
	.w8(32'hbb92be17),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90d8b8),
	.w1(32'hbc3cc4e9),
	.w2(32'h3b552694),
	.w3(32'hbaecc17a),
	.w4(32'hbb9cfdd4),
	.w5(32'h3d15449b),
	.w6(32'h3b25222f),
	.w7(32'hbbc6ac8d),
	.w8(32'h3c74db09),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb714242),
	.w1(32'hbc85ee5b),
	.w2(32'hbbdea4af),
	.w3(32'h3bd2e867),
	.w4(32'hbc09b300),
	.w5(32'h3cf792b4),
	.w6(32'hbbaf2059),
	.w7(32'h39f7db88),
	.w8(32'h3caaf431),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0a5b2),
	.w1(32'hbaeb79a3),
	.w2(32'h3b88855f),
	.w3(32'h3c2fdc24),
	.w4(32'hb9e39fd6),
	.w5(32'hbb498335),
	.w6(32'hbb850faa),
	.w7(32'h3c0eeb5c),
	.w8(32'h3bd67493),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcefa3f),
	.w1(32'h3aa2b42e),
	.w2(32'h3a11e32e),
	.w3(32'h3bf038a0),
	.w4(32'hb93a9af4),
	.w5(32'hba9191b6),
	.w6(32'h3c104980),
	.w7(32'hbabfc6ce),
	.w8(32'hb80c3791),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4c2c9),
	.w1(32'h3be189f8),
	.w2(32'h3c018db3),
	.w3(32'h3b1aa75d),
	.w4(32'h3bcbd60d),
	.w5(32'h3bf347e2),
	.w6(32'h3b9ad2f1),
	.w7(32'hbbac4767),
	.w8(32'h3b266d6a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41ae8e),
	.w1(32'h3ad8ee68),
	.w2(32'h393079ba),
	.w3(32'h3bbb7275),
	.w4(32'h3bd15236),
	.w5(32'h3c96fa24),
	.w6(32'hbb244d16),
	.w7(32'h3b34470c),
	.w8(32'h3bd919f8),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b996a7f),
	.w1(32'hbbab9f20),
	.w2(32'h3bf4e3ef),
	.w3(32'h3c248caf),
	.w4(32'hbbe070f7),
	.w5(32'h3a01a9f2),
	.w6(32'h3aea2d5d),
	.w7(32'hbc2e6252),
	.w8(32'hbb097f44),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab826d5),
	.w1(32'hbb641593),
	.w2(32'hbb8b0f59),
	.w3(32'hbaa27cd9),
	.w4(32'h3b9d8815),
	.w5(32'h3d33e0c2),
	.w6(32'hbbef1290),
	.w7(32'h3c12bdb9),
	.w8(32'h3cc435dd),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb38f29),
	.w1(32'h3ab5c446),
	.w2(32'h3bb86368),
	.w3(32'h3c9f77c7),
	.w4(32'hbbcf7708),
	.w5(32'h3b0a460a),
	.w6(32'h3bb56e8f),
	.w7(32'h3b04506b),
	.w8(32'hbbdb2ba3),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a55bd),
	.w1(32'hb9a1a10a),
	.w2(32'hbbcc8da6),
	.w3(32'hbb9b85c7),
	.w4(32'hbc314ec8),
	.w5(32'hbbe48752),
	.w6(32'hbc063a32),
	.w7(32'h37c81e30),
	.w8(32'hbb750bd8),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6de690),
	.w1(32'hbb09363f),
	.w2(32'hbb225f0e),
	.w3(32'hbbbe5b7d),
	.w4(32'hba6d0420),
	.w5(32'h3a87e8f7),
	.w6(32'h3bd068a5),
	.w7(32'h3af7f58f),
	.w8(32'h3bee0750),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a6e79),
	.w1(32'h3bc1f12b),
	.w2(32'hbb5cd302),
	.w3(32'h3bac96d4),
	.w4(32'h3b178850),
	.w5(32'hbc2736dc),
	.w6(32'h3bdbfae3),
	.w7(32'h3adfe870),
	.w8(32'hbbb3e162),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65f265),
	.w1(32'h3b43db60),
	.w2(32'hbbb0e6bb),
	.w3(32'hbba6e48f),
	.w4(32'hbadc716c),
	.w5(32'hbb885ead),
	.w6(32'h391eca4c),
	.w7(32'h3acf69a5),
	.w8(32'hb9891afb),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b205fcc),
	.w1(32'hbc4ddc47),
	.w2(32'hbc2a361e),
	.w3(32'hbb28708a),
	.w4(32'hbc5342cf),
	.w5(32'hbc987623),
	.w6(32'h3bcc47c8),
	.w7(32'hbb9287c5),
	.w8(32'hbc76e856),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c70ac),
	.w1(32'hbbf61dbe),
	.w2(32'h3b22f4b4),
	.w3(32'hbc40e569),
	.w4(32'hbc7e8534),
	.w5(32'hbc946522),
	.w6(32'hbbc3eec7),
	.w7(32'hbbbc8bb4),
	.w8(32'h3ba65bcf),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9c1be),
	.w1(32'h3b786d02),
	.w2(32'h3b5d3d48),
	.w3(32'hbc8ec14f),
	.w4(32'h3b5d5561),
	.w5(32'h3c2e1718),
	.w6(32'hbc0bd67a),
	.w7(32'h3ade4aad),
	.w8(32'h3a2d16f0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b0b5a),
	.w1(32'h3b0ffeab),
	.w2(32'hbbdc1bd5),
	.w3(32'h3b39938f),
	.w4(32'hbb99fb27),
	.w5(32'h3ab55fc7),
	.w6(32'h3bfd24c1),
	.w7(32'h3b9c35af),
	.w8(32'h3b5e9353),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b156543),
	.w1(32'hbbf63988),
	.w2(32'h3b9dc181),
	.w3(32'h3b29ad1d),
	.w4(32'h3b55ba39),
	.w5(32'h3d1a507d),
	.w6(32'hbbbbcdf1),
	.w7(32'h3b86923a),
	.w8(32'h3c45028e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b591790),
	.w1(32'hba661252),
	.w2(32'h3b56dd5e),
	.w3(32'h3baa22fd),
	.w4(32'h3ad4cf51),
	.w5(32'hbc3573d2),
	.w6(32'hbc43ae1f),
	.w7(32'h39f3af95),
	.w8(32'hbc8d2cf0),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddf04d),
	.w1(32'h3b91d68a),
	.w2(32'hbbcf006f),
	.w3(32'hbc65be07),
	.w4(32'hbbc40a71),
	.w5(32'hbb86e740),
	.w6(32'hbbc076da),
	.w7(32'hbc075de3),
	.w8(32'hbbd666ca),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd79cd),
	.w1(32'h3b5d889f),
	.w2(32'h3b0d1351),
	.w3(32'hbbb0e9a6),
	.w4(32'h3a0dbb05),
	.w5(32'hbb540329),
	.w6(32'hbbdc498a),
	.w7(32'hbbcae54b),
	.w8(32'hba20788b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc71a1),
	.w1(32'hbc03efa6),
	.w2(32'h3bee84b9),
	.w3(32'hbb838c0d),
	.w4(32'hbbb66243),
	.w5(32'hbbd914a5),
	.w6(32'hbae2c26f),
	.w7(32'h3b2abf5b),
	.w8(32'h3c514df5),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac43381),
	.w1(32'h3b838045),
	.w2(32'hbc96ba3b),
	.w3(32'hbc11eccb),
	.w4(32'hbc85a1c3),
	.w5(32'hbc923dae),
	.w6(32'hbbcb8df0),
	.w7(32'hbc274309),
	.w8(32'hbc1208e1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc153f83),
	.w1(32'hbbb2e905),
	.w2(32'h3bdde9ac),
	.w3(32'hbc63b37b),
	.w4(32'h3bc7ada8),
	.w5(32'h3ce465f3),
	.w6(32'h3b976eb1),
	.w7(32'hbb7a1a25),
	.w8(32'h3babf427),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b0ccc),
	.w1(32'h3b035560),
	.w2(32'h3b9114d8),
	.w3(32'h3c4999f3),
	.w4(32'h3be1bb6e),
	.w5(32'h3caef1a7),
	.w6(32'h3b2235fb),
	.w7(32'h39aa51c6),
	.w8(32'h3c33f44d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c094c80),
	.w1(32'h3b53af18),
	.w2(32'hb9a24ec1),
	.w3(32'h3c2bd1c7),
	.w4(32'h3b816718),
	.w5(32'hbb6dd1cc),
	.w6(32'h3a92df78),
	.w7(32'h3ba56fbb),
	.w8(32'h3ac63cf9),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad83aac),
	.w1(32'h3c05a03c),
	.w2(32'h3b2c4ee3),
	.w3(32'hbad59cbe),
	.w4(32'h3b9a0167),
	.w5(32'h3ac7b95a),
	.w6(32'hba79050b),
	.w7(32'h3a0c825c),
	.w8(32'h3c065ba3),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb109af4),
	.w1(32'hbbc2dc5b),
	.w2(32'h3b1ca520),
	.w3(32'h39bb867e),
	.w4(32'h3be91695),
	.w5(32'h3d17267d),
	.w6(32'h3bb578fa),
	.w7(32'h3b939ad5),
	.w8(32'h3c52f343),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f0c56),
	.w1(32'h3b39db08),
	.w2(32'h3c4e7d13),
	.w3(32'h3c0248fe),
	.w4(32'h3c0ab3bb),
	.w5(32'h3cb4d4ea),
	.w6(32'hbb0e0c23),
	.w7(32'h3c0b3c37),
	.w8(32'h3c238671),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7df7a),
	.w1(32'hbbcbb784),
	.w2(32'hbc4341cc),
	.w3(32'h3c27656f),
	.w4(32'hbc586f47),
	.w5(32'hbcb42d1e),
	.w6(32'h3b78b0a2),
	.w7(32'hbbdccb5a),
	.w8(32'hbc1190a2),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec1dc0),
	.w1(32'hbbc79e22),
	.w2(32'hbb8311a6),
	.w3(32'hbc5e8ea1),
	.w4(32'hbc3a0242),
	.w5(32'h3a90dc4b),
	.w6(32'hbb03b8e9),
	.w7(32'hbbf4737d),
	.w8(32'hbc318d4b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01edb4),
	.w1(32'hbc05b2b2),
	.w2(32'hbbeb2b59),
	.w3(32'hbc8c2766),
	.w4(32'hbbac3d06),
	.w5(32'h3b7d6c2c),
	.w6(32'hbc0fb06d),
	.w7(32'hbb81efca),
	.w8(32'h3b6d815f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b891b88),
	.w1(32'hbab92870),
	.w2(32'hbc143292),
	.w3(32'h3c091968),
	.w4(32'hbb8539ac),
	.w5(32'hbc84c456),
	.w6(32'h3b859d42),
	.w7(32'hbbe7c8c7),
	.w8(32'hbc128c11),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule