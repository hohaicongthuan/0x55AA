module layer_10_featuremap_168(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb514c966),
	.w1(32'hb65085cc),
	.w2(32'h35d0358d),
	.w3(32'hb3cf9257),
	.w4(32'hb5cffbd2),
	.w5(32'h363fdd0e),
	.w6(32'hb6216b98),
	.w7(32'h36132cf7),
	.w8(32'hb5272d18),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb958beeb),
	.w1(32'h388a83ae),
	.w2(32'h397ba3a9),
	.w3(32'hb9912e33),
	.w4(32'hb8bb02a3),
	.w5(32'h38d03ccd),
	.w6(32'hb8ee32db),
	.w7(32'hb8b86a71),
	.w8(32'hb7b80805),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34f58a27),
	.w1(32'h34d5c73c),
	.w2(32'h34d824bc),
	.w3(32'h3579d0e4),
	.w4(32'hb50855bf),
	.w5(32'hb484be6b),
	.w6(32'h350eb7ca),
	.w7(32'hb426b321),
	.w8(32'hb4a5a5e3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dfba23),
	.w1(32'hb89649ef),
	.w2(32'hb8c08b7a),
	.w3(32'hb8692b27),
	.w4(32'hb877b538),
	.w5(32'hb816882c),
	.w6(32'h3719eba6),
	.w7(32'h37bf766e),
	.w8(32'hb7ca5408),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5dc4f75),
	.w1(32'h373be02a),
	.w2(32'h37e91cb5),
	.w3(32'hb7b36f49),
	.w4(32'hb72e5503),
	.w5(32'h372f31d4),
	.w6(32'hb7ab3d96),
	.w7(32'hb78a2129),
	.w8(32'h374308e0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3525f545),
	.w1(32'hb5c95922),
	.w2(32'hb6cc56fd),
	.w3(32'hb4f4fd20),
	.w4(32'hb6283d2f),
	.w5(32'hb6f31b57),
	.w6(32'h35f44852),
	.w7(32'hb5b486fe),
	.w8(32'hb5e83135),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1908bf),
	.w1(32'h3916a936),
	.w2(32'hb8a19975),
	.w3(32'h3a45c513),
	.w4(32'h39df9bc8),
	.w5(32'h3a67ef7c),
	.w6(32'hb98af0a9),
	.w7(32'h38a8ea72),
	.w8(32'h3a4f20a8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95edfa),
	.w1(32'h39c6cb6e),
	.w2(32'hba04c27a),
	.w3(32'h3a13edb4),
	.w4(32'h393a308a),
	.w5(32'h3aa55fda),
	.w6(32'h397d8351),
	.w7(32'h3a0a130d),
	.w8(32'h3983ff03),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379b9373),
	.w1(32'h386071e0),
	.w2(32'h38803cd3),
	.w3(32'h387c5e78),
	.w4(32'h38e101f1),
	.w5(32'h38d6265b),
	.w6(32'h3765abd1),
	.w7(32'h38763674),
	.w8(32'h38d52684),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a1d16e),
	.w1(32'hb9bb47ed),
	.w2(32'hb99afdf9),
	.w3(32'h38d96c5d),
	.w4(32'h39183c19),
	.w5(32'h38fa3af4),
	.w6(32'h3619a7c6),
	.w7(32'h346f4102),
	.w8(32'h39813e5d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36361767),
	.w1(32'hb7a37ad4),
	.w2(32'h38441303),
	.w3(32'hb815cf16),
	.w4(32'hb863a2fc),
	.w5(32'h373b3b31),
	.w6(32'hb8181192),
	.w7(32'hb83f6e40),
	.w8(32'h3781e6b0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb962629a),
	.w1(32'hb9de989c),
	.w2(32'hb9a7e59b),
	.w3(32'h3a156c1a),
	.w4(32'h37f1ee56),
	.w5(32'h3a0e9081),
	.w6(32'hb9bb8f9a),
	.w7(32'hb88d60ab),
	.w8(32'h384e1c68),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b4190),
	.w1(32'hb959683c),
	.w2(32'hb987d915),
	.w3(32'h3996a64b),
	.w4(32'h3992e985),
	.w5(32'h380f7d57),
	.w6(32'h394b5364),
	.w7(32'h398988c4),
	.w8(32'h39c6ab16),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a007b27),
	.w1(32'h39f01f2c),
	.w2(32'h3a0c2c90),
	.w3(32'h39bf51b9),
	.w4(32'h3a1ca96d),
	.w5(32'h3a31050e),
	.w6(32'hb8b1e64e),
	.w7(32'h382483ca),
	.w8(32'h39a5732d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9419e52),
	.w1(32'h38005107),
	.w2(32'h3866c341),
	.w3(32'hb92ed842),
	.w4(32'hb8904a33),
	.w5(32'h37d7bce5),
	.w6(32'hb8f2f25c),
	.w7(32'hb791ff8d),
	.w8(32'hb71ea209),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906c088),
	.w1(32'h390cd033),
	.w2(32'h3a18907a),
	.w3(32'hba1a3eb3),
	.w4(32'h3930a0ad),
	.w5(32'h384ece57),
	.w6(32'hb9a1c0ab),
	.w7(32'h366e4638),
	.w8(32'h3846da7a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80c7fc1),
	.w1(32'hb83f5947),
	.w2(32'hb7b18177),
	.w3(32'hb7be23e7),
	.w4(32'hb83ebd04),
	.w5(32'hb81da1e4),
	.w6(32'hb7b96772),
	.w7(32'hb849c185),
	.w8(32'hb7fa1d39),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a268d99),
	.w1(32'h39415577),
	.w2(32'hb9a61e3b),
	.w3(32'h39752326),
	.w4(32'h3a2834e5),
	.w5(32'h39816571),
	.w6(32'h372ac84f),
	.w7(32'h3957c737),
	.w8(32'h39bbc8f3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3973f58e),
	.w1(32'h35c61641),
	.w2(32'hb9288b72),
	.w3(32'h39801f37),
	.w4(32'h39944725),
	.w5(32'h39469ae0),
	.w6(32'h38c083cb),
	.w7(32'h392f286b),
	.w8(32'h398596e2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60e9e64),
	.w1(32'h3614ba87),
	.w2(32'hb58c6007),
	.w3(32'hb50c09ba),
	.w4(32'h363f2c84),
	.w5(32'h34f3151f),
	.w6(32'hb53e0aaa),
	.w7(32'hb5b08995),
	.w8(32'hb60a14a4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3652dcd0),
	.w1(32'h369fb939),
	.w2(32'hb67b5969),
	.w3(32'h367076b3),
	.w4(32'h3683be83),
	.w5(32'h31734680),
	.w6(32'h36d2ab6d),
	.w7(32'h36841378),
	.w8(32'h35dc32d3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e1627f),
	.w1(32'hb87b30b3),
	.w2(32'hb6f272e5),
	.w3(32'hb8f9ce05),
	.w4(32'hb8de9cc2),
	.w5(32'hb88dcf42),
	.w6(32'hb7b5a4a7),
	.w7(32'hb76933a9),
	.w8(32'hb771d0a4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31f70e),
	.w1(32'h39f1d3af),
	.w2(32'h39c16582),
	.w3(32'hb93ca75f),
	.w4(32'hb873e629),
	.w5(32'hb918becd),
	.w6(32'hba2aa4b7),
	.w7(32'hb9493ba4),
	.w8(32'hb869432b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901e0f1),
	.w1(32'hb9166157),
	.w2(32'hb89c9f47),
	.w3(32'hb8d646e4),
	.w4(32'hb8a14d43),
	.w5(32'h380cad3a),
	.w6(32'hb9146daa),
	.w7(32'hb8c42d51),
	.w8(32'h3783dce4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c8bfd),
	.w1(32'h388d0e54),
	.w2(32'h39dfb3de),
	.w3(32'hba30cd81),
	.w4(32'hb9712bc7),
	.w5(32'h38ef8b1b),
	.w6(32'hb9b65c7c),
	.w7(32'hb929546c),
	.w8(32'h3731305a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37118299),
	.w1(32'h364ccdd5),
	.w2(32'hb7097869),
	.w3(32'h374fd0de),
	.w4(32'h37ad8b2e),
	.w5(32'h375fc1d3),
	.w6(32'h3795fe94),
	.w7(32'h380d242b),
	.w8(32'h3815ed27),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3425f4f6),
	.w1(32'h360528b1),
	.w2(32'hb595918a),
	.w3(32'hb6ef2812),
	.w4(32'hb645eb62),
	.w5(32'hb6c2bf32),
	.w6(32'h365af7e2),
	.w7(32'h34153e46),
	.w8(32'hb454851e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8939cd),
	.w1(32'hb9ad28d2),
	.w2(32'h3989d47d),
	.w3(32'hb98747a2),
	.w4(32'h392e8972),
	.w5(32'hb9856039),
	.w6(32'h39beb275),
	.w7(32'h39fcf010),
	.w8(32'h3a2f9c10),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35581baa),
	.w1(32'h37f5fe08),
	.w2(32'h389ca66a),
	.w3(32'hb88e9b08),
	.w4(32'hb872089d),
	.w5(32'hb587c0c4),
	.w6(32'hb882901c),
	.w7(32'hb88eb9e1),
	.w8(32'hb809ad1d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba502258),
	.w1(32'hb9d3750b),
	.w2(32'hb9baefc1),
	.w3(32'hb9f076d2),
	.w4(32'hb99234ad),
	.w5(32'hb9b898d7),
	.w6(32'hb88de299),
	.w7(32'h3766dd3f),
	.w8(32'h36eceb01),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb639caf5),
	.w1(32'hb633d06f),
	.w2(32'hb624f06d),
	.w3(32'hb5d5d215),
	.w4(32'hb6665586),
	.w5(32'hb66539bd),
	.w6(32'h36693d7e),
	.w7(32'hb64aa6af),
	.w8(32'h339d599e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64e1dac),
	.w1(32'hb62b1159),
	.w2(32'hb637f308),
	.w3(32'hb6914bbb),
	.w4(32'hb72bb5a5),
	.w5(32'hb724c0ef),
	.w6(32'hb6c25fd2),
	.w7(32'hb7129685),
	.w8(32'hb694c0bd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384a64fb),
	.w1(32'hb80e2ea0),
	.w2(32'hb81c6732),
	.w3(32'h385a5592),
	.w4(32'h381eb9f6),
	.w5(32'h392e5fc4),
	.w6(32'hb89ed901),
	.w7(32'h37c0c4aa),
	.w8(32'h3901261d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb890abbd),
	.w1(32'h390f0dc4),
	.w2(32'h396de583),
	.w3(32'hb98d958a),
	.w4(32'hb64230c1),
	.w5(32'h39548999),
	.w6(32'hb901bd56),
	.w7(32'hb8e76f23),
	.w8(32'hb7898202),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9369a02),
	.w1(32'hb92ea054),
	.w2(32'hb8903354),
	.w3(32'h378a4ce1),
	.w4(32'hb71990cd),
	.w5(32'h37f70e58),
	.w6(32'hb7a8369b),
	.w7(32'h3794956a),
	.w8(32'h3804cbe0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbe4d6),
	.w1(32'h391eb7e2),
	.w2(32'hb8689862),
	.w3(32'h3895affc),
	.w4(32'h374afd63),
	.w5(32'h39956966),
	.w6(32'hb80e77aa),
	.w7(32'h386dbf6a),
	.w8(32'h3934194b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904af55),
	.w1(32'h3a32fa5f),
	.w2(32'h385427aa),
	.w3(32'h3a8defab),
	.w4(32'hb8264a09),
	.w5(32'h3a40d714),
	.w6(32'hb9c1fc1a),
	.w7(32'hba2c3531),
	.w8(32'hba580511),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b4f74),
	.w1(32'h399f8b93),
	.w2(32'h3a0eb270),
	.w3(32'hba72d995),
	.w4(32'hb99c6a86),
	.w5(32'hb9934f98),
	.w6(32'hba082ee6),
	.w7(32'hb96bde20),
	.w8(32'hb9a0bdb6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba639148),
	.w1(32'h3925c6ba),
	.w2(32'h397285da),
	.w3(32'hba1fedd8),
	.w4(32'hb91888bc),
	.w5(32'hb9d12411),
	.w6(32'hb9406436),
	.w7(32'h37bdbbc0),
	.w8(32'hb8b0d3fe),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b2e25c),
	.w1(32'hb766a2ff),
	.w2(32'hb7776d8c),
	.w3(32'hb8e151c2),
	.w4(32'hb89748f4),
	.w5(32'hb81e1737),
	.w6(32'hb804e779),
	.w7(32'h374f44ea),
	.w8(32'hb69a8ca6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3614a392),
	.w1(32'hb52bd7f5),
	.w2(32'hb79bdd15),
	.w3(32'h36806581),
	.w4(32'h35f7c9e8),
	.w5(32'hb77e95ff),
	.w6(32'h3742aee2),
	.w7(32'hb65d5e38),
	.w8(32'hb6df5d36),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e6b967),
	.w1(32'hb4a6a9d8),
	.w2(32'hb6252e5f),
	.w3(32'hb71fbcc6),
	.w4(32'hb6803bee),
	.w5(32'hb6c54856),
	.w6(32'h36aeb7ab),
	.w7(32'h35f32721),
	.w8(32'hb6057628),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a5d987),
	.w1(32'hb799db4e),
	.w2(32'h388fffad),
	.w3(32'hb7a054ee),
	.w4(32'hb68e064a),
	.w5(32'h388de7cc),
	.w6(32'hb6399c71),
	.w7(32'h37d3b07b),
	.w8(32'h38bd27a7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5e3c6),
	.w1(32'hb8d3c563),
	.w2(32'h395d7df6),
	.w3(32'hb98d4b27),
	.w4(32'h39f5decc),
	.w5(32'h3818698c),
	.w6(32'hb901dcf8),
	.w7(32'h39e4f30a),
	.w8(32'h398bf104),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8f325),
	.w1(32'hb8688eb0),
	.w2(32'h38b4ed0f),
	.w3(32'hb9e728fb),
	.w4(32'hb8ef5006),
	.w5(32'h37703385),
	.w6(32'hb8c50a9f),
	.w7(32'hb748f0e2),
	.w8(32'hb7bf8f4d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9208de5),
	.w1(32'h38c587da),
	.w2(32'h390305af),
	.w3(32'hba562d65),
	.w4(32'hb991bb94),
	.w5(32'h396eba84),
	.w6(32'hb89cf412),
	.w7(32'hb8920ec7),
	.w8(32'h37ed93b3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987eacc),
	.w1(32'hb90a4071),
	.w2(32'h3879303c),
	.w3(32'hb956f127),
	.w4(32'hb85836c2),
	.w5(32'hb831790b),
	.w6(32'hb8e29b1d),
	.w7(32'hb86a38ef),
	.w8(32'hb8559025),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40ff67),
	.w1(32'h387b82a8),
	.w2(32'hb9b4e006),
	.w3(32'h3a25435c),
	.w4(32'h39a98125),
	.w5(32'h39e79475),
	.w6(32'h3890151b),
	.w7(32'h38fd72f9),
	.w8(32'h39d3e94d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a561f4),
	.w1(32'h36373d81),
	.w2(32'hb5e78222),
	.w3(32'hb781e249),
	.w4(32'h35dccdca),
	.w5(32'h372c5fcf),
	.w6(32'hb6ece81f),
	.w7(32'h36d7dde2),
	.w8(32'h372d3b35),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e381e8),
	.w1(32'h3781f047),
	.w2(32'h36212e97),
	.w3(32'h37c8e223),
	.w4(32'h3847e14d),
	.w5(32'h38090973),
	.w6(32'hb6034cd0),
	.w7(32'h37322e50),
	.w8(32'h36bb04be),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b41344),
	.w1(32'hb7c4e6bc),
	.w2(32'hb63f447e),
	.w3(32'hb7df2462),
	.w4(32'hb798f9ce),
	.w5(32'h36773d2e),
	.w6(32'hb7d66de2),
	.w7(32'hb7b5fde9),
	.w8(32'hb666fe94),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391369c4),
	.w1(32'hb6f4b4e2),
	.w2(32'h39842eaf),
	.w3(32'hb951b123),
	.w4(32'h39048c83),
	.w5(32'hb89ee284),
	.w6(32'hb8c3a5bc),
	.w7(32'h388e30fb),
	.w8(32'hb844974e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38865f36),
	.w1(32'hb767dd39),
	.w2(32'h3789d15b),
	.w3(32'hb849ec14),
	.w4(32'hb89122ad),
	.w5(32'h388cf4f4),
	.w6(32'hb893bd9b),
	.w7(32'hb88eceb3),
	.w8(32'h37bd2df3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c48df4),
	.w1(32'h38d6020a),
	.w2(32'hb9942b6f),
	.w3(32'h39a0b4cb),
	.w4(32'h39d23398),
	.w5(32'h39c6767a),
	.w6(32'hb920d0da),
	.w7(32'h3869d0df),
	.w8(32'h3960f967),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70f2146),
	.w1(32'h3584a805),
	.w2(32'h3703496f),
	.w3(32'hb949836b),
	.w4(32'hb8247506),
	.w5(32'h368b469f),
	.w6(32'h38290984),
	.w7(32'h38d6858e),
	.w8(32'h37364461),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb815ce74),
	.w1(32'hb626511f),
	.w2(32'h3713cb54),
	.w3(32'hb7f885d6),
	.w4(32'hb76939a3),
	.w5(32'h36c5c935),
	.w6(32'hb673da22),
	.w7(32'hb64628b7),
	.w8(32'h35ee95e7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb625c17f),
	.w1(32'h35544287),
	.w2(32'hb6847ce8),
	.w3(32'hb707867d),
	.w4(32'hb69fca00),
	.w5(32'hb6bbddfd),
	.w6(32'hb6486433),
	.w7(32'hb6adbe85),
	.w8(32'hb70237a2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81379c2),
	.w1(32'hb61152e2),
	.w2(32'hb81ce728),
	.w3(32'hb7a96ade),
	.w4(32'hb6f76cfe),
	.w5(32'hb72f4b79),
	.w6(32'hb699735c),
	.w7(32'hb795fe69),
	.w8(32'h37b4243b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb857a2b2),
	.w1(32'hb7a532ac),
	.w2(32'h37a5d4a5),
	.w3(32'hb8971e03),
	.w4(32'hb83995c0),
	.w5(32'hb69a150a),
	.w6(32'hb83b8ce9),
	.w7(32'hb7ce69a0),
	.w8(32'h32bfad56),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79721f9),
	.w1(32'hb7ac37f5),
	.w2(32'hb610be8e),
	.w3(32'hb7e60b5b),
	.w4(32'hb7c7e5b0),
	.w5(32'hb75ed707),
	.w6(32'h3526f38a),
	.w7(32'hb797ea3f),
	.w8(32'h374a701b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388ea17b),
	.w1(32'h3722dd0b),
	.w2(32'hb8874783),
	.w3(32'h3806de2e),
	.w4(32'h3957c741),
	.w5(32'h391297f7),
	.w6(32'hb8226589),
	.w7(32'h391f3bc3),
	.w8(32'h38d91359),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1b5a0),
	.w1(32'hb93d05a2),
	.w2(32'h38ac6aad),
	.w3(32'hb97978cd),
	.w4(32'h393fbe22),
	.w5(32'hb90e7001),
	.w6(32'h3980dc95),
	.w7(32'h39b0e2c8),
	.w8(32'h395df45e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5dabbce),
	.w1(32'hb6392085),
	.w2(32'hb49807ad),
	.w3(32'hb55a8174),
	.w4(32'hb54d6305),
	.w5(32'hb5984b27),
	.w6(32'h35f07f66),
	.w7(32'h36c0eb56),
	.w8(32'hb6821291),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e131e1),
	.w1(32'hb62538ce),
	.w2(32'hb6b8cd8e),
	.w3(32'hb67b03fa),
	.w4(32'hb58b0b11),
	.w5(32'hb697d24b),
	.w6(32'h36460e4e),
	.w7(32'h3505a3fa),
	.w8(32'hb689e45c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36686436),
	.w1(32'h343b9ac5),
	.w2(32'hb3efc5d2),
	.w3(32'h36eba050),
	.w4(32'hb62fcf4f),
	.w5(32'h34ce14ce),
	.w6(32'h36eb3c8a),
	.w7(32'hb4af6a29),
	.w8(32'h35f902f7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361d65a3),
	.w1(32'h3617c5b0),
	.w2(32'hb6be2276),
	.w3(32'h3597fb5c),
	.w4(32'h36093da4),
	.w5(32'hb6603329),
	.w6(32'h36b37d3e),
	.w7(32'h345e1c9d),
	.w8(32'hb36eed56),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba801b46),
	.w1(32'hba8e47ad),
	.w2(32'hba104230),
	.w3(32'hb93f367d),
	.w4(32'h3a126ec7),
	.w5(32'h397bb370),
	.w6(32'h398b18ae),
	.w7(32'h393dcae7),
	.w8(32'h39d07e9f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cac5f3),
	.w1(32'h3a2cac5d),
	.w2(32'h3a43850c),
	.w3(32'hba90e049),
	.w4(32'hb9b2d395),
	.w5(32'h3a6735d6),
	.w6(32'hb9c544f2),
	.w7(32'h3880deba),
	.w8(32'h3a2e65cd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990e31b),
	.w1(32'h38b9f729),
	.w2(32'h3a1a1339),
	.w3(32'hb9a01773),
	.w4(32'h38daff3c),
	.w5(32'h3991f5a2),
	.w6(32'hb9542335),
	.w7(32'h391dc0be),
	.w8(32'h38ab0970),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3be25d),
	.w1(32'h3932260e),
	.w2(32'h3a25c198),
	.w3(32'hba6e2a0d),
	.w4(32'hb96f3536),
	.w5(32'h38869042),
	.w6(32'hb9fdba6d),
	.w7(32'hb96aac92),
	.w8(32'hb821c30e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b1382c),
	.w1(32'h33a9fb70),
	.w2(32'hb6ccc269),
	.w3(32'h36cb7abb),
	.w4(32'h355c9619),
	.w5(32'hb684f5df),
	.w6(32'h36b236bb),
	.w7(32'h361ef7f9),
	.w8(32'hb600336e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363abfff),
	.w1(32'h35ba119a),
	.w2(32'hb6f96b53),
	.w3(32'hb4ea560a),
	.w4(32'h35b006ea),
	.w5(32'hb71599c3),
	.w6(32'h36c134b5),
	.w7(32'h364705c5),
	.w8(32'hb5614c99),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb484800d),
	.w1(32'hb5e2336b),
	.w2(32'hb7472840),
	.w3(32'h34eca930),
	.w4(32'h32916be8),
	.w5(32'hb764cbd1),
	.w6(32'h3737c48d),
	.w7(32'h3677bbe3),
	.w8(32'hb636a3b8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922196b),
	.w1(32'h38d45b05),
	.w2(32'h3841426e),
	.w3(32'h391ba405),
	.w4(32'h3963e588),
	.w5(32'h38e916d6),
	.w6(32'h377ee06d),
	.w7(32'h38cb6fa3),
	.w8(32'h38d1036b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36213ab6),
	.w1(32'hb5db4a0f),
	.w2(32'hb6e7aaf8),
	.w3(32'h36e2f83b),
	.w4(32'h36578e1b),
	.w5(32'hb5828f08),
	.w6(32'h3724a17e),
	.w7(32'h370b5012),
	.w8(32'h35d5a080),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939e3ac),
	.w1(32'hb8f497a5),
	.w2(32'hb967c73d),
	.w3(32'h39d7ea67),
	.w4(32'h3924cb9d),
	.w5(32'h398c21d9),
	.w6(32'h395ca482),
	.w7(32'h390d9e40),
	.w8(32'h3898a21a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a321324),
	.w1(32'h39e4400d),
	.w2(32'hb7c2ecd3),
	.w3(32'h3a0c756f),
	.w4(32'h39a5aca8),
	.w5(32'h3a315ce8),
	.w6(32'hb7cbba0a),
	.w7(32'h39367470),
	.w8(32'h3885746f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc7212),
	.w1(32'hb903171a),
	.w2(32'h39361e41),
	.w3(32'hb9faaf6d),
	.w4(32'hb92d71b7),
	.w5(32'h379511eb),
	.w6(32'hb90fda93),
	.w7(32'hb8d34b9b),
	.w8(32'h36669657),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39314472),
	.w1(32'h38e217c3),
	.w2(32'h3915ad12),
	.w3(32'h3834ffd7),
	.w4(32'h3918c0df),
	.w5(32'h3912d7c8),
	.w6(32'hb8ed00cd),
	.w7(32'h37796a0f),
	.w8(32'h38c2f9ec),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9818266),
	.w1(32'hb9442671),
	.w2(32'hb91f62a1),
	.w3(32'h392dcafb),
	.w4(32'h393f4809),
	.w5(32'h39cee4a1),
	.w6(32'hb6980bee),
	.w7(32'hb88a373c),
	.w8(32'h38f190e0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98cbd62),
	.w1(32'hb8800062),
	.w2(32'h38ea311a),
	.w3(32'hb95478eb),
	.w4(32'h390851a0),
	.w5(32'hb69ca315),
	.w6(32'hb855143f),
	.w7(32'h38c536fd),
	.w8(32'h373544f8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39698b2f),
	.w1(32'hb7800cde),
	.w2(32'hb90054bd),
	.w3(32'h397f7f88),
	.w4(32'h391494b5),
	.w5(32'h38f900a3),
	.w6(32'h38c91405),
	.w7(32'h38a61287),
	.w8(32'h391faf45),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6658f73),
	.w1(32'h359092af),
	.w2(32'h36314414),
	.w3(32'hb6f8690a),
	.w4(32'hb57a6063),
	.w5(32'h35d61227),
	.w6(32'hb64dc532),
	.w7(32'h3669c15c),
	.w8(32'h369a2b0f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h343798f0),
	.w1(32'h35d8513b),
	.w2(32'h360ed39c),
	.w3(32'h362bdc13),
	.w4(32'h363e000b),
	.w5(32'h35a8c03f),
	.w6(32'h365d22cd),
	.w7(32'h3652b69b),
	.w8(32'h35cdf858),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb573ca52),
	.w1(32'h368a98f5),
	.w2(32'hb68f3f52),
	.w3(32'h357b0b71),
	.w4(32'h365eb006),
	.w5(32'hb6adb314),
	.w6(32'h36fc1d32),
	.w7(32'hb5a652e0),
	.w8(32'hb659a289),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89588a8),
	.w1(32'hb73bc239),
	.w2(32'hb8166ecc),
	.w3(32'hb7cf4208),
	.w4(32'hb7962dd0),
	.w5(32'hb81ddb6d),
	.w6(32'h379b9acc),
	.w7(32'h37fa63cf),
	.w8(32'hb7782595),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981b742),
	.w1(32'h3904e666),
	.w2(32'h39992a07),
	.w3(32'hb9a65c54),
	.w4(32'hb8bbb7db),
	.w5(32'h387c0dc1),
	.w6(32'hb8e7cc3f),
	.w7(32'hb7818b93),
	.w8(32'hb84d6bb8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8189851),
	.w1(32'hb8327d53),
	.w2(32'hb6aac9a7),
	.w3(32'hb6a18689),
	.w4(32'hb74d4a06),
	.w5(32'h38004423),
	.w6(32'hb8382298),
	.w7(32'hb81c4950),
	.w8(32'hb7b95262),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992b1f0),
	.w1(32'h39201265),
	.w2(32'h3960d2ff),
	.w3(32'hba0caf76),
	.w4(32'hb8c98c97),
	.w5(32'h39ec14c4),
	.w6(32'hb94b182f),
	.w7(32'hb9079c94),
	.w8(32'h39605b67),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca5512),
	.w1(32'h38be5973),
	.w2(32'hb9243650),
	.w3(32'h39304146),
	.w4(32'h38e2c9bf),
	.w5(32'h39bbdf81),
	.w6(32'hb8dd96b5),
	.w7(32'h36db6d4e),
	.w8(32'h39042bef),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb46db),
	.w1(32'hb8e050d7),
	.w2(32'hb8ce85d8),
	.w3(32'hb924335b),
	.w4(32'hb85c2b6e),
	.w5(32'hb93a5bb5),
	.w6(32'hb8bef662),
	.w7(32'hb8d78e91),
	.w8(32'hb8d0fb81),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0de3b1),
	.w1(32'hb8d480cf),
	.w2(32'h399c40fa),
	.w3(32'h396f1cdc),
	.w4(32'h394e47a2),
	.w5(32'h3a0083c9),
	.w6(32'hba0ea4eb),
	.w7(32'hba7a92ff),
	.w8(32'h3835169f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98cb937),
	.w1(32'h396a3e0a),
	.w2(32'h38d47874),
	.w3(32'hb9350931),
	.w4(32'hb803e803),
	.w5(32'hb9405238),
	.w6(32'hb8a6c9ac),
	.w7(32'hb8ff7c1d),
	.w8(32'hb987e2f8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a069ca3),
	.w1(32'h394c451f),
	.w2(32'h3a1b2f70),
	.w3(32'hb8b955ca),
	.w4(32'h399290f5),
	.w5(32'h3a0cd048),
	.w6(32'hba24cadb),
	.w7(32'hb8cd675e),
	.w8(32'h3945a9f7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20cd4d),
	.w1(32'hb92cbfe2),
	.w2(32'h39622969),
	.w3(32'hb9f55c08),
	.w4(32'h389657c3),
	.w5(32'h3985fb18),
	.w6(32'hb9a28a63),
	.w7(32'hb9aa21e7),
	.w8(32'h372daac8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba185432),
	.w1(32'hb9622f51),
	.w2(32'hb8d1e7cd),
	.w3(32'hb9768d30),
	.w4(32'h37cd189d),
	.w5(32'hb8c2586e),
	.w6(32'hb7cbb944),
	.w7(32'h38b935c2),
	.w8(32'h39333422),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d18c8b),
	.w1(32'h3714956a),
	.w2(32'h378cef93),
	.w3(32'h36d611a5),
	.w4(32'h37871ac8),
	.w5(32'h36a81830),
	.w6(32'h373b18a7),
	.w7(32'h35d35610),
	.w8(32'hb70cce54),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3978b1a8),
	.w1(32'h3850e9ec),
	.w2(32'hb8adf25e),
	.w3(32'h3913c5f6),
	.w4(32'h399e1c62),
	.w5(32'h39a6e668),
	.w6(32'hb834c9d8),
	.w7(32'h38c6eb54),
	.w8(32'h396d3cbc),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f9435),
	.w1(32'hba02c771),
	.w2(32'hb9d2b4e9),
	.w3(32'h39b71c7c),
	.w4(32'h3934bee7),
	.w5(32'h398c12d5),
	.w6(32'hb9459553),
	.w7(32'hb9d925fa),
	.w8(32'hb938344a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4bbe5),
	.w1(32'h3a97872d),
	.w2(32'h3a124bfb),
	.w3(32'h3a0e27b7),
	.w4(32'h3911eb8d),
	.w5(32'h398a9b57),
	.w6(32'hb93f16f4),
	.w7(32'hb942195e),
	.w8(32'hb91b0da8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d8b0f),
	.w1(32'hb925fcb2),
	.w2(32'h391a2a6f),
	.w3(32'hba0f5387),
	.w4(32'hb97b4582),
	.w5(32'h371a9868),
	.w6(32'hb9d2e37b),
	.w7(32'hb8b1e569),
	.w8(32'hb922cba8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3e08f),
	.w1(32'hb88382f3),
	.w2(32'h38a6a4fb),
	.w3(32'hb9f8bd0e),
	.w4(32'hb9532d64),
	.w5(32'h38ac6576),
	.w6(32'hb8f280e9),
	.w7(32'hb8b3acb8),
	.w8(32'h37e3a3bf),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3931409b),
	.w1(32'h388fc0fc),
	.w2(32'hb9f14adf),
	.w3(32'h3a3a5449),
	.w4(32'h38a51d98),
	.w5(32'h3a176f18),
	.w6(32'hb9f3913a),
	.w7(32'hb9a7f299),
	.w8(32'hb9670e72),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37993697),
	.w1(32'h3785cd43),
	.w2(32'h388175d1),
	.w3(32'h3768b3d7),
	.w4(32'h38375501),
	.w5(32'h389d986d),
	.w6(32'h360548f2),
	.w7(32'h38161a75),
	.w8(32'h389ccff2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0220fe),
	.w1(32'h3a3ea195),
	.w2(32'hb865a89f),
	.w3(32'h3a7fafee),
	.w4(32'h3a146a59),
	.w5(32'h3a4b2a7e),
	.w6(32'hba63150b),
	.w7(32'hba018132),
	.w8(32'hb9f52e88),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79b9321),
	.w1(32'hb81414c3),
	.w2(32'hb8a81d84),
	.w3(32'h38432603),
	.w4(32'h391eae88),
	.w5(32'h38e91532),
	.w6(32'hb928ecd8),
	.w7(32'h3888f5fd),
	.w8(32'h38c3d305),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f28066),
	.w1(32'h37345e1f),
	.w2(32'h3825d571),
	.w3(32'hb6a8b6a9),
	.w4(32'h3719ec05),
	.w5(32'h3819a7b2),
	.w6(32'hb7a241d7),
	.w7(32'hb63b6e07),
	.w8(32'h379279d6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39202c80),
	.w1(32'h3928f809),
	.w2(32'h3a11c31a),
	.w3(32'hb9866d48),
	.w4(32'h3831a3e7),
	.w5(32'h38562372),
	.w6(32'hb8e009ab),
	.w7(32'h38678e5c),
	.w8(32'h38ba4cc7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d82c10),
	.w1(32'hb91b4454),
	.w2(32'hb9267c92),
	.w3(32'h392a29d7),
	.w4(32'h39151856),
	.w5(32'h3891ab0d),
	.w6(32'h385de9e2),
	.w7(32'h390a8280),
	.w8(32'h397920f0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf1975),
	.w1(32'hb91fc03c),
	.w2(32'hb7ebf59a),
	.w3(32'hb99450c9),
	.w4(32'hb8abe554),
	.w5(32'hb8378ed7),
	.w6(32'hb824485c),
	.w7(32'h36e7d85b),
	.w8(32'h3738662f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dcf9b1),
	.w1(32'h37436656),
	.w2(32'h385a62f6),
	.w3(32'hb95c9ffc),
	.w4(32'h37c0bff9),
	.w5(32'hb931af1a),
	.w6(32'h389ad2e2),
	.w7(32'h38e0c110),
	.w8(32'hb85057d4),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ed9092),
	.w1(32'h38d0bc06),
	.w2(32'h393ef1d0),
	.w3(32'hb8f33387),
	.w4(32'h38822896),
	.w5(32'h39082b47),
	.w6(32'hb9010fb9),
	.w7(32'hb898734b),
	.w8(32'hb8666337),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399515ec),
	.w1(32'h39cb1eb3),
	.w2(32'h397a1b6a),
	.w3(32'hba833372),
	.w4(32'hb97ca939),
	.w5(32'h3a23c32e),
	.w6(32'hba262dfc),
	.w7(32'hb971311f),
	.w8(32'h395a87f7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385610bb),
	.w1(32'h37d6caf8),
	.w2(32'h3a2187c0),
	.w3(32'hba0a58bc),
	.w4(32'h39856089),
	.w5(32'h3917a1da),
	.w6(32'hba2917d3),
	.w7(32'hb9df51e9),
	.w8(32'hb90131e6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92315f3),
	.w1(32'hb778175c),
	.w2(32'hb73ec4d5),
	.w3(32'hb95e6708),
	.w4(32'hb8a8e37b),
	.w5(32'hb791b501),
	.w6(32'hb7c46005),
	.w7(32'hb7c7f019),
	.w8(32'hb8327fa7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb711192f),
	.w1(32'hb63dcee5),
	.w2(32'hb6411088),
	.w3(32'hb724a545),
	.w4(32'hb6338a5a),
	.w5(32'hb67f5ee4),
	.w6(32'hb69cce22),
	.w7(32'hb679ab95),
	.w8(32'hb6513eee),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86ba7d4),
	.w1(32'h38c6c453),
	.w2(32'h38d9eb7e),
	.w3(32'hb94a6531),
	.w4(32'hb80d16eb),
	.w5(32'h3856c361),
	.w6(32'hb8ad6eb0),
	.w7(32'hb8b2ddb8),
	.w8(32'hb74082ec),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c932ea),
	.w1(32'h35b81e58),
	.w2(32'hb64fccdc),
	.w3(32'h357b11e7),
	.w4(32'h36175084),
	.w5(32'hb689af26),
	.w6(32'h3609a0e2),
	.w7(32'h3631c254),
	.w8(32'hb5097a0c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38067c04),
	.w1(32'h37ce741e),
	.w2(32'h37f599bb),
	.w3(32'h36655a80),
	.w4(32'hb6ce597e),
	.w5(32'h37bbc5a6),
	.w6(32'hb77b3b52),
	.w7(32'hb7683655),
	.w8(32'hb73c3bf8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944603e),
	.w1(32'hb6e79cfb),
	.w2(32'h37c444a5),
	.w3(32'hb9ab6a8d),
	.w4(32'hb8ff91e7),
	.w5(32'h378a9d68),
	.w6(32'hb753d553),
	.w7(32'hb84ca90d),
	.w8(32'hb815f886),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cde972),
	.w1(32'h37859ebd),
	.w2(32'h38931e7c),
	.w3(32'hb8b36fc3),
	.w4(32'h3784ce68),
	.w5(32'h3892b2af),
	.w6(32'hb8fe92c1),
	.w7(32'hb8582590),
	.w8(32'h382e4773),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936138c),
	.w1(32'hb9025e90),
	.w2(32'hb93e37db),
	.w3(32'h3951c386),
	.w4(32'h384f8643),
	.w5(32'h38e7723d),
	.w6(32'h38c8ec7a),
	.w7(32'hb834a6a0),
	.w8(32'h38902911),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbbe40),
	.w1(32'hb71ac8a3),
	.w2(32'h3954e111),
	.w3(32'hb9f1d163),
	.w4(32'hb92f0b9e),
	.w5(32'hb8c83b24),
	.w6(32'hb97950ce),
	.w7(32'hb91f153a),
	.w8(32'hb867b032),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363b6ae1),
	.w1(32'hb474e71f),
	.w2(32'hb5464412),
	.w3(32'hb521026e),
	.w4(32'hb4f7ae7b),
	.w5(32'h35aaa762),
	.w6(32'h366aaff5),
	.w7(32'hb5e124f3),
	.w8(32'hb59c2d01),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d392b5),
	.w1(32'hb52e93fb),
	.w2(32'h37181fd1),
	.w3(32'hb7c03252),
	.w4(32'hb6ceac95),
	.w5(32'h3705bd62),
	.w6(32'hb78caaaf),
	.w7(32'hb735c2f8),
	.w8(32'h36a8f166),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f30131),
	.w1(32'h3613bdbf),
	.w2(32'hb5ced0b5),
	.w3(32'h365351d2),
	.w4(32'h3623bee5),
	.w5(32'hb6051e94),
	.w6(32'h363c8e71),
	.w7(32'hb49ed631),
	.w8(32'hb278c1d2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb829f866),
	.w1(32'hb943dbad),
	.w2(32'hb90fb6f2),
	.w3(32'hb7f6d5e4),
	.w4(32'hb98631de),
	.w5(32'hb92e2331),
	.w6(32'hb9525679),
	.w7(32'hb98bc324),
	.w8(32'hb88ffe4b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b285bc2),
	.w1(32'h3aa6e463),
	.w2(32'h39de7368),
	.w3(32'hb90aaa95),
	.w4(32'h389ea0ae),
	.w5(32'h3aeb33a4),
	.w6(32'hbabbeddf),
	.w7(32'hba04e43c),
	.w8(32'h3a794544),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386baf9a),
	.w1(32'hb8351c3a),
	.w2(32'hb9be295c),
	.w3(32'h39170637),
	.w4(32'h3a306c3d),
	.w5(32'h39a7d41c),
	.w6(32'hb9af1431),
	.w7(32'hb9624d0c),
	.w8(32'hb95035dd),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb749733a),
	.w1(32'hb9d5feb7),
	.w2(32'hb9be760f),
	.w3(32'hb8971eec),
	.w4(32'hb986f317),
	.w5(32'hb9c18fbd),
	.w6(32'hb99064f4),
	.w7(32'hb9c9f52d),
	.w8(32'hb9a120c3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b145e),
	.w1(32'hb966a4b9),
	.w2(32'hb98701a8),
	.w3(32'hba0d9844),
	.w4(32'hb9ab083a),
	.w5(32'hb95c7b4b),
	.w6(32'hb9bb8f41),
	.w7(32'hb9d1568e),
	.w8(32'hb9ce6133),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19cc85),
	.w1(32'hba4c9691),
	.w2(32'hba39c457),
	.w3(32'hb9dbff96),
	.w4(32'hb9e6d717),
	.w5(32'hb9a3efd9),
	.w6(32'hb9b9e4d4),
	.w7(32'hb94e9998),
	.w8(32'hb94d8adc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba095306),
	.w1(32'hb97b7205),
	.w2(32'h38e9e10f),
	.w3(32'hb9bdb0dd),
	.w4(32'hb9a998f7),
	.w5(32'hb9028642),
	.w6(32'hb975ecb1),
	.w7(32'h3917c04a),
	.w8(32'h385e93e4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ca28c),
	.w1(32'hb996f922),
	.w2(32'h38ac490b),
	.w3(32'hba082b0d),
	.w4(32'h35956756),
	.w5(32'hb908c92c),
	.w6(32'hb9b18d2a),
	.w7(32'hb9928ed5),
	.w8(32'hb9477564),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ae32ec),
	.w1(32'hba1b2429),
	.w2(32'hba31519e),
	.w3(32'h39a743d8),
	.w4(32'hb7fb49a5),
	.w5(32'hb754a940),
	.w6(32'hb9587135),
	.w7(32'hb990739e),
	.w8(32'h38a025c7),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fcceb8),
	.w1(32'h37d11d1d),
	.w2(32'h38acb500),
	.w3(32'hb9b06e9c),
	.w4(32'h37bab0f7),
	.w5(32'h3850ffc3),
	.w6(32'hb8aec44a),
	.w7(32'hb8037cc4),
	.w8(32'h38c81ec8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39637ce1),
	.w1(32'hb879b10b),
	.w2(32'hb7a146a5),
	.w3(32'h38c57cf8),
	.w4(32'hb8b0033c),
	.w5(32'hb903cca8),
	.w6(32'hba12bd80),
	.w7(32'hb9edfb6c),
	.w8(32'hb83c8cea),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e72fb7),
	.w1(32'h370ff624),
	.w2(32'hb9e30fbb),
	.w3(32'h399bfb30),
	.w4(32'h38a5724b),
	.w5(32'h38f11289),
	.w6(32'hb92176af),
	.w7(32'hb946cd37),
	.w8(32'hb80d517c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a9e80),
	.w1(32'hb89dc414),
	.w2(32'hb81ff364),
	.w3(32'hba522707),
	.w4(32'hb9d96846),
	.w5(32'h395892a2),
	.w6(32'hb9afa040),
	.w7(32'hb9840396),
	.w8(32'hb991017b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb965b0d0),
	.w1(32'hb9a77b81),
	.w2(32'hb9da1c92),
	.w3(32'h399ee2ad),
	.w4(32'hb9ed33ab),
	.w5(32'hb99aefbe),
	.w6(32'hb9cc9551),
	.w7(32'hb9b582e0),
	.w8(32'hb9145792),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8da37),
	.w1(32'hb917d9c5),
	.w2(32'hb903cf42),
	.w3(32'hba222221),
	.w4(32'hb8b90878),
	.w5(32'hb8b2a052),
	.w6(32'hb92ee2fd),
	.w7(32'hb8c354ac),
	.w8(32'hb8bedf32),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba268ed8),
	.w1(32'h39ee3794),
	.w2(32'h398bf72b),
	.w3(32'hb9e9ac04),
	.w4(32'h39d3d22f),
	.w5(32'h39677e73),
	.w6(32'h390fb5ec),
	.w7(32'h3993f144),
	.w8(32'h390ec121),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f165bf),
	.w1(32'hb9a2cbf2),
	.w2(32'hba1f82f8),
	.w3(32'h3a1b043d),
	.w4(32'hb9d9e411),
	.w5(32'hb8ec516e),
	.w6(32'hba0407ec),
	.w7(32'hb8eb48a8),
	.w8(32'hb95591bf),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0fa89),
	.w1(32'hb8a6cb6d),
	.w2(32'hb903b0ae),
	.w3(32'hb9a143fe),
	.w4(32'hb871f64e),
	.w5(32'hb8ddd27f),
	.w6(32'hb8638d77),
	.w7(32'hb8d59616),
	.w8(32'h386ff781),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb800a1d0),
	.w1(32'h394c5095),
	.w2(32'h39a1a726),
	.w3(32'h376c1693),
	.w4(32'hb77ada65),
	.w5(32'h390e515d),
	.w6(32'h395807b0),
	.w7(32'h39aea9bd),
	.w8(32'h38b15c49),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f7abd7),
	.w1(32'hba3327e7),
	.w2(32'hba0c2fbd),
	.w3(32'hb85fc492),
	.w4(32'hb9d5efe0),
	.w5(32'hb9cbcaa3),
	.w6(32'hb9b26e01),
	.w7(32'hb9ca135c),
	.w8(32'hb9c337c6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1af519),
	.w1(32'hb9001ee8),
	.w2(32'h3921ea98),
	.w3(32'hba0f80a6),
	.w4(32'hb991562a),
	.w5(32'hb8169b38),
	.w6(32'hb94502f5),
	.w7(32'hb8f07a98),
	.w8(32'hb96e6938),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38674b31),
	.w1(32'hb8159007),
	.w2(32'hb960070a),
	.w3(32'h37dba628),
	.w4(32'h38c553c1),
	.w5(32'hb83fbd39),
	.w6(32'hb9164065),
	.w7(32'hb86796ce),
	.w8(32'h381ee391),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900640a),
	.w1(32'hb933bdd4),
	.w2(32'hb9138e8d),
	.w3(32'hb90ed131),
	.w4(32'hb98ef2bf),
	.w5(32'hb9a298e0),
	.w6(32'hb9751578),
	.w7(32'hb997bd58),
	.w8(32'hb80454ea),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d95467),
	.w1(32'hba124785),
	.w2(32'hba931687),
	.w3(32'hb6d9eb7d),
	.w4(32'hb88e13fb),
	.w5(32'hb93f2736),
	.w6(32'hb9eddbb2),
	.w7(32'hba246df2),
	.w8(32'hba54b9c6),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b8674),
	.w1(32'h3864da46),
	.w2(32'h38d5fb20),
	.w3(32'hb76ab26a),
	.w4(32'h38ab4c09),
	.w5(32'hb8417564),
	.w6(32'h39b0f223),
	.w7(32'h3944bfa5),
	.w8(32'h39820ee3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979ebc5),
	.w1(32'h3644ac18),
	.w2(32'hb92f36b8),
	.w3(32'h397024b4),
	.w4(32'h38e98f94),
	.w5(32'h3921aaab),
	.w6(32'hb9310355),
	.w7(32'hba0e7c80),
	.w8(32'hb8b67dc0),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba238b62),
	.w1(32'hb98c2899),
	.w2(32'h383a2cca),
	.w3(32'hb9bf9f7b),
	.w4(32'hb9b41fea),
	.w5(32'hba2be463),
	.w6(32'h37fbb642),
	.w7(32'h39c4f2fa),
	.w8(32'hb913f08c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a14079),
	.w1(32'h396b5ed5),
	.w2(32'h39b1204f),
	.w3(32'hb9eeb1ae),
	.w4(32'hb93a47fb),
	.w5(32'h38a90e21),
	.w6(32'hb99a3dd5),
	.w7(32'hb9283d17),
	.w8(32'hb8b01899),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89b6931),
	.w1(32'hb94a243b),
	.w2(32'hb933b4aa),
	.w3(32'hb9c4fb47),
	.w4(32'hb93eb04d),
	.w5(32'hb9382d38),
	.w6(32'hb95f672d),
	.w7(32'hb9567eb2),
	.w8(32'hb8d55eb9),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fcfaa4),
	.w1(32'hb9a85b65),
	.w2(32'hb9815241),
	.w3(32'hba0c02ac),
	.w4(32'hb9b159eb),
	.w5(32'hb95686f9),
	.w6(32'hb95985ef),
	.w7(32'hb8f07da4),
	.w8(32'hb8e1826a),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cab5df),
	.w1(32'hb891d091),
	.w2(32'h391900aa),
	.w3(32'hb9b8e549),
	.w4(32'hb95daba6),
	.w5(32'hb9301bfe),
	.w6(32'hb958de9e),
	.w7(32'hb8c345c7),
	.w8(32'hb973d369),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebc629),
	.w1(32'h38701f2d),
	.w2(32'h387f2473),
	.w3(32'hb9fd7d51),
	.w4(32'hb8c6bc32),
	.w5(32'hb7fcc027),
	.w6(32'h373576e3),
	.w7(32'hb8810b7e),
	.w8(32'hb901b156),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3842f3c2),
	.w1(32'hb8ab2b17),
	.w2(32'hb8fa8f29),
	.w3(32'h3786efb3),
	.w4(32'hb8a1d68f),
	.w5(32'hb9091d5b),
	.w6(32'hb90012df),
	.w7(32'hb9511e42),
	.w8(32'hb871e9f4),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82bfede),
	.w1(32'hb94d0a95),
	.w2(32'hb938749b),
	.w3(32'hb83a41c5),
	.w4(32'hb93812fc),
	.w5(32'hb95717cc),
	.w6(32'hb944693a),
	.w7(32'hb980993f),
	.w8(32'hb92e452d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b748f),
	.w1(32'h3a03a563),
	.w2(32'h3a10a17c),
	.w3(32'h37e0b160),
	.w4(32'h39d02a42),
	.w5(32'h3a113a93),
	.w6(32'hb6b776af),
	.w7(32'h394ee437),
	.w8(32'h37cfc9c3),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3851fea9),
	.w1(32'h398b95f3),
	.w2(32'h3a1bf5c4),
	.w3(32'h39585fe0),
	.w4(32'h39f2797c),
	.w5(32'h3a284897),
	.w6(32'h395c6b33),
	.w7(32'h399eb319),
	.w8(32'h38ee9bb3),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a83970),
	.w1(32'hb9f96213),
	.w2(32'hb984b628),
	.w3(32'hb9e3f0bc),
	.w4(32'hba01f4fc),
	.w5(32'hb988ca31),
	.w6(32'hb9e6efc5),
	.w7(32'hb9ad5b62),
	.w8(32'hb9cad1b5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0b9e0),
	.w1(32'hb96e2eaf),
	.w2(32'hb959bbb7),
	.w3(32'hb9f13c84),
	.w4(32'hb987f5e7),
	.w5(32'hb98239f7),
	.w6(32'hb93e32c4),
	.w7(32'hb9926f95),
	.w8(32'hb914ba64),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb976df77),
	.w1(32'hba5a4b80),
	.w2(32'hba0e4984),
	.w3(32'hb7e4160b),
	.w4(32'hba14f50d),
	.w5(32'h3629d174),
	.w6(32'hb9f4b160),
	.w7(32'hb88511a7),
	.w8(32'h39a32a9b),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9764086),
	.w1(32'hb998b357),
	.w2(32'hb98b75f7),
	.w3(32'hb9b6f4b5),
	.w4(32'hb9540238),
	.w5(32'hb9789974),
	.w6(32'hb950b821),
	.w7(32'hb9802198),
	.w8(32'hb98c9e1c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f1440),
	.w1(32'hb8a0a0fd),
	.w2(32'hb8f2ceac),
	.w3(32'hb9634d79),
	.w4(32'hb8251dc7),
	.w5(32'hb863d5a8),
	.w6(32'hb8cfe2fe),
	.w7(32'hb91d2da9),
	.w8(32'h37aee2c0),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9464d57),
	.w1(32'hb96da605),
	.w2(32'hb8992d34),
	.w3(32'hb91abf92),
	.w4(32'hb999d3bf),
	.w5(32'hb94d55ad),
	.w6(32'hb9b5d4b1),
	.w7(32'hb953f299),
	.w8(32'hb918055a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1f40f),
	.w1(32'h399dcfab),
	.w2(32'hb943b449),
	.w3(32'h38fbd770),
	.w4(32'h391e5164),
	.w5(32'h39990d55),
	.w6(32'hb8595335),
	.w7(32'h356ca1fc),
	.w8(32'h35b910cb),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab96ba),
	.w1(32'hb9323a7e),
	.w2(32'hb7d59092),
	.w3(32'hb91d893a),
	.w4(32'hb96af680),
	.w5(32'hb8b127d0),
	.w6(32'hb917741e),
	.w7(32'hb7950504),
	.w8(32'hb89fa9dd),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b6a7b),
	.w1(32'hb9badeed),
	.w2(32'hb9867a9b),
	.w3(32'hba07e396),
	.w4(32'hb97fd5cd),
	.w5(32'hb98fda4a),
	.w6(32'hb97e17e4),
	.w7(32'hb93cf1c0),
	.w8(32'hb9704ce1),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1bfb0),
	.w1(32'h39623c0b),
	.w2(32'h39289e24),
	.w3(32'hb991aecf),
	.w4(32'h3a5b72d0),
	.w5(32'h39b2c0f5),
	.w6(32'h39fe06c9),
	.w7(32'h39bd3c1d),
	.w8(32'h39b1abbc),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fdae0a),
	.w1(32'hb93d581f),
	.w2(32'h39b07a56),
	.w3(32'h38d134fc),
	.w4(32'h3a5144de),
	.w5(32'h39064cbb),
	.w6(32'h3898587f),
	.w7(32'h3a040a2f),
	.w8(32'h3739b88d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c79563),
	.w1(32'h3901bcbf),
	.w2(32'h3980b713),
	.w3(32'h39ceddb4),
	.w4(32'h39475638),
	.w5(32'h39d4b8d2),
	.w6(32'hb9a462d2),
	.w7(32'hb99ca3af),
	.w8(32'hb402b408),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3909f01f),
	.w1(32'hba0a1fcd),
	.w2(32'hba80b4ac),
	.w3(32'h399c3d5b),
	.w4(32'hb98efde2),
	.w5(32'hb98d86be),
	.w6(32'hb9bd6380),
	.w7(32'hb932493e),
	.w8(32'hb93e0d8e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39dfc7),
	.w1(32'h3889adcd),
	.w2(32'h39531e97),
	.w3(32'hba08fd60),
	.w4(32'h370fa6ce),
	.w5(32'h391013a7),
	.w6(32'h38981570),
	.w7(32'h3934f6e4),
	.w8(32'hb8adec80),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920f2b3),
	.w1(32'hb9b98cf6),
	.w2(32'hb981b00d),
	.w3(32'hb9606985),
	.w4(32'hb8b3afa4),
	.w5(32'hb93e5ac7),
	.w6(32'hb9b7225b),
	.w7(32'hb9b906ce),
	.w8(32'hb97262a3),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a09a4a),
	.w1(32'h3954af9c),
	.w2(32'h3948e651),
	.w3(32'hb98f274e),
	.w4(32'h397b0fd3),
	.w5(32'h39829433),
	.w6(32'h38e0d8f3),
	.w7(32'h38fbf2a4),
	.w8(32'h39770363),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936e014),
	.w1(32'hb92b0509),
	.w2(32'hb91714da),
	.w3(32'h39a04ec0),
	.w4(32'hb828f251),
	.w5(32'h374b39df),
	.w6(32'hb76dc793),
	.w7(32'hb80d9d7d),
	.w8(32'h3838e275),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91af028),
	.w1(32'h3993efd8),
	.w2(32'h37c934a5),
	.w3(32'h38cd0fd3),
	.w4(32'h38b807dd),
	.w5(32'hb520cffa),
	.w6(32'h39076d58),
	.w7(32'hb707f9e9),
	.w8(32'hb82e18e3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72cd7da),
	.w1(32'hb9381487),
	.w2(32'h397df933),
	.w3(32'hb967dde9),
	.w4(32'h3806126f),
	.w5(32'hb92cf325),
	.w6(32'hb957970f),
	.w7(32'hb9791f81),
	.w8(32'hb8a34ad4),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8967214),
	.w1(32'hba153a2e),
	.w2(32'hb88f8a72),
	.w3(32'hb6dbf7c0),
	.w4(32'hba2c87dd),
	.w5(32'hb99ba5b4),
	.w6(32'hb9d6ad42),
	.w7(32'hb914b7e5),
	.w8(32'hb99a9ce5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91dcce4),
	.w1(32'hb9227876),
	.w2(32'h38497e33),
	.w3(32'hb985863b),
	.w4(32'hb8d9abf1),
	.w5(32'hb832b87c),
	.w6(32'hb8e0280c),
	.w7(32'h37900b6a),
	.w8(32'hb8a5205b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97fe381),
	.w1(32'h391996ad),
	.w2(32'h39c4f232),
	.w3(32'hba03dd48),
	.w4(32'hb8cbfccf),
	.w5(32'h38149494),
	.w6(32'hb9529ffd),
	.w7(32'h39326ec3),
	.w8(32'h396cfe81),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993ecee),
	.w1(32'h3975790e),
	.w2(32'h3a47578d),
	.w3(32'h38886c09),
	.w4(32'h39f4955c),
	.w5(32'h39b1741d),
	.w6(32'hb9b4a749),
	.w7(32'hb979774c),
	.w8(32'hb88bcbaf),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15d2c9),
	.w1(32'h3990cd66),
	.w2(32'hb71c8874),
	.w3(32'h3a38510d),
	.w4(32'hb9f04511),
	.w5(32'h394af095),
	.w6(32'hb9e4e032),
	.w7(32'hb941ab22),
	.w8(32'hb9311c3e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f67050),
	.w1(32'hb9b06ded),
	.w2(32'hb970b99a),
	.w3(32'hb8f82497),
	.w4(32'hb98a5497),
	.w5(32'hb968bb87),
	.w6(32'hb9962eb8),
	.w7(32'hb98aa90f),
	.w8(32'hb98cd8be),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9083588),
	.w1(32'hb923a8bc),
	.w2(32'hb9fde817),
	.w3(32'h38b9537e),
	.w4(32'h3a11ebd0),
	.w5(32'h39c8258d),
	.w6(32'hb7dffcca),
	.w7(32'h399c8dbb),
	.w8(32'h39c2a46a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6f785),
	.w1(32'hba859638),
	.w2(32'h3850c521),
	.w3(32'hba5594d6),
	.w4(32'hb97aeb28),
	.w5(32'hba565eeb),
	.w6(32'hb9849f86),
	.w7(32'hb88737fd),
	.w8(32'hb9bcf867),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb965785a),
	.w1(32'h392c8390),
	.w2(32'h38fce05f),
	.w3(32'hb8620993),
	.w4(32'h39df0bdd),
	.w5(32'h3a0564dc),
	.w6(32'h3840c694),
	.w7(32'hb7fed2d4),
	.w8(32'h3846f7d8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396758f5),
	.w1(32'h3951a2d1),
	.w2(32'h39ce93a6),
	.w3(32'h39944f91),
	.w4(32'h39984641),
	.w5(32'h3999e9c1),
	.w6(32'hb9543ec5),
	.w7(32'h38f59c94),
	.w8(32'h35feb513),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398488d2),
	.w1(32'h3852b393),
	.w2(32'hb88cacaa),
	.w3(32'h394efdb6),
	.w4(32'h398e9a7f),
	.w5(32'h390a4701),
	.w6(32'h394d0e5b),
	.w7(32'h38caf88f),
	.w8(32'h384ce45c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88d3cb8),
	.w1(32'hb832b60f),
	.w2(32'hb93c3c37),
	.w3(32'h390e9097),
	.w4(32'hb866d624),
	.w5(32'hb8eae759),
	.w6(32'h37ee5b84),
	.w7(32'hb9009ee2),
	.w8(32'hb93b7e49),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfc599),
	.w1(32'h39d840f6),
	.w2(32'h39ce1d3a),
	.w3(32'h396a6d79),
	.w4(32'h39b420aa),
	.w5(32'h3a520337),
	.w6(32'hb6a3041f),
	.w7(32'h39dfca17),
	.w8(32'h39d4f1a6),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39942c3c),
	.w1(32'hb89b677a),
	.w2(32'hb9356dff),
	.w3(32'h3981154a),
	.w4(32'hb8eba7e8),
	.w5(32'hb8d05519),
	.w6(32'hb91afd41),
	.w7(32'hb8b6fcd9),
	.w8(32'hb8c3fbf5),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f42812),
	.w1(32'h390e13d4),
	.w2(32'h39586dd5),
	.w3(32'hba19b1c9),
	.w4(32'h3803fb5e),
	.w5(32'h3911db79),
	.w6(32'hb8fe9aa9),
	.w7(32'h37d99d02),
	.w8(32'h394901e9),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a5f5a),
	.w1(32'hb8e5ba99),
	.w2(32'hb8605994),
	.w3(32'hb99a1e87),
	.w4(32'hb846d3ae),
	.w5(32'hb7f9b6e3),
	.w6(32'hb84b9200),
	.w7(32'hb8fe543d),
	.w8(32'h38509176),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945e5bd),
	.w1(32'h39bc901b),
	.w2(32'h398273cf),
	.w3(32'h39916161),
	.w4(32'h3a043759),
	.w5(32'h3a207187),
	.w6(32'h39827624),
	.w7(32'h39cbe6bc),
	.w8(32'h3a130533),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ddd2a),
	.w1(32'hb9ae1b5a),
	.w2(32'hb97047f7),
	.w3(32'h3a07ece3),
	.w4(32'hb98386e3),
	.w5(32'hb94bae44),
	.w6(32'hb970b964),
	.w7(32'hb99a06c1),
	.w8(32'hb9a7a759),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b48361),
	.w1(32'hb90c7981),
	.w2(32'hb8d14919),
	.w3(32'hb9890710),
	.w4(32'hb8c11f65),
	.w5(32'hb8448b88),
	.w6(32'hb8df2010),
	.w7(32'hb9180609),
	.w8(32'hb816e734),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b1c7f),
	.w1(32'hb9456654),
	.w2(32'h38996712),
	.w3(32'hb9986d99),
	.w4(32'hb9c4061e),
	.w5(32'h37e4a4f7),
	.w6(32'hba53b10f),
	.w7(32'hba2596b4),
	.w8(32'hb9558496),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8977a07),
	.w1(32'hb99eb58f),
	.w2(32'hb996cf1a),
	.w3(32'hb71f7884),
	.w4(32'hb989f235),
	.w5(32'hb9a54a95),
	.w6(32'hb96976cf),
	.w7(32'hb99ff6ed),
	.w8(32'hb92b1721),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f97cb4),
	.w1(32'hb98348d9),
	.w2(32'hb993c92a),
	.w3(32'hb9133c16),
	.w4(32'hb8d3b8ae),
	.w5(32'hb937898e),
	.w6(32'hb9a660e8),
	.w7(32'hb90bc372),
	.w8(32'hb9051bf1),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba476612),
	.w1(32'hb9953857),
	.w2(32'hb84a27c9),
	.w3(32'hba623c93),
	.w4(32'hba25a4ed),
	.w5(32'hb953a063),
	.w6(32'hba1046ac),
	.w7(32'hb9b3fbe1),
	.w8(32'hb9d54bb8),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22b233),
	.w1(32'h39973f6a),
	.w2(32'h39ad1c6e),
	.w3(32'hba2a86b6),
	.w4(32'h3982731f),
	.w5(32'h39b3a40b),
	.w6(32'h3895a110),
	.w7(32'h384c95cf),
	.w8(32'h39858aaf),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d199c),
	.w1(32'hb9259c8b),
	.w2(32'hb8969963),
	.w3(32'h39b7261a),
	.w4(32'hb92b08e3),
	.w5(32'hb95752b6),
	.w6(32'hb983a318),
	.w7(32'hb92d36ff),
	.w8(32'hb9b6328a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47a051),
	.w1(32'hb81e1497),
	.w2(32'h3a193123),
	.w3(32'hba66cd73),
	.w4(32'h3838d113),
	.w5(32'h39a441cd),
	.w6(32'hb90eeb64),
	.w7(32'h399e2e68),
	.w8(32'h390a9753),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393bfba5),
	.w1(32'hb92b3248),
	.w2(32'hb92124cd),
	.w3(32'hb799a458),
	.w4(32'hb8dd94fa),
	.w5(32'hb9272152),
	.w6(32'hb997490d),
	.w7(32'hb969bf39),
	.w8(32'h383aae55),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c2900e),
	.w1(32'h36f0b6db),
	.w2(32'hb92078fc),
	.w3(32'h380c7a5d),
	.w4(32'h396a6c77),
	.w5(32'h38461c7a),
	.w6(32'h38e8091c),
	.w7(32'h384d06cc),
	.w8(32'h394745a4),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c92284),
	.w1(32'h397de9b6),
	.w2(32'h39839d42),
	.w3(32'h37305a78),
	.w4(32'h391cd409),
	.w5(32'h39139ee1),
	.w6(32'h3963e2d4),
	.w7(32'h38ddebe8),
	.w8(32'hb857f859),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65f711e),
	.w1(32'hb81ddc28),
	.w2(32'h37c27a47),
	.w3(32'hb7b1bde7),
	.w4(32'hb784ff49),
	.w5(32'hb8192fa6),
	.w6(32'h382b8b5c),
	.w7(32'h38a110d8),
	.w8(32'h3908dd1f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f779d0),
	.w1(32'h39d4e427),
	.w2(32'h39a0665b),
	.w3(32'hba000a18),
	.w4(32'hb9c74acf),
	.w5(32'h39b80625),
	.w6(32'hb9889f07),
	.w7(32'hb97e7eba),
	.w8(32'h3984feb2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83b9582),
	.w1(32'hb7eb7572),
	.w2(32'hb874a645),
	.w3(32'hb9b808ed),
	.w4(32'h3839eaf5),
	.w5(32'h3962ce6f),
	.w6(32'h38a023ae),
	.w7(32'h39112416),
	.w8(32'h3849503c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999b3fe),
	.w1(32'h3918a086),
	.w2(32'h39345f15),
	.w3(32'hba0961d1),
	.w4(32'hb902bc0d),
	.w5(32'h393868bf),
	.w6(32'hb88c745f),
	.w7(32'hb93a9ed1),
	.w8(32'hb8bf52fe),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2edbcb),
	.w1(32'hba2a4f89),
	.w2(32'hb9de7d74),
	.w3(32'h39a18d01),
	.w4(32'h3937b1c3),
	.w5(32'h3a66c53d),
	.w6(32'hb99ff51b),
	.w7(32'hba15cb27),
	.w8(32'hb842a991),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a49b22),
	.w1(32'hb8aa554c),
	.w2(32'hb6ec62e1),
	.w3(32'hb876c20d),
	.w4(32'hb900a39b),
	.w5(32'hb8b9687c),
	.w6(32'hb8dee89b),
	.w7(32'hb886c668),
	.w8(32'h39056708),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39696aec),
	.w1(32'h384b3a29),
	.w2(32'h3903fad8),
	.w3(32'hb95662b8),
	.w4(32'hb9509f32),
	.w5(32'h3883bb2a),
	.w6(32'hb98266d9),
	.w7(32'hb93dc2ed),
	.w8(32'hb920ddbd),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a7f99),
	.w1(32'h391ef72a),
	.w2(32'hba14b40e),
	.w3(32'h39856468),
	.w4(32'hb9768e80),
	.w5(32'h3948d79b),
	.w6(32'hb9582462),
	.w7(32'hb97ebed1),
	.w8(32'h399fe376),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0daf8f),
	.w1(32'h392a4e42),
	.w2(32'hb98331f0),
	.w3(32'h399b4f77),
	.w4(32'h39a6581e),
	.w5(32'h392f8b16),
	.w6(32'hb9821ac4),
	.w7(32'hb7d09a3d),
	.w8(32'h395a8b0c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19f9c4),
	.w1(32'h397d278b),
	.w2(32'hb966734f),
	.w3(32'h3a283605),
	.w4(32'h39370fe0),
	.w5(32'h37c1c969),
	.w6(32'h376f2367),
	.w7(32'hb904a080),
	.w8(32'hb8a4a454),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f21ef7),
	.w1(32'hb925a096),
	.w2(32'hb8832fa9),
	.w3(32'hb9cdf2e2),
	.w4(32'hb986fc1f),
	.w5(32'hb9a16d3d),
	.w6(32'hb9b8aa0b),
	.w7(32'hb9cc154b),
	.w8(32'hb9abdfef),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba145de5),
	.w1(32'hb82e9dd3),
	.w2(32'h39941017),
	.w3(32'hba278f03),
	.w4(32'hb907759b),
	.w5(32'hb9083375),
	.w6(32'hb8e96360),
	.w7(32'hb84f789a),
	.w8(32'h37f08430),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380262f0),
	.w1(32'hb986df56),
	.w2(32'hb92d6089),
	.w3(32'hb7d796c5),
	.w4(32'hb9a1880d),
	.w5(32'hb9a8de97),
	.w6(32'hb98d227f),
	.w7(32'hb98aa46f),
	.w8(32'hb97dc1df),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d474e),
	.w1(32'hb890ae17),
	.w2(32'hb91f7163),
	.w3(32'hb9917336),
	.w4(32'h387597e9),
	.w5(32'h3922047a),
	.w6(32'hb96534c9),
	.w7(32'hba0c0501),
	.w8(32'hba2824bd),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b81456),
	.w1(32'h389e0f34),
	.w2(32'h3807fa9b),
	.w3(32'h3786955e),
	.w4(32'h38847632),
	.w5(32'h38a6f3b7),
	.w6(32'hb84252b9),
	.w7(32'hb954503d),
	.w8(32'h39c90efb),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949ad1c),
	.w1(32'hb825d037),
	.w2(32'hb66dc081),
	.w3(32'hb80ab2b6),
	.w4(32'h3704c18a),
	.w5(32'hb7f748cf),
	.w6(32'hb8af125c),
	.w7(32'hb699d50d),
	.w8(32'h37c39107),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d82771),
	.w1(32'h3937ab54),
	.w2(32'h3932de13),
	.w3(32'h39b9762b),
	.w4(32'h399d6a77),
	.w5(32'h39f48b9b),
	.w6(32'hb8a91562),
	.w7(32'h39376e9b),
	.w8(32'h3927628b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b2f8ae),
	.w1(32'h3904d2c1),
	.w2(32'h39a77db3),
	.w3(32'hba178a9f),
	.w4(32'hb96be4c5),
	.w5(32'h39566db3),
	.w6(32'hb9fc63c1),
	.w7(32'hb91c5bd1),
	.w8(32'h396d1321),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d3e3c),
	.w1(32'hb805f015),
	.w2(32'h39391a0d),
	.w3(32'hb96afe0d),
	.w4(32'hb9acf20a),
	.w5(32'h39560d58),
	.w6(32'h38340e45),
	.w7(32'h39379d35),
	.w8(32'h39388a42),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393eaa04),
	.w1(32'hb962d386),
	.w2(32'hb9240dd1),
	.w3(32'h39807886),
	.w4(32'hb9192c51),
	.w5(32'h3710ac15),
	.w6(32'hb9930da0),
	.w7(32'hb9ad30a3),
	.w8(32'hba2ef45f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa14c34),
	.w1(32'h3a947f16),
	.w2(32'h39a56af9),
	.w3(32'h3a885351),
	.w4(32'h3a847bfe),
	.w5(32'h3a97889c),
	.w6(32'h38414c26),
	.w7(32'hb560d3c0),
	.w8(32'h39c2cce8),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8a3cb),
	.w1(32'hb9872e63),
	.w2(32'hb993bb61),
	.w3(32'h3a3b145d),
	.w4(32'hb909aecf),
	.w5(32'h37180d35),
	.w6(32'hb978e818),
	.w7(32'hb943f475),
	.w8(32'h38c83a61),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89f38d1),
	.w1(32'h3942a989),
	.w2(32'h38f7ed7a),
	.w3(32'hb789f6bd),
	.w4(32'h398e435b),
	.w5(32'h395b6401),
	.w6(32'h391cb2bd),
	.w7(32'h38d2f2fa),
	.w8(32'h395794e1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a246a67),
	.w1(32'hb8d2051c),
	.w2(32'hb928c1b1),
	.w3(32'h3a20a82a),
	.w4(32'hb840e47f),
	.w5(32'h37c0cd63),
	.w6(32'hb988ee3b),
	.w7(32'hb93ac366),
	.w8(32'h3866be5c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9186baa),
	.w1(32'hb96c489e),
	.w2(32'hb98312e3),
	.w3(32'hb91c7087),
	.w4(32'hb98598ee),
	.w5(32'hb988c5f6),
	.w6(32'hb99e5219),
	.w7(32'hb9c0961d),
	.w8(32'hb9f17891),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9a9b3),
	.w1(32'hb923aa7e),
	.w2(32'hb8c48234),
	.w3(32'hb9b0f32f),
	.w4(32'hb947463c),
	.w5(32'hb950368e),
	.w6(32'hb9338dbf),
	.w7(32'hb96ed330),
	.w8(32'hb895992b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c8d4cb),
	.w1(32'h398289a9),
	.w2(32'h393a6ff4),
	.w3(32'hb909a6b2),
	.w4(32'h39a332e1),
	.w5(32'h39891194),
	.w6(32'h394ad42b),
	.w7(32'h3910684e),
	.w8(32'h397c7b43),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961db5f),
	.w1(32'hb958f4f2),
	.w2(32'hb982928e),
	.w3(32'h39b85a06),
	.w4(32'hb8ea47f0),
	.w5(32'hb9c31d8a),
	.w6(32'hb972bd53),
	.w7(32'hb98e3a4f),
	.w8(32'hb9d60a1f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ad48c),
	.w1(32'hb93641b4),
	.w2(32'hb923d59f),
	.w3(32'hba29b470),
	.w4(32'hb987273f),
	.w5(32'hb95fc33c),
	.w6(32'hb999f02b),
	.w7(32'hb95eb0e1),
	.w8(32'hb909ef3d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13baab),
	.w1(32'hb92d6044),
	.w2(32'h39ae4b34),
	.w3(32'hb957b9a8),
	.w4(32'h3a4e9d0c),
	.w5(32'h395fab70),
	.w6(32'hb86f7860),
	.w7(32'h3960c413),
	.w8(32'h39a78c86),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45d68a),
	.w1(32'hb8fdbeb1),
	.w2(32'hb9c90c5f),
	.w3(32'h39acc428),
	.w4(32'h32d9afb6),
	.w5(32'hb8da7eaf),
	.w6(32'hb99e3760),
	.w7(32'hb8dc0e4f),
	.w8(32'h3886598f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91405b9),
	.w1(32'hba172343),
	.w2(32'hb9dca187),
	.w3(32'h3910cda4),
	.w4(32'hb8c76841),
	.w5(32'hb967e3e8),
	.w6(32'hb9be2995),
	.w7(32'hb8fe2cd8),
	.w8(32'hb8416310),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1a0f1),
	.w1(32'hb956f06b),
	.w2(32'hb85234fb),
	.w3(32'hb963f693),
	.w4(32'hb81bea8d),
	.w5(32'hb85b9392),
	.w6(32'hb995961b),
	.w7(32'hb93dc6ec),
	.w8(32'hb8f3eb49),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39183d43),
	.w1(32'h39ca84ac),
	.w2(32'h3992aadd),
	.w3(32'h389b0027),
	.w4(32'h39f676b4),
	.w5(32'h39f4bf06),
	.w6(32'h39381ac2),
	.w7(32'h391eb57f),
	.w8(32'h39d18746),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992d1b3),
	.w1(32'hb826f442),
	.w2(32'hb888bfa1),
	.w3(32'h39f98cd4),
	.w4(32'hb7e5b80e),
	.w5(32'hb86b4677),
	.w6(32'hb8390872),
	.w7(32'hb8a9ba50),
	.w8(32'hb7374e7c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8158d7a),
	.w1(32'hb8934bd1),
	.w2(32'hb8a0a462),
	.w3(32'h37469f55),
	.w4(32'hb8229079),
	.w5(32'hb86defb0),
	.w6(32'hb88b67d0),
	.w7(32'hb8b15e0a),
	.w8(32'h35b9f5b1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39107a5f),
	.w1(32'hb7c7dd0a),
	.w2(32'hb9900abd),
	.w3(32'h38399251),
	.w4(32'h39a24bd6),
	.w5(32'h38dd6f79),
	.w6(32'hba237d9e),
	.w7(32'hb9fdc478),
	.w8(32'hba29ba65),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8ed13),
	.w1(32'hb95b6fcf),
	.w2(32'hb7e3b4cb),
	.w3(32'hb8dd1109),
	.w4(32'hb90278ff),
	.w5(32'h380a77f5),
	.w6(32'hb907c6bc),
	.w7(32'h3721e6a5),
	.w8(32'hb633f676),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9726cee),
	.w1(32'hb93d1acc),
	.w2(32'hb7248b31),
	.w3(32'hb9328a1b),
	.w4(32'hb98c8e73),
	.w5(32'hb903a502),
	.w6(32'hb96eb239),
	.w7(32'hb9190c51),
	.w8(32'h370a6d2b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b64b12),
	.w1(32'h388611a8),
	.w2(32'h3968e0e5),
	.w3(32'hb8a172b0),
	.w4(32'h38a5d85a),
	.w5(32'h38963701),
	.w6(32'hb9534022),
	.w7(32'hb947f6f1),
	.w8(32'h39110100),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b45e70),
	.w1(32'hb7d02221),
	.w2(32'hb8963245),
	.w3(32'hb833916a),
	.w4(32'h3833848e),
	.w5(32'h36016444),
	.w6(32'hb878cbaa),
	.w7(32'hb9011aa1),
	.w8(32'h378f9422),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3776107e),
	.w1(32'hb989e178),
	.w2(32'hba6def58),
	.w3(32'h38e76d8e),
	.w4(32'hb6ab9880),
	.w5(32'hb95f9ede),
	.w6(32'hba0e2cbf),
	.w7(32'hba548c85),
	.w8(32'hba890817),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3486cf),
	.w1(32'hb9afa4be),
	.w2(32'hb9aef8a6),
	.w3(32'hb9bc854e),
	.w4(32'hb965f72a),
	.w5(32'hb9835323),
	.w6(32'hb901bb27),
	.w7(32'hb9b2e533),
	.w8(32'hb92cd562),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db7802),
	.w1(32'hb96b8ed7),
	.w2(32'h39e8faa8),
	.w3(32'hb9baa45d),
	.w4(32'h3a30ae1b),
	.w5(32'h38877ece),
	.w6(32'hba179060),
	.w7(32'hb7ffaee4),
	.w8(32'h395cf24d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7673666),
	.w1(32'h3bd595a1),
	.w2(32'h3b8e3fe6),
	.w3(32'hb7e3e17e),
	.w4(32'h3bff949d),
	.w5(32'h3bb1422a),
	.w6(32'h3bd7ecfd),
	.w7(32'h3ba24bd2),
	.w8(32'h3bbb3a6b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9911ee),
	.w1(32'hbc23e485),
	.w2(32'hbc3eecd8),
	.w3(32'h3bc0aa2c),
	.w4(32'hbbc9a689),
	.w5(32'hbbe18b41),
	.w6(32'hbc344e41),
	.w7(32'hbc465da2),
	.w8(32'hbc1418ce),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule