module layer_10_featuremap_336(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad5583),
	.w1(32'hbbb2ddd7),
	.w2(32'hbb9ca969),
	.w3(32'hbb900642),
	.w4(32'hbbaac38a),
	.w5(32'h3b2414ef),
	.w6(32'hbb6b824e),
	.w7(32'hbb9ce97b),
	.w8(32'h3ac5676c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c840025),
	.w1(32'h3bbc8902),
	.w2(32'h3c228cbb),
	.w3(32'h3c5088ac),
	.w4(32'hbb74f79d),
	.w5(32'hbacbb446),
	.w6(32'h3c68803a),
	.w7(32'hbb210bd7),
	.w8(32'h3bb06347),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84e0b3),
	.w1(32'hb8861188),
	.w2(32'hbaa00292),
	.w3(32'h3aac9725),
	.w4(32'h3adc6bb9),
	.w5(32'h3b8776cb),
	.w6(32'h3a7edcd1),
	.w7(32'h3a3f742a),
	.w8(32'h3b831ef7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b219b22),
	.w1(32'h3a9f3c18),
	.w2(32'hb8f80737),
	.w3(32'h3b7cf68c),
	.w4(32'h3b860dbd),
	.w5(32'h3b052faa),
	.w6(32'h3ae8c29c),
	.w7(32'h3a8e9d7e),
	.w8(32'hb9247dde),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995e58b),
	.w1(32'hbb371b12),
	.w2(32'hba6c0223),
	.w3(32'hbb6ca20d),
	.w4(32'hba091f24),
	.w5(32'h37e9a5bf),
	.w6(32'hbbaf2cd3),
	.w7(32'hbb7ba6f3),
	.w8(32'h3a7891c6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2df774),
	.w1(32'h3b3e7455),
	.w2(32'h3b007ba0),
	.w3(32'h3a08f4ce),
	.w4(32'h39256a64),
	.w5(32'h3a28e690),
	.w6(32'h3a5fe334),
	.w7(32'h3a061a70),
	.w8(32'h39dcf3c0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf9379),
	.w1(32'h3c4b4ca1),
	.w2(32'h3ca3e50e),
	.w3(32'h3b560cb4),
	.w4(32'h3c6eafb8),
	.w5(32'h3ca09d5b),
	.w6(32'hba21d5ca),
	.w7(32'h3c142abd),
	.w8(32'h3ca1e04e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c885da2),
	.w1(32'h3c1a950c),
	.w2(32'h3bb72d1d),
	.w3(32'h3ca80985),
	.w4(32'h3ca155c5),
	.w5(32'h3c73fb17),
	.w6(32'h3c95652f),
	.w7(32'h3b64113d),
	.w8(32'h3c3d1508),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ad0e4),
	.w1(32'hb9de19d3),
	.w2(32'h3a04945e),
	.w3(32'h3b539154),
	.w4(32'hba65b1d6),
	.w5(32'h3aa5aa7b),
	.w6(32'h3b971359),
	.w7(32'h3abc1251),
	.w8(32'h3b430777),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceb0b34),
	.w1(32'h3b9c8307),
	.w2(32'h3cd2f99e),
	.w3(32'h3ca4504b),
	.w4(32'hbb91fd26),
	.w5(32'h3c8f98f6),
	.w6(32'h3ca2b337),
	.w7(32'h3a7f186a),
	.w8(32'h3ccdb657),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c062f),
	.w1(32'h3b5bb650),
	.w2(32'h3aadb287),
	.w3(32'h3b7804bf),
	.w4(32'h3a0339ad),
	.w5(32'hba43d805),
	.w6(32'h3b65a533),
	.w7(32'h3a913d1c),
	.w8(32'h3a08745e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97d835),
	.w1(32'hbc3bb79a),
	.w2(32'h3beb9519),
	.w3(32'h3ba72283),
	.w4(32'hba74b572),
	.w5(32'h3c8df1d8),
	.w6(32'h3bcdef19),
	.w7(32'hbb9de20f),
	.w8(32'h3c97e7e7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb130cb),
	.w1(32'h3aab8e02),
	.w2(32'h3ce4795e),
	.w3(32'h3c4ac91e),
	.w4(32'h3b8de903),
	.w5(32'h3cb5dea2),
	.w6(32'h3bed6cc7),
	.w7(32'h3bb6166b),
	.w8(32'h3ccff234),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c309dbc),
	.w1(32'h3ba17e8a),
	.w2(32'h3bd71612),
	.w3(32'h3bb09fd6),
	.w4(32'h3ac7d163),
	.w5(32'h3bba83e6),
	.w6(32'h3b1d92a9),
	.w7(32'hbadf671f),
	.w8(32'h3be9436e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99925c),
	.w1(32'h3b825da9),
	.w2(32'h3c315f8c),
	.w3(32'h3c2ac483),
	.w4(32'hbbe68864),
	.w5(32'h399dd462),
	.w6(32'h3c8d8997),
	.w7(32'hb8d5c98f),
	.w8(32'h3c0cd9b6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc30f58),
	.w1(32'h3be28461),
	.w2(32'h3cab208c),
	.w3(32'h3c957eef),
	.w4(32'hbb929643),
	.w5(32'h3c206a3a),
	.w6(32'h3cc0b565),
	.w7(32'h3c18f545),
	.w8(32'h3cc23541),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72b95e),
	.w1(32'h3ac5830d),
	.w2(32'h3b24ceb5),
	.w3(32'h3b8e1a13),
	.w4(32'h3b2697f8),
	.w5(32'hba90ba90),
	.w6(32'h3b3b3e2b),
	.w7(32'h3a557f7e),
	.w8(32'hbb411888),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a4a3e),
	.w1(32'h3b3882e7),
	.w2(32'h3ca7f19e),
	.w3(32'h3c28c9d5),
	.w4(32'h3af1115d),
	.w5(32'h3ccb276b),
	.w6(32'h3c8096ed),
	.w7(32'h3b636a32),
	.w8(32'h3cb9c5b3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c206e3d),
	.w1(32'h3b8c0a7b),
	.w2(32'h3c7a718a),
	.w3(32'h3b63ea4b),
	.w4(32'h3b705191),
	.w5(32'h3c94be7c),
	.w6(32'h3bec7274),
	.w7(32'h3b906245),
	.w8(32'h3c90b399),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b0f5f),
	.w1(32'h3a9987ed),
	.w2(32'h3a9420f3),
	.w3(32'h389036b5),
	.w4(32'hbb370c77),
	.w5(32'h3b68e7e4),
	.w6(32'hb8bd2790),
	.w7(32'hbb2ccf2d),
	.w8(32'h3afe98d5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad448aa),
	.w1(32'h3b4d3561),
	.w2(32'hbad858f9),
	.w3(32'h3ad61d3c),
	.w4(32'hbae539dc),
	.w5(32'h3a884011),
	.w6(32'h3a6c5fe6),
	.w7(32'hbba16604),
	.w8(32'h3a80e189),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aade50b),
	.w1(32'hbbec8f90),
	.w2(32'h3b18904d),
	.w3(32'hba126848),
	.w4(32'hbc159a82),
	.w5(32'hba93de95),
	.w6(32'h3b91bc6b),
	.w7(32'hbbc6406b),
	.w8(32'h3a64dfd8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4ca822),
	.w1(32'h3bcef384),
	.w2(32'h3cb8b30b),
	.w3(32'h3d10b4c6),
	.w4(32'hbb18609a),
	.w5(32'h3c7e3d5f),
	.w6(32'h3d24b5fa),
	.w7(32'h3c5587e9),
	.w8(32'h3d2bc403),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce2e73c),
	.w1(32'hbace01cd),
	.w2(32'h3c91158b),
	.w3(32'h3c786c3c),
	.w4(32'hbc6cf600),
	.w5(32'h3c069f35),
	.w6(32'h3c9c30d1),
	.w7(32'hbbed1b78),
	.w8(32'h3c976b2b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d28d5ce),
	.w1(32'hba9d5441),
	.w2(32'h3c7b3dc5),
	.w3(32'h3d016acf),
	.w4(32'hbc61c4d7),
	.w5(32'h3b314c1c),
	.w6(32'h3d31fada),
	.w7(32'hbbb709f9),
	.w8(32'h3c47a1bf),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b518894),
	.w1(32'h3b4f91d3),
	.w2(32'h3a881914),
	.w3(32'h3b6cbe04),
	.w4(32'h3b676d85),
	.w5(32'h3b0ee257),
	.w6(32'h3b9331a5),
	.w7(32'h3b5d0093),
	.w8(32'h3b258566),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a088a5b),
	.w1(32'hba72ccc7),
	.w2(32'hba07af74),
	.w3(32'hba1bc87c),
	.w4(32'hba04b7df),
	.w5(32'hbb89742f),
	.w6(32'hb9d5ea9f),
	.w7(32'hb936fc9a),
	.w8(32'hbb8f3c24),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ff328),
	.w1(32'hbc566fd2),
	.w2(32'h3ad8f199),
	.w3(32'hbae1d568),
	.w4(32'hbc48f370),
	.w5(32'hbc514449),
	.w6(32'h3aa51af5),
	.w7(32'hbb83460b),
	.w8(32'hb9617d18),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b683bc9),
	.w1(32'hbbad0779),
	.w2(32'hbb648375),
	.w3(32'h3bfc2a4e),
	.w4(32'hbbe80522),
	.w5(32'hbbbf459c),
	.w6(32'h3c20b254),
	.w7(32'hbb8ccca5),
	.w8(32'hbb35e1bc),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c859340),
	.w1(32'hbbe0e5e1),
	.w2(32'h3bab405b),
	.w3(32'h3c88f60c),
	.w4(32'hbbd4abe7),
	.w5(32'hbae6370e),
	.w6(32'h3c9d2868),
	.w7(32'hbb5e6b60),
	.w8(32'h3c0fdcef),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00efd4),
	.w1(32'h3a3f653d),
	.w2(32'h3aa09cfd),
	.w3(32'hbb396f1a),
	.w4(32'hba925433),
	.w5(32'hb7d331d3),
	.w6(32'h370b82bc),
	.w7(32'hb909c977),
	.w8(32'h3aea06b4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a042ea7),
	.w1(32'hb9dc9544),
	.w2(32'hb971cfb0),
	.w3(32'h39e5c709),
	.w4(32'h3adb54d8),
	.w5(32'hba38ba8d),
	.w6(32'h3b1798cf),
	.w7(32'h39fe14a2),
	.w8(32'hba25a11b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff5a91),
	.w1(32'hb8c1b201),
	.w2(32'h3c111245),
	.w3(32'h3a1ca03e),
	.w4(32'hbb9649a1),
	.w5(32'h3b887fc2),
	.w6(32'h3c035b6c),
	.w7(32'hba1a501e),
	.w8(32'h3bc9ce01),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a4ccd),
	.w1(32'hba6ddf43),
	.w2(32'h3b5202f3),
	.w3(32'h3c1e375c),
	.w4(32'hbb14aa8f),
	.w5(32'hbaf287ce),
	.w6(32'h3bf98492),
	.w7(32'hba72c693),
	.w8(32'h3ada20ec),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd41e7),
	.w1(32'hb9f6f1d0),
	.w2(32'hbb29e46a),
	.w3(32'h3a37f590),
	.w4(32'hba804679),
	.w5(32'h3a397cdd),
	.w6(32'h3b359a0c),
	.w7(32'h38f0bf93),
	.w8(32'h3aefff4c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b018c9a),
	.w1(32'h3b980501),
	.w2(32'h3c18e878),
	.w3(32'hb87e97a6),
	.w4(32'h3bbf87c6),
	.w5(32'h3bfc27c8),
	.w6(32'hbb512de1),
	.w7(32'hb9d2e3a2),
	.w8(32'h3bc0a02e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb5682f),
	.w1(32'hbc4e9880),
	.w2(32'h3cb79b95),
	.w3(32'h3c2a559d),
	.w4(32'hbc77ae77),
	.w5(32'h3bf5e989),
	.w6(32'h3bc88245),
	.w7(32'hbc983459),
	.w8(32'h3c93be9f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5e63b6),
	.w1(32'hbc378768),
	.w2(32'hbbb143d1),
	.w3(32'h3d21d9d8),
	.w4(32'hbcdb67d7),
	.w5(32'hbca90e04),
	.w6(32'h3d8455fd),
	.w7(32'hbbf1faf6),
	.w8(32'h3aa87da1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfb9f80),
	.w1(32'hbc9e6b70),
	.w2(32'hbbe400e4),
	.w3(32'h3d0ba825),
	.w4(32'hbc9d3fb4),
	.w5(32'hbc664217),
	.w6(32'h3d5f2c62),
	.w7(32'hba56022a),
	.w8(32'h3c124fd7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c7c4b),
	.w1(32'hbb956217),
	.w2(32'hbb094ee1),
	.w3(32'h3b7f4ebb),
	.w4(32'hbbd895ba),
	.w5(32'hbbffa543),
	.w6(32'h3b873cb3),
	.w7(32'hbb58033f),
	.w8(32'hbb302a66),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3431ee),
	.w1(32'h3ac214eb),
	.w2(32'hbad532c4),
	.w3(32'h3a683cd7),
	.w4(32'h390664c7),
	.w5(32'h3a591d11),
	.w6(32'hb9961929),
	.w7(32'hb94ae43a),
	.w8(32'h3acf314b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2806b),
	.w1(32'h3a263670),
	.w2(32'hba8e0677),
	.w3(32'h39372595),
	.w4(32'hb9d6935f),
	.w5(32'hb802e764),
	.w6(32'h3aeed73c),
	.w7(32'hb9394f82),
	.w8(32'h3a4f1399),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c308af2),
	.w1(32'hbb53d191),
	.w2(32'hbaa62df5),
	.w3(32'h3c39c7aa),
	.w4(32'h3938a0cf),
	.w5(32'h3bd52dbf),
	.w6(32'h3c1120c6),
	.w7(32'h3b2b8e94),
	.w8(32'h3bc795a8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf124d7),
	.w1(32'h3b8d1c70),
	.w2(32'h3cce46c8),
	.w3(32'h3cd35bb0),
	.w4(32'h3bcac971),
	.w5(32'h3c998929),
	.w6(32'h3cf5191d),
	.w7(32'h3ca09979),
	.w8(32'h3d15c660),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d048351),
	.w1(32'h3ac8fd9c),
	.w2(32'h3ca07550),
	.w3(32'h3c9b5fd6),
	.w4(32'hbc3da9c5),
	.w5(32'h3bb333f3),
	.w6(32'h3cf017fb),
	.w7(32'hbb4a3319),
	.w8(32'h3c86630a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d11dd82),
	.w1(32'h3aa88e70),
	.w2(32'h3ca1ea8a),
	.w3(32'h3c96b19f),
	.w4(32'hbc63386a),
	.w5(32'h3c0cce3d),
	.w6(32'h3cf89425),
	.w7(32'hbb6c6950),
	.w8(32'h3c99973a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4641c),
	.w1(32'h3a8d58f2),
	.w2(32'h3c27b8d4),
	.w3(32'h3cafc518),
	.w4(32'hbba84d65),
	.w5(32'h3bdaec9e),
	.w6(32'h3cd31947),
	.w7(32'h3b082bb9),
	.w8(32'h3c936f5a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb6379),
	.w1(32'h3c668c14),
	.w2(32'h3ccd4a68),
	.w3(32'h3c1b013b),
	.w4(32'h3c9a400f),
	.w5(32'h3ce79e15),
	.w6(32'h3c59e170),
	.w7(32'h3c8241cf),
	.w8(32'h3cdb881a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac61a6d),
	.w1(32'hbac5a412),
	.w2(32'hba118f15),
	.w3(32'hbac7411d),
	.w4(32'hbaab114c),
	.w5(32'h38dde4ba),
	.w6(32'hbb58486e),
	.w7(32'hbae964ae),
	.w8(32'h3a8f2490),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cfb5a),
	.w1(32'hba48f7f2),
	.w2(32'hbab7424a),
	.w3(32'h3b2f4128),
	.w4(32'h3ad2f3a1),
	.w5(32'h3b234b2c),
	.w6(32'h3ba5c4d8),
	.w7(32'h3b7b35bf),
	.w8(32'h3b96061b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b953534),
	.w1(32'h39e383c5),
	.w2(32'hb9c98a9b),
	.w3(32'hbb050fd5),
	.w4(32'h3aab8882),
	.w5(32'h3a97424d),
	.w6(32'hbb1775dc),
	.w7(32'hb90c7cde),
	.w8(32'h375ea09d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cabb378),
	.w1(32'h3bf95a09),
	.w2(32'h3c81fffb),
	.w3(32'h3c6f7583),
	.w4(32'hba61c8f7),
	.w5(32'h3b9be200),
	.w6(32'h3c4dcc21),
	.w7(32'hbab14b0b),
	.w8(32'h3bc8ad4f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2df966),
	.w1(32'hb9dc3be5),
	.w2(32'h3b0b68f3),
	.w3(32'h3b4a5b1a),
	.w4(32'h3b28a499),
	.w5(32'h3b51f293),
	.w6(32'h3a9f2ebc),
	.w7(32'hb9384437),
	.w8(32'h3ae87bcf),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d6176),
	.w1(32'h3be04806),
	.w2(32'h3cbf8e8c),
	.w3(32'h3c4a20e8),
	.w4(32'h3b7604cd),
	.w5(32'h3ca3d3c0),
	.w6(32'h3c82386b),
	.w7(32'h3aa1dc5a),
	.w8(32'h3cb5d97e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21b914),
	.w1(32'h39a19776),
	.w2(32'h3b139a24),
	.w3(32'h3b56f750),
	.w4(32'h3ae41296),
	.w5(32'h3b98d356),
	.w6(32'h3bbe26e7),
	.w7(32'h3aeb700f),
	.w8(32'h3b9035c9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abae58d),
	.w1(32'h3b13dcac),
	.w2(32'h39e63f4f),
	.w3(32'h3a2f3678),
	.w4(32'hba4e6781),
	.w5(32'hb98aaeac),
	.w6(32'h3ab9b3d0),
	.w7(32'hb86c9e82),
	.w8(32'hb9d645f7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d6710),
	.w1(32'h3ae59556),
	.w2(32'hb9c4f8e2),
	.w3(32'hb919edfd),
	.w4(32'hbabf3226),
	.w5(32'hba91e3bb),
	.w6(32'h3a47a3b8),
	.w7(32'hba5abc8d),
	.w8(32'h3a1be702),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf8bbb),
	.w1(32'hba7fd2a0),
	.w2(32'hbb22b40e),
	.w3(32'h3ab39886),
	.w4(32'hbafc5694),
	.w5(32'hb9cd2d44),
	.w6(32'h3b0e41db),
	.w7(32'hbb6e150f),
	.w8(32'h3aa27b05),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6688c),
	.w1(32'hbb6c084a),
	.w2(32'hbab305c1),
	.w3(32'h3a07e9e1),
	.w4(32'hbba6bc96),
	.w5(32'hbbb8f151),
	.w6(32'h3bcea7df),
	.w7(32'hbb07a2c2),
	.w8(32'hb914f54b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a854559),
	.w1(32'h399a7833),
	.w2(32'h3a23614b),
	.w3(32'hba7ce2a5),
	.w4(32'hba82b614),
	.w5(32'h3a93389d),
	.w6(32'h3bd95ccb),
	.w7(32'h3b8c2c38),
	.w8(32'h3aa7f5c5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84b695),
	.w1(32'h3b5bd5a5),
	.w2(32'h3c33e670),
	.w3(32'h3c7aed07),
	.w4(32'h3b9f1b71),
	.w5(32'h3c594fff),
	.w6(32'h3c7a9e43),
	.w7(32'h3bbc82f1),
	.w8(32'h3c5183ec),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c832909),
	.w1(32'h3bd65d6a),
	.w2(32'h3bb8362c),
	.w3(32'h3c806b2b),
	.w4(32'h3c257d3d),
	.w5(32'h3b359f20),
	.w6(32'h3c7a3d46),
	.w7(32'h3c2b9187),
	.w8(32'h3bf7ae4e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92cb20),
	.w1(32'hbaf3a352),
	.w2(32'hbae3c8b2),
	.w3(32'hbaa9e4b2),
	.w4(32'hba3f754f),
	.w5(32'h3a78af76),
	.w6(32'hba8cfdc6),
	.w7(32'hbaa8bcc8),
	.w8(32'h3a105d87),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98601d0),
	.w1(32'h3b39015a),
	.w2(32'h3a9b5e39),
	.w3(32'h3adf635f),
	.w4(32'hb82a22a7),
	.w5(32'h3aef764f),
	.w6(32'h3abd98f1),
	.w7(32'h3a218306),
	.w8(32'h3a8aa231),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa89835),
	.w1(32'h3a61ae26),
	.w2(32'h3829f2b4),
	.w3(32'hba1621ce),
	.w4(32'h39fb8c53),
	.w5(32'hbab65d4b),
	.w6(32'hba96a7b8),
	.w7(32'hbaadbb3f),
	.w8(32'hba9dd724),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4133b4),
	.w1(32'hbae291fc),
	.w2(32'hbada278c),
	.w3(32'hbaf38c53),
	.w4(32'hb8d6c18a),
	.w5(32'hbb0cbba1),
	.w6(32'hba9921c1),
	.w7(32'hbacc770b),
	.w8(32'h3ab590f3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be98c2c),
	.w1(32'h3bf7d3bc),
	.w2(32'h3c92f903),
	.w3(32'h3c34d388),
	.w4(32'h3c2711b1),
	.w5(32'h3c883124),
	.w6(32'h3c677353),
	.w7(32'h3c54fdda),
	.w8(32'h3cea04bf),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2e392d),
	.w1(32'h3c9efd1e),
	.w2(32'h3d0f60bb),
	.w3(32'h3ced3861),
	.w4(32'h3c660faf),
	.w5(32'h3cdce4de),
	.w6(32'h3d15f99f),
	.w7(32'h3c678b05),
	.w8(32'h3cd29e54),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf6f0f8),
	.w1(32'hbb199b1a),
	.w2(32'h3c3c82a2),
	.w3(32'h3c923778),
	.w4(32'hbc09bede),
	.w5(32'h3baecebf),
	.w6(32'h3cebfa44),
	.w7(32'h3ba2f933),
	.w8(32'h3c63d059),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3b0176),
	.w1(32'hbc6a3d4c),
	.w2(32'h3cc2cc9f),
	.w3(32'h3ce27506),
	.w4(32'hbd104a69),
	.w5(32'hbb61caa5),
	.w6(32'h3d4a085f),
	.w7(32'hbcc4bb94),
	.w8(32'h3c71963d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a378dd4),
	.w1(32'h3a8cd4e1),
	.w2(32'h3a31b5f4),
	.w3(32'h3a1918d0),
	.w4(32'h3ab32f21),
	.w5(32'h3b0d90ae),
	.w6(32'h3b1e3bef),
	.w7(32'h3b09d215),
	.w8(32'h3acffb2b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cc7463),
	.w1(32'hb9b3a120),
	.w2(32'hbace2197),
	.w3(32'h3acd39b4),
	.w4(32'h3af0a7b2),
	.w5(32'h392d6be5),
	.w6(32'hba21cbb7),
	.w7(32'hbafb0ab8),
	.w8(32'hb9842380),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15b38e),
	.w1(32'hbb071f0b),
	.w2(32'hb9048ffc),
	.w3(32'h39efbcb8),
	.w4(32'h3b0500a8),
	.w5(32'h3ac9fb5a),
	.w6(32'hb8f13491),
	.w7(32'h3988cbea),
	.w8(32'hb93c8dea),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0113c6),
	.w1(32'hbb2ea3f1),
	.w2(32'h3b2c3185),
	.w3(32'h3b95d206),
	.w4(32'h3a1924bd),
	.w5(32'h3bcecabe),
	.w6(32'h3b819223),
	.w7(32'h393c1a10),
	.w8(32'h3be93de1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acde09c),
	.w1(32'h3af8bfff),
	.w2(32'h3af89dae),
	.w3(32'h3b4c12e4),
	.w4(32'h3b21e239),
	.w5(32'h39d312d9),
	.w6(32'h3aa52258),
	.w7(32'h3b248d41),
	.w8(32'hbb346d85),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaec472),
	.w1(32'h39cd4921),
	.w2(32'h3b9ced14),
	.w3(32'h3b557eda),
	.w4(32'h3c002dae),
	.w5(32'h3bc5638e),
	.w6(32'hbb42e866),
	.w7(32'h3b1b4f04),
	.w8(32'h3b872434),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98d9d0),
	.w1(32'h3ab17082),
	.w2(32'h3c065830),
	.w3(32'h3c6775e2),
	.w4(32'hbb3ecd7d),
	.w5(32'h3c567509),
	.w6(32'h3cbc2064),
	.w7(32'h3be9720d),
	.w8(32'h3c9268c9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cadf51e),
	.w1(32'h3b8a5724),
	.w2(32'h3c6bf833),
	.w3(32'h3c55d884),
	.w4(32'hbb960fb8),
	.w5(32'h3b89a0bd),
	.w6(32'h3c3dcabf),
	.w7(32'hbb7b9730),
	.w8(32'h3c1620c0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e03c0),
	.w1(32'hba99f219),
	.w2(32'h3c31ed31),
	.w3(32'h3bae6f36),
	.w4(32'hbb77272b),
	.w5(32'h3c1bce4f),
	.w6(32'h3bc44929),
	.w7(32'hbad0ea2b),
	.w8(32'h3c5d2228),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d74e9),
	.w1(32'h3b80ed00),
	.w2(32'h3c3f72a4),
	.w3(32'h3b93fab5),
	.w4(32'h3ba1bfe3),
	.w5(32'h3b5fd0c6),
	.w6(32'h3ad41b3f),
	.w7(32'h39db1222),
	.w8(32'h3bca25ed),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1485d2),
	.w1(32'hbba1cec1),
	.w2(32'h3aa1fe14),
	.w3(32'h3ba652d3),
	.w4(32'hbbd15507),
	.w5(32'h3a1bdb79),
	.w6(32'h3bd2bbcb),
	.w7(32'hbb50dd48),
	.w8(32'h3b8d61a1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a087ebb),
	.w1(32'hb99cffa3),
	.w2(32'h3c0cb886),
	.w3(32'hba7162a4),
	.w4(32'h3b044543),
	.w5(32'h3c33f4c7),
	.w6(32'hba15c829),
	.w7(32'h3874a97a),
	.w8(32'h3c290dcf),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb908ee7f),
	.w1(32'hb9717985),
	.w2(32'hba6a5cba),
	.w3(32'hba04a18d),
	.w4(32'h3a481377),
	.w5(32'h3bd8c475),
	.w6(32'hba89a240),
	.w7(32'hba338b8f),
	.w8(32'h3bb6ec59),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf725f),
	.w1(32'h3bc9fa09),
	.w2(32'h3ba4aa76),
	.w3(32'h3c0347d7),
	.w4(32'h3c113a42),
	.w5(32'hba624b9e),
	.w6(32'h3b994847),
	.w7(32'h3bb90203),
	.w8(32'hb8d737bc),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a5bc9),
	.w1(32'h37ed5df7),
	.w2(32'hb945290c),
	.w3(32'h398bf6e7),
	.w4(32'h39b8bef3),
	.w5(32'hb976dc1f),
	.w6(32'h39444343),
	.w7(32'h3891da26),
	.w8(32'h3a36d1bc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fc26a5),
	.w1(32'hb933e4cf),
	.w2(32'h384d0ef2),
	.w3(32'hba34fd13),
	.w4(32'hbac37ba0),
	.w5(32'hbb42069b),
	.w6(32'h3aa5602f),
	.w7(32'h392b0e96),
	.w8(32'hba54a4bf),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbad922),
	.w1(32'hbb32fc31),
	.w2(32'hbb751b5b),
	.w3(32'h3cabf793),
	.w4(32'hbc0473b3),
	.w5(32'hbc3065df),
	.w6(32'h3cbcfabc),
	.w7(32'hbbcb6011),
	.w8(32'hbb0335b1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef30a2),
	.w1(32'hbaaa03fc),
	.w2(32'h3a5d599f),
	.w3(32'hbb89108d),
	.w4(32'hbbadce7b),
	.w5(32'hbb3063f3),
	.w6(32'h3abf1c1c),
	.w7(32'hbada9e82),
	.w8(32'h3a36a34d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98a900),
	.w1(32'h3b81113f),
	.w2(32'h3c5b3d52),
	.w3(32'h3c0af0a0),
	.w4(32'hbb43560b),
	.w5(32'h3bfd03b1),
	.w6(32'h3c6a72be),
	.w7(32'hb9ab8b11),
	.w8(32'h3be95677),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8426a7),
	.w1(32'h3c099b8f),
	.w2(32'h3c2e488e),
	.w3(32'h3cc6d248),
	.w4(32'h3bdff1b6),
	.w5(32'h3c4a78e4),
	.w6(32'h3cdca89f),
	.w7(32'h3c7e39fc),
	.w8(32'h3c8ceebc),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21e17f),
	.w1(32'hbc2e095b),
	.w2(32'hbb39f75f),
	.w3(32'h3c56a7de),
	.w4(32'hbbef0523),
	.w5(32'hbbc8e69b),
	.w6(32'h3c790e99),
	.w7(32'hbb618de8),
	.w8(32'hbabb56fa),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e9e28),
	.w1(32'h3b8aace7),
	.w2(32'h3c693e8d),
	.w3(32'h3c1833b3),
	.w4(32'hbc0e8c32),
	.w5(32'hbad7f055),
	.w6(32'h3c358b4a),
	.w7(32'h3b814aa7),
	.w8(32'h3c6d629b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ba19c),
	.w1(32'hbc4e63a3),
	.w2(32'hbb4dc202),
	.w3(32'h3b7f7e7c),
	.w4(32'hbc49cc23),
	.w5(32'hbbdd01ae),
	.w6(32'h3bbb3113),
	.w7(32'hbc5ddf7f),
	.w8(32'hbc03bbd2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd45690),
	.w1(32'h3b932295),
	.w2(32'h3c6972b1),
	.w3(32'h3c7a44ed),
	.w4(32'hbb774901),
	.w5(32'h3b903d04),
	.w6(32'h3cb05ae8),
	.w7(32'hb9884225),
	.w8(32'h3c59d0f3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41574b),
	.w1(32'hba429eb5),
	.w2(32'h3bf92c34),
	.w3(32'h3c06db2d),
	.w4(32'hbbeff9e5),
	.w5(32'hbbb27fbe),
	.w6(32'h3bf28d4a),
	.w7(32'hbb8c8dad),
	.w8(32'h3b9cd462),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc37718),
	.w1(32'hbbe962fd),
	.w2(32'h3b334ec2),
	.w3(32'h3c80a4ae),
	.w4(32'hbc601d1a),
	.w5(32'hbb8d6119),
	.w6(32'h3cb7ab0f),
	.w7(32'hbbc1593d),
	.w8(32'h3a344aff),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe3a7e),
	.w1(32'hbb14174a),
	.w2(32'hbabd769e),
	.w3(32'hbb0a864b),
	.w4(32'hba5854f3),
	.w5(32'hb9a36729),
	.w6(32'hbba33a41),
	.w7(32'hbb3e1311),
	.w8(32'hbb98d221),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca94299),
	.w1(32'h3b4ae659),
	.w2(32'h3c85dd38),
	.w3(32'h3c3364c0),
	.w4(32'hbb9ea4a0),
	.w5(32'h3c1fdad2),
	.w6(32'h3cb21a89),
	.w7(32'h3be15a69),
	.w8(32'h3cb3d5a4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c137900),
	.w1(32'h3b13a889),
	.w2(32'h3c43a0a5),
	.w3(32'h3c0bdcae),
	.w4(32'hbb6d62fe),
	.w5(32'h3ac79ea0),
	.w6(32'h3b9436de),
	.w7(32'h3b71377b),
	.w8(32'h3c14c222),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf04ea),
	.w1(32'hba658618),
	.w2(32'h3cff6bdc),
	.w3(32'h3a57e75f),
	.w4(32'hbc8e642e),
	.w5(32'h3bdc5c85),
	.w6(32'h3b9f18af),
	.w7(32'hbc2b9f4f),
	.w8(32'h3c95edb7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d45706e),
	.w1(32'hbc911f34),
	.w2(32'hbcd5cc06),
	.w3(32'h3ceec2ef),
	.w4(32'hbd197c4c),
	.w5(32'hbd1a31ce),
	.w6(32'h3d0e6ade),
	.w7(32'hbc99574d),
	.w8(32'hbcb70dfa),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2b825),
	.w1(32'hb71261c0),
	.w2(32'h3ca2641c),
	.w3(32'h3c5845ff),
	.w4(32'hbc1ea5f5),
	.w5(32'h3c48b2ef),
	.w6(32'h3cc519af),
	.w7(32'hbb1fa84d),
	.w8(32'h3c99f9b8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62203a),
	.w1(32'h3bbad802),
	.w2(32'h3c6d0320),
	.w3(32'h3b9a481d),
	.w4(32'h3ac821ba),
	.w5(32'h3c18a145),
	.w6(32'hbb734b4e),
	.w7(32'hbbb1ab10),
	.w8(32'h3c547e29),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e218f),
	.w1(32'h3a90d3b7),
	.w2(32'hb8d5be60),
	.w3(32'h3981e54d),
	.w4(32'hb986fc2e),
	.w5(32'hb98a754d),
	.w6(32'hba213fe6),
	.w7(32'hbab08da8),
	.w8(32'hbae08c87),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d21e577),
	.w1(32'h3c7818f7),
	.w2(32'h3cf0a187),
	.w3(32'h3c695107),
	.w4(32'hbad20ed1),
	.w5(32'h3c51d119),
	.w6(32'h3b619d51),
	.w7(32'hbc173703),
	.w8(32'h3c06916d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb19cf6),
	.w1(32'hbba2cc8b),
	.w2(32'h3be15aba),
	.w3(32'h3ba98ed4),
	.w4(32'h3a435d23),
	.w5(32'h3c310b82),
	.w6(32'h3891a33a),
	.w7(32'hbba6cde4),
	.w8(32'h3bff0c7b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b1829e),
	.w1(32'hb9dada38),
	.w2(32'h3a760a2c),
	.w3(32'h37e10678),
	.w4(32'hbad56a51),
	.w5(32'hb968139c),
	.w6(32'hb9c1b83e),
	.w7(32'hbad5ee24),
	.w8(32'hba209583),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf4e68),
	.w1(32'h3af8247b),
	.w2(32'h3b550192),
	.w3(32'h3b5d0cba),
	.w4(32'h39a251e4),
	.w5(32'h39cf6c24),
	.w6(32'h3bd299d7),
	.w7(32'h3b1bbeb4),
	.w8(32'h3b20f743),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c519b07),
	.w1(32'h3b5373c8),
	.w2(32'h3c62f198),
	.w3(32'h3c0a4bca),
	.w4(32'h3b7b19cc),
	.w5(32'h3c5d1434),
	.w6(32'h3c4da5ac),
	.w7(32'h3c35bb45),
	.w8(32'h3cae2085),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6682aa),
	.w1(32'hbb428fe9),
	.w2(32'h3c079bfd),
	.w3(32'h3c1e563e),
	.w4(32'hbbdd84cb),
	.w5(32'h3b99e0dd),
	.w6(32'h3c818d71),
	.w7(32'hbb335873),
	.w8(32'h3c42b6fe),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07386c),
	.w1(32'hbb055a16),
	.w2(32'h3acbcc71),
	.w3(32'h3ba42471),
	.w4(32'hbbb7deb3),
	.w5(32'hbb52c8ca),
	.w6(32'h3c892b54),
	.w7(32'h3b42ffef),
	.w8(32'h3bb4d95a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74d51e),
	.w1(32'h3915bcfc),
	.w2(32'h3ba22836),
	.w3(32'h3c051976),
	.w4(32'hbbd3bd07),
	.w5(32'hbacfeec7),
	.w6(32'h3bf28708),
	.w7(32'hbb7d7bd3),
	.w8(32'h3ba0f91a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf2812),
	.w1(32'hbc031dfe),
	.w2(32'hbb1f5be9),
	.w3(32'h3bb7815b),
	.w4(32'hbc0d7311),
	.w5(32'h3a910c22),
	.w6(32'h3c6b56d6),
	.w7(32'hbb07efd5),
	.w8(32'h3bf53b43),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7aff6b),
	.w1(32'h3b8bd64d),
	.w2(32'h3c47ab1f),
	.w3(32'h3be8dde4),
	.w4(32'hbbe74104),
	.w5(32'hbae317da),
	.w6(32'h3c079269),
	.w7(32'h390ac460),
	.w8(32'h3bfd99ba),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5479bb),
	.w1(32'hb9d44362),
	.w2(32'h3b8c0b52),
	.w3(32'h3c1fcd6c),
	.w4(32'hbb41f268),
	.w5(32'h3b1f318d),
	.w6(32'h3c4e197d),
	.w7(32'hba636ebb),
	.w8(32'h3befe770),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35635577),
	.w1(32'h3976fafc),
	.w2(32'h3994f4f3),
	.w3(32'hb8eb8aa1),
	.w4(32'h3a127ceb),
	.w5(32'hb9b2a37e),
	.w6(32'hb9912437),
	.w7(32'h393c0caa),
	.w8(32'hb96c55fa),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8823d9),
	.w1(32'hb9cb368e),
	.w2(32'hb99a92f7),
	.w3(32'hb9600ec0),
	.w4(32'hbac7cd4a),
	.w5(32'h38389e38),
	.w6(32'h3a52691a),
	.w7(32'hb9e14b86),
	.w8(32'h3a157224),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29f3b8),
	.w1(32'h39cb0839),
	.w2(32'h3a367181),
	.w3(32'h3a3a87a7),
	.w4(32'h3a448e49),
	.w5(32'hba2a9286),
	.w6(32'h3a562ac0),
	.w7(32'hba163583),
	.w8(32'hba6731aa),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba609986),
	.w1(32'hba39ec60),
	.w2(32'hba3a89e9),
	.w3(32'h3ac0b365),
	.w4(32'hb99cf72e),
	.w5(32'hba22c90e),
	.w6(32'h3ab98668),
	.w7(32'hba396a8e),
	.w8(32'hbad299d5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c821534),
	.w1(32'hbbb1e6da),
	.w2(32'h3b8bdcb3),
	.w3(32'h3c02ba62),
	.w4(32'hbc236400),
	.w5(32'h3b5bd3e8),
	.w6(32'h3c539d2e),
	.w7(32'hbb9b461a),
	.w8(32'h3c2bbe23),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8810df),
	.w1(32'h3ae83e7d),
	.w2(32'h3b01ca73),
	.w3(32'h3b260488),
	.w4(32'h3a7ee557),
	.w5(32'h3aa2dcca),
	.w6(32'h3b38ec9e),
	.w7(32'h3a2db433),
	.w8(32'hb8f34c73),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb91b7),
	.w1(32'h3a2d5ad6),
	.w2(32'h3c09cfdc),
	.w3(32'hb980bbab),
	.w4(32'h3b45209e),
	.w5(32'h3bdc7bcd),
	.w6(32'hbb8f3b77),
	.w7(32'h3aceac48),
	.w8(32'h3bc81164),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce3f332),
	.w1(32'h3b0819de),
	.w2(32'h3bd41869),
	.w3(32'h3ca91501),
	.w4(32'hbc1acc1d),
	.w5(32'hbb88cfcd),
	.w6(32'h3ccd0966),
	.w7(32'hbb136167),
	.w8(32'h3bf0561f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0b0cf),
	.w1(32'h3a0cad80),
	.w2(32'h3a8e664e),
	.w3(32'h3932a753),
	.w4(32'h39566405),
	.w5(32'hb78c7985),
	.w6(32'h3a81ed14),
	.w7(32'h39adb143),
	.w8(32'hb99e413b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55663b),
	.w1(32'h39abe349),
	.w2(32'h3a99e6f9),
	.w3(32'hba4c5910),
	.w4(32'hba1c1b44),
	.w5(32'h39a72b19),
	.w6(32'h3a37c562),
	.w7(32'h378347e0),
	.w8(32'h3aa51429),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08c536),
	.w1(32'h3a2ca688),
	.w2(32'h3a674389),
	.w3(32'h3a0db599),
	.w4(32'h3a433705),
	.w5(32'hba27f83e),
	.w6(32'h3ab7fc4f),
	.w7(32'h3a22e10a),
	.w8(32'hb9e6359e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b55b0),
	.w1(32'hb97358e0),
	.w2(32'h3924352f),
	.w3(32'h3ac00c23),
	.w4(32'hba65bc8d),
	.w5(32'hba9e4c31),
	.w6(32'h3b3ed4b2),
	.w7(32'h3ac1f133),
	.w8(32'h3ab9c97f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1114e),
	.w1(32'h3c17359e),
	.w2(32'h3bcc54ae),
	.w3(32'hbb18b986),
	.w4(32'h3bf83efb),
	.w5(32'h3c9e3f78),
	.w6(32'h3b83f798),
	.w7(32'h3bc556bc),
	.w8(32'h3c2cc7b8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c513f6c),
	.w1(32'h3a25a62d),
	.w2(32'h3c7ecd04),
	.w3(32'h3bf63ad5),
	.w4(32'hb9026c39),
	.w5(32'h3c71edf0),
	.w6(32'h3c0efd4a),
	.w7(32'h3b8c01d1),
	.w8(32'h3ca491d4),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab246be),
	.w1(32'h3b0d627b),
	.w2(32'h3b37a251),
	.w3(32'h3a5399a2),
	.w4(32'h3a8b583c),
	.w5(32'hba3d4bc7),
	.w6(32'hba81be54),
	.w7(32'hb932b709),
	.w8(32'h3a9027e3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1c89f),
	.w1(32'h3a497a3d),
	.w2(32'h3b187b57),
	.w3(32'h3b92d70a),
	.w4(32'hb9ae3de9),
	.w5(32'h3ab1a423),
	.w6(32'h3c1aad48),
	.w7(32'h3ada7fdc),
	.w8(32'h3b7ee99d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb26ec),
	.w1(32'hb8705516),
	.w2(32'h3b57756d),
	.w3(32'h3bb812c1),
	.w4(32'hbb270a9f),
	.w5(32'hb8d3c402),
	.w6(32'h3bba402a),
	.w7(32'hbac769a8),
	.w8(32'h3ae14a63),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd87b5),
	.w1(32'hbaec4cbd),
	.w2(32'h3b830cc0),
	.w3(32'h3b237d59),
	.w4(32'hbb1b4525),
	.w5(32'h39db7c21),
	.w6(32'h3bf6c87a),
	.w7(32'h39b420be),
	.w8(32'h3b8095b9),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c692a19),
	.w1(32'h3b8ff624),
	.w2(32'h3c583ddc),
	.w3(32'h3be12f72),
	.w4(32'hbbc4a962),
	.w5(32'hb9b7946a),
	.w6(32'h3bf3b076),
	.w7(32'hbb130322),
	.w8(32'h3b720102),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5b893),
	.w1(32'h3b46f264),
	.w2(32'h3c8d2037),
	.w3(32'h3b8e5346),
	.w4(32'h3add2107),
	.w5(32'h3c60c338),
	.w6(32'h3be8a36d),
	.w7(32'h3bc2df6e),
	.w8(32'h3ca1299d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81d500),
	.w1(32'hbb3caadc),
	.w2(32'h3b8d9e87),
	.w3(32'h3c2f81df),
	.w4(32'hbc0b1b20),
	.w5(32'hba7d59a1),
	.w6(32'h3c5f7e0f),
	.w7(32'hbb8cdd6f),
	.w8(32'h3bc1a51c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e41e7),
	.w1(32'h3b9d550a),
	.w2(32'h3c0114fe),
	.w3(32'h3b8ed034),
	.w4(32'hbb916779),
	.w5(32'h3b014058),
	.w6(32'h3b917055),
	.w7(32'h3abd1bfe),
	.w8(32'h3c011e72),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a8485),
	.w1(32'h3b96f211),
	.w2(32'h3c59ecc7),
	.w3(32'h3bcf5368),
	.w4(32'h3b85c719),
	.w5(32'h3c750fab),
	.w6(32'h3bf71c06),
	.w7(32'h3b4b571f),
	.w8(32'h3c4b06df),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b791c),
	.w1(32'hba7c0e17),
	.w2(32'hba55a327),
	.w3(32'h3c29f6ab),
	.w4(32'hbbb673ca),
	.w5(32'hbb53d016),
	.w6(32'h3c883dd2),
	.w7(32'hbb31cafa),
	.w8(32'h3ae50714),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3088f8),
	.w1(32'h3b05a075),
	.w2(32'h3c0f2281),
	.w3(32'h3bd3dbda),
	.w4(32'hba3d0b9b),
	.w5(32'h3bbfd11b),
	.w6(32'h3bf7ade5),
	.w7(32'h3b5068d1),
	.w8(32'h3c57e2fa),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baabcda),
	.w1(32'hb9e052d7),
	.w2(32'h3b387498),
	.w3(32'h3b29ce89),
	.w4(32'hbb17038b),
	.w5(32'h3a836389),
	.w6(32'h3b919694),
	.w7(32'hba84ee79),
	.w8(32'h3b3c59cf),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb549d9),
	.w1(32'hbc788bc5),
	.w2(32'hbbb41da2),
	.w3(32'h3ca74371),
	.w4(32'hbc2b8556),
	.w5(32'hbafcc9c4),
	.w6(32'h3cb350fa),
	.w7(32'hbbd99b33),
	.w8(32'h3bcff565),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e18ef),
	.w1(32'hba4e930d),
	.w2(32'hba2d6683),
	.w3(32'h3c0b7a6e),
	.w4(32'hbb1be112),
	.w5(32'hbb24bc5e),
	.w6(32'h3c5b5ede),
	.w7(32'h3abe8145),
	.w8(32'h3b734ae8),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39944c53),
	.w1(32'hb8fff5f9),
	.w2(32'h3995c3bd),
	.w3(32'h3898151d),
	.w4(32'h3a3878cc),
	.w5(32'hb90fc29b),
	.w6(32'hb9de62b1),
	.w7(32'h39127c9e),
	.w8(32'hb9b4b6d2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9597a91),
	.w1(32'hba1f262a),
	.w2(32'hb9d06a76),
	.w3(32'hba03d373),
	.w4(32'hb7966fa7),
	.w5(32'h38653ee3),
	.w6(32'hb9deba70),
	.w7(32'hb9fcbdf7),
	.w8(32'h381953fd),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb060f7),
	.w1(32'h39b9c914),
	.w2(32'h3b19d818),
	.w3(32'h3bbcda8f),
	.w4(32'hbab84602),
	.w5(32'hba917ddc),
	.w6(32'h3bb8ba67),
	.w7(32'hbaf657f9),
	.w8(32'h3a1e0152),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4b5ab),
	.w1(32'hbb33ad51),
	.w2(32'h3b4aeaca),
	.w3(32'h3c0b876f),
	.w4(32'hbc2f6c58),
	.w5(32'hbbb6e55f),
	.w6(32'h3c86007c),
	.w7(32'hbb795cc3),
	.w8(32'h3bda68ea),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cabf828),
	.w1(32'h3af9c4f0),
	.w2(32'h3caba619),
	.w3(32'h3c9e0e35),
	.w4(32'hbaa459cb),
	.w5(32'h3c8045df),
	.w6(32'h3c8d23f8),
	.w7(32'hba75b13d),
	.w8(32'h3c842da2),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a4c2c6),
	.w1(32'hb99fb4d4),
	.w2(32'hb847c19c),
	.w3(32'hba13245e),
	.w4(32'h39e0b470),
	.w5(32'h3714f783),
	.w6(32'hba807909),
	.w7(32'hb8282cf0),
	.w8(32'h382427d7),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c835f4b),
	.w1(32'h3aeefdc9),
	.w2(32'h3c89c65c),
	.w3(32'h3c33a51d),
	.w4(32'hba97fa8b),
	.w5(32'h3c610f0f),
	.w6(32'h3c6859b7),
	.w7(32'h3b914dc8),
	.w8(32'h3ca3d388),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a6637),
	.w1(32'h3aad1d9c),
	.w2(32'h3c0ac908),
	.w3(32'h3bf04b68),
	.w4(32'hbb55ca6b),
	.w5(32'h3ab5757a),
	.w6(32'h3c12d156),
	.w7(32'h3ac00922),
	.w8(32'h3c14f79e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9272ba),
	.w1(32'h3be814dd),
	.w2(32'h3c9bdb00),
	.w3(32'h3b08f255),
	.w4(32'h3b32c0f8),
	.w5(32'h3c46fb86),
	.w6(32'hbba78d3b),
	.w7(32'h3b0f38d2),
	.w8(32'h3c7186a4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4a9ce),
	.w1(32'hbc485c13),
	.w2(32'h3c283c94),
	.w3(32'h3ba06d10),
	.w4(32'hbc810d63),
	.w5(32'hb9d9198a),
	.w6(32'h3c881df8),
	.w7(32'hbc165b99),
	.w8(32'h3bd17986),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c394890),
	.w1(32'h3b4f033e),
	.w2(32'h3a884ba7),
	.w3(32'h3bf76dee),
	.w4(32'h3b1b13c0),
	.w5(32'h39c19b64),
	.w6(32'h3c1a8ff1),
	.w7(32'h3ac78ef9),
	.w8(32'h3b06bdfa),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09c6da),
	.w1(32'hbadb8ad4),
	.w2(32'hbb2d2007),
	.w3(32'hba4f4c6e),
	.w4(32'hb9fba77a),
	.w5(32'hbaffafd2),
	.w6(32'hba8ff884),
	.w7(32'hbaffc426),
	.w8(32'hbb813cdd),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50dd47),
	.w1(32'hbc123c8e),
	.w2(32'hbbd07138),
	.w3(32'h3c042118),
	.w4(32'hbc22dfb5),
	.w5(32'hbb9bb752),
	.w6(32'h3c8c59e9),
	.w7(32'hbb638c52),
	.w8(32'h3b90cce1),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad654d),
	.w1(32'hbb469de3),
	.w2(32'hbb387ef7),
	.w3(32'h3c4fbbae),
	.w4(32'hbc3c8baa),
	.w5(32'hbb5b34fe),
	.w6(32'h3c99e094),
	.w7(32'hbb5112a0),
	.w8(32'h3b8a9af0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad43b4),
	.w1(32'hbc3b9557),
	.w2(32'hbb160841),
	.w3(32'h3ba14458),
	.w4(32'hbc5d5ea0),
	.w5(32'hbbc2e266),
	.w6(32'h3c34f3fc),
	.w7(32'hbc08310c),
	.w8(32'hb9eec7e4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966d864),
	.w1(32'h3a892136),
	.w2(32'h3b18f268),
	.w3(32'h3aff7e3c),
	.w4(32'h3b26959e),
	.w5(32'h3b6b5c30),
	.w6(32'h3ad756cd),
	.w7(32'h3abd78d6),
	.w8(32'h3bb1bbc0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af769aa),
	.w1(32'h3b0ebe45),
	.w2(32'h3ac8c26b),
	.w3(32'h3aec2f92),
	.w4(32'h3a47d765),
	.w5(32'hb9c9f660),
	.w6(32'h3b2d78ab),
	.w7(32'h3ab23d69),
	.w8(32'h3a5ba48f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6cdc86),
	.w1(32'h3bab36fd),
	.w2(32'h3c2ad0a2),
	.w3(32'h3be2ad60),
	.w4(32'h39ad3cb9),
	.w5(32'h3c0d04f6),
	.w6(32'h3c1369be),
	.w7(32'h3b9d8e75),
	.w8(32'h3c332f66),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf46450),
	.w1(32'hb9fc774d),
	.w2(32'h3b06453f),
	.w3(32'hba255784),
	.w4(32'h398b5ec4),
	.w5(32'h3b1ed638),
	.w6(32'hbad98535),
	.w7(32'hba3fd89f),
	.w8(32'h3a65481c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20713d),
	.w1(32'hbb5484ab),
	.w2(32'h3a71b972),
	.w3(32'h3bef754c),
	.w4(32'hbafaa362),
	.w5(32'h3a222008),
	.w6(32'h3c3a18b1),
	.w7(32'hba5a4aea),
	.w8(32'h3b836781),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a22a63),
	.w1(32'h38b12308),
	.w2(32'h3a3ccc94),
	.w3(32'hba04fbba),
	.w4(32'hb9a8a0e9),
	.w5(32'h3996306f),
	.w6(32'h394412d9),
	.w7(32'hb920770a),
	.w8(32'hb9892425),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7554c7),
	.w1(32'hbb8d2d4b),
	.w2(32'h3b80f648),
	.w3(32'h3bee52d4),
	.w4(32'hba6eed50),
	.w5(32'h3b6de43f),
	.w6(32'h3c24d371),
	.w7(32'hbb34a737),
	.w8(32'h3b541e95),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374d9973),
	.w1(32'hba6624eb),
	.w2(32'hb8e50f9b),
	.w3(32'hba69ba80),
	.w4(32'h38dc85c6),
	.w5(32'h3a6569d2),
	.w6(32'hbab2af08),
	.w7(32'hb9b64b48),
	.w8(32'h398ceacf),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa88d93),
	.w1(32'h3a74f1ca),
	.w2(32'h3ac5d13a),
	.w3(32'h3b1207f5),
	.w4(32'h3ab4b5f2),
	.w5(32'h3aabf207),
	.w6(32'h3b6c1400),
	.w7(32'h3b07edb9),
	.w8(32'h3a93c086),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ff948),
	.w1(32'h3ab5d285),
	.w2(32'h3b88d527),
	.w3(32'h3c12527a),
	.w4(32'hbb919202),
	.w5(32'h3aedf733),
	.w6(32'h3c667940),
	.w7(32'hb8c1f66b),
	.w8(32'h3bdd3139),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdc2346),
	.w1(32'h3a993fdc),
	.w2(32'h3c6f5f46),
	.w3(32'h3cae44cf),
	.w4(32'h3af0db1c),
	.w5(32'h3cde566d),
	.w6(32'h3cc100d6),
	.w7(32'h3b60de84),
	.w8(32'h3cef40cb),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babe1dc),
	.w1(32'hbbf0692c),
	.w2(32'hbb26ae97),
	.w3(32'h3b597220),
	.w4(32'hbc056818),
	.w5(32'hbb23c06c),
	.w6(32'h3c073209),
	.w7(32'hbba69eaf),
	.w8(32'h399d417c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9eae46),
	.w1(32'h39dcf40c),
	.w2(32'h3c435a97),
	.w3(32'h3c27bf3f),
	.w4(32'hbbbe69c2),
	.w5(32'h3bf9cc73),
	.w6(32'h3c4bea7d),
	.w7(32'hbb5c05dd),
	.w8(32'h3c3827f1),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7bf5a),
	.w1(32'hb8485ec9),
	.w2(32'h3b395dfe),
	.w3(32'h3b994059),
	.w4(32'h3a8e0f70),
	.w5(32'hba1aeb71),
	.w6(32'h3ad1caac),
	.w7(32'hbaa0e4c0),
	.w8(32'hb96aa6aa),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc19b09),
	.w1(32'hbb43a315),
	.w2(32'h3cd9bc35),
	.w3(32'h3c83105e),
	.w4(32'hbc27e89a),
	.w5(32'h3c7bfd7c),
	.w6(32'h3cc37055),
	.w7(32'h3c175783),
	.w8(32'h3ce45720),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9730c9),
	.w1(32'h3aa45bb2),
	.w2(32'h3c68d939),
	.w3(32'h3c47d01e),
	.w4(32'hbbd5fab6),
	.w5(32'h3b80b6e6),
	.w6(32'h3c93fb0c),
	.w7(32'hbae64cf5),
	.w8(32'h3c084992),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29dd1a),
	.w1(32'hb99702a4),
	.w2(32'h3c856f46),
	.w3(32'h3bad4eeb),
	.w4(32'hbacd0234),
	.w5(32'h3c80c7e2),
	.w6(32'h3c14779a),
	.w7(32'h3b0a4296),
	.w8(32'h3ca2f74c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38860ebb),
	.w1(32'hb9cf3c0b),
	.w2(32'hba33e4bf),
	.w3(32'hb9c839bd),
	.w4(32'hba62ea0b),
	.w5(32'hba48972a),
	.w6(32'hba01f402),
	.w7(32'hb9fa6e04),
	.w8(32'hba3efcda),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c020d34),
	.w1(32'h3b3309c5),
	.w2(32'h3c0977e5),
	.w3(32'h3b8b1fb0),
	.w4(32'hbaf8da37),
	.w5(32'h3b86ac8b),
	.w6(32'h3b49d041),
	.w7(32'hbb022597),
	.w8(32'h3b8c0fcb),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba726e77),
	.w1(32'hba8dfe11),
	.w2(32'hb9a0c51a),
	.w3(32'hba808799),
	.w4(32'hb91fd890),
	.w5(32'hba5ba859),
	.w6(32'hba96596e),
	.w7(32'hb977cedc),
	.w8(32'hba8a4e4f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ecfa8b),
	.w1(32'h3a2396af),
	.w2(32'h3bf935a8),
	.w3(32'hb988c6f5),
	.w4(32'h39315cef),
	.w5(32'h3b31686a),
	.w6(32'h3a769ba7),
	.w7(32'h39949d10),
	.w8(32'h3b9cb1d0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d4cad),
	.w1(32'h393f4702),
	.w2(32'h3adb7e2a),
	.w3(32'h3bc0af8c),
	.w4(32'h39971408),
	.w5(32'h397a7eb9),
	.w6(32'h3ba3e1ec),
	.w7(32'hba59fbae),
	.w8(32'h3aa2a000),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e9950),
	.w1(32'hbab5de5b),
	.w2(32'h3c2f5c8d),
	.w3(32'h3be29081),
	.w4(32'hbbcc9b57),
	.w5(32'h3adb670e),
	.w6(32'h3c381118),
	.w7(32'hba5618a7),
	.w8(32'h3c23797e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00756e),
	.w1(32'hb9c528ed),
	.w2(32'hba5e1950),
	.w3(32'hb9b0859d),
	.w4(32'hb9b26a4d),
	.w5(32'hba371aa5),
	.w6(32'hba5bbea8),
	.w7(32'hba1d83b6),
	.w8(32'hba07a004),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3729191b),
	.w1(32'h393085b8),
	.w2(32'h3a0dee16),
	.w3(32'h375a22d0),
	.w4(32'h3a2540ae),
	.w5(32'h3a5233b6),
	.w6(32'hb90ef81d),
	.w7(32'hb6cdcfb6),
	.w8(32'h39c44117),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6425c),
	.w1(32'hbb0bbfcf),
	.w2(32'hbaf13efe),
	.w3(32'h3b8cb374),
	.w4(32'hbb8ea922),
	.w5(32'hbb3fdb60),
	.w6(32'h3bf22c56),
	.w7(32'hbb096cf7),
	.w8(32'hba4c4f44),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8791d7),
	.w1(32'h3add708d),
	.w2(32'h3bc9ddf9),
	.w3(32'h3c797abd),
	.w4(32'hbaa8f029),
	.w5(32'hba4227ac),
	.w6(32'h3c7e8cb0),
	.w7(32'h3b9ebe0e),
	.w8(32'h3bac3918),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8e9ce),
	.w1(32'hbb832725),
	.w2(32'h3b6538eb),
	.w3(32'h3c028bf9),
	.w4(32'hbb0d6ae9),
	.w5(32'h3b706472),
	.w6(32'hbb574b34),
	.w7(32'hbc22990b),
	.w8(32'h3b8bfece),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05bb74),
	.w1(32'hbb01b795),
	.w2(32'h39c0747e),
	.w3(32'h3b3af738),
	.w4(32'hba666704),
	.w5(32'h3acc5010),
	.w6(32'h3b3da4ba),
	.w7(32'hb95c32d5),
	.w8(32'h3b7c8458),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2a27a1),
	.w1(32'h3c79fd0f),
	.w2(32'h3d42fee5),
	.w3(32'h3d0d6ee0),
	.w4(32'h3c3ad8f4),
	.w5(32'h3d3a96a3),
	.w6(32'h3cfa2b61),
	.w7(32'h3c9d97fb),
	.w8(32'h3d3582fa),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1c6afa),
	.w1(32'hbb2af0f0),
	.w2(32'h3c2fe1ab),
	.w3(32'h3d0b7dd7),
	.w4(32'hbc477744),
	.w5(32'hbc03fa85),
	.w6(32'h3d16be1b),
	.w7(32'hbc1f4d2c),
	.w8(32'h3ba37de0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15f93d),
	.w1(32'hb953ec14),
	.w2(32'h3af4ffdc),
	.w3(32'hba77f795),
	.w4(32'h3b305292),
	.w5(32'h3b998a70),
	.w6(32'hbaa72447),
	.w7(32'h3a607279),
	.w8(32'h3b8140ba),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f26b7),
	.w1(32'hba43c133),
	.w2(32'hb89941dc),
	.w3(32'h38c70ae9),
	.w4(32'h3a582122),
	.w5(32'h3a611ba8),
	.w6(32'h3986b9ab),
	.w7(32'h391ba854),
	.w8(32'hb9172c69),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8b34a),
	.w1(32'h3a35d970),
	.w2(32'h3a8b8081),
	.w3(32'h3a1dc822),
	.w4(32'h3ac47513),
	.w5(32'h3aa811fd),
	.w6(32'h39781539),
	.w7(32'h3acc212e),
	.w8(32'h3a0ead28),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba562da7),
	.w1(32'h38a6ec69),
	.w2(32'h3a2a364f),
	.w3(32'h39b80167),
	.w4(32'h3a8a44da),
	.w5(32'hb9d75aa4),
	.w6(32'h39935246),
	.w7(32'h3aa371e4),
	.w8(32'h398b33b2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb853a829),
	.w1(32'h3b5ca37e),
	.w2(32'h3bdf69b2),
	.w3(32'h39c12cae),
	.w4(32'h3b9e9932),
	.w5(32'h3bb44433),
	.w6(32'hb9a21466),
	.w7(32'h3b4c7b68),
	.w8(32'h3bdb0189),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5afb4a),
	.w1(32'h3a335e73),
	.w2(32'h3b5276a4),
	.w3(32'h3b9753b0),
	.w4(32'hbbefadc2),
	.w5(32'hbabe0100),
	.w6(32'h3c58578c),
	.w7(32'h3ac949f2),
	.w8(32'h3c30d16f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd40535),
	.w1(32'h3b324f7f),
	.w2(32'h3ca91fa7),
	.w3(32'h3c862f95),
	.w4(32'hbc26936a),
	.w5(32'h3bf0ed56),
	.w6(32'h3caae2ee),
	.w7(32'hbba110a3),
	.w8(32'h3c254afb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c65b4),
	.w1(32'hbb62c541),
	.w2(32'h38d5c0b4),
	.w3(32'h3b5222e2),
	.w4(32'hbafe845c),
	.w5(32'hba0a50cd),
	.w6(32'h3bae528d),
	.w7(32'h3a3c0992),
	.w8(32'h3b3046a0),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ba56c),
	.w1(32'h3bf1148b),
	.w2(32'h3c9fada7),
	.w3(32'h3bec09af),
	.w4(32'h39e85d7a),
	.w5(32'h3c573a1f),
	.w6(32'h3c72ad98),
	.w7(32'h3bfd53ae),
	.w8(32'h3cac3377),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8549d1),
	.w1(32'hbaa96cba),
	.w2(32'h3b0a1648),
	.w3(32'h3ae206d6),
	.w4(32'hb942ed7d),
	.w5(32'h3b3add4b),
	.w6(32'h3a7f87b9),
	.w7(32'hba8e2824),
	.w8(32'h3b13a2ce),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba969410),
	.w1(32'hba02e1e1),
	.w2(32'hba1bed16),
	.w3(32'hba1b160d),
	.w4(32'hb85061fb),
	.w5(32'hba0ab8d1),
	.w6(32'hba727f3d),
	.w7(32'hba042032),
	.w8(32'h39c5773d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c4b92),
	.w1(32'h3b11859a),
	.w2(32'h3a01b1e7),
	.w3(32'h3ab636f0),
	.w4(32'h37a9d2ea),
	.w5(32'hbad325ed),
	.w6(32'h3b3872df),
	.w7(32'h3a815c45),
	.w8(32'hbace88e1),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa46ee),
	.w1(32'hb503db78),
	.w2(32'hb9489690),
	.w3(32'hba867506),
	.w4(32'h37d60149),
	.w5(32'hba684d6f),
	.w6(32'hba6b8717),
	.w7(32'hb93fc349),
	.w8(32'hbab0badc),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7bfd8d),
	.w1(32'hbaab2fd9),
	.w2(32'h3b19ffe3),
	.w3(32'h3c4bb529),
	.w4(32'hbbec45e6),
	.w5(32'hbb8c2748),
	.w6(32'h3c84f850),
	.w7(32'hbb20d17a),
	.w8(32'h3bfb0c96),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb28270),
	.w1(32'hbbc38a34),
	.w2(32'h3a8ac52d),
	.w3(32'h3c417aed),
	.w4(32'hbc7d31d3),
	.w5(32'hbbd64a60),
	.w6(32'h3cdf5e0f),
	.w7(32'hbb9a01de),
	.w8(32'h3bcb5ef5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca746d6),
	.w1(32'h3b1c3a05),
	.w2(32'h3c451e34),
	.w3(32'h3c5784f4),
	.w4(32'hbbb12f25),
	.w5(32'h3b84120c),
	.w6(32'h3c9d611f),
	.w7(32'h3a87ea7b),
	.w8(32'h3c56d044),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59252e),
	.w1(32'hbacb3712),
	.w2(32'hbb89bf0d),
	.w3(32'h3b5c592b),
	.w4(32'hbab3075d),
	.w5(32'hbb2938e2),
	.w6(32'h3bc6c3ce),
	.w7(32'hb8c64ba0),
	.w8(32'hba780b69),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc8f1e),
	.w1(32'h3a86d7fe),
	.w2(32'h3c473753),
	.w3(32'h3c6103dd),
	.w4(32'hbc270d04),
	.w5(32'hbad715b0),
	.w6(32'h3ca40fc9),
	.w7(32'hbaddf912),
	.w8(32'h3c31e1bb),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c152ec9),
	.w1(32'hbaa3f917),
	.w2(32'h3bec7928),
	.w3(32'h3bcf0777),
	.w4(32'hbad641d5),
	.w5(32'h3ba32ed7),
	.w6(32'h3c23f165),
	.w7(32'h3b117020),
	.w8(32'h3c22027a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb07803),
	.w1(32'hbb674a20),
	.w2(32'h3c979eec),
	.w3(32'h3c88c384),
	.w4(32'hbc3daa96),
	.w5(32'h3c3e8473),
	.w6(32'h3c75daa4),
	.w7(32'hbbebff9f),
	.w8(32'h3c826cfb),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b11b7),
	.w1(32'h388b4ff7),
	.w2(32'hb9b5931a),
	.w3(32'hb9833386),
	.w4(32'hb8dda871),
	.w5(32'h37c84c0e),
	.w6(32'h3898dbc2),
	.w7(32'h3906c483),
	.w8(32'hb98e1ab9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35fc0e),
	.w1(32'hb96bb27a),
	.w2(32'h3a1711b3),
	.w3(32'hb8a30164),
	.w4(32'h39b97639),
	.w5(32'h3a045a51),
	.w6(32'hb9acecd9),
	.w7(32'h37f24d86),
	.w8(32'h39a5b2dc),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5dc35),
	.w1(32'hbadadbb2),
	.w2(32'h3c103daf),
	.w3(32'h3c3283fc),
	.w4(32'hbb7616b8),
	.w5(32'h3c202fd3),
	.w6(32'h3c96f88d),
	.w7(32'h3ab1e6b6),
	.w8(32'h3c3e63cd),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae60e2),
	.w1(32'hbb31746a),
	.w2(32'h3c7256d7),
	.w3(32'h3c5c9611),
	.w4(32'hbba7f717),
	.w5(32'h3c92d2ef),
	.w6(32'h3c9dcf49),
	.w7(32'h3a485b99),
	.w8(32'h3ca2dbc3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cca304e),
	.w1(32'h3a8c3187),
	.w2(32'h3c3862c7),
	.w3(32'h3c58c2c7),
	.w4(32'hbc2b223e),
	.w5(32'h3b5c1d19),
	.w6(32'h3cbc8203),
	.w7(32'hbb2becf9),
	.w8(32'h3c2ad0cc),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e0532),
	.w1(32'h3a826448),
	.w2(32'h3aa81563),
	.w3(32'h3bba1efe),
	.w4(32'h3c0fbd83),
	.w5(32'h3b811d3b),
	.w6(32'hbbe368db),
	.w7(32'h3a3bdc71),
	.w8(32'h3bfdff35),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca67ad),
	.w1(32'h3a103a56),
	.w2(32'h3aa6d5be),
	.w3(32'hb7500057),
	.w4(32'h3a3b4c97),
	.w5(32'hb8b8ec38),
	.w6(32'h3a2c5671),
	.w7(32'h3a65e6d7),
	.w8(32'hb92970f5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a984a),
	.w1(32'h3a310929),
	.w2(32'hba1fd6e7),
	.w3(32'h3a739e18),
	.w4(32'h3a739eaa),
	.w5(32'h3a89d05f),
	.w6(32'h3a1db7a4),
	.w7(32'h39acf152),
	.w8(32'h3945d3ec),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd79c0b),
	.w1(32'hbbc8cb3d),
	.w2(32'h3c6527cc),
	.w3(32'h39b34446),
	.w4(32'h3c22841b),
	.w5(32'h3cbe0b0f),
	.w6(32'hbb7b202f),
	.w7(32'h3ad56406),
	.w8(32'h3c9085c1),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9acfc5),
	.w1(32'h3b3406cd),
	.w2(32'h3c967c16),
	.w3(32'h3c89637b),
	.w4(32'h3acca6eb),
	.w5(32'h3c91d075),
	.w6(32'h3c8f91af),
	.w7(32'h3c03de6d),
	.w8(32'h3ccc25d9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2fa67),
	.w1(32'h3aed5880),
	.w2(32'h3c09c4b6),
	.w3(32'hba6cc327),
	.w4(32'h3b2fe215),
	.w5(32'h3c3019d6),
	.w6(32'hbb5fe82f),
	.w7(32'h3abd8af4),
	.w8(32'h3c438497),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c464549),
	.w1(32'hbc3bc8ab),
	.w2(32'hbb4e091f),
	.w3(32'h3c2cabc6),
	.w4(32'hbc4f4aff),
	.w5(32'hbbc8087f),
	.w6(32'h3c966c6a),
	.w7(32'hbbbc531c),
	.w8(32'h390b806d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb0123c),
	.w1(32'h3af36ae9),
	.w2(32'h3c1bea1d),
	.w3(32'h3c8bbe48),
	.w4(32'hbc2c7db1),
	.w5(32'hbb96e011),
	.w6(32'h3cbdfa3c),
	.w7(32'hbb1456c2),
	.w8(32'h3be8e5b4),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba383ed2),
	.w1(32'hba4a15c2),
	.w2(32'hb9cfcdc5),
	.w3(32'hba8677d7),
	.w4(32'hb9d63f65),
	.w5(32'h38be9252),
	.w6(32'hbaa5be13),
	.w7(32'hb9997892),
	.w8(32'h3a0db30e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e092ea),
	.w1(32'hb8c744eb),
	.w2(32'hb915e1e3),
	.w3(32'h39c3c912),
	.w4(32'h39d6ccd4),
	.w5(32'h3a4e46a2),
	.w6(32'hb8cc0c6d),
	.w7(32'hb6f8cd45),
	.w8(32'h3a273e2b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e5275),
	.w1(32'hb917aaec),
	.w2(32'hbad1135e),
	.w3(32'hb9b57287),
	.w4(32'h3b3019b1),
	.w5(32'h3ae75f71),
	.w6(32'h3ac0cde9),
	.w7(32'h3b2a4654),
	.w8(32'h3a7ccb2c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b2a4a4),
	.w1(32'hba334230),
	.w2(32'hba295b24),
	.w3(32'hba07db8d),
	.w4(32'hba37167c),
	.w5(32'h3b84de78),
	.w6(32'hbae249c7),
	.w7(32'hbaba89c3),
	.w8(32'h3b6314da),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bb9be),
	.w1(32'h3c0bb2e0),
	.w2(32'h3c115e58),
	.w3(32'h3b58ac1e),
	.w4(32'h3c0e760b),
	.w5(32'h3997d55f),
	.w6(32'h3b59a2d6),
	.w7(32'h3b8022e7),
	.w8(32'hba549137),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3eebfb),
	.w1(32'h3ad3caf5),
	.w2(32'h3b5dfcf2),
	.w3(32'h3aecde86),
	.w4(32'hbc1e052d),
	.w5(32'h3bc4c4e0),
	.w6(32'h3c10f26e),
	.w7(32'hbb527daf),
	.w8(32'h3c77b396),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91184c),
	.w1(32'hb85dbb42),
	.w2(32'hb981234d),
	.w3(32'h3c27aeea),
	.w4(32'hbb94057d),
	.w5(32'hbc254526),
	.w6(32'h3c5a6f39),
	.w7(32'hbb29e024),
	.w8(32'h3b910434),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c9e03),
	.w1(32'hb9e6098d),
	.w2(32'hbc129c1e),
	.w3(32'hba5b3fb0),
	.w4(32'h3bd02ca4),
	.w5(32'h3b493c88),
	.w6(32'hbb8cdc91),
	.w7(32'hbb4e30e9),
	.w8(32'hbaadf525),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4fd3a),
	.w1(32'h3b9921fb),
	.w2(32'h3c9d5c40),
	.w3(32'h3b85ed1d),
	.w4(32'h3b8f21ef),
	.w5(32'h3c0bb061),
	.w6(32'h3b740cd1),
	.w7(32'hbb171edd),
	.w8(32'h3c877424),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd7680),
	.w1(32'hbc44fec9),
	.w2(32'hbbc0d23d),
	.w3(32'hbc25ebbb),
	.w4(32'hbc5771da),
	.w5(32'h3bc3697f),
	.w6(32'hbb4dc19a),
	.w7(32'hbc2366b5),
	.w8(32'h3c371048),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391935d7),
	.w1(32'h3b80180b),
	.w2(32'h3abd1378),
	.w3(32'h3afa09fe),
	.w4(32'h3b2c5422),
	.w5(32'hbb12940c),
	.w6(32'h3bd7dd15),
	.w7(32'h3a746c9c),
	.w8(32'hb8df0771),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00ef03),
	.w1(32'hb9e40fed),
	.w2(32'h3bbb1637),
	.w3(32'hba27f6d5),
	.w4(32'h3b87fa2f),
	.w5(32'h3b2cafc1),
	.w6(32'h3adffd24),
	.w7(32'h3bfcf8ed),
	.w8(32'h3ab4fe51),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc971c8),
	.w1(32'hbc2ca753),
	.w2(32'hbc0e4d87),
	.w3(32'hbbc9ecdf),
	.w4(32'hbbfa61d5),
	.w5(32'hbc395e72),
	.w6(32'hbc0e5b76),
	.w7(32'hbbf5a518),
	.w8(32'hbbda2435),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb23376),
	.w1(32'h3b357164),
	.w2(32'hbaf66b51),
	.w3(32'h3b54d0f5),
	.w4(32'hbb045cb6),
	.w5(32'h3b8e3244),
	.w6(32'h3c021fc7),
	.w7(32'hb81a8e5f),
	.w8(32'h3bb250e6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9af635),
	.w1(32'h3aec1393),
	.w2(32'hba28cdb9),
	.w3(32'h3acaeee0),
	.w4(32'hba73b17d),
	.w5(32'hba9e34b4),
	.w6(32'h3a838911),
	.w7(32'hbb3e5172),
	.w8(32'hba919e7a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6441dd),
	.w1(32'h3c120f50),
	.w2(32'h3b8c1b93),
	.w3(32'h3b958455),
	.w4(32'h3bb1f199),
	.w5(32'hbb109c96),
	.w6(32'h3b32715a),
	.w7(32'h3bae81ab),
	.w8(32'hbbbde6a6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b866e67),
	.w1(32'h3b5a13c8),
	.w2(32'hbabccef9),
	.w3(32'h3bb4904a),
	.w4(32'h3a3efca1),
	.w5(32'hb9231fcb),
	.w6(32'h3c5adfd4),
	.w7(32'h3b21f803),
	.w8(32'h3b9af772),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55ff2e),
	.w1(32'hbb8b377e),
	.w2(32'h3c6b8ca6),
	.w3(32'h3c04b71d),
	.w4(32'hbbf07d41),
	.w5(32'h3c10a6ac),
	.w6(32'h3b80cbad),
	.w7(32'h3b5e43c1),
	.w8(32'h3c92ea61),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c237250),
	.w1(32'h3be675fc),
	.w2(32'h3c327e3b),
	.w3(32'h3b8379f1),
	.w4(32'h3b2abd14),
	.w5(32'h3bb9ad18),
	.w6(32'h3bfad202),
	.w7(32'h3b5c3a01),
	.w8(32'h3c11308a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ac277),
	.w1(32'h3c061ac5),
	.w2(32'h3cbd5116),
	.w3(32'h3c2830af),
	.w4(32'h3bd563c6),
	.w5(32'h3c553753),
	.w6(32'h3c20638c),
	.w7(32'h3bbfc599),
	.w8(32'h3c978281),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45b52d),
	.w1(32'h3b21309f),
	.w2(32'h3b4c9699),
	.w3(32'h3b6fb4f8),
	.w4(32'hbba9adaf),
	.w5(32'hbc0e8aed),
	.w6(32'h3bb38a61),
	.w7(32'hba6fed16),
	.w8(32'hbba1ad21),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba312f),
	.w1(32'hbbe1856c),
	.w2(32'hbbe6c520),
	.w3(32'hba3a1ac1),
	.w4(32'hbaa66bbe),
	.w5(32'h3c06cd90),
	.w6(32'hbbf073f6),
	.w7(32'hbb3ee278),
	.w8(32'h3c229908),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1e5fa),
	.w1(32'hba7389df),
	.w2(32'h3a0369db),
	.w3(32'h3b7f6730),
	.w4(32'h3ae17380),
	.w5(32'hba96a810),
	.w6(32'h3a97f090),
	.w7(32'hba8fd248),
	.w8(32'hb9359436),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38dece),
	.w1(32'hba1ebcb8),
	.w2(32'hbb082b36),
	.w3(32'hba1b85a4),
	.w4(32'h3abc9117),
	.w5(32'hba3e2d17),
	.w6(32'hbae0398a),
	.w7(32'hbaa86c2b),
	.w8(32'hbb393a5b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d07b1),
	.w1(32'h3a8721df),
	.w2(32'h3c130444),
	.w3(32'h3b969ea3),
	.w4(32'hbb8395b4),
	.w5(32'hba2ae5a2),
	.w6(32'h3be9f328),
	.w7(32'hbb97216e),
	.w8(32'h3b0fd604),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbead5d4),
	.w1(32'hbbd07dc2),
	.w2(32'hbb4f3c34),
	.w3(32'hbbc5f767),
	.w4(32'hbb81d3ed),
	.w5(32'hbb199f9e),
	.w6(32'hbba9e705),
	.w7(32'hbb698eea),
	.w8(32'hbaa3b2c8),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2caa33),
	.w1(32'hbb409220),
	.w2(32'h3b5097d0),
	.w3(32'h3add7706),
	.w4(32'hbabb689e),
	.w5(32'hbb21d2e6),
	.w6(32'h3bb0f36f),
	.w7(32'h3aa7fd4b),
	.w8(32'hbad30de5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc9f39),
	.w1(32'h3bb00a40),
	.w2(32'h3c19e88e),
	.w3(32'hba1c479d),
	.w4(32'h3a8ddd8f),
	.w5(32'hbb9be8cd),
	.w6(32'hbb8749cb),
	.w7(32'h3c2fd4d5),
	.w8(32'hbba206e4),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc41ca6),
	.w1(32'h3b8d65d3),
	.w2(32'hbbfd7100),
	.w3(32'hbb7abb54),
	.w4(32'h3ba8889f),
	.w5(32'h3a1f1bbb),
	.w6(32'hbaad294f),
	.w7(32'h3b42de46),
	.w8(32'hbb681712),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39b56c),
	.w1(32'hba96989d),
	.w2(32'h3c12427d),
	.w3(32'h3bd19a26),
	.w4(32'h398b80a9),
	.w5(32'h3bb2484d),
	.w6(32'h3bc0677f),
	.w7(32'h3c54bfc4),
	.w8(32'h3b2569c4),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb12f85),
	.w1(32'h3c1061d6),
	.w2(32'h3a372f2e),
	.w3(32'h3a6a97da),
	.w4(32'h3b89a5d2),
	.w5(32'hbb4afd9e),
	.w6(32'hba8f8867),
	.w7(32'h3b09bcff),
	.w8(32'hb9d0302d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cacf595),
	.w1(32'h3c6188a7),
	.w2(32'h3cefff3b),
	.w3(32'h3c1a26ad),
	.w4(32'h3bb25443),
	.w5(32'h3b522327),
	.w6(32'h3c6f47fe),
	.w7(32'h3c68ecf1),
	.w8(32'h3c78ef7b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ff58f),
	.w1(32'h3b4b8c78),
	.w2(32'hbac29fdb),
	.w3(32'h3b96470d),
	.w4(32'h3b134b53),
	.w5(32'h3b12a637),
	.w6(32'h3a9c1f57),
	.w7(32'hba8e8fe9),
	.w8(32'h3ab096f9),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44f0ad),
	.w1(32'hbc40f622),
	.w2(32'hbc4107d5),
	.w3(32'h3c3bd9f7),
	.w4(32'hbb7374e3),
	.w5(32'hbc6d79eb),
	.w6(32'h3ca51d01),
	.w7(32'hbaf3fe34),
	.w8(32'hbcabc808),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule