module layer_10_featuremap_313(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02f0ac),
	.w1(32'h3b4ce0fc),
	.w2(32'hb9ca970b),
	.w3(32'h3858c2a8),
	.w4(32'hbb861ed5),
	.w5(32'h3afe6c1d),
	.w6(32'h3b4a79ef),
	.w7(32'hbacad98e),
	.w8(32'h3b77613d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e57f0),
	.w1(32'h3ae4c56b),
	.w2(32'h3ba4eb74),
	.w3(32'hb87f815d),
	.w4(32'h3ab15d6f),
	.w5(32'hba6d0294),
	.w6(32'h3a8c542e),
	.w7(32'h3b5c5a58),
	.w8(32'hbb42cd59),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3c2f2),
	.w1(32'h3b1c2955),
	.w2(32'hba197297),
	.w3(32'h3b271cdf),
	.w4(32'h3a96a86e),
	.w5(32'h39693e9a),
	.w6(32'h3aa05933),
	.w7(32'h3a972d23),
	.w8(32'h3a5f2173),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af55b5f),
	.w1(32'h3aa0f087),
	.w2(32'h3b5b7cc3),
	.w3(32'h3a8ad428),
	.w4(32'h39739d6a),
	.w5(32'h3b8162c3),
	.w6(32'h38b10090),
	.w7(32'h3a856969),
	.w8(32'hbbc56b57),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abda33e),
	.w1(32'h3ad31dd0),
	.w2(32'h3ab6344e),
	.w3(32'h3baaac03),
	.w4(32'h3b36536f),
	.w5(32'hbac5708f),
	.w6(32'hbbf561d0),
	.w7(32'hbc08b4a3),
	.w8(32'hbb56f93b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb491d1d),
	.w1(32'hba0e4fd9),
	.w2(32'hbafd0cb0),
	.w3(32'h3a5c3e6f),
	.w4(32'hbb0aa5ae),
	.w5(32'h3b856ff2),
	.w6(32'hbb443402),
	.w7(32'hbb241d21),
	.w8(32'hba04e0dd),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fea21),
	.w1(32'h3bc264dd),
	.w2(32'h3bcedabd),
	.w3(32'h3bc4e322),
	.w4(32'h3b80412d),
	.w5(32'h3b2751e9),
	.w6(32'h3aabf2fc),
	.w7(32'h3b2421e1),
	.w8(32'h3b61aeb9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb20aec),
	.w1(32'h3be03872),
	.w2(32'h3bae6f9f),
	.w3(32'h3b8ff4b6),
	.w4(32'h3a4de928),
	.w5(32'h3a05d45a),
	.w6(32'h3ba508eb),
	.w7(32'h3b25400d),
	.w8(32'hba8936ed),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b02aa5),
	.w1(32'h3b17b06c),
	.w2(32'h3b0b9e38),
	.w3(32'h3b26804d),
	.w4(32'h398df6c2),
	.w5(32'hbaef44d1),
	.w6(32'h3ae52446),
	.w7(32'h3ac5e865),
	.w8(32'hbb53b161),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb466ca8),
	.w1(32'hb9f0ba33),
	.w2(32'hba89f390),
	.w3(32'hb62f78ec),
	.w4(32'hbb5fc0ab),
	.w5(32'hbb794de4),
	.w6(32'hbb610d79),
	.w7(32'hbb5bddee),
	.w8(32'hbb77e8e3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a01d8),
	.w1(32'hba7ea381),
	.w2(32'hbaf36a4d),
	.w3(32'hbaa9c22f),
	.w4(32'hbb99c6f3),
	.w5(32'hbad56709),
	.w6(32'hbb816291),
	.w7(32'hbb696ed2),
	.w8(32'hbb3b5692),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ddfe4),
	.w1(32'h3b863361),
	.w2(32'hba91ab7b),
	.w3(32'hbb16502c),
	.w4(32'hbb220100),
	.w5(32'hbba26ca4),
	.w6(32'h39ac30cb),
	.w7(32'h3a02b159),
	.w8(32'hbb34c123),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380030b8),
	.w1(32'hbb62f08d),
	.w2(32'hbb5a45f3),
	.w3(32'hbba72962),
	.w4(32'hbba3dbee),
	.w5(32'hba82f93f),
	.w6(32'hbb2b3f6e),
	.w7(32'hbb456b2d),
	.w8(32'hb9d17280),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39452f2a),
	.w1(32'hba8b71a8),
	.w2(32'hb9a4a42a),
	.w3(32'hbb5a2a1a),
	.w4(32'hbb610542),
	.w5(32'h3a92efc5),
	.w6(32'hbafbe852),
	.w7(32'hbb29454c),
	.w8(32'h3aeead0c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a9320),
	.w1(32'h3b6ae2cb),
	.w2(32'h3b09b30f),
	.w3(32'h3aefb413),
	.w4(32'h3acbb800),
	.w5(32'hbb3727b4),
	.w6(32'h3aec2484),
	.w7(32'h3a9bd8b3),
	.w8(32'hbaf91bc6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f91f1),
	.w1(32'h3a085c61),
	.w2(32'hbaf412d0),
	.w3(32'hbb88084b),
	.w4(32'hbbabfd92),
	.w5(32'hb9233d98),
	.w6(32'hba046e1d),
	.w7(32'hbb0c6d0e),
	.w8(32'hb9c7278f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b248cfb),
	.w1(32'h3abb67a0),
	.w2(32'h3b2e4a6a),
	.w3(32'hb998ed0b),
	.w4(32'h3ab78d23),
	.w5(32'hb96e9273),
	.w6(32'hba972897),
	.w7(32'h3af8cb99),
	.w8(32'hba70fca4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae3448),
	.w1(32'hbae086d1),
	.w2(32'hba84cdfc),
	.w3(32'hb9618553),
	.w4(32'hba7cfdf5),
	.w5(32'hbb5866d9),
	.w6(32'hba70016e),
	.w7(32'hba794cce),
	.w8(32'h3abddd31),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba073437),
	.w1(32'hbb5bf301),
	.w2(32'hbb6e0693),
	.w3(32'hbaa79f38),
	.w4(32'h3aba7465),
	.w5(32'h398938cc),
	.w6(32'h3b1204b5),
	.w7(32'h3a80b397),
	.w8(32'hb918dd8f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf983a),
	.w1(32'hb99e216c),
	.w2(32'hbb9a63b7),
	.w3(32'hbb38e960),
	.w4(32'hbb35a817),
	.w5(32'hbad5addb),
	.w6(32'hbb2c8ffe),
	.w7(32'hbb9c671f),
	.w8(32'hb8a4462e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae64fb0),
	.w1(32'hb9e17402),
	.w2(32'hbb6d7674),
	.w3(32'hbb8274e2),
	.w4(32'hbbd216ac),
	.w5(32'h3b61e47d),
	.w6(32'hb8a36551),
	.w7(32'hbb9ca7a8),
	.w8(32'h3b160d5d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32b7eb),
	.w1(32'h3bad0f8d),
	.w2(32'h3beafafb),
	.w3(32'h3bbd96d8),
	.w4(32'h3ba67dc6),
	.w5(32'hba870761),
	.w6(32'h3b89a86b),
	.w7(32'h3b9c651a),
	.w8(32'hbac55436),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b394c11),
	.w1(32'h3b3f445b),
	.w2(32'h3b3393f4),
	.w3(32'hba9d014b),
	.w4(32'hbac56589),
	.w5(32'hbb44f3aa),
	.w6(32'h3a9bab39),
	.w7(32'h39af08ee),
	.w8(32'h3a3e9fb7),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb042058),
	.w1(32'hbb453dc8),
	.w2(32'hbb7cdbaa),
	.w3(32'hbba036ec),
	.w4(32'hbc022050),
	.w5(32'h3b359462),
	.w6(32'hbb3fcbb1),
	.w7(32'hbb9eebe2),
	.w8(32'h3a074cc5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa7032),
	.w1(32'hba599a0f),
	.w2(32'hba30f0ef),
	.w3(32'h3bb594ca),
	.w4(32'h3b9ddc53),
	.w5(32'hb991087e),
	.w6(32'h3968bb39),
	.w7(32'hbabab032),
	.w8(32'h3a1f5722),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cbf554),
	.w1(32'h3aa5042a),
	.w2(32'hb975b4b9),
	.w3(32'h3a878098),
	.w4(32'h3a0f3d73),
	.w5(32'h3b6a296e),
	.w6(32'h3aa57a84),
	.w7(32'h3972a8db),
	.w8(32'h3b2138e5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27b8b5),
	.w1(32'h3baae795),
	.w2(32'h3b36c72c),
	.w3(32'h3b97c3c9),
	.w4(32'h3b8c9202),
	.w5(32'hb7bedc35),
	.w6(32'h3bacbc3d),
	.w7(32'h3bb9d34d),
	.w8(32'hbb558f19),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0aa217),
	.w1(32'h3afe4c7e),
	.w2(32'h3aae810d),
	.w3(32'h3b0eab58),
	.w4(32'hba5241f1),
	.w5(32'h3b5f304d),
	.w6(32'hb9096928),
	.w7(32'hba66cfe4),
	.w8(32'h3991601b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba112955),
	.w1(32'hb787e529),
	.w2(32'hb9058743),
	.w3(32'h39330ee6),
	.w4(32'h3a6ee7f3),
	.w5(32'h3ab8a7fb),
	.w6(32'hbb12c205),
	.w7(32'hbb61f9eb),
	.w8(32'h3a9dd275),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b086d),
	.w1(32'h39cad7a9),
	.w2(32'hb9ce4b57),
	.w3(32'hba3c416d),
	.w4(32'hba94797d),
	.w5(32'hbb2dc1f4),
	.w6(32'hb9518b01),
	.w7(32'hb9f019e5),
	.w8(32'hbb425c25),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf23ff2),
	.w1(32'hbc0bf46b),
	.w2(32'hbbd01182),
	.w3(32'h36b0c31c),
	.w4(32'h3ab88a5c),
	.w5(32'hbb988896),
	.w6(32'hbbe43876),
	.w7(32'hbb9be97b),
	.w8(32'hbb4f0ac1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf062d8),
	.w1(32'hbb88e673),
	.w2(32'hb9fe1308),
	.w3(32'hbb8c81e8),
	.w4(32'hbb247bd2),
	.w5(32'h3a820585),
	.w6(32'hbb39558f),
	.w7(32'hbb0b8774),
	.w8(32'h3b612110),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb975b0d),
	.w1(32'hbbd54586),
	.w2(32'hbaaf05d2),
	.w3(32'h3b263537),
	.w4(32'h3ba60cf0),
	.w5(32'hb9a8c3fa),
	.w6(32'hbaf76411),
	.w7(32'h37e8424f),
	.w8(32'hbad9af44),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb252eef),
	.w1(32'hbaefeba2),
	.w2(32'hbafa81d6),
	.w3(32'hbaaa8d8e),
	.w4(32'hbb19de59),
	.w5(32'h3b79ecdf),
	.w6(32'hbadda787),
	.w7(32'hbb1fd29d),
	.w8(32'h3abdcb0c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed1f5a),
	.w1(32'hb90f8a94),
	.w2(32'h3929046a),
	.w3(32'h3b1cfb6d),
	.w4(32'h3a737359),
	.w5(32'hbb79176b),
	.w6(32'h3ae31cc2),
	.w7(32'h3b025bd9),
	.w8(32'hbb90c181),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49a598),
	.w1(32'hbb21311e),
	.w2(32'hbb045ea0),
	.w3(32'hbaca444e),
	.w4(32'hbab43bc0),
	.w5(32'h3ad7c155),
	.w6(32'hbb49325c),
	.w7(32'hbb368ce5),
	.w8(32'h3ab31c04),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4d279),
	.w1(32'hba947b05),
	.w2(32'hbad7924f),
	.w3(32'h3b56c531),
	.w4(32'h3b22b39a),
	.w5(32'hbaf44997),
	.w6(32'hba9b0244),
	.w7(32'h391a6092),
	.w8(32'h3ab95e85),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fcdb5),
	.w1(32'h3b741501),
	.w2(32'hbaaef29a),
	.w3(32'h3ac0a3fa),
	.w4(32'hbb1aa587),
	.w5(32'hbb9566bd),
	.w6(32'h3bb22233),
	.w7(32'h3ae3e325),
	.w8(32'hbbae9bb9),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63dbdb),
	.w1(32'hba1d5489),
	.w2(32'hba10a210),
	.w3(32'hbb4fbd6d),
	.w4(32'hbb3524bc),
	.w5(32'h3a93e10d),
	.w6(32'hbbe1984b),
	.w7(32'hbba20f9c),
	.w8(32'h3b52dd64),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9660e),
	.w1(32'h3b91674d),
	.w2(32'h3b3fff83),
	.w3(32'h3b1fea07),
	.w4(32'hbafad2a7),
	.w5(32'hbae605fb),
	.w6(32'h3b599c8e),
	.w7(32'h3b26bb2a),
	.w8(32'hbb33660c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b2e68),
	.w1(32'hbb106f5f),
	.w2(32'hba9476d6),
	.w3(32'hbabf3db3),
	.w4(32'hba8069bd),
	.w5(32'h3b5b4169),
	.w6(32'hbada16b4),
	.w7(32'hba9bd53e),
	.w8(32'h39143b87),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dee4f),
	.w1(32'h3bce86ed),
	.w2(32'h3bd270c0),
	.w3(32'h3b91f6d8),
	.w4(32'h3b8a36af),
	.w5(32'hbbbbd1eb),
	.w6(32'h3b168279),
	.w7(32'h3b42b5cc),
	.w8(32'hbb11c293),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dece4),
	.w1(32'hbb5b9337),
	.w2(32'hbb79446a),
	.w3(32'hbb93c030),
	.w4(32'hbbb34487),
	.w5(32'hbb17a656),
	.w6(32'h39e7b0c5),
	.w7(32'hba78097f),
	.w8(32'hbb20dc36),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab25cdb),
	.w1(32'hbb61bd5f),
	.w2(32'hb90d9739),
	.w3(32'h3a12e844),
	.w4(32'h3b0f8782),
	.w5(32'h3a05284c),
	.w6(32'hba434cdd),
	.w7(32'h3b0f73f8),
	.w8(32'hbad1a637),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66f309),
	.w1(32'h39d6309c),
	.w2(32'h3b9ff417),
	.w3(32'h3abcbadf),
	.w4(32'h3a8158b5),
	.w5(32'hbb1b5d15),
	.w6(32'hba901384),
	.w7(32'h3a5ce4a3),
	.w8(32'hbaca4ebf),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41af82),
	.w1(32'hbada447a),
	.w2(32'hbaad50fb),
	.w3(32'hbbce54e5),
	.w4(32'hbb4119af),
	.w5(32'h3a22a60b),
	.w6(32'hbbbbb721),
	.w7(32'hbb3be1cd),
	.w8(32'hba272103),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61237a),
	.w1(32'hba136a29),
	.w2(32'hbb073d45),
	.w3(32'hba5390dc),
	.w4(32'hba38a90c),
	.w5(32'h3ae2f688),
	.w6(32'hbb22625f),
	.w7(32'hbb42b829),
	.w8(32'h3a85e19f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ea87d),
	.w1(32'h3b63db9e),
	.w2(32'h3b8d828e),
	.w3(32'h3b58081d),
	.w4(32'h3b2a5af4),
	.w5(32'hbb5ff6f3),
	.w6(32'h3b23be94),
	.w7(32'h3b212d50),
	.w8(32'hbb0a86e0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb008347),
	.w1(32'hbb20d4e2),
	.w2(32'hbb17a7dc),
	.w3(32'hbae56ca6),
	.w4(32'hbb15f787),
	.w5(32'h3ba60b8d),
	.w6(32'hba8396c5),
	.w7(32'hbadbcb24),
	.w8(32'h3af7a893),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fc772),
	.w1(32'h3c0317fc),
	.w2(32'h3bff575f),
	.w3(32'h3bff26f3),
	.w4(32'h3b9633b5),
	.w5(32'h3bbcf084),
	.w6(32'h3bc4ed63),
	.w7(32'h3b57f199),
	.w8(32'h3bcd863b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1adf20),
	.w1(32'h38cec929),
	.w2(32'hb91e55bb),
	.w3(32'h3bf93ad2),
	.w4(32'h3b9c9a79),
	.w5(32'h38f7fc53),
	.w6(32'h3b415a4e),
	.w7(32'h3a34c55c),
	.w8(32'h3a8b8ced),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9365b65),
	.w1(32'hba9fa6b5),
	.w2(32'h3aadcb02),
	.w3(32'hba475f59),
	.w4(32'hba228fb3),
	.w5(32'hba450fe9),
	.w6(32'hb94b841f),
	.w7(32'h3a1e2268),
	.w8(32'hb96e5f57),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5691ec),
	.w1(32'hbb1c5b11),
	.w2(32'hbb038291),
	.w3(32'hbab8ca87),
	.w4(32'hba169ed5),
	.w5(32'h3bb14043),
	.w6(32'hba5b21ef),
	.w7(32'hba540bde),
	.w8(32'h3b2cba02),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e7c27),
	.w1(32'h3ba35f79),
	.w2(32'hbb59a6ab),
	.w3(32'hba11a897),
	.w4(32'hbb946a8c),
	.w5(32'hba4f07f0),
	.w6(32'h399c351c),
	.w7(32'hbbd3b954),
	.w8(32'hba89759f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab60e9e),
	.w1(32'hbac70117),
	.w2(32'hbb3e1b9d),
	.w3(32'hbb22fd6f),
	.w4(32'hbaaff307),
	.w5(32'h3aaed917),
	.w6(32'hbb10ab90),
	.w7(32'hbb08040c),
	.w8(32'hbaf1e606),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57739c),
	.w1(32'hbb58ae60),
	.w2(32'hbb038f96),
	.w3(32'h371ec43d),
	.w4(32'hba7204cb),
	.w5(32'hbae3d712),
	.w6(32'hbb2f8129),
	.w7(32'hbab3517c),
	.w8(32'hbacd83c3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae21a1e),
	.w1(32'hbb2a60ab),
	.w2(32'hbb2f5f7e),
	.w3(32'hbb28abb4),
	.w4(32'hbb153715),
	.w5(32'h3b5774bb),
	.w6(32'hbad750a3),
	.w7(32'hbb1af6dd),
	.w8(32'h3b64c7ba),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a5293),
	.w1(32'h3b1e51b4),
	.w2(32'hbb74a140),
	.w3(32'hba456f79),
	.w4(32'hbb8073b3),
	.w5(32'h3bc74e80),
	.w6(32'h38958075),
	.w7(32'hbb5c9c56),
	.w8(32'h3abfca9e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b715aa1),
	.w1(32'h3c12f4ed),
	.w2(32'h3c0f212a),
	.w3(32'h3c0dcef7),
	.w4(32'h3b94bf20),
	.w5(32'h3b8847f1),
	.w6(32'h3be72c92),
	.w7(32'h3b89410a),
	.w8(32'hba0c85f7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7808c14),
	.w1(32'h38052ee2),
	.w2(32'h3b5b8c4b),
	.w3(32'h3c03b2b3),
	.w4(32'h3c33fc99),
	.w5(32'hbb04fae4),
	.w6(32'h3a8332ff),
	.w7(32'h3b5307b8),
	.w8(32'hbae72ff7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e0644),
	.w1(32'h3b12ce2e),
	.w2(32'h3a5541ad),
	.w3(32'hba8e8e40),
	.w4(32'h393b71a8),
	.w5(32'h39be36f5),
	.w6(32'hbb2f8f08),
	.w7(32'hbb05a526),
	.w8(32'hb9ed77b1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8095cb),
	.w1(32'h3a5a4fa1),
	.w2(32'h3a6465ff),
	.w3(32'h3a21efb9),
	.w4(32'hb9cb5994),
	.w5(32'h3ba36a19),
	.w6(32'hbade3a40),
	.w7(32'hbb1c7c80),
	.w8(32'h39a23374),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82eea1),
	.w1(32'h39ea1ad0),
	.w2(32'h392430d6),
	.w3(32'h3be4bd0e),
	.w4(32'h3bc3b193),
	.w5(32'h3a738680),
	.w6(32'h3af20349),
	.w7(32'h3a5fa6ea),
	.w8(32'hb8fc271f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902e696),
	.w1(32'hb9c8aca1),
	.w2(32'hb9e8436c),
	.w3(32'hb967ee97),
	.w4(32'hbabb5a18),
	.w5(32'h3aff2c74),
	.w6(32'hb9236502),
	.w7(32'hba4d0ddb),
	.w8(32'h3b1c0d77),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac441f9),
	.w1(32'hba2826d8),
	.w2(32'hbb19a84c),
	.w3(32'hbae52b57),
	.w4(32'hbaeeef66),
	.w5(32'hba313188),
	.w6(32'hba9d5027),
	.w7(32'hbadd2e2d),
	.w8(32'hbb86aba6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bf575),
	.w1(32'hbb8c27f7),
	.w2(32'hbbc0aaab),
	.w3(32'h38ea4286),
	.w4(32'h39a2f302),
	.w5(32'hba1c9593),
	.w6(32'hbb2f4f05),
	.w7(32'hbb8af9c9),
	.w8(32'h3a5d38c4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7852a9),
	.w1(32'h3b82fc28),
	.w2(32'hb908b44f),
	.w3(32'hba5c1c7b),
	.w4(32'hbb07fa41),
	.w5(32'h3b40bfdd),
	.w6(32'h3a8ee25f),
	.w7(32'hba0537c9),
	.w8(32'h3b4094e0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83689b),
	.w1(32'h3ba205b7),
	.w2(32'h3bd0f510),
	.w3(32'h3b83b54a),
	.w4(32'h3bc891de),
	.w5(32'h3b4dc9e7),
	.w6(32'h3bb85fcb),
	.w7(32'h3bf38124),
	.w8(32'h3b993c43),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06931b),
	.w1(32'h3b074ee3),
	.w2(32'h3b22d4a3),
	.w3(32'h3aab2e49),
	.w4(32'h390bab95),
	.w5(32'hbb41a50d),
	.w6(32'h3ac08124),
	.w7(32'h3959b994),
	.w8(32'hbb889772),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37b2b4),
	.w1(32'hbb405024),
	.w2(32'hba6380c1),
	.w3(32'hbb1ed85c),
	.w4(32'hbb1611cf),
	.w5(32'hba587186),
	.w6(32'hbb51edf0),
	.w7(32'hba514abc),
	.w8(32'h3a39acc5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a92aa),
	.w1(32'hb9bdc197),
	.w2(32'hb9c9346c),
	.w3(32'h3a861d97),
	.w4(32'h3aba426f),
	.w5(32'hbaf92447),
	.w6(32'h3af56fff),
	.w7(32'h3aee14a1),
	.w8(32'h3aaee46e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadfa27),
	.w1(32'h3b1f5033),
	.w2(32'hbaaf9886),
	.w3(32'hba958d3f),
	.w4(32'hbabf35cc),
	.w5(32'hbb2dfe17),
	.w6(32'h3a3cffbb),
	.w7(32'hbb196ca4),
	.w8(32'hbb00e9fe),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb351bc5),
	.w1(32'hbb54e22b),
	.w2(32'hbb5cd85a),
	.w3(32'hb9d92a9e),
	.w4(32'hbad31418),
	.w5(32'h3828474f),
	.w6(32'hba73728c),
	.w7(32'hbaa1875c),
	.w8(32'h39e4f15c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e9bc7),
	.w1(32'hba5a8931),
	.w2(32'hba2245e0),
	.w3(32'hbaa8c4e7),
	.w4(32'hba5cea56),
	.w5(32'hbb0f0f94),
	.w6(32'hbae27e3f),
	.w7(32'hba4da2ee),
	.w8(32'h3873320c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e8bc5),
	.w1(32'h3b8a5403),
	.w2(32'hbb070efd),
	.w3(32'hbb4ee310),
	.w4(32'hbbbf5687),
	.w5(32'hbb604fe9),
	.w6(32'h3a2601b0),
	.w7(32'hbabe0a1f),
	.w8(32'hbad177fb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bca72),
	.w1(32'hbb832d79),
	.w2(32'hbb5a8938),
	.w3(32'hbb551ecc),
	.w4(32'hbb2d2c4e),
	.w5(32'hbb31a555),
	.w6(32'hbb0b833b),
	.w7(32'hbafde204),
	.w8(32'hbb7f179f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35e404),
	.w1(32'hbb4a9bc5),
	.w2(32'hbb436512),
	.w3(32'hba851e07),
	.w4(32'hba36106e),
	.w5(32'hb9f7e14a),
	.w6(32'hbad319eb),
	.w7(32'hbb21d161),
	.w8(32'hbb6d7bbd),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb021022),
	.w1(32'hbac6aeae),
	.w2(32'hb9949e94),
	.w3(32'hba9f3734),
	.w4(32'hba969b65),
	.w5(32'hbb616f33),
	.w6(32'hbb9c4bf2),
	.w7(32'hbb872314),
	.w8(32'hbb02cd27),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dadd8),
	.w1(32'hbb2a2fc1),
	.w2(32'hbb6961dc),
	.w3(32'hbb5c437e),
	.w4(32'hbb09f57a),
	.w5(32'h39cae35a),
	.w6(32'hbb1fbafb),
	.w7(32'hbb013541),
	.w8(32'hbadfd9f3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932ad9b),
	.w1(32'h3a848669),
	.w2(32'h39edcad2),
	.w3(32'h3ac45249),
	.w4(32'h3a48549d),
	.w5(32'h3ad434c9),
	.w6(32'hbb6e3f7f),
	.w7(32'hbae3c891),
	.w8(32'h3b4f0fd1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9dba4d),
	.w1(32'h3b7cb837),
	.w2(32'h3a8fb1d4),
	.w3(32'h3aa67224),
	.w4(32'hbaa5a91a),
	.w5(32'hbac12da2),
	.w6(32'h3b90d195),
	.w7(32'h39e60143),
	.w8(32'hbb0f958d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3046df),
	.w1(32'hbb2b1d4a),
	.w2(32'hbb4131d8),
	.w3(32'hba90b9dd),
	.w4(32'hbadb9141),
	.w5(32'hba44571e),
	.w6(32'hbb0503e2),
	.w7(32'hbb186490),
	.w8(32'hbab49c56),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28538c),
	.w1(32'hba5065a7),
	.w2(32'hbac3e0c0),
	.w3(32'hb9858b27),
	.w4(32'hbb248098),
	.w5(32'h3afc1119),
	.w6(32'hbb163c5d),
	.w7(32'hbb17531d),
	.w8(32'h3b5f9234),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13ba4d),
	.w1(32'h3bcb0452),
	.w2(32'h3b842378),
	.w3(32'hbb41af6c),
	.w4(32'hb8a0072e),
	.w5(32'hbb0181e0),
	.w6(32'h3af8dd07),
	.w7(32'h3bcf74da),
	.w8(32'hbb525770),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5dedb4),
	.w1(32'hb9ffc70d),
	.w2(32'hbaa28ec4),
	.w3(32'hbb08803b),
	.w4(32'hbb0573d4),
	.w5(32'hbbaa9ad6),
	.w6(32'hbb1129d7),
	.w7(32'hbb104320),
	.w8(32'hbbbfe287),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb820e8d),
	.w1(32'hbb88508d),
	.w2(32'hbb8afe0f),
	.w3(32'hbb926e64),
	.w4(32'hbb80a2e7),
	.w5(32'h3bd2faac),
	.w6(32'hbbb80ae7),
	.w7(32'hbb8d4cc1),
	.w8(32'h3b016e3d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b768438),
	.w1(32'h3c1dc8a0),
	.w2(32'h3a7b4b7e),
	.w3(32'h3b899963),
	.w4(32'hb998b556),
	.w5(32'h3b27a1d7),
	.w6(32'h3b1b8ffa),
	.w7(32'h39b86324),
	.w8(32'hb9c90345),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fa531),
	.w1(32'hba1d2da9),
	.w2(32'hbab71bc8),
	.w3(32'h3b5489cd),
	.w4(32'h3b42d61e),
	.w5(32'h3b8f00c6),
	.w6(32'h38765e75),
	.w7(32'hba7d18b8),
	.w8(32'h3a2c2039),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b220542),
	.w1(32'h3b985919),
	.w2(32'h3ba919ca),
	.w3(32'h3bbc782a),
	.w4(32'h3b9e9497),
	.w5(32'hbad5608c),
	.w6(32'h3ae5b7bc),
	.w7(32'h3b2c0b66),
	.w8(32'hba0b5a8a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb015ac3),
	.w1(32'hbb42ba2b),
	.w2(32'h3a926789),
	.w3(32'hbaac0b22),
	.w4(32'hbab6d992),
	.w5(32'hbb4c0133),
	.w6(32'hbb0a976c),
	.w7(32'h3a9133b8),
	.w8(32'h38ee4ad4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a887c),
	.w1(32'hb8fb7020),
	.w2(32'h3911471b),
	.w3(32'hbb5a65be),
	.w4(32'hbbba84b2),
	.w5(32'h3acfb829),
	.w6(32'hbaea4be1),
	.w7(32'hbb029ae7),
	.w8(32'h39b00870),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd5218),
	.w1(32'hbb53f10c),
	.w2(32'h38f7183d),
	.w3(32'h386b7d6f),
	.w4(32'hbad72712),
	.w5(32'hb9f5dbad),
	.w6(32'hbb2a430e),
	.w7(32'hbaf4e47c),
	.w8(32'hbb8fa4ec),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd8787),
	.w1(32'h39de2f10),
	.w2(32'h3be70ceb),
	.w3(32'h397cefc6),
	.w4(32'h3b379455),
	.w5(32'h3a838ff8),
	.w6(32'hbb749046),
	.w7(32'hba769277),
	.w8(32'h3b5df376),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3796b2b4),
	.w1(32'h3a922267),
	.w2(32'h39a96c8b),
	.w3(32'h39e4f32f),
	.w4(32'hb83f6345),
	.w5(32'hbb53d96a),
	.w6(32'h3b404dcd),
	.w7(32'h3ae9b9c2),
	.w8(32'hba3cdaa6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6977d9),
	.w1(32'h3a92ac6a),
	.w2(32'hbaa26b0c),
	.w3(32'hbab65c6b),
	.w4(32'hbb959cbd),
	.w5(32'hbb654759),
	.w6(32'hb9169a1b),
	.w7(32'hbb0d931b),
	.w8(32'h39e44a85),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95afd9),
	.w1(32'h3bbc705a),
	.w2(32'h3a22d7e2),
	.w3(32'hbaeb4c00),
	.w4(32'h39c2f73b),
	.w5(32'hba99c020),
	.w6(32'h3ba2307b),
	.w7(32'h3bb17606),
	.w8(32'hbac3a6ea),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb90f6),
	.w1(32'hba2b2f97),
	.w2(32'h3aca79ec),
	.w3(32'h37723a4d),
	.w4(32'hba3ada71),
	.w5(32'hbb826876),
	.w6(32'hbac02e4c),
	.w7(32'h398129da),
	.w8(32'hbb47c492),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacdcff),
	.w1(32'hbbb4a93d),
	.w2(32'h3ad1d861),
	.w3(32'h3ab835c5),
	.w4(32'h3b833552),
	.w5(32'h3b048410),
	.w6(32'hbb016b48),
	.w7(32'h3af4c5aa),
	.w8(32'h3aa49536),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fa1c5),
	.w1(32'h3a746089),
	.w2(32'h3a87e02f),
	.w3(32'h3a5a9b03),
	.w4(32'hbaade921),
	.w5(32'hba3fc14e),
	.w6(32'h3ace974b),
	.w7(32'h3917e4d1),
	.w8(32'h3ab51df4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5a726),
	.w1(32'hba081bce),
	.w2(32'hbb0d3a8b),
	.w3(32'hba3c6aa2),
	.w4(32'hbad73a99),
	.w5(32'hbba05688),
	.w6(32'h39c95c9d),
	.w7(32'hbb23c552),
	.w8(32'hbb1fa05c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6492c4),
	.w1(32'hbb1c070c),
	.w2(32'hbb2542b4),
	.w3(32'hbb8dfb78),
	.w4(32'hbb8b3d75),
	.w5(32'hbc08b8bd),
	.w6(32'hbabdba9b),
	.w7(32'hbb25fd05),
	.w8(32'hbb83de84),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4f483),
	.w1(32'h3b6e9063),
	.w2(32'h3aa077b1),
	.w3(32'hbb88e115),
	.w4(32'hbb112da7),
	.w5(32'h3b36ffe3),
	.w6(32'h3b097abb),
	.w7(32'h3bb4a681),
	.w8(32'h3b59cfb4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b941b82),
	.w1(32'h3b0d573e),
	.w2(32'hbac914ec),
	.w3(32'h3b3e20f7),
	.w4(32'hbaedcac1),
	.w5(32'hbb8db714),
	.w6(32'h3b66331a),
	.w7(32'hba9e7f04),
	.w8(32'hbba1fab8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c8142),
	.w1(32'hbb3c2f94),
	.w2(32'hbaa91719),
	.w3(32'hbb8b0d25),
	.w4(32'hbbbf1472),
	.w5(32'h3923e812),
	.w6(32'hbb870ad2),
	.w7(32'hbb2e0864),
	.w8(32'h39af3983),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c1ae9),
	.w1(32'hbad6cd1e),
	.w2(32'hbb510c48),
	.w3(32'hbac5a024),
	.w4(32'hbb1f64da),
	.w5(32'h399815b3),
	.w6(32'hba1cd579),
	.w7(32'hbb2586ce),
	.w8(32'h3a124186),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e3b99),
	.w1(32'hba5fb7d6),
	.w2(32'hb95d913a),
	.w3(32'h3a2d7389),
	.w4(32'h3af62265),
	.w5(32'hbab4987c),
	.w6(32'hba7ebaa4),
	.w7(32'h3a937054),
	.w8(32'hbab11820),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2c138),
	.w1(32'hb8c412bb),
	.w2(32'hba1026ff),
	.w3(32'hb958dd77),
	.w4(32'hbae9103a),
	.w5(32'hbb02d25e),
	.w6(32'h3aeef457),
	.w7(32'h39aeae3d),
	.w8(32'h3ab0fb37),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab30b24),
	.w1(32'h3af83dc0),
	.w2(32'hb977f900),
	.w3(32'hbb28e1b0),
	.w4(32'hbb31bfa5),
	.w5(32'hb9b2fe48),
	.w6(32'h3b808c91),
	.w7(32'h3a37a6e4),
	.w8(32'hba4d6fae),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a663db2),
	.w1(32'h398e27c3),
	.w2(32'h399060b5),
	.w3(32'hbaa395ef),
	.w4(32'hbb3f5f9a),
	.w5(32'hbb0f9cf8),
	.w6(32'hba59f546),
	.w7(32'hba9733ed),
	.w8(32'h388c9461),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b059fb3),
	.w1(32'h39b24e3e),
	.w2(32'h3ac24222),
	.w3(32'hbad373bc),
	.w4(32'hbb8aa0ee),
	.w5(32'hbb4d40cc),
	.w6(32'h3b25e1e4),
	.w7(32'h3b6e9ba5),
	.w8(32'hbad74079),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983d273),
	.w1(32'h3a3d97bb),
	.w2(32'h3a5aa41b),
	.w3(32'hbb0a642c),
	.w4(32'hba8f44c8),
	.w5(32'h3b839511),
	.w6(32'h3b5e2343),
	.w7(32'h3b45e5c0),
	.w8(32'h3b36d434),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a1b7d),
	.w1(32'h3b5b83bd),
	.w2(32'h3a9f43f0),
	.w3(32'hbaa8a469),
	.w4(32'hbaf3ec80),
	.w5(32'h3bda4dca),
	.w6(32'h3ac57d3f),
	.w7(32'hb94b57c0),
	.w8(32'h3b3683e9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba63b5e),
	.w1(32'h3b232c1b),
	.w2(32'h3b663856),
	.w3(32'h3bf84011),
	.w4(32'h3bc3c50b),
	.w5(32'h39e7615d),
	.w6(32'h3ab06b90),
	.w7(32'h3b8de0cb),
	.w8(32'h3b0713eb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05d732),
	.w1(32'h3b7bf6fc),
	.w2(32'h3ba735db),
	.w3(32'hbaeefb3c),
	.w4(32'h3a4182eb),
	.w5(32'hbad8eea0),
	.w6(32'h3ab7618e),
	.w7(32'h35f78a83),
	.w8(32'hba93f291),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c7cc7),
	.w1(32'hbabbeb7c),
	.w2(32'h3ab2c90f),
	.w3(32'hbb40fdb4),
	.w4(32'hb9e6b4d1),
	.w5(32'h3b4c5cf2),
	.w6(32'hba8fd418),
	.w7(32'hbb4a2042),
	.w8(32'h3b59b9f0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8289c),
	.w1(32'h3b333b74),
	.w2(32'h3b0c22ca),
	.w3(32'hbae7907f),
	.w4(32'hbb36889c),
	.w5(32'h3b131b00),
	.w6(32'h3a88739e),
	.w7(32'h3a82c999),
	.w8(32'h3b394a3e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a833c3d),
	.w1(32'h3b95e3e1),
	.w2(32'h3b9f5159),
	.w3(32'h3b63151c),
	.w4(32'h3b90742d),
	.w5(32'hb8a05323),
	.w6(32'h3b7cafec),
	.w7(32'h3b4fd50c),
	.w8(32'h3abea571),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39672d1a),
	.w1(32'h3ad8fd64),
	.w2(32'h398f70f8),
	.w3(32'hbb02a72a),
	.w4(32'hbb2acaca),
	.w5(32'h3b79b981),
	.w6(32'hb98c9dea),
	.w7(32'hbb272918),
	.w8(32'h38320343),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97e6ac),
	.w1(32'h3afd0d86),
	.w2(32'hba6905cb),
	.w3(32'h3b812cfc),
	.w4(32'h3aab5ef3),
	.w5(32'hbb286622),
	.w6(32'h3ac1a557),
	.w7(32'hba73e2d4),
	.w8(32'hbb9a25d0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb52f6),
	.w1(32'hbb29e219),
	.w2(32'h39bcfe96),
	.w3(32'hbb78b94e),
	.w4(32'hbb1c9f5b),
	.w5(32'h3c22f34e),
	.w6(32'hbb6c8a77),
	.w7(32'hb9a468f8),
	.w8(32'h3ba0ff2a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dc3e3),
	.w1(32'h3ade304c),
	.w2(32'hb9f8dd63),
	.w3(32'h3a8fb0e8),
	.w4(32'hbb684b46),
	.w5(32'h3b3f0f42),
	.w6(32'hb9cb29e6),
	.w7(32'hbb476ad6),
	.w8(32'h3ac4a5a3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06b4e4),
	.w1(32'h3a81644e),
	.w2(32'hbbbcd56b),
	.w3(32'h3b92aceb),
	.w4(32'h3af87521),
	.w5(32'hba5beb33),
	.w6(32'hbb1e421b),
	.w7(32'hbb393afb),
	.w8(32'hbbbfb812),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33e280),
	.w1(32'hba75775f),
	.w2(32'h3bbaddb7),
	.w3(32'h3b410212),
	.w4(32'hbb89ab23),
	.w5(32'h3b49edc5),
	.w6(32'h3ba714b0),
	.w7(32'h3c0c8b9a),
	.w8(32'h3ae9cf9f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa471f5),
	.w1(32'hbba52c14),
	.w2(32'h3ad70831),
	.w3(32'h3b56412f),
	.w4(32'h3baf298d),
	.w5(32'hba8d8311),
	.w6(32'h3b3d0d22),
	.w7(32'h3c170f41),
	.w8(32'hbb7661e8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfc7f5),
	.w1(32'h3b5564fd),
	.w2(32'h3bcbff5d),
	.w3(32'h3afd0e5e),
	.w4(32'hbad8fa49),
	.w5(32'h3a059974),
	.w6(32'h3b9c6d11),
	.w7(32'h3a7427a3),
	.w8(32'h3aef1d74),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b335bfb),
	.w1(32'hba9c1ab5),
	.w2(32'hbac9b6a3),
	.w3(32'h3a97d985),
	.w4(32'h39d9014a),
	.w5(32'hbb3ea270),
	.w6(32'h3ba47de0),
	.w7(32'h3b806042),
	.w8(32'h3acfeb11),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84247b),
	.w1(32'hbb0aad1d),
	.w2(32'h3a35fb58),
	.w3(32'hbb0ebe85),
	.w4(32'hbb9802a1),
	.w5(32'hbaa17a32),
	.w6(32'h3bbafe9f),
	.w7(32'h3b6d5c72),
	.w8(32'hbb46801d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96e3c3),
	.w1(32'hbb201cb6),
	.w2(32'hba8d3840),
	.w3(32'hbae63c2b),
	.w4(32'hba2069f9),
	.w5(32'h3b51f2ed),
	.w6(32'hba9da122),
	.w7(32'hbb8421a5),
	.w8(32'h3b383f31),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddbf0f),
	.w1(32'h3b1ca8ed),
	.w2(32'h3b9369f0),
	.w3(32'h3b81e0d3),
	.w4(32'hbac554bc),
	.w5(32'h3bbf6c81),
	.w6(32'hb943476b),
	.w7(32'h3b351c66),
	.w8(32'hb900f451),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813e1d),
	.w1(32'hbac4aae1),
	.w2(32'h3b5e06d5),
	.w3(32'h3ba9b7f9),
	.w4(32'h3bda27fd),
	.w5(32'hb8bd06d9),
	.w6(32'h3baef17a),
	.w7(32'h3b66b653),
	.w8(32'h3b8290e8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb777d477),
	.w1(32'h3aed28d6),
	.w2(32'h3ad0375e),
	.w3(32'h3a21327e),
	.w4(32'hbb3be809),
	.w5(32'hbaf2ba29),
	.w6(32'h3b900452),
	.w7(32'h3aa03394),
	.w8(32'h3a5ba38a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a184800),
	.w1(32'h37877c01),
	.w2(32'hb8232741),
	.w3(32'hbb4eb23b),
	.w4(32'hbb003c5a),
	.w5(32'hbba84ab9),
	.w6(32'h3a3e68cc),
	.w7(32'h3a11471f),
	.w8(32'hbc267dae),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc0847),
	.w1(32'hbaf73c44),
	.w2(32'h3a3869c5),
	.w3(32'hbb789c47),
	.w4(32'hbc03b839),
	.w5(32'hbb18ad37),
	.w6(32'hbb67e15d),
	.w7(32'h39938982),
	.w8(32'h3a8625cb),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53d057),
	.w1(32'h3b233eec),
	.w2(32'h3a9a6457),
	.w3(32'hba8f8416),
	.w4(32'hbb9def69),
	.w5(32'hbb0b2584),
	.w6(32'h3baaf034),
	.w7(32'h3b09b30b),
	.w8(32'h3aac3766),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9a12a),
	.w1(32'h3aed178a),
	.w2(32'h3b7f5fde),
	.w3(32'hbb41bbb3),
	.w4(32'h3a11bf93),
	.w5(32'hba388fc0),
	.w6(32'h3b3e9470),
	.w7(32'h3b088262),
	.w8(32'h3b9c61cd),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d805f),
	.w1(32'h3c380669),
	.w2(32'h3b493d3b),
	.w3(32'hbadd6d2c),
	.w4(32'hbbbe6b2a),
	.w5(32'h3b98e8e1),
	.w6(32'h3b248bb0),
	.w7(32'hba55b16b),
	.w8(32'h3b9cb5a6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be124e2),
	.w1(32'h3bdd909d),
	.w2(32'h3c060c02),
	.w3(32'h3b8822dd),
	.w4(32'h3bd910fe),
	.w5(32'hbb1a5aed),
	.w6(32'h3b7f8f61),
	.w7(32'h3bd40caa),
	.w8(32'h38a5700a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f449e9),
	.w1(32'hba207019),
	.w2(32'h399f911a),
	.w3(32'hba960c46),
	.w4(32'hbb7b9b74),
	.w5(32'hbb24123f),
	.w6(32'h3b7bda1a),
	.w7(32'h3b893ea1),
	.w8(32'h38a5b654),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b318aa6),
	.w1(32'h3b2d9f09),
	.w2(32'h3a628fba),
	.w3(32'hbaff5fad),
	.w4(32'hbb810a9a),
	.w5(32'h3adf07ab),
	.w6(32'h3ba3d60b),
	.w7(32'h3b1acc6a),
	.w8(32'hba752d2a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafbee1),
	.w1(32'h3a61309d),
	.w2(32'hba88777b),
	.w3(32'hba665b61),
	.w4(32'hbb272f88),
	.w5(32'hba6a3de3),
	.w6(32'hba85b9d4),
	.w7(32'hbb8464a4),
	.w8(32'hbba06e6b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0eae4),
	.w1(32'hbc075da8),
	.w2(32'hbbb97d3c),
	.w3(32'h39eb6fcd),
	.w4(32'hb9c822b0),
	.w5(32'h3c2a637f),
	.w6(32'hbb978a43),
	.w7(32'hba59d5a9),
	.w8(32'h3ba1a895),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16af32),
	.w1(32'hbabd95fb),
	.w2(32'hbb2403c2),
	.w3(32'h3bd95224),
	.w4(32'h3b236ae3),
	.w5(32'hbb81789b),
	.w6(32'h3b8f6b2a),
	.w7(32'h3a010cbc),
	.w8(32'hbb109b76),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cfd59),
	.w1(32'hbae10b4b),
	.w2(32'hba970624),
	.w3(32'hbb65ba44),
	.w4(32'hbaa2cd54),
	.w5(32'hbae78654),
	.w6(32'h39febe29),
	.w7(32'h3aa2205f),
	.w8(32'hbb19c9b1),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8de359),
	.w1(32'hbc0f9400),
	.w2(32'hba80181d),
	.w3(32'h3b00bfd8),
	.w4(32'h39d05a46),
	.w5(32'hb9c030a1),
	.w6(32'hbb81cc31),
	.w7(32'h3b3fa7ab),
	.w8(32'h3b5e131a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c2f6f),
	.w1(32'h3b2d89ea),
	.w2(32'h3a53a204),
	.w3(32'hb8decf44),
	.w4(32'h3aa62a11),
	.w5(32'hbac156f1),
	.w6(32'h3bc3ad97),
	.w7(32'h3a494b95),
	.w8(32'hbad7cd86),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab99658),
	.w1(32'hba5c41ba),
	.w2(32'hbb05e81e),
	.w3(32'hba183249),
	.w4(32'hba0b40f6),
	.w5(32'hbb211125),
	.w6(32'h399664ce),
	.w7(32'hba3a48c9),
	.w8(32'hbb3e4258),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfd0fc),
	.w1(32'hbaf97044),
	.w2(32'hba80145a),
	.w3(32'hbaf735a6),
	.w4(32'hba9150cc),
	.w5(32'h3bb37ea6),
	.w6(32'hbb1d54ba),
	.w7(32'hbacdf370),
	.w8(32'h3b11aea4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43407d),
	.w1(32'hb94104de),
	.w2(32'hba0d68fe),
	.w3(32'h3b593d66),
	.w4(32'h3a663923),
	.w5(32'h3ab64a23),
	.w6(32'h3b52aeb5),
	.w7(32'h3b35dcd9),
	.w8(32'hb965b03c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46cabe),
	.w1(32'hbbee2e9b),
	.w2(32'h3b61caf5),
	.w3(32'h3b7cd10a),
	.w4(32'h3bd550f2),
	.w5(32'h3aa17595),
	.w6(32'hbb81088e),
	.w7(32'h3bea998e),
	.w8(32'h3af43150),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3c0d7),
	.w1(32'h3acbe01d),
	.w2(32'hbb00f5fa),
	.w3(32'h3b30ced3),
	.w4(32'h3947d443),
	.w5(32'h3a9fc7bb),
	.w6(32'h3ada2d93),
	.w7(32'hbb123cd0),
	.w8(32'h3b07601f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6767fb),
	.w1(32'h3b7913c9),
	.w2(32'h3a885fcb),
	.w3(32'h3ac140db),
	.w4(32'hba8c6fcf),
	.w5(32'hbb36b195),
	.w6(32'h3b0f97d4),
	.w7(32'hba50b7a5),
	.w8(32'hbb16b485),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3910fc8a),
	.w1(32'h3a4018bd),
	.w2(32'h3b8922b5),
	.w3(32'h3a8c2f80),
	.w4(32'h3acd0ad7),
	.w5(32'hbb6305cf),
	.w6(32'h3a29ad57),
	.w7(32'h3bdee667),
	.w8(32'hb9ef0a71),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2a561),
	.w1(32'h3a95c619),
	.w2(32'hb8854aed),
	.w3(32'hbae0a0d1),
	.w4(32'h3a5a703f),
	.w5(32'hbb2db737),
	.w6(32'h3b1ac59e),
	.w7(32'h3ba91fc4),
	.w8(32'h3a53e2ab),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bdb35),
	.w1(32'hbb5c424e),
	.w2(32'h39facd1f),
	.w3(32'hbb876ce7),
	.w4(32'h3ab3f5e1),
	.w5(32'hbabfd350),
	.w6(32'h3a4e8287),
	.w7(32'h3b921af1),
	.w8(32'hb96f17ea),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab73017),
	.w1(32'h399e456f),
	.w2(32'h3804ce18),
	.w3(32'hba953e5e),
	.w4(32'hba8271a4),
	.w5(32'h3a7f8669),
	.w6(32'h39602eb6),
	.w7(32'hba448847),
	.w8(32'h3ad128bd),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d0f1e),
	.w1(32'h3889eac8),
	.w2(32'h3b9272b1),
	.w3(32'h3b222172),
	.w4(32'h3a2e5c37),
	.w5(32'h3ad68442),
	.w6(32'h3b532d1c),
	.w7(32'h3c0cced0),
	.w8(32'h3b3eff9c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392511e1),
	.w1(32'h39ba9743),
	.w2(32'hba73e9f9),
	.w3(32'h3bafec87),
	.w4(32'h3b737453),
	.w5(32'h3bd98378),
	.w6(32'h3bc5d771),
	.w7(32'h3ba083ee),
	.w8(32'h3b9f9467),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b40c2),
	.w1(32'hbb2f40e9),
	.w2(32'hba1735b9),
	.w3(32'h3b6989ad),
	.w4(32'h3b7f50d8),
	.w5(32'hbaf20283),
	.w6(32'hba4572e7),
	.w7(32'h3add1928),
	.w8(32'h3af55e34),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71c010),
	.w1(32'h3be83809),
	.w2(32'h3b5217ad),
	.w3(32'hbb957a00),
	.w4(32'h3946971e),
	.w5(32'h3baf84df),
	.w6(32'hba97380b),
	.w7(32'h3bcca5af),
	.w8(32'h3b05037d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc158bc8),
	.w1(32'hb79120f0),
	.w2(32'h3be2aab6),
	.w3(32'h3bc779b1),
	.w4(32'h3b82022c),
	.w5(32'hbb8e78d5),
	.w6(32'h3bd71303),
	.w7(32'h3ad5cbd6),
	.w8(32'hbaea1491),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17871b),
	.w1(32'hbb2291d0),
	.w2(32'hbb809a4d),
	.w3(32'hbb4c10bc),
	.w4(32'hbb473ca4),
	.w5(32'hba13f505),
	.w6(32'hbb4e5737),
	.w7(32'hbbab5566),
	.w8(32'hb99862fb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0198b2),
	.w1(32'hba733b87),
	.w2(32'hb84a3b32),
	.w3(32'h3b0237b1),
	.w4(32'h3a6437ad),
	.w5(32'h3a1d978b),
	.w6(32'h3b4d0e5d),
	.w7(32'h3b2609aa),
	.w8(32'hba0eaf7f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00eeff),
	.w1(32'h3b85a5de),
	.w2(32'h3b90c257),
	.w3(32'h3b7387e2),
	.w4(32'h39d628bf),
	.w5(32'hba977465),
	.w6(32'h3b47a32b),
	.w7(32'h3b250258),
	.w8(32'h3a45f471),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f3812),
	.w1(32'h3856d9fd),
	.w2(32'h39d1e105),
	.w3(32'hbaec3642),
	.w4(32'hbac6fe4f),
	.w5(32'h393571b4),
	.w6(32'hbaa4eb57),
	.w7(32'hbac37889),
	.w8(32'h391afcdb),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca8e1e),
	.w1(32'h3b04f6d3),
	.w2(32'hbb198dea),
	.w3(32'hbab6eeeb),
	.w4(32'h3a5f369a),
	.w5(32'hbb819845),
	.w6(32'hba4de504),
	.w7(32'h3909bbba),
	.w8(32'hba4d3a46),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86c197),
	.w1(32'hba3f2078),
	.w2(32'h3bb9a663),
	.w3(32'hbb84c3a1),
	.w4(32'hba8d8020),
	.w5(32'hbba59daf),
	.w6(32'hbb31cf7d),
	.w7(32'h3ae05e93),
	.w8(32'hbaced84b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4673bd),
	.w1(32'hba679adb),
	.w2(32'hb942650a),
	.w3(32'hba27d6b5),
	.w4(32'h39dff7d7),
	.w5(32'h3bc43cd1),
	.w6(32'h3ba5572e),
	.w7(32'h3c36f536),
	.w8(32'h3ace4c07),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60c5ef),
	.w1(32'hb93169c4),
	.w2(32'hbbb4d092),
	.w3(32'h3b865bd0),
	.w4(32'hbabc356c),
	.w5(32'h3ad09d02),
	.w6(32'hbadbce3e),
	.w7(32'hbbb9eff3),
	.w8(32'hbb29c1bd),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc6d65),
	.w1(32'h3b409089),
	.w2(32'hbb32f32b),
	.w3(32'h3b17876c),
	.w4(32'hb99e792b),
	.w5(32'hbb82b53a),
	.w6(32'hba99bf44),
	.w7(32'hbb7b4ba7),
	.w8(32'hba021220),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38de63),
	.w1(32'hbb3994b2),
	.w2(32'hbb8ce580),
	.w3(32'hbb9f5863),
	.w4(32'hbb5eb79d),
	.w5(32'h3b1db774),
	.w6(32'hba963277),
	.w7(32'hba548b83),
	.w8(32'hba73048f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98409a),
	.w1(32'hba87c7f3),
	.w2(32'h3b0b4868),
	.w3(32'hbaf29c6b),
	.w4(32'hbaabf8a4),
	.w5(32'hbb2f5b2f),
	.w6(32'hbbbc6019),
	.w7(32'h3ac4d750),
	.w8(32'hbb5ed34d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37e60a),
	.w1(32'h393b6a9e),
	.w2(32'hbad92ac0),
	.w3(32'hbbbb30f7),
	.w4(32'hbbc93e48),
	.w5(32'hbb710f5c),
	.w6(32'h39b5d406),
	.w7(32'hbb8bbfc5),
	.w8(32'hbb41b738),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9bdef),
	.w1(32'hbb13182f),
	.w2(32'hb9f1d3e0),
	.w3(32'hbae639fe),
	.w4(32'hbb216e81),
	.w5(32'h3b6add2b),
	.w6(32'hbaa24d2b),
	.w7(32'h3a4e457a),
	.w8(32'h3c5f34b9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20ed94),
	.w1(32'h3bae225f),
	.w2(32'hbb88e3ad),
	.w3(32'hba06d065),
	.w4(32'hbbb48b03),
	.w5(32'hb9910196),
	.w6(32'h3c4337a2),
	.w7(32'hba3a3d80),
	.w8(32'h3a34c8f9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9581c00),
	.w1(32'h3a9187d5),
	.w2(32'hb99df6f6),
	.w3(32'hbaa2de81),
	.w4(32'hb9247e59),
	.w5(32'h3b8c1777),
	.w6(32'h3b4294f9),
	.w7(32'h3ac92243),
	.w8(32'h3b55904f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adee237),
	.w1(32'h3b8c92f6),
	.w2(32'h3b8967d5),
	.w3(32'h3bc30046),
	.w4(32'h3bfae937),
	.w5(32'hbb4c503a),
	.w6(32'h3b4a17b6),
	.w7(32'h3b7f0b79),
	.w8(32'hbbae8963),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73b7ab),
	.w1(32'hbb499e10),
	.w2(32'hba4e3b81),
	.w3(32'h39867a56),
	.w4(32'h3a5d7c82),
	.w5(32'h3b0bf0c0),
	.w6(32'hbb0578ae),
	.w7(32'h3b38c15b),
	.w8(32'h3b0bb290),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af38a90),
	.w1(32'h3a9f0a30),
	.w2(32'h39706a58),
	.w3(32'h3b22227f),
	.w4(32'h3a8b05fd),
	.w5(32'h3b762cd2),
	.w6(32'h3b3f9440),
	.w7(32'h39c4fbbc),
	.w8(32'h3afd5a77),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae03175),
	.w1(32'h3991737f),
	.w2(32'hb9fa0c57),
	.w3(32'hbad56a56),
	.w4(32'h3a273782),
	.w5(32'hbb16c18f),
	.w6(32'hba946ad8),
	.w7(32'hbb0f1fdf),
	.w8(32'hba12a1f1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a51a5),
	.w1(32'h3a8e2ccb),
	.w2(32'h3a8be639),
	.w3(32'hbb7bd8b0),
	.w4(32'hbb31f8d9),
	.w5(32'h3b975138),
	.w6(32'hbb2c7e37),
	.w7(32'hbb3eb418),
	.w8(32'h385b128f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19476f),
	.w1(32'h3bb1de87),
	.w2(32'h3a66cb8e),
	.w3(32'hbb28322a),
	.w4(32'hbbb0ba1d),
	.w5(32'h3ab3f70c),
	.w6(32'h3a707adb),
	.w7(32'hb9157421),
	.w8(32'hba98ead1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b8008),
	.w1(32'h3a625505),
	.w2(32'hbb6c77b5),
	.w3(32'h39ab421e),
	.w4(32'h3a55eb4f),
	.w5(32'hb99e2bd5),
	.w6(32'hba62f0a2),
	.w7(32'hbad10aec),
	.w8(32'hbb0a60f5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa23d5),
	.w1(32'hb969eecc),
	.w2(32'hb9e28df2),
	.w3(32'h39c5db96),
	.w4(32'hbb0c3108),
	.w5(32'hbb17fa60),
	.w6(32'h3b1fa473),
	.w7(32'hba1f24fb),
	.w8(32'hbb899bc6),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb942ee7),
	.w1(32'hbb757bf9),
	.w2(32'h39d3e2f2),
	.w3(32'h3b702fd5),
	.w4(32'hb77ba90b),
	.w5(32'hb937f792),
	.w6(32'h3aaa13a6),
	.w7(32'hb9ad57e2),
	.w8(32'hbabd3c9c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fc56f),
	.w1(32'hb9537ca2),
	.w2(32'hba536f57),
	.w3(32'h387bde44),
	.w4(32'h3a889f68),
	.w5(32'h3b8cc7bf),
	.w6(32'hbaf4eafb),
	.w7(32'hbafcb10f),
	.w8(32'h3b377983),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b862510),
	.w1(32'h3a1e3866),
	.w2(32'hbaec1316),
	.w3(32'h3b92ca46),
	.w4(32'hb88d01fb),
	.w5(32'h3b4d205a),
	.w6(32'h3a3f9901),
	.w7(32'h3939c689),
	.w8(32'h3b5ed4e2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ff669),
	.w1(32'h3b2ca259),
	.w2(32'h3bb695ef),
	.w3(32'h3a94e6f4),
	.w4(32'h3b8b3149),
	.w5(32'hb9ec4f12),
	.w6(32'h3b3c631c),
	.w7(32'h3b97e6ac),
	.w8(32'h3c342dbc),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc37ba4),
	.w1(32'h3c74d0bf),
	.w2(32'h3a226d19),
	.w3(32'h3ae64e97),
	.w4(32'hbba30c46),
	.w5(32'hba188e89),
	.w6(32'h3c80232e),
	.w7(32'hbacc246c),
	.w8(32'h3ac22ae8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eac273),
	.w1(32'h3a06ba8a),
	.w2(32'hbac1d68b),
	.w3(32'h3affda66),
	.w4(32'h3a99f9d0),
	.w5(32'hbb440080),
	.w6(32'h3b886fa9),
	.w7(32'h3be0023f),
	.w8(32'h3b21e2bf),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba3e1d),
	.w1(32'hbb402d1c),
	.w2(32'hbb2a51ce),
	.w3(32'hbb8a8216),
	.w4(32'hbbe5cc4b),
	.w5(32'hbb684ee4),
	.w6(32'h3bca2c6f),
	.w7(32'h3ae352b3),
	.w8(32'hbbbb5373),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a4a4a),
	.w1(32'h3a99372b),
	.w2(32'h3b10d8c4),
	.w3(32'hbb7a5c18),
	.w4(32'hbb76fd3c),
	.w5(32'h3a4b1910),
	.w6(32'hbb53a89a),
	.w7(32'hbac62392),
	.w8(32'hba2d0d8c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfc7ad),
	.w1(32'hba2a6441),
	.w2(32'hbad351dc),
	.w3(32'h3b612334),
	.w4(32'hba8805af),
	.w5(32'h3b071cc9),
	.w6(32'hb9e982d9),
	.w7(32'hbb214175),
	.w8(32'hba16cd7e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1bd78),
	.w1(32'h3ac16409),
	.w2(32'h3b65f90d),
	.w3(32'h3b693b88),
	.w4(32'hbb21bfad),
	.w5(32'hba74ea28),
	.w6(32'h3b4a6b5c),
	.w7(32'h3b55aa6b),
	.w8(32'hbbffd249),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40ec05),
	.w1(32'h3a9d676d),
	.w2(32'h3b8da8df),
	.w3(32'hbb02b54b),
	.w4(32'hbb43ec50),
	.w5(32'hbab01aa4),
	.w6(32'h389c457c),
	.w7(32'h3b0f032c),
	.w8(32'h38307932),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc206d1),
	.w1(32'hba472383),
	.w2(32'hbba67a18),
	.w3(32'hbb0daf95),
	.w4(32'hbc143c35),
	.w5(32'hb9c3d65b),
	.w6(32'h38830765),
	.w7(32'hbbb5092a),
	.w8(32'hbab55820),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb122e14),
	.w1(32'hbb477b32),
	.w2(32'hbb24bc7e),
	.w3(32'hbbd097d8),
	.w4(32'hbb239c2b),
	.w5(32'h3ac519b9),
	.w6(32'hbbc5a7af),
	.w7(32'hbb2f07d0),
	.w8(32'h3b37a74d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f4706),
	.w1(32'h3b52e795),
	.w2(32'h3ae27677),
	.w3(32'h3b2b9a75),
	.w4(32'h394d471a),
	.w5(32'hba55ae4a),
	.w6(32'h3b90a18a),
	.w7(32'h3af04541),
	.w8(32'h3b7da720),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9afa22),
	.w1(32'h3b70f3b4),
	.w2(32'hba91d983),
	.w3(32'hbabab2d9),
	.w4(32'hbb12f399),
	.w5(32'hba7e6553),
	.w6(32'h391ae01a),
	.w7(32'hbb9e5e85),
	.w8(32'hba361fbd),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c00b0),
	.w1(32'hba30beef),
	.w2(32'h394157f1),
	.w3(32'hbafe4cf5),
	.w4(32'hbabfe05c),
	.w5(32'hbb32a5f2),
	.w6(32'hbaff9967),
	.w7(32'hba9451c9),
	.w8(32'hbb53b331),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51770c),
	.w1(32'hbb05f36b),
	.w2(32'hbaa0cda5),
	.w3(32'hbb810ca5),
	.w4(32'hbad652c3),
	.w5(32'hbbb0c453),
	.w6(32'hbba1507f),
	.w7(32'hba24078d),
	.w8(32'hbb85c2dd),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6be610),
	.w1(32'h3b916836),
	.w2(32'h3bb21020),
	.w3(32'hbb5eb894),
	.w4(32'hbad1c82b),
	.w5(32'h3a1e62a4),
	.w6(32'hba6c8340),
	.w7(32'h3ae53919),
	.w8(32'h36d16710),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11a64b),
	.w1(32'hbac04264),
	.w2(32'hbae07b01),
	.w3(32'h3a10924d),
	.w4(32'h3b2dc547),
	.w5(32'hbaac5961),
	.w6(32'hbb41f12c),
	.w7(32'h3aa2f61a),
	.w8(32'hba4b0a5f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98bc7e),
	.w1(32'hbaded0a7),
	.w2(32'hbb6bf31d),
	.w3(32'h3a7a531c),
	.w4(32'hbc057f28),
	.w5(32'hbaf2574a),
	.w6(32'h3a92a89b),
	.w7(32'hbb45c5e0),
	.w8(32'hbbc19ed5),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb16693),
	.w1(32'hbb5cfddc),
	.w2(32'h3ab626ad),
	.w3(32'h3ad4771f),
	.w4(32'h3b7491c9),
	.w5(32'h3a237cfa),
	.w6(32'hbb13bf47),
	.w7(32'h3aff819d),
	.w8(32'hba8bf18b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e839f),
	.w1(32'h3b9c3bc1),
	.w2(32'h3b35b95f),
	.w3(32'hb9bb7782),
	.w4(32'hbb4d11f7),
	.w5(32'hbadad9e8),
	.w6(32'hb9971e68),
	.w7(32'hbab4f5b5),
	.w8(32'h3a5018b9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af154fa),
	.w1(32'h3ac5a3fb),
	.w2(32'h3a780e99),
	.w3(32'hbaea97d1),
	.w4(32'hba90b401),
	.w5(32'h38ecba7e),
	.w6(32'h3a366ca0),
	.w7(32'h3a2a7d3e),
	.w8(32'hb9e9fc8b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c81e5e),
	.w1(32'h3a25b082),
	.w2(32'hb8b2e7fe),
	.w3(32'hba213361),
	.w4(32'hbb560b87),
	.w5(32'hbba743e0),
	.w6(32'h38d9286d),
	.w7(32'hba4b2293),
	.w8(32'hba9eb2d1),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee4d9f),
	.w1(32'h3a90f4ab),
	.w2(32'hbb0eca98),
	.w3(32'hbb91a7e9),
	.w4(32'hbb916b6a),
	.w5(32'h3b6627be),
	.w6(32'h3ae0f536),
	.w7(32'hb84cd862),
	.w8(32'hbb5eda3d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eee045),
	.w1(32'hba61493e),
	.w2(32'h3aa66ea6),
	.w3(32'h3b50a8b6),
	.w4(32'h3a3b0617),
	.w5(32'hbabcea79),
	.w6(32'hbbb3c838),
	.w7(32'hbaa5ea76),
	.w8(32'hbb13395d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab69a69),
	.w1(32'hb95e9e95),
	.w2(32'hba045331),
	.w3(32'hb94468b2),
	.w4(32'h3a2561cf),
	.w5(32'h392087ee),
	.w6(32'hbb17f2b2),
	.w7(32'h3a912771),
	.w8(32'h3b8cb6d5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e3486),
	.w1(32'h3b87c430),
	.w2(32'hb97dd98c),
	.w3(32'h3b318a96),
	.w4(32'hbabfd454),
	.w5(32'hbbc3a5d5),
	.w6(32'h3bc3d2d9),
	.w7(32'h3a92eeea),
	.w8(32'hbbdf5f50),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba96594),
	.w1(32'hbb1c3db2),
	.w2(32'hbb466d60),
	.w3(32'hbb27308f),
	.w4(32'hbb9d19f5),
	.w5(32'h3b0d540c),
	.w6(32'hba9ef847),
	.w7(32'hbb2bf9f2),
	.w8(32'h3b9402d7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6302b),
	.w1(32'h3af1d247),
	.w2(32'h3aa7ac01),
	.w3(32'h3b7d0e72),
	.w4(32'h3b5bf2a2),
	.w5(32'hbac8591d),
	.w6(32'h3bbe5655),
	.w7(32'h3b63f80e),
	.w8(32'h3b9a0757),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84abf2),
	.w1(32'h3bcf6d07),
	.w2(32'h3bd87a3d),
	.w3(32'hb918bed7),
	.w4(32'hbb9acd0b),
	.w5(32'hbacf54cc),
	.w6(32'h3c6e2860),
	.w7(32'h3c3cbb37),
	.w8(32'h3a30ab5d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbdefc),
	.w1(32'hba050009),
	.w2(32'hbb5822eb),
	.w3(32'hba5cdf30),
	.w4(32'hbb6abb75),
	.w5(32'h3a794a82),
	.w6(32'h3b54cefd),
	.w7(32'hbb1058e8),
	.w8(32'h38cb5a40),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b329c75),
	.w1(32'h3a9dd57d),
	.w2(32'h3b24a93d),
	.w3(32'h3abcb137),
	.w4(32'h39b91c94),
	.w5(32'hbb1f3a4e),
	.w6(32'h3b45a707),
	.w7(32'h3b751627),
	.w8(32'h3a7fd1a5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7fd07e),
	.w1(32'h3a835daa),
	.w2(32'hba331f77),
	.w3(32'hbb0c6a1e),
	.w4(32'hba292edc),
	.w5(32'h3bdf624f),
	.w6(32'h3ac5c4d5),
	.w7(32'hbaa3e075),
	.w8(32'h3b6d604b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd03c00),
	.w1(32'hbbd3a2f5),
	.w2(32'h3a3a4257),
	.w3(32'hbb7f8e5e),
	.w4(32'h3b91d06c),
	.w5(32'h39f151c9),
	.w6(32'hbc1eae85),
	.w7(32'hb9abb4af),
	.w8(32'hbb9535da),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dc97d),
	.w1(32'h3ab2c832),
	.w2(32'hba1c5735),
	.w3(32'h3bad8c6b),
	.w4(32'h3b427c12),
	.w5(32'hba5842f6),
	.w6(32'h3babbd82),
	.w7(32'hba2b1e0b),
	.w8(32'h3a3530cd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a758225),
	.w1(32'hbafc8eec),
	.w2(32'hbb84c327),
	.w3(32'h3a6a1d8e),
	.w4(32'h399a846e),
	.w5(32'hbaef517d),
	.w6(32'hb9869d75),
	.w7(32'hb9ba6a8a),
	.w8(32'hba9e4c88),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4bc8c),
	.w1(32'hbb101591),
	.w2(32'h3add6863),
	.w3(32'hbb3939e7),
	.w4(32'h3a7c107b),
	.w5(32'hba92832f),
	.w6(32'h3a1b5680),
	.w7(32'hb99ea516),
	.w8(32'hbad030c9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60d1ac),
	.w1(32'hba58be75),
	.w2(32'hbb69b5e1),
	.w3(32'h3b0d6959),
	.w4(32'hba676256),
	.w5(32'hbb669ad1),
	.w6(32'h390a7e79),
	.w7(32'hba7c62fb),
	.w8(32'hbb10546b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95e6b8),
	.w1(32'hbb8ea5de),
	.w2(32'h3b3e05b2),
	.w3(32'hbbe6b679),
	.w4(32'hbab2ed44),
	.w5(32'hbb821df4),
	.w6(32'hbbe1f99a),
	.w7(32'h3a8d039c),
	.w8(32'hb89d3955),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d5187),
	.w1(32'hb92694d0),
	.w2(32'h3bb0c053),
	.w3(32'hbc00e4aa),
	.w4(32'hbbe02221),
	.w5(32'h3ad82a86),
	.w6(32'hbb3a49c4),
	.w7(32'h38d43f33),
	.w8(32'hbb0ecf1f),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61aae8),
	.w1(32'hba1ad8fe),
	.w2(32'h3b7f4c9f),
	.w3(32'h3b3f4886),
	.w4(32'h3ae230cc),
	.w5(32'hbb1d56b9),
	.w6(32'h3b55ebd5),
	.w7(32'h3b42dd3d),
	.w8(32'h3a748656),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05fc0f),
	.w1(32'h3ba6fd31),
	.w2(32'h39db729a),
	.w3(32'hbb33e707),
	.w4(32'h3b46da3f),
	.w5(32'hbb020e01),
	.w6(32'h3b051def),
	.w7(32'h3aa0c461),
	.w8(32'hbb3cb6de),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70dd7b),
	.w1(32'hba9133d9),
	.w2(32'hb91b26eb),
	.w3(32'h3b45c535),
	.w4(32'h3b2d2054),
	.w5(32'h3b91b9bc),
	.w6(32'h3b6eb3e7),
	.w7(32'h3b89dc99),
	.w8(32'h3b1ab526),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa3f53),
	.w1(32'h39f395fd),
	.w2(32'hbafcb543),
	.w3(32'h3b8d1d99),
	.w4(32'h3a8806c5),
	.w5(32'hbb434676),
	.w6(32'h3c0bb207),
	.w7(32'hbb42c521),
	.w8(32'h3b1a75a3),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a0f1a),
	.w1(32'hbab5db0f),
	.w2(32'h3b85fd67),
	.w3(32'h3be3c59d),
	.w4(32'h3b7ab0e2),
	.w5(32'hba8abdc1),
	.w6(32'h3c41a209),
	.w7(32'h3c213dd7),
	.w8(32'hbb4f9e80),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb150ad9),
	.w1(32'h3b635a81),
	.w2(32'h3b24b8d6),
	.w3(32'hb9ee40e4),
	.w4(32'hbaf1d2ac),
	.w5(32'hbab923ce),
	.w6(32'hbb3652dd),
	.w7(32'hba3941e1),
	.w8(32'hba90f84d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56e01e),
	.w1(32'hba3140bb),
	.w2(32'h3b81cc0b),
	.w3(32'hba9777a2),
	.w4(32'h3aaef825),
	.w5(32'hbb72d96e),
	.w6(32'hbb387ca5),
	.w7(32'h3b34010d),
	.w8(32'hbb46f0f1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6f97f),
	.w1(32'h3a81fc60),
	.w2(32'hb934e501),
	.w3(32'h3b245c7c),
	.w4(32'hb9003056),
	.w5(32'hba8ac2f0),
	.w6(32'hba5b38dc),
	.w7(32'hbb68d733),
	.w8(32'h3ba378db),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb170383),
	.w1(32'h3bfa3c62),
	.w2(32'h3c09fbe8),
	.w3(32'h3c498276),
	.w4(32'h3bf40379),
	.w5(32'h3ac2f514),
	.w6(32'h3bfa60fb),
	.w7(32'h3c1cdcc6),
	.w8(32'h3b8df244),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3c316),
	.w1(32'h3bba76ac),
	.w2(32'h3ac17d1e),
	.w3(32'h3b2b63da),
	.w4(32'h3be6aca2),
	.w5(32'h3b688263),
	.w6(32'h3bc8c6e7),
	.w7(32'h3bac1296),
	.w8(32'h3b54863e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e830e5),
	.w1(32'h3aa71871),
	.w2(32'h3a8de760),
	.w3(32'h3afb27c3),
	.w4(32'h3b04fdf9),
	.w5(32'h3ac85015),
	.w6(32'h38e8daf7),
	.w7(32'h3bfd5e27),
	.w8(32'h39348f83),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d013f),
	.w1(32'hbaa02b8b),
	.w2(32'hb85c7ab9),
	.w3(32'h3be7e26f),
	.w4(32'h3b9d79e8),
	.w5(32'hbbd9fdd6),
	.w6(32'h3b9bf891),
	.w7(32'h3ba4f1f0),
	.w8(32'hbbca54d2),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d9ae2),
	.w1(32'hbb8ae2a2),
	.w2(32'hbaee5b1f),
	.w3(32'hbb9ffe43),
	.w4(32'h39e37ac1),
	.w5(32'h3a980481),
	.w6(32'hbb4da470),
	.w7(32'h3a7fb71e),
	.w8(32'hba348ff7),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb559a7f),
	.w1(32'hb9ac1088),
	.w2(32'hbb07fe2c),
	.w3(32'h3b5aeafc),
	.w4(32'h3ae98eef),
	.w5(32'h3b8df32d),
	.w6(32'h3ad0c46f),
	.w7(32'h3aa90638),
	.w8(32'h3a8ed4a5),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad16e23),
	.w1(32'hba3f0173),
	.w2(32'h3bb16a4b),
	.w3(32'h3b4a7698),
	.w4(32'h3b86f66c),
	.w5(32'h3b2b177e),
	.w6(32'h3b6a18b5),
	.w7(32'h3b882da5),
	.w8(32'h3b183143),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1814d),
	.w1(32'hb9599694),
	.w2(32'h3a01fda5),
	.w3(32'h3b027aa1),
	.w4(32'hbae938cc),
	.w5(32'hb93c9217),
	.w6(32'hbb0dbe96),
	.w7(32'h399f734c),
	.w8(32'hba051065),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05f2f2),
	.w1(32'h3a85af72),
	.w2(32'h3a7056a6),
	.w3(32'hba20e622),
	.w4(32'h39d108e9),
	.w5(32'hba871a39),
	.w6(32'hb9e29f4b),
	.w7(32'h3aae7f36),
	.w8(32'hbb380d31),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98bddcc),
	.w1(32'hbb1c5ec0),
	.w2(32'hbb6ef681),
	.w3(32'hbb2a72c5),
	.w4(32'hba91c356),
	.w5(32'h3b1ee82b),
	.w6(32'hbba1ac58),
	.w7(32'hbb65bc0d),
	.w8(32'h3b49708f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95a39f),
	.w1(32'h3aa5ba66),
	.w2(32'hbbc456b0),
	.w3(32'h3c500706),
	.w4(32'h3be079a7),
	.w5(32'h3a7d8478),
	.w6(32'h3cdc8364),
	.w7(32'h3b3f88b1),
	.w8(32'hba1c31bd),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45c935),
	.w1(32'hba9f3811),
	.w2(32'h39b98ee2),
	.w3(32'hba93535e),
	.w4(32'hbbb77cb9),
	.w5(32'h39eaf5eb),
	.w6(32'hbbc52d00),
	.w7(32'hba5c2230),
	.w8(32'hba5b13a2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80a7c4a),
	.w1(32'h3a83d205),
	.w2(32'h3a3e7cc5),
	.w3(32'hba2a11c2),
	.w4(32'hbaad3222),
	.w5(32'h3a0206d2),
	.w6(32'hbaf82f44),
	.w7(32'hba97555b),
	.w8(32'h3ba4b0a2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81107a),
	.w1(32'h3b923ae8),
	.w2(32'hba8a18a8),
	.w3(32'h3bcb3070),
	.w4(32'h3b7b144e),
	.w5(32'h3b2b1106),
	.w6(32'hbb86d386),
	.w7(32'h3c41c379),
	.w8(32'h3b93c363),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35be1cd8),
	.w1(32'h3a8f52ad),
	.w2(32'hbb440ea7),
	.w3(32'h3bae7411),
	.w4(32'h3a8617d2),
	.w5(32'h3bb83c88),
	.w6(32'h3be73264),
	.w7(32'h3b393bbd),
	.w8(32'h3b85f642),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5b55d),
	.w1(32'h3ba1900b),
	.w2(32'h3baaf9bf),
	.w3(32'h3c6c8482),
	.w4(32'h3b98379d),
	.w5(32'hb9130455),
	.w6(32'h3c1b12ef),
	.w7(32'h3bb43832),
	.w8(32'h39fce25b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc7f7f),
	.w1(32'h3b3c8866),
	.w2(32'h3a908143),
	.w3(32'h3adf9a15),
	.w4(32'hba38f8ac),
	.w5(32'h3ad5e7bd),
	.w6(32'hbb552806),
	.w7(32'hb7d53b86),
	.w8(32'h3acb8aac),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65e384),
	.w1(32'hbb202d04),
	.w2(32'hb98fcd18),
	.w3(32'h3ab68a1d),
	.w4(32'h39a72983),
	.w5(32'hbb27d05f),
	.w6(32'hba6694c0),
	.w7(32'h37c5a6e0),
	.w8(32'h39605272),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e6db5),
	.w1(32'h3a7a9bf2),
	.w2(32'hbaaaf146),
	.w3(32'hbbed64d4),
	.w4(32'hbbc17c0e),
	.w5(32'hbb0eac9c),
	.w6(32'hbb5c10d1),
	.w7(32'hbbe098c0),
	.w8(32'hbad91733),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a945372),
	.w1(32'hbb40db1b),
	.w2(32'hbb3d1c8a),
	.w3(32'hbbb45223),
	.w4(32'hbb6a9e1e),
	.w5(32'hb7102c01),
	.w6(32'hbb496c5c),
	.w7(32'hbb8b6a6c),
	.w8(32'hb9afd3d6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b641c67),
	.w1(32'h3af0bea1),
	.w2(32'h38a256df),
	.w3(32'hbb825317),
	.w4(32'hba8e0142),
	.w5(32'hbb2e82e1),
	.w6(32'hbb2a9e4b),
	.w7(32'hbb937bbe),
	.w8(32'hbb3798c5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae10ba),
	.w1(32'hb89dd4e1),
	.w2(32'hbb19eb66),
	.w3(32'h3a9d31d6),
	.w4(32'h3b0c7bc3),
	.w5(32'h3ac496ba),
	.w6(32'hbadabbbd),
	.w7(32'hbb28147f),
	.w8(32'hbb391bc3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f8383),
	.w1(32'hbb4108cb),
	.w2(32'hba32f0ed),
	.w3(32'h3b2c7c0d),
	.w4(32'h39fb28f0),
	.w5(32'hbbf4a1a4),
	.w6(32'h3b019bd9),
	.w7(32'h3a5d4f30),
	.w8(32'hbbe67c3b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe59e06),
	.w1(32'hbc08f3e4),
	.w2(32'hbbb41504),
	.w3(32'hbba1fff1),
	.w4(32'hbbbdc13d),
	.w5(32'h3a337737),
	.w6(32'hbbb034ac),
	.w7(32'hbb8dbb16),
	.w8(32'hba6ee5f6),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule