module layer_10_featuremap_242(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2feee6),
	.w1(32'h3bc759f5),
	.w2(32'h3b5555d9),
	.w3(32'h3c3c607a),
	.w4(32'h3bb10801),
	.w5(32'h3bac3fd8),
	.w6(32'h3c865b92),
	.w7(32'h3b59f07e),
	.w8(32'h38780d60),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdb5ad),
	.w1(32'h3c0f6c28),
	.w2(32'h3c87c4ee),
	.w3(32'h3c141eb1),
	.w4(32'h3c12c630),
	.w5(32'h391aec61),
	.w6(32'h3c00bd22),
	.w7(32'h3c0b1d3b),
	.w8(32'h3a9c704f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30f015),
	.w1(32'h39a0c4a5),
	.w2(32'hba8deda2),
	.w3(32'h3a57294d),
	.w4(32'h3afe5506),
	.w5(32'hbaa806db),
	.w6(32'h3a6b34fd),
	.w7(32'hbad40e8f),
	.w8(32'h39890545),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a3ce2e),
	.w1(32'hb9c5ba26),
	.w2(32'hbadc3ecb),
	.w3(32'hba91b30c),
	.w4(32'hbb09b494),
	.w5(32'hbaf51bb4),
	.w6(32'h3a97452b),
	.w7(32'hba84fcbf),
	.w8(32'hbb3ff855),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b61ca),
	.w1(32'hb8c59eff),
	.w2(32'h3a9dbbf6),
	.w3(32'hbb62f04b),
	.w4(32'hba608ab6),
	.w5(32'hbb203c0c),
	.w6(32'hbb19d497),
	.w7(32'hb9d2a033),
	.w8(32'hba415178),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933c57c),
	.w1(32'h3b31d678),
	.w2(32'h398225e6),
	.w3(32'h3a72b0e6),
	.w4(32'hbb37b9f8),
	.w5(32'h3afab7b3),
	.w6(32'h3b8a8d98),
	.w7(32'hb9e92512),
	.w8(32'h3afc2a6d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a980182),
	.w1(32'h3b8de2a0),
	.w2(32'h3b389035),
	.w3(32'h3b2e6025),
	.w4(32'h3b6b1dc3),
	.w5(32'h3b8916a4),
	.w6(32'h3bcc7828),
	.w7(32'h3b47eaea),
	.w8(32'h3bbf7362),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8048f),
	.w1(32'hbc2fed11),
	.w2(32'hbc2c3349),
	.w3(32'hbc162756),
	.w4(32'hbba0f7ba),
	.w5(32'h3b7dbe72),
	.w6(32'hbc1c3b7b),
	.w7(32'hbc08ce5a),
	.w8(32'hba668ec7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20c724),
	.w1(32'h3afb980f),
	.w2(32'h3b260a5c),
	.w3(32'h3b449bbf),
	.w4(32'h3b190be3),
	.w5(32'hbb59ea1d),
	.w6(32'h3b8a96a0),
	.w7(32'h3b0f5cf7),
	.w8(32'hbaaa92fb),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380813e6),
	.w1(32'h3ba27bea),
	.w2(32'h3b6f4d97),
	.w3(32'h3b98a3f2),
	.w4(32'h3adbd0db),
	.w5(32'hbb88b43b),
	.w6(32'h3bf0b688),
	.w7(32'h3b1ea6bc),
	.w8(32'hbb40602e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe6cae),
	.w1(32'hb927edfc),
	.w2(32'hbb36d283),
	.w3(32'hbad62cef),
	.w4(32'hbb66997e),
	.w5(32'h3ae8449d),
	.w6(32'h3ad9ee3b),
	.w7(32'hbb99eb5b),
	.w8(32'h3af1edd1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5460d0),
	.w1(32'hbb904c31),
	.w2(32'hbc0f55bb),
	.w3(32'hb81fbed2),
	.w4(32'h3a8c67b9),
	.w5(32'hbb963804),
	.w6(32'hbb35a068),
	.w7(32'hbb8486df),
	.w8(32'hbbf7c1c6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba44c4b),
	.w1(32'hbbf2160e),
	.w2(32'hbaa5780f),
	.w3(32'hbb04699b),
	.w4(32'hbbc22ff1),
	.w5(32'h3aca5b38),
	.w6(32'hbb87660e),
	.w7(32'hbba5cea8),
	.w8(32'h3af6c671),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f3b7f),
	.w1(32'hbba3d5e9),
	.w2(32'hbbadcf5e),
	.w3(32'hbb79a9c6),
	.w4(32'hbbd89f3f),
	.w5(32'hbb9d9c44),
	.w6(32'hbac94695),
	.w7(32'hbbbae722),
	.w8(32'hb91fe183),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bf625),
	.w1(32'h3bdc7940),
	.w2(32'h38004b4d),
	.w3(32'h3b0c2e0c),
	.w4(32'h3a09c277),
	.w5(32'hb8b856f2),
	.w6(32'h3bbcb3cf),
	.w7(32'h3abe24de),
	.w8(32'hbb077986),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77f0df2),
	.w1(32'hbb2667fa),
	.w2(32'hbae816cf),
	.w3(32'h3a907f6a),
	.w4(32'hbb903590),
	.w5(32'hbb19ebae),
	.w6(32'hb87285a6),
	.w7(32'hbbcc2088),
	.w8(32'hbb505ab6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb696ffd),
	.w1(32'h39e95d63),
	.w2(32'h3a2be023),
	.w3(32'h389ea993),
	.w4(32'hbaa03c62),
	.w5(32'hba840117),
	.w6(32'h3b933c9a),
	.w7(32'h39ee5fad),
	.w8(32'h3a88e0cc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc396e78),
	.w1(32'hbc6cd101),
	.w2(32'hbc781cc0),
	.w3(32'hbc99bdd3),
	.w4(32'hbc77b96b),
	.w5(32'hbb84ac85),
	.w6(32'hbc446186),
	.w7(32'hbc3db102),
	.w8(32'hbab527fb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53dc8e),
	.w1(32'hbb9c1df5),
	.w2(32'hbb93b1d8),
	.w3(32'hbb75c99d),
	.w4(32'hbb623989),
	.w5(32'hbb7f6f6e),
	.w6(32'hbb0d24ef),
	.w7(32'hbb2af482),
	.w8(32'hbb85145c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66550d9),
	.w1(32'h39c095b3),
	.w2(32'h3a1a2cc9),
	.w3(32'hbb5eed4f),
	.w4(32'hb92d8316),
	.w5(32'h3aaae61a),
	.w6(32'hba75d2b2),
	.w7(32'h3a60b059),
	.w8(32'hbaf329b0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74e1f2),
	.w1(32'hbaaf0a80),
	.w2(32'h3b4cdb2b),
	.w3(32'h3b275c46),
	.w4(32'hb9be44b2),
	.w5(32'h3b0dd87d),
	.w6(32'h3b81e154),
	.w7(32'h3b2d31ff),
	.w8(32'h3b4f40b1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3b7dc),
	.w1(32'h3bb9465e),
	.w2(32'h3b519de3),
	.w3(32'h3bd15fe1),
	.w4(32'h3bd0dfbe),
	.w5(32'h3b17181a),
	.w6(32'h3bf87447),
	.w7(32'h3bdd1eeb),
	.w8(32'h3b50d2d8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3eda71),
	.w1(32'hbcc9594e),
	.w2(32'hbcb903bb),
	.w3(32'hbcc10033),
	.w4(32'hbc92af3b),
	.w5(32'hbbb321a7),
	.w6(32'hbcdf5c50),
	.w7(32'hbc836050),
	.w8(32'hbadbc138),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b933ce5),
	.w1(32'h3abaf82b),
	.w2(32'h3af07bea),
	.w3(32'h3b7875d3),
	.w4(32'hbb389551),
	.w5(32'hbaa5d5c8),
	.w6(32'h3c07ff41),
	.w7(32'hbb626d7a),
	.w8(32'hbb7b1aaf),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5659f),
	.w1(32'h3b9fb08e),
	.w2(32'h3a5eab2e),
	.w3(32'h3b6510b2),
	.w4(32'h3b908f63),
	.w5(32'hbb884312),
	.w6(32'h3b47ed28),
	.w7(32'hbb8f9e78),
	.w8(32'hbb5b3e50),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb029b67),
	.w1(32'h3af10582),
	.w2(32'hbb1a08ef),
	.w3(32'hbb361866),
	.w4(32'hbae28ba4),
	.w5(32'h39a75e22),
	.w6(32'h3b8f164e),
	.w7(32'h3af155ee),
	.w8(32'h3a1c1723),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e66f4b),
	.w1(32'h39214cb6),
	.w2(32'hbbba8e46),
	.w3(32'h39c6a990),
	.w4(32'hbb7e4926),
	.w5(32'h3bf32118),
	.w6(32'h3ab804b4),
	.w7(32'hbb761eab),
	.w8(32'h3baf7363),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc781b),
	.w1(32'h3c2cec81),
	.w2(32'h3c22b51d),
	.w3(32'h3c2cba9f),
	.w4(32'h3c0ed202),
	.w5(32'hb9b6d994),
	.w6(32'h3c6fdbfb),
	.w7(32'h3c322b29),
	.w8(32'h3981449e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97a047),
	.w1(32'h3bb3b735),
	.w2(32'h3b2c9429),
	.w3(32'h3a8f8958),
	.w4(32'hba66769a),
	.w5(32'hb992dd90),
	.w6(32'h3ba8d224),
	.w7(32'hb9b51b9e),
	.w8(32'hb93926e0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14bf2a),
	.w1(32'h3b5daf7a),
	.w2(32'h39400da1),
	.w3(32'h3b9ca40a),
	.w4(32'h3bdc36d1),
	.w5(32'hbb471b4f),
	.w6(32'h3bb1485b),
	.w7(32'h3afd9f9b),
	.w8(32'hbb1ff708),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04eccc),
	.w1(32'hbac623bd),
	.w2(32'h3a848745),
	.w3(32'hbb342de4),
	.w4(32'hbb2079df),
	.w5(32'h3b85b8bf),
	.w6(32'hbbc179d8),
	.w7(32'h3b3ee23b),
	.w8(32'hbb312a58),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f5d1a),
	.w1(32'hbb7a78ea),
	.w2(32'h3a17f8d0),
	.w3(32'h3bc77217),
	.w4(32'h3c3a8e71),
	.w5(32'hbc044c5b),
	.w6(32'h3ab2acf0),
	.w7(32'h3b269763),
	.w8(32'hbb8d380d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0280c),
	.w1(32'hba9a9cf5),
	.w2(32'h3a8bfe40),
	.w3(32'hbb88b2e5),
	.w4(32'h39379400),
	.w5(32'hba471e6f),
	.w6(32'h39554d8a),
	.w7(32'h3b6d3851),
	.w8(32'h399e8597),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2820a1),
	.w1(32'h3b1e50c6),
	.w2(32'h3b312643),
	.w3(32'h3b13d933),
	.w4(32'hbaec51b9),
	.w5(32'h39da2b70),
	.w6(32'h3b8f1d9b),
	.w7(32'hba5013cc),
	.w8(32'hb9c40c10),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6324a),
	.w1(32'hba08afc3),
	.w2(32'hbaa230ec),
	.w3(32'hba3e2531),
	.w4(32'h3a998245),
	.w5(32'h3976b370),
	.w6(32'hb90497f7),
	.w7(32'hbaca371a),
	.w8(32'hbb0b9156),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b71b7),
	.w1(32'hbbc7e9f9),
	.w2(32'hbbfc25eb),
	.w3(32'hbb17d8e5),
	.w4(32'hbbbe5746),
	.w5(32'hbba8c6b7),
	.w6(32'hbb11f85b),
	.w7(32'hbbc9294f),
	.w8(32'hbb08b773),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9a93f),
	.w1(32'hbad06d40),
	.w2(32'hbae1ffbe),
	.w3(32'hbbe05a0e),
	.w4(32'hbc06e00d),
	.w5(32'hbbf456f2),
	.w6(32'hbc146f9a),
	.w7(32'hb9d8e06a),
	.w8(32'hbbf29681),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f23b5f),
	.w1(32'h3c86596e),
	.w2(32'h37bbc1b7),
	.w3(32'h3c30c9f4),
	.w4(32'h3bff02f1),
	.w5(32'h3ac49406),
	.w6(32'h3c310632),
	.w7(32'hbb48fc87),
	.w8(32'hbbc9f197),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd59b16),
	.w1(32'h3c4a68fd),
	.w2(32'h3be6885e),
	.w3(32'h3c1439a8),
	.w4(32'h3c21241b),
	.w5(32'h3b46258a),
	.w6(32'h3bd4cf30),
	.w7(32'h3b6ceff1),
	.w8(32'h3b45c947),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86a8ec),
	.w1(32'h3ae6df7e),
	.w2(32'hbb36996e),
	.w3(32'h3bc7c8ff),
	.w4(32'hb998fe40),
	.w5(32'hbb3d3449),
	.w6(32'h3bf0e10f),
	.w7(32'h3b48ea13),
	.w8(32'hbb324693),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84541c),
	.w1(32'hbb20e7b4),
	.w2(32'hbaa6f533),
	.w3(32'hbb53e239),
	.w4(32'hbb152024),
	.w5(32'hbb7a617a),
	.w6(32'hbb988946),
	.w7(32'hbb014479),
	.w8(32'hbaab05f1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87cd28),
	.w1(32'hba96367a),
	.w2(32'hbb9e2bdf),
	.w3(32'hba0a44e1),
	.w4(32'hba4a8881),
	.w5(32'hbbdc60e3),
	.w6(32'h3b35800e),
	.w7(32'h3abb9d98),
	.w8(32'hbc44d39c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf33759),
	.w1(32'hbc081c5d),
	.w2(32'hbc10eb71),
	.w3(32'hbbb9c6f6),
	.w4(32'hbb765449),
	.w5(32'hbb0d75fe),
	.w6(32'hbc136827),
	.w7(32'hbbf5e2c5),
	.w8(32'hbbad7b52),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77ca38),
	.w1(32'hbbc259d8),
	.w2(32'hbb840507),
	.w3(32'hbbcd438d),
	.w4(32'hbb904c7d),
	.w5(32'hbb8146b5),
	.w6(32'hbbbde184),
	.w7(32'hbbe9fc28),
	.w8(32'h3ac2fb92),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05614d),
	.w1(32'h3c03a28a),
	.w2(32'h3b1bdd3d),
	.w3(32'h3c187974),
	.w4(32'h3bf4b5a9),
	.w5(32'h37ef0b18),
	.w6(32'h3c57ca75),
	.w7(32'h3c14fecc),
	.w8(32'h3a8efa57),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a309c06),
	.w1(32'hbb160535),
	.w2(32'hba845561),
	.w3(32'hbac5e864),
	.w4(32'h3afaaa23),
	.w5(32'hbb70ba1f),
	.w6(32'h3aa88004),
	.w7(32'h3b6aee0c),
	.w8(32'hbb4bb191),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb506188),
	.w1(32'hbb64e5c5),
	.w2(32'hbbbe5f39),
	.w3(32'hbb3c673d),
	.w4(32'hbb8dd1f1),
	.w5(32'h3b1cb5f5),
	.w6(32'hbbabe529),
	.w7(32'hbbac90ca),
	.w8(32'hbad002ae),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6228a5),
	.w1(32'hbc909a00),
	.w2(32'hbc6c8a2b),
	.w3(32'hbc916a45),
	.w4(32'hbc913d3c),
	.w5(32'hbc5fd248),
	.w6(32'hbcb0e2b1),
	.w7(32'hbc70a47d),
	.w8(32'hbc35ddaf),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d5a59d),
	.w1(32'hbb79abce),
	.w2(32'h3869d46e),
	.w3(32'hba4f9651),
	.w4(32'hbad4985c),
	.w5(32'h3bdc19b6),
	.w6(32'h3a84fff0),
	.w7(32'hb92b0216),
	.w8(32'h3be82afc),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b374fe3),
	.w1(32'h3b8c8f02),
	.w2(32'h3a412a72),
	.w3(32'h3be74aa0),
	.w4(32'h3bf6548b),
	.w5(32'h3b1270f9),
	.w6(32'h3c08ae2b),
	.w7(32'h3bbef8bf),
	.w8(32'h3b132c13),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0419b6),
	.w1(32'h3b13cac8),
	.w2(32'h3b166e2e),
	.w3(32'hba697d51),
	.w4(32'hba89ff44),
	.w5(32'hba9ef2eb),
	.w6(32'h3a85d2da),
	.w7(32'h3a9018e0),
	.w8(32'hbaa29ba1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae357ca),
	.w1(32'hbabe2602),
	.w2(32'hba804980),
	.w3(32'hbb10f46b),
	.w4(32'h3985b1b1),
	.w5(32'h3aba582a),
	.w6(32'h3ab9f19a),
	.w7(32'h3a7f5491),
	.w8(32'h393adf35),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb679891),
	.w1(32'hbb9e1041),
	.w2(32'hbbfa1f0a),
	.w3(32'hb7a8a01f),
	.w4(32'hbb4e37e1),
	.w5(32'hbb0ca46a),
	.w6(32'hbb02d62f),
	.w7(32'hbbd776ea),
	.w8(32'h3b30b0f1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb922f4e),
	.w1(32'hbc7113fc),
	.w2(32'hbc883e0d),
	.w3(32'hbc801a5d),
	.w4(32'hbc957c2e),
	.w5(32'hbc0ab4ca),
	.w6(32'hbc6b5504),
	.w7(32'hbc4cfbf2),
	.w8(32'hbc06290b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdad74),
	.w1(32'hbb83d314),
	.w2(32'hbb9cb0bd),
	.w3(32'hbbe42421),
	.w4(32'hbb9ad58d),
	.w5(32'h3a2d788d),
	.w6(32'hbb93ac43),
	.w7(32'hbb84982b),
	.w8(32'hbb0a49fd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17e226),
	.w1(32'h39b6f3cf),
	.w2(32'h39048884),
	.w3(32'hbb1cf382),
	.w4(32'hba990338),
	.w5(32'hbb17650a),
	.w6(32'hb59bb788),
	.w7(32'hbb5ee389),
	.w8(32'hbb19b5c6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb7071),
	.w1(32'hbb1c17a1),
	.w2(32'hb795b3ef),
	.w3(32'hbb56f887),
	.w4(32'h3a79f48e),
	.w5(32'hbb2f84a1),
	.w6(32'hbbb68d2f),
	.w7(32'hba3a192f),
	.w8(32'hbac60198),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade996f),
	.w1(32'hbbe0dbf9),
	.w2(32'hbbcd7f4c),
	.w3(32'hbb6d53a3),
	.w4(32'hbbb333be),
	.w5(32'h3bb9bd3b),
	.w6(32'hbba97f28),
	.w7(32'hbbcb0697),
	.w8(32'h3bd053a2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f08f2),
	.w1(32'h3bc45e2d),
	.w2(32'h3a8bd628),
	.w3(32'h3be71790),
	.w4(32'h3c0a8fd8),
	.w5(32'hbbbadeaa),
	.w6(32'h3c127fb6),
	.w7(32'h3bc4c75e),
	.w8(32'hbbb5f9ab),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8db70),
	.w1(32'hbb829aca),
	.w2(32'hbbe407d8),
	.w3(32'hbbf91bb6),
	.w4(32'hbb11a1a8),
	.w5(32'h3a8cff04),
	.w6(32'hbc199659),
	.w7(32'hbbae6569),
	.w8(32'h3a584064),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5c957),
	.w1(32'hbb783915),
	.w2(32'hba6dfc5a),
	.w3(32'hbb31e138),
	.w4(32'hb9cb4320),
	.w5(32'h3b07a519),
	.w6(32'hbb87448f),
	.w7(32'hb98c6dbb),
	.w8(32'h3ae3d774),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26a81c),
	.w1(32'hbbd7dac4),
	.w2(32'hba121e45),
	.w3(32'hbc16b60f),
	.w4(32'hb8883531),
	.w5(32'hbb5b4964),
	.w6(32'hbba9d455),
	.w7(32'hb951623e),
	.w8(32'hbb8f2ac0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a470cdb),
	.w1(32'hb9222a40),
	.w2(32'hb8c4d3e8),
	.w3(32'h3a457804),
	.w4(32'h3ac2f9fd),
	.w5(32'hba6163c0),
	.w6(32'h3a2d9bad),
	.w7(32'h3a54a7ee),
	.w8(32'hba867b55),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39964838),
	.w1(32'hbb4ae301),
	.w2(32'hbb12e4ee),
	.w3(32'hbb138f8d),
	.w4(32'hbb4ba891),
	.w5(32'hbb2438b9),
	.w6(32'hbb1652e6),
	.w7(32'hbb210a61),
	.w8(32'hbb6db5bc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba926c35),
	.w1(32'hbb0bfd15),
	.w2(32'hba7fc760),
	.w3(32'hba9b4893),
	.w4(32'h3afccffb),
	.w5(32'hba76ff7c),
	.w6(32'hb92845ec),
	.w7(32'h3a111563),
	.w8(32'hbb29880d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15727a),
	.w1(32'hb9484509),
	.w2(32'hbb1e61ba),
	.w3(32'h3a313d67),
	.w4(32'h39dd162d),
	.w5(32'h3bbfdf42),
	.w6(32'h39a999b1),
	.w7(32'hbab649ee),
	.w8(32'h3c192cc2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd41639),
	.w1(32'hb9d88e94),
	.w2(32'hbb7b779a),
	.w3(32'h3a33a67b),
	.w4(32'hbaa27d8a),
	.w5(32'hbbdaf863),
	.w6(32'hbaa69e41),
	.w7(32'hbbe3e47a),
	.w8(32'hbbbba295),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb171579),
	.w1(32'h3b850433),
	.w2(32'hba1a9682),
	.w3(32'hbb79dc08),
	.w4(32'hbbf0f59d),
	.w5(32'hbb9bcb02),
	.w6(32'hbb993605),
	.w7(32'hbbe34b36),
	.w8(32'hbbe4963e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61af29),
	.w1(32'hbc384a7a),
	.w2(32'hbc347abd),
	.w3(32'hbc7a1a96),
	.w4(32'hbbec3975),
	.w5(32'hbb25f954),
	.w6(32'hbc3161c5),
	.w7(32'hbbe8803a),
	.w8(32'hbb5fa55c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc51084),
	.w1(32'h3c12692e),
	.w2(32'h3ae5825c),
	.w3(32'h3c3f280f),
	.w4(32'h3bd558c3),
	.w5(32'hbb7d86b0),
	.w6(32'h3bea9394),
	.w7(32'hb95a0748),
	.w8(32'hbbe43a54),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f9fa8),
	.w1(32'hbb01e45b),
	.w2(32'hbb89c334),
	.w3(32'hbb666a47),
	.w4(32'hbb975ab0),
	.w5(32'h3b062c2b),
	.w6(32'hbaea039c),
	.w7(32'hbb66d87a),
	.w8(32'h3a99ca56),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c53ac),
	.w1(32'h3b80aac0),
	.w2(32'h3ae147af),
	.w3(32'h3b43e3b1),
	.w4(32'hbb1bc2c7),
	.w5(32'h3b595a1c),
	.w6(32'h3bd55915),
	.w7(32'hbb0c5f57),
	.w8(32'hba88caee),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381019b5),
	.w1(32'hbaf13868),
	.w2(32'hbb5ab17d),
	.w3(32'h3b3f91f5),
	.w4(32'h3b089bf6),
	.w5(32'hbb312b60),
	.w6(32'hb9d6f648),
	.w7(32'hbb80c7b9),
	.w8(32'hbb3fd9af),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11d52a),
	.w1(32'hbb9bb85f),
	.w2(32'h3af612a1),
	.w3(32'h3a25757e),
	.w4(32'hb91c9542),
	.w5(32'h3b49159c),
	.w6(32'hbba3e581),
	.w7(32'h3ba66b14),
	.w8(32'h3b98fd55),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ca6f2),
	.w1(32'hb920006e),
	.w2(32'hbbacdaaf),
	.w3(32'h3b496efb),
	.w4(32'hbb1f3605),
	.w5(32'hbac8bade),
	.w6(32'h3b68deed),
	.w7(32'hbbd7aebe),
	.w8(32'hbb04d46c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9876f4),
	.w1(32'hbc2f0295),
	.w2(32'hb9988d84),
	.w3(32'hbbfa95ab),
	.w4(32'hbc25cda2),
	.w5(32'hb90cbf79),
	.w6(32'hbc38c626),
	.w7(32'hbb020508),
	.w8(32'h3b192cc9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012828),
	.w1(32'hbc48a925),
	.w2(32'hbc565ac2),
	.w3(32'hbc35801d),
	.w4(32'hbc984590),
	.w5(32'hbb43bd9f),
	.w6(32'hbcaa5360),
	.w7(32'hbc667292),
	.w8(32'hb90c2c9b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06be29),
	.w1(32'h3bc0b15b),
	.w2(32'h3a4ba29d),
	.w3(32'h3b84b7ec),
	.w4(32'h3a58a3fc),
	.w5(32'hbb54f367),
	.w6(32'h3b72de2e),
	.w7(32'hbab8846f),
	.w8(32'h3b3185b1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99864d),
	.w1(32'h3af22c11),
	.w2(32'h3a818f17),
	.w3(32'h3aa389a2),
	.w4(32'h3b20c4ec),
	.w5(32'h3ab60f28),
	.w6(32'h3ac292bf),
	.w7(32'h39fc53a7),
	.w8(32'h3b42faca),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f59fe),
	.w1(32'h3a665f49),
	.w2(32'h3b928b57),
	.w3(32'hbaef221a),
	.w4(32'hbb4dd20b),
	.w5(32'h3bd52c7e),
	.w6(32'h3a2c6db2),
	.w7(32'h39fe5f3e),
	.w8(32'h3bbcef08),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c027b2b),
	.w1(32'h3be684f2),
	.w2(32'h3bbf7907),
	.w3(32'h3c0de77a),
	.w4(32'h3c193869),
	.w5(32'h3a9466de),
	.w6(32'h3b951cb8),
	.w7(32'h3b9d7cef),
	.w8(32'h3a6ce5df),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb706f6a),
	.w1(32'hbc0d7dd2),
	.w2(32'hbbf7bcde),
	.w3(32'hbb604a40),
	.w4(32'hbbaf8304),
	.w5(32'hbb6a56ca),
	.w6(32'hbba253b1),
	.w7(32'hbb45a048),
	.w8(32'hbb00bf27),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87d973e),
	.w1(32'hba9d9ccc),
	.w2(32'hba9097f7),
	.w3(32'hba5ea855),
	.w4(32'hbb11a720),
	.w5(32'hbc116e12),
	.w6(32'hbb00bf0b),
	.w7(32'hbb46e755),
	.w8(32'hbc077979),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6b8ce),
	.w1(32'hbb989ea3),
	.w2(32'hbc3c8224),
	.w3(32'hbbe263d1),
	.w4(32'hbc4f8c6c),
	.w5(32'hba85d75a),
	.w6(32'hbbb77c51),
	.w7(32'hbc4b0339),
	.w8(32'hbaa2555a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39336354),
	.w1(32'h3a05f0bb),
	.w2(32'h39f9883d),
	.w3(32'hb9ad4b6e),
	.w4(32'hbac3f426),
	.w5(32'h3ab9e228),
	.w6(32'hbaa26e9a),
	.w7(32'hbb2e2bb9),
	.w8(32'h3b0d9821),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b134266),
	.w1(32'hba7a71d1),
	.w2(32'h3b827848),
	.w3(32'hbb1d66e2),
	.w4(32'h3b852bc1),
	.w5(32'h3b530a77),
	.w6(32'h39be7514),
	.w7(32'h3b810fac),
	.w8(32'h3ba40f3f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93f75a),
	.w1(32'h3b1c63fd),
	.w2(32'hbb0b6638),
	.w3(32'h3bc029a2),
	.w4(32'h3bbd2fc7),
	.w5(32'h3b692194),
	.w6(32'h3b306d29),
	.w7(32'hba9dc293),
	.w8(32'hb9985f19),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a3f84),
	.w1(32'h3aad7e21),
	.w2(32'h3ab41c0a),
	.w3(32'h3a271949),
	.w4(32'hbab42b2d),
	.w5(32'h3b0bf04b),
	.w6(32'h3a6c230f),
	.w7(32'h3a018083),
	.w8(32'h3a84dbc5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a744718),
	.w1(32'h3b03aafa),
	.w2(32'h3aee1c75),
	.w3(32'h3b80952e),
	.w4(32'h3b28594d),
	.w5(32'hbaef10e1),
	.w6(32'h3b9f8042),
	.w7(32'h3aa8b692),
	.w8(32'h3b75de40),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7dea3f),
	.w1(32'hbc698ea7),
	.w2(32'hbbc9099d),
	.w3(32'hbca89a74),
	.w4(32'hbc7816f7),
	.w5(32'h3bd268d5),
	.w6(32'hbca9673a),
	.w7(32'hbbab8529),
	.w8(32'h3bcdcd55),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c002316),
	.w1(32'h3c5ad9fc),
	.w2(32'h3bde4483),
	.w3(32'h3bfac8ec),
	.w4(32'h3a858f51),
	.w5(32'hbb7d4edc),
	.w6(32'h3c3ae0e2),
	.w7(32'h3b94b984),
	.w8(32'hbb975fff),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b69f6),
	.w1(32'hbb629489),
	.w2(32'hbb2bfb76),
	.w3(32'hbc0b72f8),
	.w4(32'hbb310cf5),
	.w5(32'hbadc4eb6),
	.w6(32'hbbd47852),
	.w7(32'hbabf1619),
	.w8(32'hbb856552),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7973b8),
	.w1(32'h3af3a5d8),
	.w2(32'h3b1bc49c),
	.w3(32'h3a504294),
	.w4(32'h3c1a8590),
	.w5(32'hbb91a6d5),
	.w6(32'h3a521bb1),
	.w7(32'h3b188eba),
	.w8(32'hbba92e7c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e96b3),
	.w1(32'hbb945b0f),
	.w2(32'hbb1fa4ce),
	.w3(32'hbb422c46),
	.w4(32'h3b2a3e4a),
	.w5(32'h3a22f0a7),
	.w6(32'hbaea0fea),
	.w7(32'h3b0c2db8),
	.w8(32'h3aa9abd9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915c26b),
	.w1(32'h3bc9fd4e),
	.w2(32'h3ad422d3),
	.w3(32'h3bd94124),
	.w4(32'h3b2fcdd1),
	.w5(32'hbaa9bad8),
	.w6(32'h3bf71acc),
	.w7(32'h38520c17),
	.w8(32'hbb90af14),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb371693),
	.w1(32'h3aeb2e03),
	.w2(32'hbbad4aea),
	.w3(32'h3b8c5934),
	.w4(32'h3957a706),
	.w5(32'h3b78e070),
	.w6(32'h3b5ab9da),
	.w7(32'hbbba7630),
	.w8(32'h3a9411ee),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eabe5),
	.w1(32'h3b2e66bb),
	.w2(32'h3c12b93c),
	.w3(32'h3ba9e2e5),
	.w4(32'h3bd671d0),
	.w5(32'hbbce223f),
	.w6(32'h3b42d153),
	.w7(32'h3c17e842),
	.w8(32'hbb79a485),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3041c),
	.w1(32'hbb0278fa),
	.w2(32'hb9b2080a),
	.w3(32'hbbe907f7),
	.w4(32'hbb727ed1),
	.w5(32'h3b2e9d9e),
	.w6(32'hbb3fbddf),
	.w7(32'h3acd5a80),
	.w8(32'h3ab0bac5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1795a),
	.w1(32'hbb3ad2df),
	.w2(32'hbbf57a24),
	.w3(32'h3b5d2078),
	.w4(32'h3bdbe0d9),
	.w5(32'hbb04d3e8),
	.w6(32'hbb6eacaa),
	.w7(32'hba40f044),
	.w8(32'hbb80a3fd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c073e7f),
	.w1(32'h3d2f3223),
	.w2(32'h3b628aa0),
	.w3(32'hbd3df255),
	.w4(32'hbd01d44f),
	.w5(32'hba916f64),
	.w6(32'hbd16698e),
	.w7(32'hbca44c56),
	.w8(32'hbaf35ba2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34166b),
	.w1(32'h3c6999a5),
	.w2(32'h3bb6d489),
	.w3(32'h3c15a5c2),
	.w4(32'h3c5691b3),
	.w5(32'h3b3988ea),
	.w6(32'h3c2ce33e),
	.w7(32'h3c5120d0),
	.w8(32'hbbda5dbb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c244395),
	.w1(32'h3cd46cb6),
	.w2(32'h3c27fc41),
	.w3(32'h3bc7eae9),
	.w4(32'h3c00a772),
	.w5(32'h3b62d5fc),
	.w6(32'hbba50369),
	.w7(32'hbba319b9),
	.w8(32'h3ab17f8a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b139d13),
	.w1(32'h399efbc4),
	.w2(32'hba699714),
	.w3(32'hbb5ea652),
	.w4(32'hbb88013e),
	.w5(32'h3c179641),
	.w6(32'hbb8e7463),
	.w7(32'h3a920f0f),
	.w8(32'hb8d9e7bb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae83a2),
	.w1(32'hbc20ef50),
	.w2(32'hb8da4724),
	.w3(32'h3ca584f8),
	.w4(32'h3c461086),
	.w5(32'hbc139a07),
	.w6(32'h3b0609a8),
	.w7(32'h3b80cc7d),
	.w8(32'hbc230651),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f100d),
	.w1(32'hbca893dd),
	.w2(32'hbc8b32ba),
	.w3(32'hbcc2e937),
	.w4(32'hbd1c72a6),
	.w5(32'hbcafde65),
	.w6(32'hbd354cc0),
	.w7(32'hbca385a5),
	.w8(32'hbc3beb06),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1157cd),
	.w1(32'h3d2fa114),
	.w2(32'h3bec87a0),
	.w3(32'hbce4aeef),
	.w4(32'hbcb7bdf2),
	.w5(32'hbc017c82),
	.w6(32'hbc877b82),
	.w7(32'hbc829156),
	.w8(32'hbc5d14f2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d23b80),
	.w1(32'h3cadeb78),
	.w2(32'h3c8a9382),
	.w3(32'hbc68aacb),
	.w4(32'hbb64d648),
	.w5(32'h3b56e4da),
	.w6(32'hbbe49281),
	.w7(32'hbc506a32),
	.w8(32'h3bacf32c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3881d559),
	.w1(32'h3c621db8),
	.w2(32'hba3c81e4),
	.w3(32'hbb6e1ecf),
	.w4(32'hbb31951c),
	.w5(32'h3be66fe1),
	.w6(32'h3b30fce0),
	.w7(32'hba9af692),
	.w8(32'h3b89acfd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fd6a5),
	.w1(32'hbbecb1c4),
	.w2(32'hbc00a448),
	.w3(32'hb9e5f030),
	.w4(32'h3baa63f1),
	.w5(32'hbaaabb5b),
	.w6(32'hbb92266b),
	.w7(32'hbaafc0fc),
	.w8(32'hbad4e982),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90cd85),
	.w1(32'hbb919bf9),
	.w2(32'hbb530905),
	.w3(32'h3c28354b),
	.w4(32'h3c0eff20),
	.w5(32'hbbcaa42d),
	.w6(32'h3bbe5389),
	.w7(32'hb9fe7f28),
	.w8(32'hbb27125a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b25cd),
	.w1(32'h3c0db31a),
	.w2(32'h3bff886d),
	.w3(32'hbc01470c),
	.w4(32'hbbb684fd),
	.w5(32'hb9c5da83),
	.w6(32'hbbb0063c),
	.w7(32'hbb868e57),
	.w8(32'hbb7a102a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e4c31),
	.w1(32'hbb74fbdd),
	.w2(32'h3a3011b0),
	.w3(32'h3a312512),
	.w4(32'hbb31f76f),
	.w5(32'hba1a83b0),
	.w6(32'hbb18003f),
	.w7(32'h3a306f6d),
	.w8(32'h3b39b76c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8ab50),
	.w1(32'h3add1723),
	.w2(32'h39c809e7),
	.w3(32'h3a016c03),
	.w4(32'h3b993794),
	.w5(32'hba1aac97),
	.w6(32'h3b0eef04),
	.w7(32'h3a633e06),
	.w8(32'hb9975bb8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafe864),
	.w1(32'h3bd007ec),
	.w2(32'h3b3fb636),
	.w3(32'hba004c09),
	.w4(32'hbb85099d),
	.w5(32'hbac576fb),
	.w6(32'h3bae147a),
	.w7(32'h38ce003f),
	.w8(32'hbbd10ef6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1c50d),
	.w1(32'h3d1a4b8b),
	.w2(32'hbc010917),
	.w3(32'hbb789710),
	.w4(32'h3baffba0),
	.w5(32'hbb5b8e74),
	.w6(32'hbbca9e76),
	.w7(32'h3b3dea15),
	.w8(32'hbba65811),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba202c3f),
	.w1(32'h3a8fd665),
	.w2(32'h3bb849f3),
	.w3(32'hbb22897d),
	.w4(32'hbb73974e),
	.w5(32'hbaf0e3a4),
	.w6(32'hbb93aff8),
	.w7(32'hba53fd98),
	.w8(32'hbb115e6e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcdac1),
	.w1(32'hbbbd8e9f),
	.w2(32'hbc2000c4),
	.w3(32'hbb8e614d),
	.w4(32'hbc11fc82),
	.w5(32'hbbb889e5),
	.w6(32'hbb2433c0),
	.w7(32'hbbf1ec53),
	.w8(32'hbbba7e49),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4af760),
	.w1(32'h3bd432c9),
	.w2(32'h3b6c4c35),
	.w3(32'hb9952e9e),
	.w4(32'h3bbee05b),
	.w5(32'h3c2d9b3d),
	.w6(32'hbc2c41d5),
	.w7(32'hbc2e8426),
	.w8(32'h3be120cc),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb329e),
	.w1(32'hbb6ffd40),
	.w2(32'hbbc3d80c),
	.w3(32'hbb0dfe5c),
	.w4(32'h3b68f579),
	.w5(32'h3a8494f3),
	.w6(32'hb92f948e),
	.w7(32'h3b101191),
	.w8(32'hbc0db5a4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb999e82),
	.w1(32'hbbd578d5),
	.w2(32'hbb951114),
	.w3(32'h3c0c08a3),
	.w4(32'h3be1d6a3),
	.w5(32'h3b8b2292),
	.w6(32'hbbd32316),
	.w7(32'hbb956452),
	.w8(32'h3b6656a2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c237ff5),
	.w1(32'h3c5d57a7),
	.w2(32'h3bdb8a99),
	.w3(32'h3bca5ed2),
	.w4(32'h3b57f911),
	.w5(32'h3b329637),
	.w6(32'h3c12b081),
	.w7(32'h3b8f8c09),
	.w8(32'hbad0bacf),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1898c6),
	.w1(32'hbc3569fd),
	.w2(32'hbb1f5035),
	.w3(32'hbabe4885),
	.w4(32'hbb40379c),
	.w5(32'hbc0f5422),
	.w6(32'hbbb749cf),
	.w7(32'h3b931143),
	.w8(32'hbbf6cc52),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8fb2a),
	.w1(32'h3bf34ed0),
	.w2(32'h3bb5c941),
	.w3(32'hbb7bfdf6),
	.w4(32'h3b9cec7d),
	.w5(32'h39024f7f),
	.w6(32'hbc091570),
	.w7(32'hbc2f8a62),
	.w8(32'hba953051),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc57027),
	.w1(32'h3bb484bd),
	.w2(32'hb9ef845d),
	.w3(32'h3b7e00e9),
	.w4(32'h3b1e4580),
	.w5(32'hbb871a3d),
	.w6(32'h3bf5f5eb),
	.w7(32'h3b0c9e6e),
	.w8(32'hbac095da),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad9d81),
	.w1(32'hbbf23041),
	.w2(32'hbbd88ca1),
	.w3(32'h3983dfce),
	.w4(32'hbb2d5953),
	.w5(32'h3ae596af),
	.w6(32'hbae9cb46),
	.w7(32'hbb50eeec),
	.w8(32'hbb04d264),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbad73a),
	.w1(32'h3a9685d0),
	.w2(32'hbadbb3e9),
	.w3(32'h3abfaa32),
	.w4(32'h3b18c9a9),
	.w5(32'h3b32297a),
	.w6(32'h3bae3e2c),
	.w7(32'h3a8eaab3),
	.w8(32'hba565cb8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcdfff),
	.w1(32'h3b5b1937),
	.w2(32'hb7499838),
	.w3(32'h3c275f31),
	.w4(32'h3b413e8d),
	.w5(32'hbc011ce4),
	.w6(32'hb931632c),
	.w7(32'hbb12e7fe),
	.w8(32'hbac238aa),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c233ac3),
	.w1(32'h3c63e9e0),
	.w2(32'hbb9d1b5a),
	.w3(32'hbba2e5e0),
	.w4(32'h3b310ae2),
	.w5(32'hbba540ff),
	.w6(32'h3a97b7a6),
	.w7(32'h3befa771),
	.w8(32'hbb2e406a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa93cf6),
	.w1(32'hba8e2d14),
	.w2(32'h3b8dde57),
	.w3(32'hbb4a9211),
	.w4(32'hba67fd92),
	.w5(32'h3b10911b),
	.w6(32'h3ab107da),
	.w7(32'h3abcaa07),
	.w8(32'h3acb8464),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2fa27),
	.w1(32'h3b9e574c),
	.w2(32'hbb488d38),
	.w3(32'h3beb0282),
	.w4(32'h39d8e6b8),
	.w5(32'h3b8ee3a3),
	.w6(32'hbace31d1),
	.w7(32'hbc012fa2),
	.w8(32'hbbd10d0d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb256c1c),
	.w1(32'hbae19041),
	.w2(32'hba25f5cf),
	.w3(32'hba6bae6a),
	.w4(32'hbb518fe6),
	.w5(32'h393fea89),
	.w6(32'hbbca84cd),
	.w7(32'hbb2e22b2),
	.w8(32'h3b485d76),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb146817),
	.w1(32'hbc23e886),
	.w2(32'hbc047c1d),
	.w3(32'h3baab9d7),
	.w4(32'h3b1a5d56),
	.w5(32'hb97172fc),
	.w6(32'hb984b73f),
	.w7(32'h39253ce1),
	.w8(32'hbc9cd4f8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6599e8),
	.w1(32'h3c0ce99b),
	.w2(32'h39f41a46),
	.w3(32'h3b43b9ee),
	.w4(32'h3c286715),
	.w5(32'h3ace5fe4),
	.w6(32'hbc2476bf),
	.w7(32'hbc2c9614),
	.w8(32'h3ac7b764),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2816c6),
	.w1(32'h3b814d35),
	.w2(32'hb7e9046e),
	.w3(32'h3bdb12ad),
	.w4(32'h3be3bcd1),
	.w5(32'h3ac6ab71),
	.w6(32'h3b5b4c02),
	.w7(32'h3a61f211),
	.w8(32'h3b695111),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71a61a),
	.w1(32'hb9e11648),
	.w2(32'hbb8400fc),
	.w3(32'hbc710615),
	.w4(32'hbc03dd61),
	.w5(32'hbb99140c),
	.w6(32'hbc5be127),
	.w7(32'hbbef82cd),
	.w8(32'hbba25af9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa34d28),
	.w1(32'hbab8710e),
	.w2(32'hbc25c87a),
	.w3(32'h3c15c2c2),
	.w4(32'h3b8acc99),
	.w5(32'h3aee53cb),
	.w6(32'h3b15cfd5),
	.w7(32'hbafcc1cc),
	.w8(32'h3ba33e4d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7922c),
	.w1(32'h3b2f07b3),
	.w2(32'hb8d6188c),
	.w3(32'h3b089d7d),
	.w4(32'h3b94ab99),
	.w5(32'hbaca4622),
	.w6(32'h3b3a6022),
	.w7(32'h3b2f28cd),
	.w8(32'hbaad2e38),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56412f),
	.w1(32'hbc4d6b41),
	.w2(32'hbc1dc9e6),
	.w3(32'hbb64d05f),
	.w4(32'hbb7275bf),
	.w5(32'h3abcb05b),
	.w6(32'hbc167025),
	.w7(32'hbbc66593),
	.w8(32'hbaca6f08),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb820872),
	.w1(32'h3afe4e76),
	.w2(32'h39d03c76),
	.w3(32'h3b89ac8c),
	.w4(32'h3aa58188),
	.w5(32'hbb99f129),
	.w6(32'hba208022),
	.w7(32'hbb968a23),
	.w8(32'hbbc619f4),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3f7d6),
	.w1(32'h3a89983d),
	.w2(32'h3c115eff),
	.w3(32'hbbacf9ff),
	.w4(32'hbbdb54f8),
	.w5(32'hbc334aef),
	.w6(32'h3b150165),
	.w7(32'hbad4f913),
	.w8(32'hbc0d16c7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5213e),
	.w1(32'h3c1576b4),
	.w2(32'h3bbc5667),
	.w3(32'hbc6e9ffd),
	.w4(32'hbbec6d1e),
	.w5(32'hbbc35e52),
	.w6(32'hbbd957ff),
	.w7(32'hbab63d09),
	.w8(32'hba81fdc1),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0473c6),
	.w1(32'h3b82fd26),
	.w2(32'hbb88eeb1),
	.w3(32'h3b1f68ef),
	.w4(32'h3bfd13e3),
	.w5(32'hbb8cfaa6),
	.w6(32'h3c3ee12d),
	.w7(32'h3ba1e5c0),
	.w8(32'hba6949f7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15db75),
	.w1(32'h3a9136e8),
	.w2(32'h3b8c6ff9),
	.w3(32'hbb907555),
	.w4(32'h3a1de5dd),
	.w5(32'hbb97bfb6),
	.w6(32'hbb12b858),
	.w7(32'hbb188921),
	.w8(32'h3b1e6746),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0a1b3),
	.w1(32'h3b57828d),
	.w2(32'h3a250db3),
	.w3(32'hbb609867),
	.w4(32'h3af9ded8),
	.w5(32'hbab661e0),
	.w6(32'hbb6d8371),
	.w7(32'h3b87b790),
	.w8(32'h382b90a4),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39471bb2),
	.w1(32'h3c6959af),
	.w2(32'h3b7979bc),
	.w3(32'hbbf79b10),
	.w4(32'h3aae06b9),
	.w5(32'hbc26e744),
	.w6(32'h39b7a4ad),
	.w7(32'hba9a1e3a),
	.w8(32'hbbfa8f4a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b983a62),
	.w1(32'h3cc0d0fd),
	.w2(32'h3c4da10c),
	.w3(32'hbc7d33e0),
	.w4(32'hbc07c177),
	.w5(32'hbaaa70f9),
	.w6(32'hbc379a35),
	.w7(32'hbbc9afae),
	.w8(32'hbadcb66f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66f58a),
	.w1(32'h3c40875a),
	.w2(32'h3b9e428f),
	.w3(32'h3b6dbc99),
	.w4(32'h3a9814dd),
	.w5(32'hbbdec102),
	.w6(32'hbc006634),
	.w7(32'hbbc286d2),
	.w8(32'hbbfaa9ec),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ca2b0),
	.w1(32'hbb3538f1),
	.w2(32'h3bd3fc16),
	.w3(32'hbc2d4cb3),
	.w4(32'hbc00a2d0),
	.w5(32'h3a938da8),
	.w6(32'hbbf1ac93),
	.w7(32'h3aa6fd7c),
	.w8(32'h39e912f6),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76ea55),
	.w1(32'hbaadd5be),
	.w2(32'hbb6d474a),
	.w3(32'h3b8975bf),
	.w4(32'h3be06b2b),
	.w5(32'h3bf3aa12),
	.w6(32'hbb38f81b),
	.w7(32'h3b89a09e),
	.w8(32'h3b157157),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3afcc3),
	.w1(32'hbc986590),
	.w2(32'hbc8c5dcc),
	.w3(32'h3c2b2626),
	.w4(32'h3b92fea7),
	.w5(32'hba13dbda),
	.w6(32'hb9899035),
	.w7(32'hbb8e4a43),
	.w8(32'hba5c5650),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe25f0),
	.w1(32'h3c0e7f8a),
	.w2(32'h3ba0caf3),
	.w3(32'h3bdc8d1e),
	.w4(32'hba5bd21b),
	.w5(32'hbb24646d),
	.w6(32'h3c482844),
	.w7(32'hba85de11),
	.w8(32'h3b17c152),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56315f),
	.w1(32'h3b885211),
	.w2(32'hbba2f52f),
	.w3(32'hbb53a69a),
	.w4(32'hb8c1ceda),
	.w5(32'hbbebebe7),
	.w6(32'hbc564011),
	.w7(32'h3b7f0424),
	.w8(32'hbc4ded56),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6455af),
	.w1(32'h3cb0960f),
	.w2(32'h3bee9628),
	.w3(32'hbb0d0fca),
	.w4(32'h3bc5c2bb),
	.w5(32'hbb582973),
	.w6(32'h3bd4d909),
	.w7(32'h3bdab3c5),
	.w8(32'hbb1be2e1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d6eb8),
	.w1(32'h3c3e35f8),
	.w2(32'h3bc97bd0),
	.w3(32'hbb258cc4),
	.w4(32'h3acfbe41),
	.w5(32'h3aeb2c1a),
	.w6(32'h396037f8),
	.w7(32'h3a538c45),
	.w8(32'hb96030b1),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2602b3),
	.w1(32'hbb566d7b),
	.w2(32'hb996860e),
	.w3(32'hbb878332),
	.w4(32'h3a7943db),
	.w5(32'hbb38e43e),
	.w6(32'hbb464499),
	.w7(32'hbada76e6),
	.w8(32'hbba22025),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20cbb4),
	.w1(32'hbb13b722),
	.w2(32'hbb04c622),
	.w3(32'hba635f89),
	.w4(32'h3b49778b),
	.w5(32'hb79ca1e2),
	.w6(32'hbaa3e5e5),
	.w7(32'hb8c8b250),
	.w8(32'h3b95441e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ba650),
	.w1(32'h3c8538d2),
	.w2(32'h3c2be5de),
	.w3(32'h3a8b446d),
	.w4(32'h3bc0c834),
	.w5(32'h3be47745),
	.w6(32'h3b533afc),
	.w7(32'h3aa73d74),
	.w8(32'h3b98e5d5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ad8f5),
	.w1(32'h3a93bfa8),
	.w2(32'h3a7a628b),
	.w3(32'h39b5b4bd),
	.w4(32'hbaafeaa7),
	.w5(32'hbb238a86),
	.w6(32'h3b48dbfa),
	.w7(32'h3bac2b88),
	.w8(32'hbb26387c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58fce4),
	.w1(32'h3b8fef1a),
	.w2(32'h3ad485e3),
	.w3(32'hbc1ef14e),
	.w4(32'hbcad8eeb),
	.w5(32'hbbaa1688),
	.w6(32'h3907a6a1),
	.w7(32'hbb222458),
	.w8(32'h3b510308),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c3c33),
	.w1(32'h3b781520),
	.w2(32'hb9ef3621),
	.w3(32'hb91965ba),
	.w4(32'hbba4ab32),
	.w5(32'h3b8afe96),
	.w6(32'h3ba03572),
	.w7(32'hba71e3c5),
	.w8(32'hbbcd4f61),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dc93d),
	.w1(32'h3c6d6a67),
	.w2(32'hbbec9565),
	.w3(32'hbc25d251),
	.w4(32'hbc187db1),
	.w5(32'hbc964a01),
	.w6(32'hbc874ec4),
	.w7(32'h3aeaa205),
	.w8(32'hb99a39e8),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00b8d5),
	.w1(32'h3d1d122c),
	.w2(32'h3c8cc700),
	.w3(32'hbcd03ae4),
	.w4(32'hbc3071d3),
	.w5(32'hbb827e4a),
	.w6(32'hbbe86fa8),
	.w7(32'hbb8fcf20),
	.w8(32'hbbaa8e62),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5995e),
	.w1(32'hba9ee9d0),
	.w2(32'hbac2310b),
	.w3(32'hbb5ae5b9),
	.w4(32'h3bda2fb2),
	.w5(32'hbc207e7f),
	.w6(32'h3c173c10),
	.w7(32'h3c0019c1),
	.w8(32'hbbbdebc7),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca076e3),
	.w1(32'h3d2cb7d9),
	.w2(32'h3c83404e),
	.w3(32'hbcd6b147),
	.w4(32'hbc3e5f3d),
	.w5(32'hbbd02bcc),
	.w6(32'hbc22ebd7),
	.w7(32'h3a5334e0),
	.w8(32'hb9ccecf6),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf4775),
	.w1(32'h3c6f7a9e),
	.w2(32'h3bc86bfe),
	.w3(32'hbbd55e9e),
	.w4(32'hbc451d9e),
	.w5(32'hbbbe12e7),
	.w6(32'h3c1d306f),
	.w7(32'h3af7ea5b),
	.w8(32'h3a9cd322),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fc0fb),
	.w1(32'h3bd25b06),
	.w2(32'h3b85af40),
	.w3(32'hbaf0bb19),
	.w4(32'h3a345f23),
	.w5(32'hbb53ddfd),
	.w6(32'h3a0f70e2),
	.w7(32'h3a550b1b),
	.w8(32'h3a07eb8c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e6eba),
	.w1(32'h3c7ab119),
	.w2(32'h3c742f45),
	.w3(32'hbb36306c),
	.w4(32'hbb5d98f5),
	.w5(32'h3c23f06c),
	.w6(32'h3be101ef),
	.w7(32'h3b632315),
	.w8(32'h3b4cbb06),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc72cb3),
	.w1(32'hbcf9b877),
	.w2(32'hbc3f8161),
	.w3(32'h3c9f2e55),
	.w4(32'h3cb96ebe),
	.w5(32'hbb9022e6),
	.w6(32'h3c051089),
	.w7(32'h3c088cd3),
	.w8(32'hbb55a4b4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d3977),
	.w1(32'hba9d3707),
	.w2(32'h3b8b9035),
	.w3(32'hbc1a2940),
	.w4(32'hbc64c012),
	.w5(32'hbb4aed8b),
	.w6(32'hbc5f53a4),
	.w7(32'hbc53975d),
	.w8(32'hbb733651),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf6f0f),
	.w1(32'h3b934874),
	.w2(32'hbaeaf1be),
	.w3(32'hb9040aeb),
	.w4(32'h3a91ea6a),
	.w5(32'hbbb2620c),
	.w6(32'hbaf2e437),
	.w7(32'hbb63914c),
	.w8(32'hbbb2b9d2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c169c01),
	.w1(32'h3ca058a7),
	.w2(32'h3bee3d64),
	.w3(32'hba03d77d),
	.w4(32'hba288bef),
	.w5(32'hbc409f54),
	.w6(32'hbc6210e7),
	.w7(32'hbc99249f),
	.w8(32'hbc19c30c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c244767),
	.w1(32'h3cee1c95),
	.w2(32'h3b0217ee),
	.w3(32'hbcdb12b6),
	.w4(32'hbc5aed41),
	.w5(32'h3b2eb5e4),
	.w6(32'hbc532eb1),
	.w7(32'hbc3eb5b1),
	.w8(32'hba3bbc27),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88b21d),
	.w1(32'hbc188143),
	.w2(32'hbc2e42ac),
	.w3(32'h3bbb2e99),
	.w4(32'h3c16af74),
	.w5(32'h3b709398),
	.w6(32'hbc0b1e7c),
	.w7(32'hbb3c65e7),
	.w8(32'h39b62096),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33ada6),
	.w1(32'hbb62824c),
	.w2(32'h3a4c4fe0),
	.w3(32'h3bba3c0c),
	.w4(32'hbb0a34c7),
	.w5(32'h3ba8a140),
	.w6(32'h3b29683e),
	.w7(32'h3ad8f75d),
	.w8(32'h3b400879),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6a741),
	.w1(32'hbb9dba08),
	.w2(32'hba9a6a9f),
	.w3(32'h3b6a5b6d),
	.w4(32'h3bee2a2d),
	.w5(32'h3c04cb0b),
	.w6(32'hbaa03580),
	.w7(32'h38b6517f),
	.w8(32'h3b3a8dc1),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ddb26),
	.w1(32'hbca91aa2),
	.w2(32'hbc367507),
	.w3(32'h3c5ba64f),
	.w4(32'h3c02a589),
	.w5(32'hbc382406),
	.w6(32'h3b044d4f),
	.w7(32'h3aa5f752),
	.w8(32'hbb17fdfc),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c1ec3),
	.w1(32'h3c2c3844),
	.w2(32'h3bbc8197),
	.w3(32'hbc181866),
	.w4(32'hbbdd3854),
	.w5(32'h3b13f85f),
	.w6(32'hbbb87c8d),
	.w7(32'hba25366b),
	.w8(32'h398cb62c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0a263),
	.w1(32'hbc89b278),
	.w2(32'hbc412d59),
	.w3(32'h3bc54b05),
	.w4(32'h3b85a186),
	.w5(32'h3b91c694),
	.w6(32'hb9d8fc4e),
	.w7(32'hba9692a6),
	.w8(32'hbc162548),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35df78),
	.w1(32'h3c4e7387),
	.w2(32'h3b0fe71d),
	.w3(32'hb9b68c2b),
	.w4(32'hbc098340),
	.w5(32'hbbc5c463),
	.w6(32'hbc8d88a3),
	.w7(32'hbbb3f0a4),
	.w8(32'hbbf997bd),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba802fb),
	.w1(32'h3c44efe8),
	.w2(32'hb9ec2cd3),
	.w3(32'h3a533027),
	.w4(32'h3b32dc76),
	.w5(32'hbb03ee87),
	.w6(32'hbc19149f),
	.w7(32'hbc239301),
	.w8(32'hbb92e846),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf28af1),
	.w1(32'hb987931c),
	.w2(32'h3a955736),
	.w3(32'hbbfe88a7),
	.w4(32'hbc46445f),
	.w5(32'hbb8f2cd7),
	.w6(32'hbb9dd56c),
	.w7(32'hbc2fc4bf),
	.w8(32'hbb57862a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a086361),
	.w1(32'h3bc0c2e3),
	.w2(32'h3cbbb65f),
	.w3(32'hbc79c295),
	.w4(32'hbc826b8c),
	.w5(32'hbb88878d),
	.w6(32'h3b89e954),
	.w7(32'hbbe4668c),
	.w8(32'hbb2feb27),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbf24c),
	.w1(32'h3c44d414),
	.w2(32'h3b2e8cee),
	.w3(32'hbbafadd8),
	.w4(32'hbb8b239d),
	.w5(32'hbb2760a0),
	.w6(32'hbb8dce6a),
	.w7(32'h3a499d94),
	.w8(32'hbc1b7f2a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5a401),
	.w1(32'h3bf93f9e),
	.w2(32'hbbd57515),
	.w3(32'hbaac3e41),
	.w4(32'h3ad83c6f),
	.w5(32'hbbea3c89),
	.w6(32'hbbed685a),
	.w7(32'hbb26e61d),
	.w8(32'hbc0c9983),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8aaf4d),
	.w1(32'hbae2dafe),
	.w2(32'hba454f76),
	.w3(32'hbba94d8d),
	.w4(32'hbbde7f5a),
	.w5(32'hba167d38),
	.w6(32'hbbb3d765),
	.w7(32'hbb94f1ce),
	.w8(32'h3b10c1f1),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa937c),
	.w1(32'h3b808379),
	.w2(32'h3855d9a6),
	.w3(32'hbb94e563),
	.w4(32'hbbaa1805),
	.w5(32'hbb8baf60),
	.w6(32'hbb25617e),
	.w7(32'hbbd110e1),
	.w8(32'h39289dac),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe69a71),
	.w1(32'hbbea9f7b),
	.w2(32'hbb7231ae),
	.w3(32'hbc1aea66),
	.w4(32'hbbad9d7e),
	.w5(32'h3c087dfd),
	.w6(32'hbb0a00b9),
	.w7(32'hba805c93),
	.w8(32'h3aae3556),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b701c),
	.w1(32'hbd02437c),
	.w2(32'hbc9ffaff),
	.w3(32'h3bce37e3),
	.w4(32'h3af66bb6),
	.w5(32'h3b005340),
	.w6(32'h3c0f0a63),
	.w7(32'h3ac4c919),
	.w8(32'h3bd74cd2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b494b),
	.w1(32'h3c3ad9d8),
	.w2(32'h3c494aee),
	.w3(32'h3c0606ff),
	.w4(32'h3c400a4c),
	.w5(32'h3a81d092),
	.w6(32'h3c3ebf66),
	.w7(32'h3c0b49b8),
	.w8(32'hbab87495),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95e7ac),
	.w1(32'h3c2f84f7),
	.w2(32'h3bc0994e),
	.w3(32'h3b8db01a),
	.w4(32'h3a7b70f6),
	.w5(32'h3af84388),
	.w6(32'hbb9670e6),
	.w7(32'hbb67dca1),
	.w8(32'hbc24ee24),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb336871),
	.w1(32'h3b8c4f4b),
	.w2(32'h3b07e50d),
	.w3(32'hb7b14828),
	.w4(32'h3bce95ee),
	.w5(32'hbb96fd01),
	.w6(32'h3c3156f4),
	.w7(32'hbba11b31),
	.w8(32'hbb955885),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb142ec),
	.w1(32'h3be32b88),
	.w2(32'h3bdad0b4),
	.w3(32'hbb7b30ac),
	.w4(32'h3a011d37),
	.w5(32'h3b48b2a4),
	.w6(32'h3acc7ac3),
	.w7(32'h3a020064),
	.w8(32'h3b06a823),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f99bb),
	.w1(32'h3b3c3713),
	.w2(32'hb98ebb22),
	.w3(32'hb8ce1555),
	.w4(32'h3b6a0b83),
	.w5(32'hbb9b64d5),
	.w6(32'h3ba72731),
	.w7(32'h3ba7eb49),
	.w8(32'hbc2b237b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48f664),
	.w1(32'h3c0a3936),
	.w2(32'h3bca2d8e),
	.w3(32'hbb18f065),
	.w4(32'hbb8c9e17),
	.w5(32'hba35a6d5),
	.w6(32'hbb42501f),
	.w7(32'hbc5c4ff4),
	.w8(32'hbb5f26a0),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aee15),
	.w1(32'hbb98316f),
	.w2(32'hbc1733f3),
	.w3(32'h3c0a6ec5),
	.w4(32'h3c1fe3d9),
	.w5(32'h3c3f6168),
	.w6(32'h3aeb0603),
	.w7(32'hbb0439f8),
	.w8(32'h3be21981),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1d163),
	.w1(32'hbccca9f2),
	.w2(32'hbbc1bc42),
	.w3(32'h3c8e115a),
	.w4(32'h3c810a05),
	.w5(32'h3b90bda1),
	.w6(32'h3b8041bd),
	.w7(32'h3be7b366),
	.w8(32'h3b6e1ede),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb85a07),
	.w1(32'h3c8086dc),
	.w2(32'h3b770e42),
	.w3(32'hbb62baa4),
	.w4(32'h3bddd9fe),
	.w5(32'hbb470702),
	.w6(32'hbb44dd55),
	.w7(32'h3c8716e5),
	.w8(32'h3887b206),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d7eed),
	.w1(32'h3d49fd58),
	.w2(32'h3c87aaa1),
	.w3(32'hbcf91a4b),
	.w4(32'hbc55230a),
	.w5(32'hbbb706e4),
	.w6(32'hbc6c4b3d),
	.w7(32'hbc1c6110),
	.w8(32'hbbc3447d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7366b),
	.w1(32'h390ea6fd),
	.w2(32'h3a631ed3),
	.w3(32'hbba1225f),
	.w4(32'hbc2b01e1),
	.w5(32'h3a54045c),
	.w6(32'hbc509b6b),
	.w7(32'hbbf891a2),
	.w8(32'hbb8316d6),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd37347),
	.w1(32'hbbebe418),
	.w2(32'h3ab3f66c),
	.w3(32'h3be0fe31),
	.w4(32'h3b4b3af0),
	.w5(32'hbbfd324d),
	.w6(32'h3b7b6646),
	.w7(32'h3b9f245a),
	.w8(32'hbba1a8cc),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d7c56),
	.w1(32'h3af69edc),
	.w2(32'h3bb63046),
	.w3(32'hbbd6e074),
	.w4(32'hbc0f50fe),
	.w5(32'hbc43590f),
	.w6(32'hbc088898),
	.w7(32'hbb50b1c0),
	.w8(32'h3a743e66),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69b20d),
	.w1(32'h3cad692d),
	.w2(32'h3c50d78b),
	.w3(32'hbc89e98c),
	.w4(32'hbc22e853),
	.w5(32'hba7f295b),
	.w6(32'hba01cea9),
	.w7(32'hbc0a14e8),
	.w8(32'h3b2a8096),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5369b3),
	.w1(32'h3bc52356),
	.w2(32'hb890a3e0),
	.w3(32'hbb07b08b),
	.w4(32'h3b87e931),
	.w5(32'hbc1ba19e),
	.w6(32'h3b45c095),
	.w7(32'h3b39a751),
	.w8(32'hbb80c147),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6915ef),
	.w1(32'h3ce218a1),
	.w2(32'h3c582fe0),
	.w3(32'hbb5cfa6d),
	.w4(32'hbb2ca748),
	.w5(32'h3a2c618b),
	.w6(32'hbb049ccb),
	.w7(32'hbbcaf19b),
	.w8(32'hb8f5e1ef),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b947cf2),
	.w1(32'h3bc2ed90),
	.w2(32'h3c0212c0),
	.w3(32'h3ba4414f),
	.w4(32'hbb2c0cc7),
	.w5(32'hbb850888),
	.w6(32'h3b6b0aff),
	.w7(32'hbbab5e0c),
	.w8(32'hbbea4b94),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a310c76),
	.w1(32'h3caada9b),
	.w2(32'hb9f01c48),
	.w3(32'hbbcab22c),
	.w4(32'hb99ec629),
	.w5(32'h3a8f43df),
	.w6(32'hbc068485),
	.w7(32'hbb7b6886),
	.w8(32'h3bc401c9),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc1d4e),
	.w1(32'hbc6ad2b2),
	.w2(32'hbc27056f),
	.w3(32'h3cae15be),
	.w4(32'h3c5eb1d3),
	.w5(32'h3a7bbc6c),
	.w6(32'h3bab179c),
	.w7(32'h3bbe21a6),
	.w8(32'hbaabae24),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba116214),
	.w1(32'h3c075fad),
	.w2(32'h3b64bd6d),
	.w3(32'h3b740305),
	.w4(32'h3c04c397),
	.w5(32'h3c3b5e9c),
	.w6(32'hbb884c21),
	.w7(32'hbb959bff),
	.w8(32'h3c08134d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc766498),
	.w1(32'hbce6d8ec),
	.w2(32'hbc8cca1b),
	.w3(32'h3cb56b2e),
	.w4(32'h3c20acb9),
	.w5(32'hbc97af88),
	.w6(32'h3c124822),
	.w7(32'h3b21e434),
	.w8(32'hbafe17e2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60a3af),
	.w1(32'h3d06f060),
	.w2(32'h3c848791),
	.w3(32'hbc988a43),
	.w4(32'hbc9499af),
	.w5(32'h3c013d2b),
	.w6(32'hba2641fd),
	.w7(32'hbbcba9f7),
	.w8(32'hbb3a0f54),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a919dc8),
	.w1(32'h3b63a803),
	.w2(32'hbaf9bd11),
	.w3(32'h3b7fa570),
	.w4(32'hbbb39c2f),
	.w5(32'h3c077ff4),
	.w6(32'hbb3623b3),
	.w7(32'hbbb980ce),
	.w8(32'h3bb87a86),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ad270),
	.w1(32'hbca2b0a0),
	.w2(32'hbc0b060e),
	.w3(32'h3c6a6ae6),
	.w4(32'h3c2561b8),
	.w5(32'h38d2221e),
	.w6(32'h3b7ecc38),
	.w7(32'h3bee42c1),
	.w8(32'hbbb33dd7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb735aaf),
	.w1(32'h3b0c531c),
	.w2(32'hbb41ce51),
	.w3(32'hbbb66c6d),
	.w4(32'hbbf38223),
	.w5(32'hbb11b91c),
	.w6(32'hbbda1d62),
	.w7(32'hbbf4ff56),
	.w8(32'hbbc1c38b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b321163),
	.w1(32'h3c501774),
	.w2(32'h3abb52d0),
	.w3(32'h3ba2c7ca),
	.w4(32'h3b85667f),
	.w5(32'hbb928c48),
	.w6(32'hbacc43f7),
	.w7(32'hbc01381c),
	.w8(32'hbba4433a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1564c),
	.w1(32'h3c2118c4),
	.w2(32'h3b48874d),
	.w3(32'hbc5d3511),
	.w4(32'hbc46b219),
	.w5(32'h3b224e74),
	.w6(32'hbb72f6f7),
	.w7(32'hbbab0db6),
	.w8(32'h3b068173),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb139195),
	.w1(32'h3adba5ff),
	.w2(32'h3a4a002a),
	.w3(32'h3a87c8c5),
	.w4(32'hbb8cc477),
	.w5(32'hbadccb91),
	.w6(32'h3c562288),
	.w7(32'h3b19861e),
	.w8(32'h3873a72c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1ddf9),
	.w1(32'h3c1ee16e),
	.w2(32'h3bbe3a56),
	.w3(32'hbb850fc0),
	.w4(32'h3b186809),
	.w5(32'h3b2951b6),
	.w6(32'h39ce44fa),
	.w7(32'h3a9a2f63),
	.w8(32'hbb4ab516),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d6014),
	.w1(32'hbb9bba46),
	.w2(32'hbb8966c5),
	.w3(32'h3b7e5768),
	.w4(32'h3bae7617),
	.w5(32'hb9d61d9a),
	.w6(32'hbc2557e3),
	.w7(32'hbb20637c),
	.w8(32'hbb0c7455),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20e48a),
	.w1(32'hbc1b5f26),
	.w2(32'hbc06e31a),
	.w3(32'hbc2a3e81),
	.w4(32'hbafee61e),
	.w5(32'h3807894c),
	.w6(32'hbc9075df),
	.w7(32'hbbc5156c),
	.w8(32'hbbda2e70),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c82e3),
	.w1(32'hb9f3762f),
	.w2(32'h3a2109cf),
	.w3(32'hbc9d0f7a),
	.w4(32'hbc88c0f4),
	.w5(32'hbc907e3d),
	.w6(32'hbcc28844),
	.w7(32'hbbfd037f),
	.w8(32'hbc5f4d9e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0b774),
	.w1(32'h3ccbb246),
	.w2(32'h3ba7617c),
	.w3(32'hbc96de3b),
	.w4(32'h3b220951),
	.w5(32'h3c2dc0c5),
	.w6(32'hbbfd6bb1),
	.w7(32'h3b35f855),
	.w8(32'h3b5dde44),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e4fe6),
	.w1(32'hbc01bb66),
	.w2(32'hbbea11c8),
	.w3(32'h3c4af8b3),
	.w4(32'h3c5299f3),
	.w5(32'h3b16e018),
	.w6(32'h3c05ed4c),
	.w7(32'h3ba29449),
	.w8(32'h3b8ed323),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d2821),
	.w1(32'h3b7e8a3d),
	.w2(32'h3bd9ec38),
	.w3(32'h3b77d800),
	.w4(32'h3bbc15df),
	.w5(32'hba4666c3),
	.w6(32'h3aa01beb),
	.w7(32'h3bbb2600),
	.w8(32'hbc38cb2e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab441e),
	.w1(32'h3b44aad2),
	.w2(32'h3bd38553),
	.w3(32'hbc02f1f9),
	.w4(32'hbb389b9c),
	.w5(32'h3c69e3a4),
	.w6(32'hbc245263),
	.w7(32'hbc1f081b),
	.w8(32'h3c16e267),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2274b5),
	.w1(32'hbd1e5b1b),
	.w2(32'hbcb54e9b),
	.w3(32'h3cf33e17),
	.w4(32'h3c59b05a),
	.w5(32'h3b80fe8e),
	.w6(32'h3c1d3eba),
	.w7(32'h3bd3f96a),
	.w8(32'h3b84bed0),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8065e4),
	.w1(32'h3c7de64d),
	.w2(32'hbb5086d6),
	.w3(32'hbc1566f2),
	.w4(32'hbc852cca),
	.w5(32'hbb6dbb37),
	.w6(32'hbc7dd1ed),
	.w7(32'hbb267184),
	.w8(32'hbb405255),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95be7d0),
	.w1(32'hbb259a07),
	.w2(32'hbb940c75),
	.w3(32'hbb49e41f),
	.w4(32'hbb841256),
	.w5(32'h394bd000),
	.w6(32'hbb823cfe),
	.w7(32'hbb99a243),
	.w8(32'hb94fe698),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dacc8b),
	.w1(32'hbaff00f8),
	.w2(32'hbbcfbdd4),
	.w3(32'hbb19dc65),
	.w4(32'hbb4a1c0b),
	.w5(32'h3ba4f076),
	.w6(32'hbafc2c1e),
	.w7(32'hbb25b697),
	.w8(32'h3b1db8cd),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba956c5),
	.w1(32'h3bbb7dc1),
	.w2(32'hbb55110a),
	.w3(32'h3bfbe817),
	.w4(32'h3affe135),
	.w5(32'hbba2f633),
	.w6(32'h3bdbcb6a),
	.w7(32'hbac31bb6),
	.w8(32'hbbfc8d28),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe4449),
	.w1(32'h3a20ec5c),
	.w2(32'h3b027955),
	.w3(32'hbb751a3d),
	.w4(32'hbbb45818),
	.w5(32'h39940c8b),
	.w6(32'hbbc1d9f8),
	.w7(32'hbb01dc21),
	.w8(32'h3a450fe3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b9fc4),
	.w1(32'hbc33ec91),
	.w2(32'hbc36b3fe),
	.w3(32'hbc88b765),
	.w4(32'hbc41f9d9),
	.w5(32'hbc0f8b1d),
	.w6(32'hbc80a814),
	.w7(32'hbc16c66c),
	.w8(32'hbc3371f1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7e530),
	.w1(32'hbba6878e),
	.w2(32'hb92625d0),
	.w3(32'hbbf72337),
	.w4(32'hbb9b1dfe),
	.w5(32'h37e06d3d),
	.w6(32'hbc223123),
	.w7(32'hbb45a831),
	.w8(32'hba9107c8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf523e3),
	.w1(32'hbbb50b5c),
	.w2(32'hbbc7d702),
	.w3(32'h3b2bb2b4),
	.w4(32'hbb2dadec),
	.w5(32'hbada38be),
	.w6(32'h3ad3537a),
	.w7(32'hba6f803e),
	.w8(32'hbaee1d7c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2a38e),
	.w1(32'hbbaf9889),
	.w2(32'hbacfe360),
	.w3(32'hbbb4edef),
	.w4(32'hbb973e48),
	.w5(32'hba947124),
	.w6(32'hbba93a87),
	.w7(32'hbb1832c8),
	.w8(32'h3a7fe72a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51e9a3),
	.w1(32'hba36de32),
	.w2(32'hbb803a2f),
	.w3(32'hbb384204),
	.w4(32'hbc08e723),
	.w5(32'h39cbf68e),
	.w6(32'hba5f963c),
	.w7(32'hbc1b363a),
	.w8(32'hb9fe1636),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c16501),
	.w1(32'hbb14709b),
	.w2(32'hbb9da8eb),
	.w3(32'hbb249f85),
	.w4(32'hbb5da2b0),
	.w5(32'hbb9a6b56),
	.w6(32'hbb5ae409),
	.w7(32'hbb8f6120),
	.w8(32'hbb26959c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32fce2),
	.w1(32'hbb5f1545),
	.w2(32'hbbbfd947),
	.w3(32'hbbb38de1),
	.w4(32'hbbeb4822),
	.w5(32'h3b98891b),
	.w6(32'hbba0843d),
	.w7(32'hbbee9747),
	.w8(32'h3b503387),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ce210),
	.w1(32'h3b01f7ac),
	.w2(32'h39fa7b61),
	.w3(32'h3b3c9997),
	.w4(32'h3b870f2f),
	.w5(32'hbb9f8d2c),
	.w6(32'hba14452e),
	.w7(32'h3a9f4064),
	.w8(32'hbbaa0083),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ed22f),
	.w1(32'hbb53c024),
	.w2(32'hbb95aa18),
	.w3(32'hbb8beac4),
	.w4(32'hbb30670e),
	.w5(32'h3b378c78),
	.w6(32'hbb54840e),
	.w7(32'hbb683db8),
	.w8(32'h3abe4982),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba806b9c),
	.w1(32'h3a932c6e),
	.w2(32'h3b1d5f2a),
	.w3(32'h3adc20ae),
	.w4(32'h3ba084e0),
	.w5(32'h3a0eef64),
	.w6(32'h3b2b16a9),
	.w7(32'h3b8b2ba3),
	.w8(32'hbac30f22),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba958be1),
	.w1(32'hbae18551),
	.w2(32'h3ab005e3),
	.w3(32'h3b1cfe09),
	.w4(32'h3ba5d579),
	.w5(32'hbb69636b),
	.w6(32'h3a28d430),
	.w7(32'h3b7f189a),
	.w8(32'hba9b8468),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe76b6),
	.w1(32'hbba8bb83),
	.w2(32'hbb3efc4a),
	.w3(32'hbb80c6ce),
	.w4(32'hbb9d3936),
	.w5(32'hbab6fc87),
	.w6(32'hbac53294),
	.w7(32'hbad81a1a),
	.w8(32'hbb085bf5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96e99d),
	.w1(32'h3797300a),
	.w2(32'hbb2c3eab),
	.w3(32'hbb8a1d11),
	.w4(32'hbbf2a74e),
	.w5(32'hbb58113c),
	.w6(32'hbb2d6fde),
	.w7(32'hbbe2207b),
	.w8(32'hbb8694d6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90b108),
	.w1(32'hbaa35cb0),
	.w2(32'h3aa92de1),
	.w3(32'hbb9f9e5d),
	.w4(32'hbacf160a),
	.w5(32'h3ba20720),
	.w6(32'hbb738d80),
	.w7(32'h39eb2cf7),
	.w8(32'h3b88672a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8b53e),
	.w1(32'h3b9a5e0a),
	.w2(32'h3b6f1584),
	.w3(32'h3b865efd),
	.w4(32'h3b95f94d),
	.w5(32'hbaa9c9aa),
	.w6(32'h3b526dea),
	.w7(32'h3b67986a),
	.w8(32'h3986b741),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28a806),
	.w1(32'hbb1a9a76),
	.w2(32'hbaace3e6),
	.w3(32'hbb557d7d),
	.w4(32'hbbb7bf46),
	.w5(32'hbb4687ee),
	.w6(32'hba30fc39),
	.w7(32'hbb606c3b),
	.w8(32'hbb65f656),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0b3a2),
	.w1(32'hbbc92a5b),
	.w2(32'hbb822875),
	.w3(32'hbbc596e1),
	.w4(32'hbb572ffd),
	.w5(32'hbb7d43fa),
	.w6(32'hbbeedad2),
	.w7(32'hbb0b1ed1),
	.w8(32'hbb4c897a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08ba27),
	.w1(32'h395cd552),
	.w2(32'hbb4c8a58),
	.w3(32'hbb57338d),
	.w4(32'hbbe936d5),
	.w5(32'hbaa5ce5c),
	.w6(32'hbb9b9a06),
	.w7(32'hbbd99c44),
	.w8(32'h38efa5ee),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee2516),
	.w1(32'h3b086eaf),
	.w2(32'h3b09147a),
	.w3(32'h3a26d5ce),
	.w4(32'h3aa893fe),
	.w5(32'h3aae7c80),
	.w6(32'h3a4e1138),
	.w7(32'h3b4bf292),
	.w8(32'h3aca3b8a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49efbf),
	.w1(32'hba069fac),
	.w2(32'h3b2a1be3),
	.w3(32'h3a6ce243),
	.w4(32'h3b49ddd0),
	.w5(32'h3b6dad5d),
	.w6(32'h3a9bc6b4),
	.w7(32'h3aabfbcd),
	.w8(32'hb9d928e1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2effb),
	.w1(32'hba1c646c),
	.w2(32'h3b267fa9),
	.w3(32'h3b67ff12),
	.w4(32'hbacca27a),
	.w5(32'hbb63471a),
	.w6(32'hbb225c64),
	.w7(32'h399bf4fb),
	.w8(32'h3a96a455),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a4b6a2),
	.w1(32'hbaeb8df4),
	.w2(32'hbb0a8601),
	.w3(32'hbb587019),
	.w4(32'h3b72d4dd),
	.w5(32'hbb0e9105),
	.w6(32'hbbb1bd63),
	.w7(32'h3a058655),
	.w8(32'hbb9e06b2),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62cb2b),
	.w1(32'hbb1ecfb2),
	.w2(32'hba9a915d),
	.w3(32'hb9085eef),
	.w4(32'hbb59d162),
	.w5(32'hbabb3365),
	.w6(32'hbb7f9549),
	.w7(32'hbb6918db),
	.w8(32'hba58f932),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe551c3),
	.w1(32'hbc2dd4ba),
	.w2(32'hbbd79856),
	.w3(32'hbc0a4a49),
	.w4(32'hbbba3907),
	.w5(32'h390a6a87),
	.w6(32'hbc08d8f6),
	.w7(32'hbb986189),
	.w8(32'h3a3b2bdb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e8c545),
	.w1(32'hbb2c1c5e),
	.w2(32'hbb9205bd),
	.w3(32'hba4f6c9e),
	.w4(32'hbaed64a1),
	.w5(32'hbac220fe),
	.w6(32'hbb6cdb33),
	.w7(32'hbb451b0d),
	.w8(32'hb9dfe921),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78fb8a),
	.w1(32'hba8bb91e),
	.w2(32'hb9f2e8cc),
	.w3(32'hbbd3b7bd),
	.w4(32'hbb29a394),
	.w5(32'h3b9ec22f),
	.w6(32'hbab10070),
	.w7(32'hbb022276),
	.w8(32'hbaa81865),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule