module layer_10_featuremap_271(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc379fc),
	.w1(32'hbc2f87f6),
	.w2(32'hbbfb6aed),
	.w3(32'h3a863c25),
	.w4(32'h3b19ccb5),
	.w5(32'hbbcbea52),
	.w6(32'hbb55d5f5),
	.w7(32'hbba6b954),
	.w8(32'hbbf696e6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac7759),
	.w1(32'hbb218750),
	.w2(32'hbb9e6207),
	.w3(32'h3b3c7dcf),
	.w4(32'hbb784d65),
	.w5(32'h3c0f9e8b),
	.w6(32'h3ac8c9e7),
	.w7(32'hbb534175),
	.w8(32'h3bc048d8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe58db),
	.w1(32'hbc977182),
	.w2(32'hbc2f36f7),
	.w3(32'h3ba4236e),
	.w4(32'h3c183c78),
	.w5(32'hbb2b5407),
	.w6(32'h3c27bebe),
	.w7(32'h3a965ed0),
	.w8(32'h3b2eb7e2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dd533),
	.w1(32'h3bba5965),
	.w2(32'h3c058db4),
	.w3(32'hbb4f6b2a),
	.w4(32'h3ae2013a),
	.w5(32'hbb6ac711),
	.w6(32'hb99eda0f),
	.w7(32'h3a6aea3a),
	.w8(32'hbc4425fa),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b856f),
	.w1(32'hbbacfd96),
	.w2(32'h39e8fbed),
	.w3(32'h3b4652c3),
	.w4(32'hba280800),
	.w5(32'hb9d6d3a4),
	.w6(32'hbc41d663),
	.w7(32'hbb62c45f),
	.w8(32'h3b3fd612),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09d50d),
	.w1(32'h3b319937),
	.w2(32'h3b758fd4),
	.w3(32'h3991a65d),
	.w4(32'hbaac43fd),
	.w5(32'hbbe18d00),
	.w6(32'hb7e0e0b9),
	.w7(32'h3a608c00),
	.w8(32'hbbae7e5d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81ce7d),
	.w1(32'hba9b6bc0),
	.w2(32'h3b02e3d1),
	.w3(32'hbba31b4a),
	.w4(32'hba890c13),
	.w5(32'hba62b4ef),
	.w6(32'hba3bd714),
	.w7(32'hba4cc428),
	.w8(32'h3b5b76f7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa78d54),
	.w1(32'h3b875252),
	.w2(32'h3ba921c1),
	.w3(32'hbb6c0d97),
	.w4(32'hbb5f1104),
	.w5(32'h3b615960),
	.w6(32'hbb4aa10f),
	.w7(32'hbb1ace19),
	.w8(32'h3bec9c40),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5f7aa),
	.w1(32'h3b0e46e9),
	.w2(32'h3a7abc1a),
	.w3(32'h3b216f13),
	.w4(32'h3b8dc674),
	.w5(32'hbb130d2b),
	.w6(32'h3b6f2954),
	.w7(32'h3b964e9f),
	.w8(32'h3aa94e7c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f9183),
	.w1(32'h3b30e9be),
	.w2(32'h3b842f8f),
	.w3(32'hba9066ca),
	.w4(32'hbb0a7371),
	.w5(32'h3900135a),
	.w6(32'hbb742c18),
	.w7(32'h3973d1e0),
	.w8(32'hbb3a1856),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb098d1c),
	.w1(32'hbb407a99),
	.w2(32'h3b2043af),
	.w3(32'h3ba42d0a),
	.w4(32'h3bb51206),
	.w5(32'h3be4c267),
	.w6(32'hbb1027a2),
	.w7(32'h3a1a5b36),
	.w8(32'h3b049897),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb648751),
	.w1(32'hbc4d18ab),
	.w2(32'hbba354df),
	.w3(32'h3b995249),
	.w4(32'h3b9013d9),
	.w5(32'h3c784a78),
	.w6(32'h3c47eb28),
	.w7(32'h3bb2821a),
	.w8(32'hba22a3c4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf2857),
	.w1(32'hbbe86021),
	.w2(32'hbc103696),
	.w3(32'h3cb3d736),
	.w4(32'h3c8112b8),
	.w5(32'hba39f364),
	.w6(32'hbb8a1761),
	.w7(32'hbc073850),
	.w8(32'hbba71b08),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff5774),
	.w1(32'hbbeee1b9),
	.w2(32'h3a8a5dd2),
	.w3(32'h3b42fa6c),
	.w4(32'h3b5137ad),
	.w5(32'h3aca6260),
	.w6(32'hbb56b93a),
	.w7(32'h36eecae1),
	.w8(32'h3a7d876b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b391302),
	.w1(32'h3b2bd29d),
	.w2(32'hba3e9e73),
	.w3(32'hbac347c6),
	.w4(32'h3a9077cd),
	.w5(32'h398b37ce),
	.w6(32'hbb0afb41),
	.w7(32'hbb967a20),
	.w8(32'hbb13cdff),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94bd04),
	.w1(32'hbab8143d),
	.w2(32'h3b13f566),
	.w3(32'h3ba1b536),
	.w4(32'hbb0ec15f),
	.w5(32'h3b6cb978),
	.w6(32'h39258d6f),
	.w7(32'h3a86179a),
	.w8(32'hba9b8d38),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a11096),
	.w1(32'h3a3e9dfb),
	.w2(32'h3a6f69cb),
	.w3(32'h3c37b65b),
	.w4(32'h3ba8b01a),
	.w5(32'h3c4df3e1),
	.w6(32'h3b7c3da7),
	.w7(32'h3ad5a701),
	.w8(32'hbac8f1f4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc537ab5),
	.w1(32'hbc60a522),
	.w2(32'hbc27583f),
	.w3(32'h3c8e64bc),
	.w4(32'h3c660267),
	.w5(32'hbbb92b88),
	.w6(32'hbc0734ec),
	.w7(32'hbc186c6c),
	.w8(32'hbbdaa6ea),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefb473),
	.w1(32'hb9f1e4e5),
	.w2(32'hbae58ffa),
	.w3(32'hbb8a3fa2),
	.w4(32'hbbab8e46),
	.w5(32'h399f22a6),
	.w6(32'hbbcea2cd),
	.w7(32'hbb97db80),
	.w8(32'hbbc5a7d5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43d8af),
	.w1(32'hbc0b6a04),
	.w2(32'hbc485e55),
	.w3(32'h3be56125),
	.w4(32'h3b66d01a),
	.w5(32'hba928d44),
	.w6(32'hbbffea3f),
	.w7(32'hba9b6b18),
	.w8(32'hbb184e61),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b054a14),
	.w1(32'h387a764b),
	.w2(32'h3afdd0b2),
	.w3(32'h3c471b82),
	.w4(32'h3b41f69d),
	.w5(32'hbc7f5114),
	.w6(32'h3b8877d0),
	.w7(32'h3b38f99d),
	.w8(32'h3b7a8914),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53bfaa),
	.w1(32'h3ca39066),
	.w2(32'h3c828b8b),
	.w3(32'hbca0bd0a),
	.w4(32'hbc7219f5),
	.w5(32'h3a0f705e),
	.w6(32'h3b92049f),
	.w7(32'h3bc38cda),
	.w8(32'h3b0b7c4e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc506858),
	.w1(32'hbc5379f3),
	.w2(32'hbc14767e),
	.w3(32'h3b8fce03),
	.w4(32'h3ba0a954),
	.w5(32'hbb9ad531),
	.w6(32'h3ad94e74),
	.w7(32'hbbb31115),
	.w8(32'hbc93e040),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35ae79),
	.w1(32'hbb9cc43e),
	.w2(32'hba971ccd),
	.w3(32'hbaec093d),
	.w4(32'h3ae70d57),
	.w5(32'h3bc80830),
	.w6(32'hbc5d77c3),
	.w7(32'h3af6bb2a),
	.w8(32'hbb96b67d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a6147),
	.w1(32'hbba15d3c),
	.w2(32'hbc144d2d),
	.w3(32'h3c1bcf50),
	.w4(32'h3c24d6f6),
	.w5(32'hbbf91446),
	.w6(32'h3afd61cf),
	.w7(32'hbb972260),
	.w8(32'hbb882d45),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44e642),
	.w1(32'h3b5b7253),
	.w2(32'h3b113432),
	.w3(32'h3ae19d89),
	.w4(32'hbab6a46b),
	.w5(32'hbc00e099),
	.w6(32'h3bb6d32b),
	.w7(32'h3aa90a4b),
	.w8(32'h38ce071d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e00f1),
	.w1(32'h3b7abb13),
	.w2(32'hbaec2464),
	.w3(32'hbc2b388d),
	.w4(32'hbbcea1b5),
	.w5(32'h3ad9b7e9),
	.w6(32'h3b8f6b98),
	.w7(32'h3afd406e),
	.w8(32'h3b2aa7e2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f5853),
	.w1(32'h3a13b86f),
	.w2(32'hb9845d95),
	.w3(32'h3b10e487),
	.w4(32'hb9cd8c90),
	.w5(32'h39fc0e7f),
	.w6(32'h3b678dd6),
	.w7(32'h3b93419f),
	.w8(32'h3a2aaa55),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a5d62),
	.w1(32'hbbdb8e7b),
	.w2(32'hbc02c07a),
	.w3(32'h3bc7024c),
	.w4(32'h3b9eacd9),
	.w5(32'h3b3485fd),
	.w6(32'h3af23ed2),
	.w7(32'hb9d6c321),
	.w8(32'h3b827aff),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f3178e),
	.w1(32'hbc3b5882),
	.w2(32'hbc1de07d),
	.w3(32'h3bd49394),
	.w4(32'hba60f50b),
	.w5(32'hbb16a444),
	.w6(32'hbb1e2678),
	.w7(32'hb9029f71),
	.w8(32'hbc2fd5f7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc385c76),
	.w1(32'hbc448956),
	.w2(32'hbb9cf14f),
	.w3(32'hbbd4243e),
	.w4(32'hbba988d6),
	.w5(32'h3c376d72),
	.w6(32'hbbdba2c7),
	.w7(32'hbc05875a),
	.w8(32'h3bede531),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc246dca),
	.w1(32'hbc5e11b0),
	.w2(32'hbbea34fc),
	.w3(32'h3c26c163),
	.w4(32'h3be26368),
	.w5(32'h3ac17c01),
	.w6(32'h3c5278b0),
	.w7(32'hbb3ce31a),
	.w8(32'hbb05ef24),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9158b8),
	.w1(32'h3ad22623),
	.w2(32'h3c099dd4),
	.w3(32'h3af32b17),
	.w4(32'hbb7c3def),
	.w5(32'h3c9147fd),
	.w6(32'h3ab57905),
	.w7(32'hbb9f6ad8),
	.w8(32'hbb03fde9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27ee20),
	.w1(32'hbca2057c),
	.w2(32'hbc4d69aa),
	.w3(32'h3cee3744),
	.w4(32'h3c13ca8d),
	.w5(32'h3b821f3b),
	.w6(32'hbbd6a38e),
	.w7(32'hbc2529ad),
	.w8(32'hbb6560b9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cdb2b1),
	.w1(32'hbbebf6ba),
	.w2(32'hbbfed1a1),
	.w3(32'h3beeaa76),
	.w4(32'h37f596e1),
	.w5(32'h3c3ca753),
	.w6(32'hb9f1ac4f),
	.w7(32'hbb52f93a),
	.w8(32'hbba1d930),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e775b),
	.w1(32'hbc79b2b7),
	.w2(32'hbc360656),
	.w3(32'h3c9b3191),
	.w4(32'h3b86ff93),
	.w5(32'hbbc130e7),
	.w6(32'hbc3b54c8),
	.w7(32'hbbe13a59),
	.w8(32'hbc0e6708),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30f1b1),
	.w1(32'hbb6716f6),
	.w2(32'hbb8e97a7),
	.w3(32'hbbd83e80),
	.w4(32'hbb621cf0),
	.w5(32'hbb4e1ee3),
	.w6(32'hbbe74e03),
	.w7(32'hbc25ce2f),
	.w8(32'h3b798755),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a9954),
	.w1(32'h3b0b4a2a),
	.w2(32'h3b31e0eb),
	.w3(32'hba9f28fe),
	.w4(32'hbbd2b2c3),
	.w5(32'h3b8a286e),
	.w6(32'h3bd4426f),
	.w7(32'h3bb369f7),
	.w8(32'hbc2bdf46),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5637c),
	.w1(32'hbacc5941),
	.w2(32'hbbe6c1a1),
	.w3(32'h3c04563b),
	.w4(32'h3af73aaf),
	.w5(32'hbcb83e27),
	.w6(32'hbbe464dd),
	.w7(32'hbb399d02),
	.w8(32'h3bb7624f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a82ce),
	.w1(32'h3c9e6eca),
	.w2(32'h3c8972d4),
	.w3(32'hbcb2509c),
	.w4(32'hbca37c1d),
	.w5(32'h3bed8f43),
	.w6(32'h3b11c287),
	.w7(32'h3b8803d6),
	.w8(32'h3b62c9e4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb21e19),
	.w1(32'hbc17d1e3),
	.w2(32'hbbbd7871),
	.w3(32'h3c0426e6),
	.w4(32'h3c149015),
	.w5(32'hbbebb9ee),
	.w6(32'hbac427b3),
	.w7(32'hbb491d40),
	.w8(32'hbb26d538),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13a128),
	.w1(32'h3b74b122),
	.w2(32'h3b5c0e31),
	.w3(32'hba7904fb),
	.w4(32'hbb5e8ef8),
	.w5(32'h3bf39494),
	.w6(32'h3b77d109),
	.w7(32'h38ee0760),
	.w8(32'hbaaf64fe),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d3c85),
	.w1(32'hbc3fb3ad),
	.w2(32'hbc40a7e1),
	.w3(32'h3c15e6a9),
	.w4(32'h3b363eac),
	.w5(32'h3c04d318),
	.w6(32'hbbe8072c),
	.w7(32'hbb9fed03),
	.w8(32'hbc2542cc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46705d),
	.w1(32'hbc92d23e),
	.w2(32'hbc9a721d),
	.w3(32'h3c86ab2a),
	.w4(32'h3bd8744b),
	.w5(32'hbba3239d),
	.w6(32'hbc50c737),
	.w7(32'hbc516657),
	.w8(32'h3b040db4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40f842),
	.w1(32'h3c4b6e94),
	.w2(32'h3c124e0b),
	.w3(32'hbbcd9170),
	.w4(32'hbbfd58b1),
	.w5(32'hbc141482),
	.w6(32'h3aa83e35),
	.w7(32'h3bba4c47),
	.w8(32'hbb07b12f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2ddf1),
	.w1(32'hb9a844d2),
	.w2(32'hbadc4ca6),
	.w3(32'hbc34a21d),
	.w4(32'hbbaf317a),
	.w5(32'hbbecac38),
	.w6(32'h39be81aa),
	.w7(32'hbabebd59),
	.w8(32'hbb82bf06),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29d349),
	.w1(32'h399d7aec),
	.w2(32'hba147441),
	.w3(32'hbc2780e1),
	.w4(32'hbc071382),
	.w5(32'hbc1d447b),
	.w6(32'hbaa2e6db),
	.w7(32'hbbac8ff1),
	.w8(32'hbb006d6a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58c4b5),
	.w1(32'h3c043d3a),
	.w2(32'h3bafb0da),
	.w3(32'hbc97f253),
	.w4(32'hbc140830),
	.w5(32'h3bbaacc7),
	.w6(32'hbbc8ac93),
	.w7(32'hbbbcebf8),
	.w8(32'hbc64c150),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc583aa1),
	.w1(32'hbc6cef78),
	.w2(32'hbc47688b),
	.w3(32'h3c5d029c),
	.w4(32'h3c49dd79),
	.w5(32'hbc5218a0),
	.w6(32'hbbba79e0),
	.w7(32'hbc20f5c5),
	.w8(32'h3b8fa0cd),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d0b2f),
	.w1(32'h3c6c682b),
	.w2(32'h3c30f470),
	.w3(32'hbc6f4d6e),
	.w4(32'hbc621aca),
	.w5(32'hba9056cf),
	.w6(32'h3bed5464),
	.w7(32'h3b7784de),
	.w8(32'hbadd09e3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b301c0d),
	.w1(32'hbbec9c5a),
	.w2(32'hbb357e01),
	.w3(32'hb8f89542),
	.w4(32'hbc210c7e),
	.w5(32'h3b12fe6c),
	.w6(32'hbb9c6813),
	.w7(32'h3acc5975),
	.w8(32'hbb93080c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb592280),
	.w1(32'hbb849967),
	.w2(32'hbbbef7c9),
	.w3(32'h3b89b4f3),
	.w4(32'hbbb6c648),
	.w5(32'h3c0b316e),
	.w6(32'hbb69737f),
	.w7(32'hbbaea75c),
	.w8(32'hbaf77fa0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba11afe),
	.w1(32'hbc104230),
	.w2(32'hbae9e2b8),
	.w3(32'h3c0aa9f1),
	.w4(32'h3bff7dde),
	.w5(32'h3a8b5d33),
	.w6(32'hb93e9a07),
	.w7(32'hbb3297de),
	.w8(32'h3c1a5294),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29255e),
	.w1(32'hbbf26464),
	.w2(32'hbc421088),
	.w3(32'h3bbc492a),
	.w4(32'h3c239b47),
	.w5(32'h3bb40887),
	.w6(32'h39d2e26d),
	.w7(32'hbc0a6798),
	.w8(32'hb9fedf7c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1ca59),
	.w1(32'hbbdd6522),
	.w2(32'hbc0f78a7),
	.w3(32'h3c5feac9),
	.w4(32'h3bf81838),
	.w5(32'h3c25d719),
	.w6(32'hba7d8b59),
	.w7(32'hb9d6a3a1),
	.w8(32'hbac07fb5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a129430),
	.w1(32'hbb796e6c),
	.w2(32'hbbe8aafa),
	.w3(32'h3c729d1c),
	.w4(32'h3b8da035),
	.w5(32'h3b67e53c),
	.w6(32'h3b886729),
	.w7(32'h3b180c68),
	.w8(32'h3b53f842),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3613e),
	.w1(32'hbb3197cf),
	.w2(32'hbb8595a0),
	.w3(32'h39d8a627),
	.w4(32'h3b0a63eb),
	.w5(32'h3acf5a69),
	.w6(32'h3a876269),
	.w7(32'hba52059c),
	.w8(32'h3c52014d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20bc5a),
	.w1(32'hbbb7936b),
	.w2(32'hbbb2062d),
	.w3(32'h3c7520a2),
	.w4(32'h3b03f74e),
	.w5(32'hbc2ef44c),
	.w6(32'h3aff5c97),
	.w7(32'hbb184dc6),
	.w8(32'h3b030df4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf70217),
	.w1(32'h3bdbf13d),
	.w2(32'h3bd462e7),
	.w3(32'hbc183b6e),
	.w4(32'hbbd81753),
	.w5(32'hbc671011),
	.w6(32'h3bd7c68f),
	.w7(32'h3b99419b),
	.w8(32'h3b677e26),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e5bf5),
	.w1(32'h3cca33f3),
	.w2(32'h3c721b1e),
	.w3(32'hbcd41199),
	.w4(32'hbc8fdb78),
	.w5(32'hbb311edb),
	.w6(32'h3c65dfc9),
	.w7(32'h3bdfcf8c),
	.w8(32'hbb1809f0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de4571),
	.w1(32'hbb220baf),
	.w2(32'hbbcc4468),
	.w3(32'hbb3d769a),
	.w4(32'h3a534f84),
	.w5(32'hbbcd862a),
	.w6(32'hbc125d61),
	.w7(32'hbbe2fd51),
	.w8(32'hbb8063de),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba025633),
	.w1(32'h3bf2f090),
	.w2(32'h3ba81d4c),
	.w3(32'h3a81e453),
	.w4(32'h3aa49898),
	.w5(32'hbb49d758),
	.w6(32'h3b7a0ac9),
	.w7(32'h3b0bfce4),
	.w8(32'hbb82d448),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67cd2e),
	.w1(32'hbb8bc00b),
	.w2(32'h3aad0fbd),
	.w3(32'h3ba5ca4c),
	.w4(32'h3af77202),
	.w5(32'h374ef538),
	.w6(32'h3b6ea68c),
	.w7(32'h3ba799b0),
	.w8(32'hbad9dca1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cc5ae),
	.w1(32'hbbddf972),
	.w2(32'hbbd63a84),
	.w3(32'h3befb96e),
	.w4(32'h3a2bb40b),
	.w5(32'h3b0d7531),
	.w6(32'hbb7c734c),
	.w7(32'hbbd5d89f),
	.w8(32'hbb81bad5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf47d2),
	.w1(32'hbb92fe96),
	.w2(32'hbb1c76ae),
	.w3(32'h3c1f7c79),
	.w4(32'h3b9e0989),
	.w5(32'h3b6c4508),
	.w6(32'h3a834042),
	.w7(32'h3b220a50),
	.w8(32'hba727b54),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa72176),
	.w1(32'hbbcb6a14),
	.w2(32'hbaed4831),
	.w3(32'h3c8c543c),
	.w4(32'h3c36b25b),
	.w5(32'h3afdeb5f),
	.w6(32'hba4ed59a),
	.w7(32'hbb196ee4),
	.w8(32'h3ba97185),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb0361),
	.w1(32'hbb3ad9de),
	.w2(32'h3bc0c363),
	.w3(32'h39e5ef0e),
	.w4(32'h3a75e624),
	.w5(32'hbb46d9cf),
	.w6(32'hbaaf0bdc),
	.w7(32'h3a31d694),
	.w8(32'h3bc12c7a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3daa17),
	.w1(32'h3af46722),
	.w2(32'hbb16a712),
	.w3(32'hbbb32b0d),
	.w4(32'h3b01c52f),
	.w5(32'h3bcd2d9a),
	.w6(32'hbb527aa2),
	.w7(32'hbb516069),
	.w8(32'hbb0721c2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba3758),
	.w1(32'hbc4acc56),
	.w2(32'hbbfa8015),
	.w3(32'h3c4c76e8),
	.w4(32'h3c074bcc),
	.w5(32'h3c079bfe),
	.w6(32'hbb0f1dfc),
	.w7(32'h3b7f6f11),
	.w8(32'hbbc0cb1d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29d5bd),
	.w1(32'hbca39d03),
	.w2(32'hbc909020),
	.w3(32'h3cc3dec2),
	.w4(32'h3c171571),
	.w5(32'hbb423ace),
	.w6(32'hbc24c394),
	.w7(32'hbc3d9149),
	.w8(32'hb9e4de85),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a043e76),
	.w1(32'hb7e42998),
	.w2(32'hbad3982b),
	.w3(32'hb9239ec4),
	.w4(32'hbb00ed07),
	.w5(32'hbb807c3c),
	.w6(32'h3a8ef659),
	.w7(32'hb91c5794),
	.w8(32'hbb807fed),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb503727),
	.w1(32'hbc0973be),
	.w2(32'hba43fe5e),
	.w3(32'h3bfc26c4),
	.w4(32'hbb6dc040),
	.w5(32'h3ba1e708),
	.w6(32'hbb7da799),
	.w7(32'hbc2ddafb),
	.w8(32'hbbfbc7a0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1daa1f),
	.w1(32'hbbe0bedd),
	.w2(32'hbb691850),
	.w3(32'h3b3123c6),
	.w4(32'h3bcce467),
	.w5(32'hb9ab255c),
	.w6(32'hbb983af5),
	.w7(32'hbbb714ca),
	.w8(32'hbb6d54a4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c822c),
	.w1(32'hbc313561),
	.w2(32'hbc582d82),
	.w3(32'h3c819b73),
	.w4(32'h3b7fd2bb),
	.w5(32'h3bdc0704),
	.w6(32'hbbe8b366),
	.w7(32'hbc66bfda),
	.w8(32'h3b2a8f31),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39a613),
	.w1(32'hbbcd28db),
	.w2(32'hb98c7988),
	.w3(32'h3be4536d),
	.w4(32'h3b042c92),
	.w5(32'h3cbdb439),
	.w6(32'hbadafb66),
	.w7(32'hbb1cd068),
	.w8(32'hbaf5cae2),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f8976),
	.w1(32'hbca38911),
	.w2(32'hbc575f59),
	.w3(32'h3cf368bc),
	.w4(32'h3caef587),
	.w5(32'h3a9ff0a8),
	.w6(32'hba792a14),
	.w7(32'hbbecfa6b),
	.w8(32'h3aaadd20),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe62552),
	.w1(32'hbc261379),
	.w2(32'hb881cf2a),
	.w3(32'h3b969df5),
	.w4(32'h3ba6a197),
	.w5(32'h3bc2f9fc),
	.w6(32'hb9751e3f),
	.w7(32'hbbb9cd48),
	.w8(32'hbb086cd7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36edcb01),
	.w1(32'hbba67a46),
	.w2(32'hbaeaab50),
	.w3(32'h3c43f6e0),
	.w4(32'h3b04cc7b),
	.w5(32'hbbe759a9),
	.w6(32'hbb69ff8a),
	.w7(32'hbb5a95ff),
	.w8(32'hbbae746c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9ea79),
	.w1(32'h3a8ffe7f),
	.w2(32'hbae1fae8),
	.w3(32'hbc336bc9),
	.w4(32'hbafb83ec),
	.w5(32'h3b8b1687),
	.w6(32'h3b6eafc2),
	.w7(32'hbac2dd5f),
	.w8(32'h3b3599c9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22375b),
	.w1(32'h3b366c0d),
	.w2(32'h3b943fa0),
	.w3(32'h3c026e75),
	.w4(32'h3b7738b6),
	.w5(32'hbbb25a46),
	.w6(32'h3adb06d8),
	.w7(32'h3aa9c9ed),
	.w8(32'h3bdd6cd5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f39ed),
	.w1(32'h3c0dfa6d),
	.w2(32'h3bb6f054),
	.w3(32'hbc236fda),
	.w4(32'hbc26754c),
	.w5(32'h3c277f4e),
	.w6(32'h3c1e5ebb),
	.w7(32'h3a77a66c),
	.w8(32'hbbc13795),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc622c6f),
	.w1(32'hbc867bc4),
	.w2(32'hbc46b815),
	.w3(32'h3c909398),
	.w4(32'h3c1bad24),
	.w5(32'h3b8b98f2),
	.w6(32'hbc1ba2f9),
	.w7(32'hbc4f8d57),
	.w8(32'hbabd1951),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43c596),
	.w1(32'hbbb6cb51),
	.w2(32'hba4cbfcb),
	.w3(32'h3c0f766a),
	.w4(32'h3c1adade),
	.w5(32'hbc1fddd9),
	.w6(32'h3ba3efff),
	.w7(32'h3aae2d86),
	.w8(32'hbac17bde),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59782d),
	.w1(32'h3bc88a47),
	.w2(32'hbabde82f),
	.w3(32'hbc4ff5c9),
	.w4(32'hbc28e6b6),
	.w5(32'h3add0daf),
	.w6(32'h3a1199cd),
	.w7(32'hba45f247),
	.w8(32'h3be59b1f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1291c2),
	.w1(32'hbb9f5645),
	.w2(32'hbbeef348),
	.w3(32'h3b7be2c6),
	.w4(32'h3b912630),
	.w5(32'h3ac5e4b7),
	.w6(32'h3c84b158),
	.w7(32'h3ba1ac22),
	.w8(32'hbb65992c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09d1d2),
	.w1(32'hbb7b6ec5),
	.w2(32'hbb055f76),
	.w3(32'h3b2526a9),
	.w4(32'h3bd3f968),
	.w5(32'h3a938d4c),
	.w6(32'hbad55425),
	.w7(32'hbb18fea3),
	.w8(32'h3babc4ac),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b987acd),
	.w1(32'hbc2c971f),
	.w2(32'hbbb17583),
	.w3(32'h3b9d99e3),
	.w4(32'h3ad0287d),
	.w5(32'hbb72858c),
	.w6(32'hbab8f68c),
	.w7(32'hb93ea991),
	.w8(32'hbb190d7a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26e9c3),
	.w1(32'hbb378899),
	.w2(32'hbb465882),
	.w3(32'h3b2009b2),
	.w4(32'hba971b6d),
	.w5(32'hbb92123a),
	.w6(32'hb9a678e0),
	.w7(32'hbb0a42f7),
	.w8(32'h3aa5b036),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1e733),
	.w1(32'h3bf83190),
	.w2(32'h3bcce884),
	.w3(32'hb82573fd),
	.w4(32'h3a35c61c),
	.w5(32'h3ab3b1c0),
	.w6(32'h3b8e847f),
	.w7(32'h3b313f95),
	.w8(32'hbb361653),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8bbad),
	.w1(32'hbc2ef08d),
	.w2(32'h3b291987),
	.w3(32'h3c32f04c),
	.w4(32'h3beda49e),
	.w5(32'hbaedb8d7),
	.w6(32'hbc04c947),
	.w7(32'h3b456b50),
	.w8(32'hbc065e1a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c71df),
	.w1(32'hbaf9cf6f),
	.w2(32'hbb634929),
	.w3(32'h3a32b3b0),
	.w4(32'h3b425811),
	.w5(32'hbb986b4d),
	.w6(32'hbb1c412d),
	.w7(32'h3b671f63),
	.w8(32'hbc06f8ef),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1b8e9),
	.w1(32'hbc51bd3f),
	.w2(32'hba961ce9),
	.w3(32'h3c18b62c),
	.w4(32'h3c2ebb6c),
	.w5(32'h3bcac857),
	.w6(32'hbc123bcb),
	.w7(32'h3c0ab5bf),
	.w8(32'hbb68ffa2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39215901),
	.w1(32'hbc0b0f6f),
	.w2(32'h3abf1790),
	.w3(32'h3bf43868),
	.w4(32'h3bcd576d),
	.w5(32'hbc260f15),
	.w6(32'h3a9cc452),
	.w7(32'h3b4e7ae5),
	.w8(32'hba160de1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cadca),
	.w1(32'h3babae76),
	.w2(32'h3c502cab),
	.w3(32'hbba374a7),
	.w4(32'hbb0dc1e8),
	.w5(32'hbbe036da),
	.w6(32'h3b782d51),
	.w7(32'h3c2d229a),
	.w8(32'hbad5515d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b3c7d),
	.w1(32'hbb1ef526),
	.w2(32'h37276113),
	.w3(32'hb9b94b4c),
	.w4(32'hbb4bad3c),
	.w5(32'h3be5b801),
	.w6(32'hb92b28e0),
	.w7(32'h3b11ce2d),
	.w8(32'h3bdc9c0c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb30003),
	.w1(32'hbc19011f),
	.w2(32'hbbf9d3fd),
	.w3(32'h3af1b7c5),
	.w4(32'h3ab98d60),
	.w5(32'hbc5a6117),
	.w6(32'h3b80499b),
	.w7(32'h3bba59a4),
	.w8(32'h3b610175),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb343f5),
	.w1(32'h3c6cfb5e),
	.w2(32'h3c227777),
	.w3(32'hbcc921b5),
	.w4(32'hbc5ae7bc),
	.w5(32'hbbb1785e),
	.w6(32'h3c32577c),
	.w7(32'h3c03ac20),
	.w8(32'hbba15a35),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99eb8a),
	.w1(32'h39b9eacf),
	.w2(32'h3ab30412),
	.w3(32'h3b01bbf2),
	.w4(32'hbb642179),
	.w5(32'hb99a248a),
	.w6(32'h3b54fb8c),
	.w7(32'hbaf6a9f0),
	.w8(32'hbb03191f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa9a3e),
	.w1(32'h3969e8f4),
	.w2(32'h3c13ca2f),
	.w3(32'hbae746ee),
	.w4(32'h3b977a44),
	.w5(32'hbb0c1484),
	.w6(32'hbabe1de8),
	.w7(32'h3c285a7e),
	.w8(32'hbc144ad0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68b71b),
	.w1(32'h3b7377f6),
	.w2(32'h3a430b20),
	.w3(32'h3b16ef17),
	.w4(32'hbac539d9),
	.w5(32'h3b86d06d),
	.w6(32'h3be61bf6),
	.w7(32'hbb07827c),
	.w8(32'hbb04f161),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90d413),
	.w1(32'hbb66caab),
	.w2(32'h3aec9b68),
	.w3(32'hbbb3c25b),
	.w4(32'hb9d14850),
	.w5(32'hbbb9119b),
	.w6(32'h3b7b5d5c),
	.w7(32'h3b71ceea),
	.w8(32'hbae13e87),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58b3f7),
	.w1(32'h3a16e6a5),
	.w2(32'hbb6e81cb),
	.w3(32'h3b907ca3),
	.w4(32'h3ae933b2),
	.w5(32'hbba6db31),
	.w6(32'h3c95bc63),
	.w7(32'h398b22ac),
	.w8(32'hbb9eee6d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf9723),
	.w1(32'h3abe0136),
	.w2(32'hba1582bd),
	.w3(32'h3a0f59ec),
	.w4(32'hbbd72128),
	.w5(32'hbbb02727),
	.w6(32'h3b8353ae),
	.w7(32'hbbd4c268),
	.w8(32'hbbdbf782),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb092df),
	.w1(32'hba1b62b6),
	.w2(32'hb8d97bc6),
	.w3(32'hbad693fe),
	.w4(32'h3c03cc05),
	.w5(32'hbb97f69a),
	.w6(32'hbba28b24),
	.w7(32'h3ba03dfc),
	.w8(32'h3ae54263),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2dbe),
	.w1(32'hbbff8c8f),
	.w2(32'hbb0d8c34),
	.w3(32'hbb1c8d3e),
	.w4(32'h3b903e63),
	.w5(32'h3b2d0875),
	.w6(32'hbb5e86cb),
	.w7(32'hbb8a0804),
	.w8(32'h3ab48afc),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c61216),
	.w1(32'h3a753de3),
	.w2(32'h3b8bb89d),
	.w3(32'h3b8699f4),
	.w4(32'h3b7d57c3),
	.w5(32'hbbca6941),
	.w6(32'hbb0993c9),
	.w7(32'hb97d9dc5),
	.w8(32'hbbe4a011),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd857b),
	.w1(32'hbc281ed2),
	.w2(32'h3bb02715),
	.w3(32'hbb4e3894),
	.w4(32'h3a8bacb2),
	.w5(32'h3b9bf1af),
	.w6(32'hbc5ef078),
	.w7(32'hbad90afb),
	.w8(32'h3a00ceb5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11d35e),
	.w1(32'h3aa380c8),
	.w2(32'hb87ff882),
	.w3(32'h3a10763f),
	.w4(32'hbaaa6a6e),
	.w5(32'h3b04bf3f),
	.w6(32'h3ba58214),
	.w7(32'h3b3ca5f1),
	.w8(32'hbb93ebc8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9084e),
	.w1(32'hbba8723e),
	.w2(32'h3bce40e0),
	.w3(32'hbc0e13de),
	.w4(32'h3b88e9cd),
	.w5(32'hbae6a224),
	.w6(32'hbc40b30e),
	.w7(32'h3bae9e82),
	.w8(32'hbb05c063),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56d35b),
	.w1(32'hbb5a77c6),
	.w2(32'hbc031132),
	.w3(32'hba9c2b86),
	.w4(32'hbbdbb4e6),
	.w5(32'hbb978bb4),
	.w6(32'hbaf794f4),
	.w7(32'hbba271ff),
	.w8(32'hbc02fcf1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb880cdf),
	.w1(32'hbba7bfd6),
	.w2(32'h39c9ec6f),
	.w3(32'hbba51d7f),
	.w4(32'hbb84e45d),
	.w5(32'hbba95d0d),
	.w6(32'h3b04ab79),
	.w7(32'h3b7386f6),
	.w8(32'hbbf9a39e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0719c8),
	.w1(32'h3a27286b),
	.w2(32'h3a04169e),
	.w3(32'hbb62e498),
	.w4(32'hbb458c76),
	.w5(32'hbbbfb212),
	.w6(32'h3b3c1f0c),
	.w7(32'hbb4122c6),
	.w8(32'hbbbd7a28),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb957b5e),
	.w1(32'hbbca30fa),
	.w2(32'hbbbd8e17),
	.w3(32'hbb841632),
	.w4(32'hbbe3c01a),
	.w5(32'h3ab95861),
	.w6(32'hbb60ba60),
	.w7(32'hbc1dc970),
	.w8(32'h3959fef0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a9daa),
	.w1(32'h3b0f9312),
	.w2(32'h3bcac908),
	.w3(32'hbb50dcbc),
	.w4(32'hbb9ff1c7),
	.w5(32'h3c2977cb),
	.w6(32'hbb5ba1e8),
	.w7(32'hbb408a4c),
	.w8(32'hbab6feb0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6417ab),
	.w1(32'h3c48e991),
	.w2(32'h3c1ded40),
	.w3(32'h3c67c03a),
	.w4(32'h3b429957),
	.w5(32'hbbe7ea1a),
	.w6(32'h3c1d6c18),
	.w7(32'h3c57fbb2),
	.w8(32'hbbbcb29d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1e187),
	.w1(32'hba9ff459),
	.w2(32'h3b3a1beb),
	.w3(32'h3b437758),
	.w4(32'hbb0b86de),
	.w5(32'h3b61fe43),
	.w6(32'h3c8665c7),
	.w7(32'hba7eb4ab),
	.w8(32'h3ac8c1e2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b2aff),
	.w1(32'h3ac6e295),
	.w2(32'h3b828776),
	.w3(32'h3af97f2c),
	.w4(32'h3b79da2a),
	.w5(32'hbbd2161c),
	.w6(32'hba0dc4d4),
	.w7(32'h3b930f04),
	.w8(32'hbbaa6dbd),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc044020),
	.w1(32'hbb7ac72d),
	.w2(32'hbbddca10),
	.w3(32'hbb4a0cfa),
	.w4(32'hbb7a7300),
	.w5(32'h3b3397fa),
	.w6(32'hbb62ee3c),
	.w7(32'h3b0be03b),
	.w8(32'h3aa8e4cb),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1021a),
	.w1(32'h3c2a4e08),
	.w2(32'h3b105be1),
	.w3(32'h3c9068ac),
	.w4(32'h3b793e51),
	.w5(32'hbc1a4d1c),
	.w6(32'h3c4a46d1),
	.w7(32'h3b0dd4e0),
	.w8(32'hb97b9c16),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1862f),
	.w1(32'hba38e13d),
	.w2(32'hbb9284bd),
	.w3(32'hbb4ed498),
	.w4(32'h39e66cdf),
	.w5(32'h3aaf8595),
	.w6(32'hbba53bcd),
	.w7(32'hba5a4a31),
	.w8(32'h3957ff85),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b122350),
	.w1(32'hbb14e124),
	.w2(32'h3aa5b9e0),
	.w3(32'hbb0d9e21),
	.w4(32'hbb77cdff),
	.w5(32'h3bdf8b59),
	.w6(32'hbaea0653),
	.w7(32'hbb701ad4),
	.w8(32'h3c5da930),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a78e7),
	.w1(32'hbbfa15f1),
	.w2(32'hbaa9a2f5),
	.w3(32'hbbeba6b6),
	.w4(32'h3a6a6ff5),
	.w5(32'h3b9de25a),
	.w6(32'hbc1c7c1e),
	.w7(32'hb9c38c8b),
	.w8(32'hbc30a6a8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba34171),
	.w1(32'hbbafc14e),
	.w2(32'hbb894290),
	.w3(32'hbaaa0004),
	.w4(32'hbbe4d229),
	.w5(32'hbc16330f),
	.w6(32'hbb26a178),
	.w7(32'hbb19806a),
	.w8(32'hbb0fd8b1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe60ac),
	.w1(32'hbacc3e3a),
	.w2(32'h3a472fb7),
	.w3(32'hbb4fa42d),
	.w4(32'h3ab0cd43),
	.w5(32'h3b1da294),
	.w6(32'hbb3ac516),
	.w7(32'h3b6383cf),
	.w8(32'h390f6ccb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc536f42),
	.w1(32'hba043105),
	.w2(32'h392c9cf8),
	.w3(32'hbb6f7d8d),
	.w4(32'hbafb0184),
	.w5(32'h3bbbc0ab),
	.w6(32'h3952edf8),
	.w7(32'hba09e630),
	.w8(32'h3bc60815),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8738d4),
	.w1(32'hb9581381),
	.w2(32'hbb40353b),
	.w3(32'hba89a016),
	.w4(32'h3b3b6320),
	.w5(32'h3aa8a8fe),
	.w6(32'hbb5c9d91),
	.w7(32'hbc08584e),
	.w8(32'hbb175ae1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9d6f4),
	.w1(32'hb96c384e),
	.w2(32'h3a7db2b5),
	.w3(32'hba64f150),
	.w4(32'h3b362f32),
	.w5(32'h3c5bfffb),
	.w6(32'h3bb392f1),
	.w7(32'h3b0fdc0f),
	.w8(32'h3cbd5b1e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e663c),
	.w1(32'hba0583d6),
	.w2(32'h3be1c03b),
	.w3(32'hba519ff1),
	.w4(32'h3ba6710e),
	.w5(32'hbbc7901c),
	.w6(32'hbc42eb59),
	.w7(32'hba904731),
	.w8(32'hbb0c23b5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0d186),
	.w1(32'h3b3d7505),
	.w2(32'hbb2716a5),
	.w3(32'h3bc85b26),
	.w4(32'hbbbafc50),
	.w5(32'hbb2136e3),
	.w6(32'h3b1589f7),
	.w7(32'hbbd32f20),
	.w8(32'h3a174b32),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ef362),
	.w1(32'hbaffb239),
	.w2(32'h3a5447a3),
	.w3(32'hbaa37cb9),
	.w4(32'h3ae239fa),
	.w5(32'hbbc8f307),
	.w6(32'h3b4fc5a7),
	.w7(32'h3bac630a),
	.w8(32'hbc2c33b0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcccbd),
	.w1(32'hbc888a47),
	.w2(32'hbbb01bbb),
	.w3(32'hbb164a91),
	.w4(32'hbc283759),
	.w5(32'h3a3ec68e),
	.w6(32'hbb082977),
	.w7(32'hbc8f0979),
	.w8(32'hbbf7c77d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e3487),
	.w1(32'h3a2a0f95),
	.w2(32'h3b3b6f48),
	.w3(32'h3961ca8d),
	.w4(32'h3a729e50),
	.w5(32'h3b3dcf6c),
	.w6(32'h3c0de574),
	.w7(32'h3bd77b21),
	.w8(32'hbaf48c7b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d14e4),
	.w1(32'hbb29887f),
	.w2(32'hbb3d0ea5),
	.w3(32'h3b9f6308),
	.w4(32'h3b9988d4),
	.w5(32'h3afaf371),
	.w6(32'h3ba7b0b3),
	.w7(32'h3bd7e3e3),
	.w8(32'h3b112428),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f4503),
	.w1(32'h3a8f071c),
	.w2(32'h3a0b00df),
	.w3(32'hb9d7cd66),
	.w4(32'h398c5bdf),
	.w5(32'h3c0e8d12),
	.w6(32'h3b78f881),
	.w7(32'h3aa37b70),
	.w8(32'h3c35a6e0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6e8fb),
	.w1(32'h3c0d5bf0),
	.w2(32'h3ba8aeac),
	.w3(32'h3be5929d),
	.w4(32'h3b9f6c95),
	.w5(32'hbb5cd2e2),
	.w6(32'h3c2b067d),
	.w7(32'h3b8ddc41),
	.w8(32'hbbb6446c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b2448),
	.w1(32'hbbae7ada),
	.w2(32'hbb0ac4f6),
	.w3(32'hba9ea0a4),
	.w4(32'hbb5c8ca0),
	.w5(32'hba3ceb19),
	.w6(32'h3aeec526),
	.w7(32'hbb22555a),
	.w8(32'hbb008f9d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81fdb7e),
	.w1(32'h3a39585e),
	.w2(32'hbb263ad2),
	.w3(32'h3a23a484),
	.w4(32'hbaa679d1),
	.w5(32'h39e348d5),
	.w6(32'h3b05397f),
	.w7(32'hbaa6d031),
	.w8(32'hb954223e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb887e1ed),
	.w1(32'hb9b8966e),
	.w2(32'h3991f38f),
	.w3(32'hba8680be),
	.w4(32'hbab33ead),
	.w5(32'h3b46676b),
	.w6(32'h3a22c364),
	.w7(32'hba0fab62),
	.w8(32'h3b1b377b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68455d),
	.w1(32'h3a6fb2f8),
	.w2(32'h3a492863),
	.w3(32'h39157b8f),
	.w4(32'hbb34dcd2),
	.w5(32'h3c1352a0),
	.w6(32'h3be6862f),
	.w7(32'hba101dd1),
	.w8(32'h3c0dd26e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5c71d),
	.w1(32'hbaa8f060),
	.w2(32'h3b282768),
	.w3(32'hbb46f77c),
	.w4(32'hbb2285af),
	.w5(32'hbb393e46),
	.w6(32'hbbef3597),
	.w7(32'hb86b0417),
	.w8(32'hbb573688),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a7760),
	.w1(32'hbadd9cc8),
	.w2(32'h3bc89a33),
	.w3(32'h3b45d582),
	.w4(32'h3b043265),
	.w5(32'h39e8b8fb),
	.w6(32'hbb1d7ca3),
	.w7(32'h3ba9e5ba),
	.w8(32'hbb0d5efc),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399feed5),
	.w1(32'h3c1679b3),
	.w2(32'h3b17a979),
	.w3(32'h3b71acf5),
	.w4(32'h3b757a70),
	.w5(32'h3ac9e212),
	.w6(32'h3b1b78a8),
	.w7(32'h3b52f1fe),
	.w8(32'h3b923c22),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add15dc),
	.w1(32'h3b8d13b6),
	.w2(32'h3b9eced0),
	.w3(32'hb9e40e86),
	.w4(32'hba1533eb),
	.w5(32'hbb31c9ff),
	.w6(32'h3bb659c5),
	.w7(32'h3b88c896),
	.w8(32'hbb881595),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6fb2b),
	.w1(32'h3b3a2882),
	.w2(32'h39d235c2),
	.w3(32'h3bd37893),
	.w4(32'hbb0f66ce),
	.w5(32'h3b852182),
	.w6(32'h3c6b8fc1),
	.w7(32'h3b0ccf3e),
	.w8(32'h3b838106),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f9d83),
	.w1(32'hbb1b0ca3),
	.w2(32'hba5a341a),
	.w3(32'h3bc9ea88),
	.w4(32'h3ac7fa08),
	.w5(32'h391b55fa),
	.w6(32'h3c19fa79),
	.w7(32'h3ae37b1a),
	.w8(32'h3bc14a0b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5a720),
	.w1(32'hbb42c4c2),
	.w2(32'hbafbdd36),
	.w3(32'h3ab3bbfb),
	.w4(32'hbab44a0b),
	.w5(32'hbbae7ebb),
	.w6(32'hbbcbfcd2),
	.w7(32'h3a5f2953),
	.w8(32'hbbbaaada),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ecdb4),
	.w1(32'hb9b08c1a),
	.w2(32'hbb48546f),
	.w3(32'h3b9f775b),
	.w4(32'h3b632498),
	.w5(32'h3acff647),
	.w6(32'h3bab1994),
	.w7(32'h3bffbc14),
	.w8(32'hbba7e129),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfadf00),
	.w1(32'h3bafe89c),
	.w2(32'hbb473e98),
	.w3(32'hbb0c2d69),
	.w4(32'hbb813cd4),
	.w5(32'hbb663c14),
	.w6(32'h39540e14),
	.w7(32'hbbec45fb),
	.w8(32'hbc08866a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb38d60),
	.w1(32'h3c46634b),
	.w2(32'h3b9cda38),
	.w3(32'h3c6cc32a),
	.w4(32'hb915cfd2),
	.w5(32'h3b326502),
	.w6(32'h3cdd01c9),
	.w7(32'h3b101fec),
	.w8(32'h390d6699),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c95db),
	.w1(32'hba484a18),
	.w2(32'h3ae85f3c),
	.w3(32'hba613fae),
	.w4(32'h3b003ec6),
	.w5(32'hbb28c53e),
	.w6(32'hbb6cd3de),
	.w7(32'h3983c548),
	.w8(32'hbaec4f4f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b667bd),
	.w1(32'h3b9318ba),
	.w2(32'h3b4a7428),
	.w3(32'h3af7b4ba),
	.w4(32'hbb598207),
	.w5(32'h3b9aa19f),
	.w6(32'hba81b1c2),
	.w7(32'hbae678ba),
	.w8(32'h3c124ad4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a295b),
	.w1(32'h3bdb07bf),
	.w2(32'h3a9e154f),
	.w3(32'h3c0f17b7),
	.w4(32'h3ab094f7),
	.w5(32'hbc09bf42),
	.w6(32'h3bdc5825),
	.w7(32'h3ba2fb17),
	.w8(32'hbb1d60f8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0311ae),
	.w1(32'hbbdf5c3b),
	.w2(32'hbbd4fe85),
	.w3(32'h3b1f85d3),
	.w4(32'hbb921c5e),
	.w5(32'hba909b54),
	.w6(32'h3b2ce905),
	.w7(32'hbb698f39),
	.w8(32'hbb9f2d6d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a60c6a),
	.w1(32'h3b4fd7a0),
	.w2(32'h3c0b5b75),
	.w3(32'h3bb47801),
	.w4(32'h3b926e2e),
	.w5(32'h3ac6c989),
	.w6(32'h3c3efdac),
	.w7(32'h3bc154cf),
	.w8(32'h3abf4d5e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab55dcd),
	.w1(32'hbbf1d6bb),
	.w2(32'hbaa21348),
	.w3(32'hbbbf4961),
	.w4(32'h3aaecb4e),
	.w5(32'hbb06835f),
	.w6(32'h3a6651ee),
	.w7(32'h3b4f925d),
	.w8(32'hb9f1b15b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebaa86),
	.w1(32'hbb3de1da),
	.w2(32'hbc367f87),
	.w3(32'hba10e38f),
	.w4(32'hbc3596de),
	.w5(32'hbb23835a),
	.w6(32'hbb8b99cb),
	.w7(32'hbc44ce5a),
	.w8(32'hbb2a76b8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19ed52),
	.w1(32'hbb24968e),
	.w2(32'hb9ea233c),
	.w3(32'hbb2b721b),
	.w4(32'h3bc0529d),
	.w5(32'h39f2c916),
	.w6(32'hbb515883),
	.w7(32'h37a73ff4),
	.w8(32'h3ae57c24),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1cab8),
	.w1(32'hbc37d84f),
	.w2(32'h3bd914f8),
	.w3(32'hbbc0722b),
	.w4(32'h3b8c6ad9),
	.w5(32'hbae6aa5c),
	.w6(32'hbbe923b7),
	.w7(32'h3aade32e),
	.w8(32'h3bee46b0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe4f31),
	.w1(32'hb9fe246f),
	.w2(32'h3a28ec1a),
	.w3(32'hbac225fd),
	.w4(32'hbb8d6707),
	.w5(32'h3bada96a),
	.w6(32'h3a053991),
	.w7(32'h3a1e9c83),
	.w8(32'h3c1813e8),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0693a5),
	.w1(32'hbae4f4ae),
	.w2(32'h3bbc3d57),
	.w3(32'h3b941a3e),
	.w4(32'h3a316cdb),
	.w5(32'hb9425a3c),
	.w6(32'hba6e929a),
	.w7(32'h3b451fc1),
	.w8(32'h3c9715ae),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c449fb3),
	.w1(32'hbb076802),
	.w2(32'h3ba2f94d),
	.w3(32'h3b90e8aa),
	.w4(32'h3c27cebd),
	.w5(32'h3abe3718),
	.w6(32'h3c0c4049),
	.w7(32'h3c0bba20),
	.w8(32'h3c1fcac4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26ace6),
	.w1(32'hba84da2e),
	.w2(32'h3a15f853),
	.w3(32'hbb435d11),
	.w4(32'hba748f92),
	.w5(32'hb9ff2521),
	.w6(32'hbc249d5a),
	.w7(32'h3af8525d),
	.w8(32'h3b9fea6a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19cf58),
	.w1(32'hb9374eec),
	.w2(32'hbbd4c761),
	.w3(32'h3b0950aa),
	.w4(32'hbadc45b4),
	.w5(32'h3b9c6215),
	.w6(32'hbaebedf8),
	.w7(32'hbbfb2ef1),
	.w8(32'h3af789d2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c603e16),
	.w1(32'h3c6ef32d),
	.w2(32'h3be4c92b),
	.w3(32'h3c7dcff7),
	.w4(32'h3a904a09),
	.w5(32'hbb4d402b),
	.w6(32'h3c8cc997),
	.w7(32'h3bccc2b7),
	.w8(32'h3c4f51f0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c3224),
	.w1(32'hbb67be07),
	.w2(32'hbbcf9044),
	.w3(32'h3aabdc54),
	.w4(32'hbaa68408),
	.w5(32'hbb38524d),
	.w6(32'hbb48b8a5),
	.w7(32'hbb843bdf),
	.w8(32'hbb4948a9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18b076),
	.w1(32'hbb351190),
	.w2(32'h39cf38c0),
	.w3(32'hbbd07ff4),
	.w4(32'hba3d96c9),
	.w5(32'hbc0cbbb1),
	.w6(32'h3ac2776b),
	.w7(32'h3a9fbfd3),
	.w8(32'h3b8ecdad),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f6651),
	.w1(32'h3b7f824a),
	.w2(32'hba96cf9f),
	.w3(32'hb98df9f7),
	.w4(32'hba10ad60),
	.w5(32'h3b1dc31b),
	.w6(32'h3ba45ba9),
	.w7(32'h3b3c4411),
	.w8(32'hb80653a2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ce49c),
	.w1(32'hba088e31),
	.w2(32'hbb07380e),
	.w3(32'h3b2bd82c),
	.w4(32'h3b8a85d5),
	.w5(32'hbab22dbb),
	.w6(32'hb9f469d7),
	.w7(32'h3b7da95a),
	.w8(32'h3b0265a3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d5852),
	.w1(32'hbb318dfa),
	.w2(32'h3b44e407),
	.w3(32'hbbbf0d4e),
	.w4(32'hbb977fde),
	.w5(32'h3b393e0a),
	.w6(32'hbbd7bdb7),
	.w7(32'hbbaf7a4d),
	.w8(32'hbb35b2c4),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b194948),
	.w1(32'h3b8f940d),
	.w2(32'h3bbd733e),
	.w3(32'h3ab6d2a9),
	.w4(32'h3bc5c57e),
	.w5(32'hbbe34570),
	.w6(32'h3c25924f),
	.w7(32'h3bc58114),
	.w8(32'hbc04010d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb948a50),
	.w1(32'hb8dfe7d9),
	.w2(32'h3ac59507),
	.w3(32'hbabeda12),
	.w4(32'h3b9c3360),
	.w5(32'h3afc5759),
	.w6(32'h3abd6ca6),
	.w7(32'h3bb6a9ac),
	.w8(32'h3a169046),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98e767),
	.w1(32'h3a6ac724),
	.w2(32'h3b0c2587),
	.w3(32'h3b28581f),
	.w4(32'hbb12bead),
	.w5(32'hbb99bd0d),
	.w6(32'h3c379b00),
	.w7(32'h3c0b8e94),
	.w8(32'h3b363211),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a3b4d),
	.w1(32'h3b8f3b86),
	.w2(32'h3ba83082),
	.w3(32'h3b124e00),
	.w4(32'h3ad148f5),
	.w5(32'hbb0dd3fd),
	.w6(32'h3bca3ff8),
	.w7(32'h3b92aef0),
	.w8(32'hbbeeb2ba),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d78c0),
	.w1(32'hbbffda6a),
	.w2(32'h3b09d249),
	.w3(32'hbc0f79e6),
	.w4(32'hbb4430f3),
	.w5(32'hbb7da277),
	.w6(32'hbbee0e26),
	.w7(32'hb88a78f8),
	.w8(32'hbb83927c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc146aa6),
	.w1(32'hbbeeb2c3),
	.w2(32'h3b7e05c9),
	.w3(32'hbc0ebf52),
	.w4(32'hbada05d4),
	.w5(32'hbaa40da7),
	.w6(32'hbb5a9735),
	.w7(32'h3b380879),
	.w8(32'h38d8c0fe),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b060b15),
	.w1(32'h3afc011c),
	.w2(32'hbb41c716),
	.w3(32'h3afb8ead),
	.w4(32'hba258877),
	.w5(32'hbb38bcd9),
	.w6(32'h3b73e883),
	.w7(32'h3a117b7e),
	.w8(32'h3b29e521),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1e6ab),
	.w1(32'h3b3af6f0),
	.w2(32'h3c02ab43),
	.w3(32'h3ab0527f),
	.w4(32'h3ac8cbbc),
	.w5(32'h3a82146c),
	.w6(32'h3b37eddf),
	.w7(32'h3c0b1196),
	.w8(32'h39088f89),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eb726),
	.w1(32'hbaca18a7),
	.w2(32'hb931f593),
	.w3(32'hbb392442),
	.w4(32'h3ab99664),
	.w5(32'hbba5378f),
	.w6(32'h3b285b88),
	.w7(32'hb9a9eddb),
	.w8(32'hbc678f88),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a2471),
	.w1(32'h3c8f99f9),
	.w2(32'hbaa351a2),
	.w3(32'h3bb2058d),
	.w4(32'h3b9c70e6),
	.w5(32'h39077491),
	.w6(32'h3d12f68f),
	.w7(32'h3a27f801),
	.w8(32'hbc081acd),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde28ad),
	.w1(32'h3b07df08),
	.w2(32'h3a9e3fe6),
	.w3(32'h3bd0e3ba),
	.w4(32'h39c943d6),
	.w5(32'h3c0f22d3),
	.w6(32'h3b8e6517),
	.w7(32'h3b819dd0),
	.w8(32'h3a833c84),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8797690),
	.w1(32'h3b951350),
	.w2(32'h3b6b3fe7),
	.w3(32'h3a6c2d84),
	.w4(32'hbaf5c67c),
	.w5(32'h3be60fdc),
	.w6(32'h3b87983f),
	.w7(32'h3af841cb),
	.w8(32'h3c2c20d1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd827a2),
	.w1(32'hbbd46bf3),
	.w2(32'hbb52e5ea),
	.w3(32'hbb836df0),
	.w4(32'h3a83bc86),
	.w5(32'h3bed1ba4),
	.w6(32'hbc031798),
	.w7(32'hbc47775b),
	.w8(32'hba352134),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c0064),
	.w1(32'h3bf9d004),
	.w2(32'hb9ec1904),
	.w3(32'h3ac7c370),
	.w4(32'hba2ed250),
	.w5(32'hbb945635),
	.w6(32'h3b9537cf),
	.w7(32'hbb26e33a),
	.w8(32'hbba44dbb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda0a4c),
	.w1(32'hba60e473),
	.w2(32'hbb9a5c64),
	.w3(32'hbb72f508),
	.w4(32'hba8b6eb5),
	.w5(32'hbabc2b94),
	.w6(32'hbabaac5d),
	.w7(32'hbb1f25f7),
	.w8(32'hbb06e6bf),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ecda2),
	.w1(32'h39976e90),
	.w2(32'h3af0a9f9),
	.w3(32'hb998b2bd),
	.w4(32'hbaf7717f),
	.w5(32'hbb7844e6),
	.w6(32'hbadb41de),
	.w7(32'h3a7d104f),
	.w8(32'hbc051f50),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc582f),
	.w1(32'hbbabddfd),
	.w2(32'h3a09893c),
	.w3(32'hbc0340b7),
	.w4(32'h3b597994),
	.w5(32'h3ac2425b),
	.w6(32'hbb41bc23),
	.w7(32'hbb9083bb),
	.w8(32'h3a803714),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae505bd),
	.w1(32'h3a35f159),
	.w2(32'hb9a5d727),
	.w3(32'h3ab1ac9a),
	.w4(32'h3a434529),
	.w5(32'h3b5e59c4),
	.w6(32'h3b365b2c),
	.w7(32'hbaa263c0),
	.w8(32'hbb1fc3b3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba96ec8),
	.w1(32'hbbf1f28c),
	.w2(32'hbbb5d230),
	.w3(32'hbbd6cd01),
	.w4(32'h3b490bee),
	.w5(32'hbc3aa946),
	.w6(32'hbbf05702),
	.w7(32'hbad9c6ec),
	.w8(32'hbb12a3a3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6093ec),
	.w1(32'hbab4a796),
	.w2(32'h3a4b2b32),
	.w3(32'hbb95e609),
	.w4(32'h3a88f664),
	.w5(32'h3a6a43b0),
	.w6(32'h3b21bafc),
	.w7(32'h3b042f94),
	.w8(32'hbbca267a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5854b),
	.w1(32'hbb8fcbc8),
	.w2(32'h3b1eb3c4),
	.w3(32'hbb2eb687),
	.w4(32'hbb273ef6),
	.w5(32'h39769eb2),
	.w6(32'h3b55ac88),
	.w7(32'hba038f58),
	.w8(32'h3a7b0bfe),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cea7e6),
	.w1(32'h3a8b866e),
	.w2(32'h39b1f0ee),
	.w3(32'hbbdb6728),
	.w4(32'hbb85f86b),
	.w5(32'hbb86467b),
	.w6(32'hbbcdb4f5),
	.w7(32'hbb258338),
	.w8(32'hba640445),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8caf9),
	.w1(32'h3a2f77b5),
	.w2(32'hbb5a511b),
	.w3(32'hbaa310e6),
	.w4(32'hbbdff35e),
	.w5(32'h3b8895ad),
	.w6(32'hbab2e163),
	.w7(32'hbb495b67),
	.w8(32'hbad902b5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe04a54),
	.w1(32'h3b10a56e),
	.w2(32'hbb3e1c89),
	.w3(32'h3b93b009),
	.w4(32'h3a6891f2),
	.w5(32'h3c19e65c),
	.w6(32'h3bd3d998),
	.w7(32'hbb668efb),
	.w8(32'hba5a13ba),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb987e43),
	.w1(32'h3a904d55),
	.w2(32'hb895f9e3),
	.w3(32'hbbacc08a),
	.w4(32'hbb2b0004),
	.w5(32'h3b3163eb),
	.w6(32'hbbe086d2),
	.w7(32'hb799d6aa),
	.w8(32'hbad93c18),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bf087),
	.w1(32'h3a113cf6),
	.w2(32'hbb455c0a),
	.w3(32'hb7baa944),
	.w4(32'hba9cd24b),
	.w5(32'hbbe01957),
	.w6(32'h3b031145),
	.w7(32'hbb64ea9f),
	.w8(32'hbbcacf7d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba32132),
	.w1(32'hba979ddf),
	.w2(32'h3a8bddfc),
	.w3(32'hbc309c92),
	.w4(32'hbbdd00a9),
	.w5(32'h3c007fc1),
	.w6(32'hbb60a236),
	.w7(32'hba368d73),
	.w8(32'h3c352739),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0ac41),
	.w1(32'h3c0f9e72),
	.w2(32'h3be02c79),
	.w3(32'h3c51e91a),
	.w4(32'h3be505de),
	.w5(32'h3a63a127),
	.w6(32'h3cb6153e),
	.w7(32'h3729b0a9),
	.w8(32'h394eae45),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a601b9),
	.w1(32'h39d6e514),
	.w2(32'h3ace3989),
	.w3(32'h3b987944),
	.w4(32'h3a3dda4c),
	.w5(32'hbbe46184),
	.w6(32'hbb509828),
	.w7(32'h3b92feef),
	.w8(32'hbbe0c3e0),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb6025),
	.w1(32'hbb237132),
	.w2(32'h39594d15),
	.w3(32'h39daed71),
	.w4(32'h39478e47),
	.w5(32'hbbd078dc),
	.w6(32'h3b310728),
	.w7(32'h3aae1024),
	.w8(32'hbbf8c2ad),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9a1ca),
	.w1(32'h3c0d04f7),
	.w2(32'hb8f5fd52),
	.w3(32'h3bcf2d1a),
	.w4(32'h3a6762f9),
	.w5(32'hbbbb077e),
	.w6(32'h3ccba3e5),
	.w7(32'h3adbeb5a),
	.w8(32'hbc023eed),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0986fb),
	.w1(32'hbb0f6938),
	.w2(32'hbb637a39),
	.w3(32'hbb89381f),
	.w4(32'hbb905726),
	.w5(32'hbb144038),
	.w6(32'hbbda9595),
	.w7(32'hba973e32),
	.w8(32'hba65d0a3),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba13766),
	.w1(32'h3ad4cd0e),
	.w2(32'h3b3d836e),
	.w3(32'h3b6a7b64),
	.w4(32'hba0e8796),
	.w5(32'h3a867188),
	.w6(32'h3a9a1dce),
	.w7(32'hbbc31fd8),
	.w8(32'h3b858449),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccb058),
	.w1(32'hbb494355),
	.w2(32'hbb8f4a6d),
	.w3(32'hbb2afab6),
	.w4(32'hbb934c52),
	.w5(32'hbb2f6615),
	.w6(32'hbba1e8ba),
	.w7(32'hbba047e9),
	.w8(32'hba8c6aa3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab11bce),
	.w1(32'h3b639c96),
	.w2(32'h3980db05),
	.w3(32'h3abdc621),
	.w4(32'h39c0d2f7),
	.w5(32'hbb370926),
	.w6(32'hba04488c),
	.w7(32'h3b1d75ff),
	.w8(32'hb9d88678),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb5427),
	.w1(32'h3b435f36),
	.w2(32'h3aa6cb37),
	.w3(32'h3b661dda),
	.w4(32'hbbde512c),
	.w5(32'hba966960),
	.w6(32'h3b1c9413),
	.w7(32'hbab27da2),
	.w8(32'hbaf53cc0),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c0a4e),
	.w1(32'hba5d3360),
	.w2(32'h3bb2d5e7),
	.w3(32'hba0819ee),
	.w4(32'hba0b075f),
	.w5(32'hbb367d81),
	.w6(32'h3b196d48),
	.w7(32'h3bfde237),
	.w8(32'hbbaebd34),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86d359),
	.w1(32'h3a102aae),
	.w2(32'h3bf632ad),
	.w3(32'h3b359c07),
	.w4(32'h3bc1c98e),
	.w5(32'h3afbaa6f),
	.w6(32'h3bded7dc),
	.w7(32'h3c1771c6),
	.w8(32'h3b9151d5),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4830d9),
	.w1(32'h3a249e67),
	.w2(32'hba9bb893),
	.w3(32'hbad9696c),
	.w4(32'hbae1aa35),
	.w5(32'h3934105b),
	.w6(32'h3b849d50),
	.w7(32'h3a4d072d),
	.w8(32'hbb9703d7),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1925c0),
	.w1(32'h3a321615),
	.w2(32'hbba7f279),
	.w3(32'hbb8975ce),
	.w4(32'h3b08f7e3),
	.w5(32'hbbcc0858),
	.w6(32'hba264ed4),
	.w7(32'hbb8a58d9),
	.w8(32'hbb0f41ed),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a92cc),
	.w1(32'h3b8ffae2),
	.w2(32'h3b6054e6),
	.w3(32'h3b8c403e),
	.w4(32'h3b42b5f8),
	.w5(32'hbbcbf8ed),
	.w6(32'h3b26924d),
	.w7(32'h3b0f5885),
	.w8(32'h3abd89c2),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfda03),
	.w1(32'h3b6863a3),
	.w2(32'h3b75b3d8),
	.w3(32'h3bffea28),
	.w4(32'hb8346156),
	.w5(32'h3bd3c17f),
	.w6(32'h3ca48704),
	.w7(32'hbb16d15a),
	.w8(32'h3b52bfa2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa30bd6),
	.w1(32'hbb3d8591),
	.w2(32'h3a81e5c2),
	.w3(32'h3adddb31),
	.w4(32'h3b759f9a),
	.w5(32'hbbb825c3),
	.w6(32'h3b1b6be2),
	.w7(32'h3b15be89),
	.w8(32'hbb0e1cee),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9572c5e),
	.w1(32'hbb3851ea),
	.w2(32'hbbb0ddf1),
	.w3(32'h3bc45467),
	.w4(32'hbba9f9c4),
	.w5(32'h3af3da8c),
	.w6(32'h3bdadbd6),
	.w7(32'hbc5f0ad6),
	.w8(32'hbc33ece6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabb290),
	.w1(32'hbb5ca438),
	.w2(32'h3a583b65),
	.w3(32'hbb82a62a),
	.w4(32'hbbe88296),
	.w5(32'hbb1e8652),
	.w6(32'h3b735d97),
	.w7(32'h3a5f6385),
	.w8(32'h399f660c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb841509),
	.w1(32'hbc1431c5),
	.w2(32'h39f719b3),
	.w3(32'hba3225b5),
	.w4(32'hbba16e44),
	.w5(32'hbb7ae7a6),
	.w6(32'h3b26ca92),
	.w7(32'hbb0eae46),
	.w8(32'hb7b2b29e),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb560732),
	.w1(32'hbbbb42bb),
	.w2(32'hbb4aca5b),
	.w3(32'hbb4e0b77),
	.w4(32'h3b60f913),
	.w5(32'h3b94e327),
	.w6(32'hbbdee5d2),
	.w7(32'hbb95d85b),
	.w8(32'h3bbc6ead),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee7e7e),
	.w1(32'h3aa885e5),
	.w2(32'h3b597f01),
	.w3(32'h3bad8c44),
	.w4(32'h3b9d4636),
	.w5(32'hb9a5f8a8),
	.w6(32'h3bf42fa8),
	.w7(32'h3b81fa82),
	.w8(32'hba923e8d),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e707f),
	.w1(32'hbc2d3df1),
	.w2(32'h3c74f515),
	.w3(32'hbc393db0),
	.w4(32'h3c0ad9d5),
	.w5(32'h3c4de7ca),
	.w6(32'hbbd9005b),
	.w7(32'h3c2b3596),
	.w8(32'h3c7550d3),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd64cd),
	.w1(32'h3a06684c),
	.w2(32'hbb5fa2da),
	.w3(32'h3a5bc7d5),
	.w4(32'hbb5693f4),
	.w5(32'hbb0d3e89),
	.w6(32'hbc00d9e9),
	.w7(32'hba6004f2),
	.w8(32'hbc8028f8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12f855),
	.w1(32'hbb309e3a),
	.w2(32'h3c215e48),
	.w3(32'h3aa2b320),
	.w4(32'h3c01af00),
	.w5(32'h3bdb3f46),
	.w6(32'h3c9b7a54),
	.w7(32'hbb01260c),
	.w8(32'h3c76be94),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9219b0),
	.w1(32'hbacec860),
	.w2(32'h3b55b0f7),
	.w3(32'h3be586dd),
	.w4(32'h3a69d1f6),
	.w5(32'hbba0afd1),
	.w6(32'h3b80c19c),
	.w7(32'h3ba6fe6f),
	.w8(32'hbbff0d21),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd28f1d),
	.w1(32'hbb8e2edd),
	.w2(32'hbbfddcf1),
	.w3(32'h3a94f9fa),
	.w4(32'hbbf4060d),
	.w5(32'hbbef4d03),
	.w6(32'h3bbd458c),
	.w7(32'hbbdf9910),
	.w8(32'hbc1fd2b3),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaab197),
	.w1(32'h3a3c847b),
	.w2(32'h3b47f7a2),
	.w3(32'h3af48337),
	.w4(32'h3a99e451),
	.w5(32'hbba1aa55),
	.w6(32'h3bf2a64f),
	.w7(32'h3b17ac46),
	.w8(32'hbbeee6a5),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3750b17c),
	.w1(32'h3b8435d6),
	.w2(32'h3ba0d662),
	.w3(32'h3ad72f73),
	.w4(32'h3b11f92e),
	.w5(32'hbbfd6f4f),
	.w6(32'h3ac70b43),
	.w7(32'h3ae25163),
	.w8(32'hbc38ad6e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1de1e4),
	.w1(32'h3bb2b88d),
	.w2(32'h3b6af446),
	.w3(32'h3ab8dedf),
	.w4(32'h3be6f89e),
	.w5(32'hbbb3fc79),
	.w6(32'h3af49b7f),
	.w7(32'h3bf71cc1),
	.w8(32'hb9c40b9b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93de3b),
	.w1(32'h3b3c5290),
	.w2(32'h3b2ee1d1),
	.w3(32'h3b4d7eb2),
	.w4(32'hbb597082),
	.w5(32'hbaab46c6),
	.w6(32'h3b4ccab1),
	.w7(32'h39d86224),
	.w8(32'hbade9931),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393613eb),
	.w1(32'hbb1907b5),
	.w2(32'h3a62b5b2),
	.w3(32'hbb0e9759),
	.w4(32'h3b399906),
	.w5(32'hbb6d2131),
	.w6(32'hbb873e18),
	.w7(32'h3b0ddcc3),
	.w8(32'hbb850ca7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb25e1),
	.w1(32'hbb31595d),
	.w2(32'h3ac77d5b),
	.w3(32'hb84a0dbc),
	.w4(32'h3badfe1c),
	.w5(32'hbbbf6de0),
	.w6(32'h385768dc),
	.w7(32'h3aaf570f),
	.w8(32'hbbe07cb0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb838a7c),
	.w1(32'h3b86b1ea),
	.w2(32'hbb86810f),
	.w3(32'h39d4e624),
	.w4(32'hbbeefc2e),
	.w5(32'hbae32347),
	.w6(32'h3b53420d),
	.w7(32'hbbb43bb5),
	.w8(32'hbb1a296c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb840880),
	.w1(32'hbbf6813e),
	.w2(32'hbaf58f4d),
	.w3(32'hbaf12ddd),
	.w4(32'hbba68901),
	.w5(32'hba99fec5),
	.w6(32'hbbe27232),
	.w7(32'hbbe32cb4),
	.w8(32'hba4ffc24),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34f5a0),
	.w1(32'hbb472341),
	.w2(32'hba64276a),
	.w3(32'hba8fadcd),
	.w4(32'hba13c904),
	.w5(32'hbb45fe8c),
	.w6(32'hba1c6a77),
	.w7(32'hbbded22f),
	.w8(32'hbc047dd6),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8db1f3),
	.w1(32'hbb9365b3),
	.w2(32'hbb2f0ee7),
	.w3(32'hbb08b09c),
	.w4(32'hb908dd63),
	.w5(32'hbac24d94),
	.w6(32'hbb6e2610),
	.w7(32'hbafcc433),
	.w8(32'h3b6237ef),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0cfef),
	.w1(32'h3b8050fb),
	.w2(32'hbaa810b7),
	.w3(32'hbb08efba),
	.w4(32'hbadd7683),
	.w5(32'hb925aa2b),
	.w6(32'h3b99f829),
	.w7(32'h3b71a22b),
	.w8(32'h3a532ebd),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc838c),
	.w1(32'hba06fe1c),
	.w2(32'h39e81109),
	.w3(32'hb91ae6e2),
	.w4(32'h3a5cf123),
	.w5(32'hbb3f151c),
	.w6(32'h3b2cc8ab),
	.w7(32'hba7ffc36),
	.w8(32'hbb296b8c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70dd65),
	.w1(32'hbac8ee0f),
	.w2(32'h3a9e1ab0),
	.w3(32'hba99fa4c),
	.w4(32'h3b766edb),
	.w5(32'h3aba45c5),
	.w6(32'hbb6c8b01),
	.w7(32'h3656c4e0),
	.w8(32'h37911754),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e22763),
	.w1(32'hbac145f0),
	.w2(32'h3b52944e),
	.w3(32'hba086d14),
	.w4(32'h3a8af782),
	.w5(32'h39ef3bc3),
	.w6(32'hbc001f43),
	.w7(32'hba516d9d),
	.w8(32'hb8697591),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08e039),
	.w1(32'h39083e23),
	.w2(32'h3b8cc73c),
	.w3(32'h38e0b443),
	.w4(32'h3bca569a),
	.w5(32'h3c55f9d6),
	.w6(32'hbb05b137),
	.w7(32'h3b95cbd8),
	.w8(32'h3c404795),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c498ebb),
	.w1(32'h3ad0adce),
	.w2(32'h3bad2fd5),
	.w3(32'h3adb474e),
	.w4(32'h3bca3685),
	.w5(32'hbb548e1c),
	.w6(32'h3b4fe7b4),
	.w7(32'h3b6e29bd),
	.w8(32'hbac89e08),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dc8f6),
	.w1(32'hb9828ba1),
	.w2(32'hbb152c92),
	.w3(32'h3a0804ed),
	.w4(32'hba4041c7),
	.w5(32'h3ac9245d),
	.w6(32'h3b2f2fcc),
	.w7(32'hbabfc419),
	.w8(32'h3b37775a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab92302),
	.w1(32'hbb0eb771),
	.w2(32'hba9ef063),
	.w3(32'h3ae4c6eb),
	.w4(32'hbb1f5fa1),
	.w5(32'h3b90a501),
	.w6(32'h3ac73b1c),
	.w7(32'hbb81527a),
	.w8(32'h3bc276d2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d378d),
	.w1(32'hba80e2ae),
	.w2(32'h3a5e65d9),
	.w3(32'h3b438e44),
	.w4(32'h3b941db2),
	.w5(32'hbad45985),
	.w6(32'h3b9ba54f),
	.w7(32'h3bafeae3),
	.w8(32'h3ae59a11),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb312b9d),
	.w1(32'hba782ec1),
	.w2(32'hba6561bb),
	.w3(32'hbb39454b),
	.w4(32'h3b403c34),
	.w5(32'hbb1bb6fb),
	.w6(32'hbb8f30b5),
	.w7(32'hb91e70c0),
	.w8(32'hbb9e40b8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb558311),
	.w1(32'hbb80b4cb),
	.w2(32'hb733a442),
	.w3(32'h3abb965b),
	.w4(32'h3baba662),
	.w5(32'h3b6db6b6),
	.w6(32'h3977b9ed),
	.w7(32'h3b467c1b),
	.w8(32'h3b1710c4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87d73c),
	.w1(32'h3a08cc07),
	.w2(32'h3a4f3db2),
	.w3(32'h3b30e235),
	.w4(32'h399c4df9),
	.w5(32'h3a651156),
	.w6(32'h3b6c08b4),
	.w7(32'hbb583382),
	.w8(32'h39b3b71d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ee399),
	.w1(32'h3c112781),
	.w2(32'h3bdb3c8a),
	.w3(32'hbaf263de),
	.w4(32'hba928236),
	.w5(32'hbb8b8589),
	.w6(32'h3b28cb5b),
	.w7(32'h3b96ca36),
	.w8(32'hbaf68975),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18bcf2),
	.w1(32'hbb58f92f),
	.w2(32'hbb914607),
	.w3(32'hbbb0e3b8),
	.w4(32'hbb8118db),
	.w5(32'hbb3a9c96),
	.w6(32'hbb2ae69c),
	.w7(32'hbb48ae18),
	.w8(32'hbadcdd92),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b247c2c),
	.w1(32'hbaffa56e),
	.w2(32'h3adfcdff),
	.w3(32'hbbb2df01),
	.w4(32'h3bec76da),
	.w5(32'hbb30536e),
	.w6(32'hbbb97451),
	.w7(32'h3bcc7a82),
	.w8(32'hbb7cd34f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb558dbe),
	.w1(32'hbbbd823e),
	.w2(32'hbbaa8415),
	.w3(32'hbba2f572),
	.w4(32'hbaafbd25),
	.w5(32'hbbfb4e81),
	.w6(32'hbb578e99),
	.w7(32'hbb850c65),
	.w8(32'hbb8a4c90),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a88b97),
	.w1(32'h39dca938),
	.w2(32'h39154280),
	.w3(32'hb9c22133),
	.w4(32'h3af027bf),
	.w5(32'hbbd6b9b0),
	.w6(32'h3804bb56),
	.w7(32'hba035bf4),
	.w8(32'hbb6b7cc7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb890db7),
	.w1(32'hbbae69a5),
	.w2(32'hbb924777),
	.w3(32'h3bb8f82e),
	.w4(32'h3b123e27),
	.w5(32'hb9c9b14e),
	.w6(32'h3c59dc7a),
	.w7(32'h3b974270),
	.w8(32'h3b970f34),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ac8a1),
	.w1(32'hbc506800),
	.w2(32'hbc3a86c1),
	.w3(32'hbc06742d),
	.w4(32'hbb1897e4),
	.w5(32'hbb483dd9),
	.w6(32'hbbce02b5),
	.w7(32'hbc62afad),
	.w8(32'hbb971fb0),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ea182),
	.w1(32'hbb22e50c),
	.w2(32'hbbb7b30a),
	.w3(32'h3ba198f1),
	.w4(32'hbba2c3d5),
	.w5(32'h3a505d7b),
	.w6(32'h3bce8ebb),
	.w7(32'hbbb9d293),
	.w8(32'h3ae8f978),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acafe6e),
	.w1(32'hbb9897ff),
	.w2(32'hbc0835bb),
	.w3(32'hbb73daab),
	.w4(32'h3903a35a),
	.w5(32'hbaa419b6),
	.w6(32'hbc13c44f),
	.w7(32'hbc3df26d),
	.w8(32'hba97a76b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5f919),
	.w1(32'hb995f355),
	.w2(32'hba339077),
	.w3(32'h39c68970),
	.w4(32'h3b4073cb),
	.w5(32'h3ae3327f),
	.w6(32'hbb5f6233),
	.w7(32'h39f55400),
	.w8(32'h389be81a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba609395),
	.w1(32'hbb6aa351),
	.w2(32'hbbb3adc8),
	.w3(32'h39371a58),
	.w4(32'hb98f1989),
	.w5(32'h3b814e85),
	.w6(32'hbbe59ce4),
	.w7(32'hbbfbcb8a),
	.w8(32'h3acb467e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba657314),
	.w1(32'hbb1d689f),
	.w2(32'h3b245034),
	.w3(32'hba16d094),
	.w4(32'h3b65f7ba),
	.w5(32'h3bb7ea86),
	.w6(32'hbb3d458c),
	.w7(32'h3b178b83),
	.w8(32'hba8eeb4a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule