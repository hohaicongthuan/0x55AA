module layer_10_featuremap_142(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a45e64),
	.w1(32'hbb7faf2a),
	.w2(32'hbb084b18),
	.w3(32'hb7763661),
	.w4(32'hb8aae1b6),
	.w5(32'hba14e92b),
	.w6(32'hbafc4834),
	.w7(32'hb97742a5),
	.w8(32'h3a8e07e7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01a6d8),
	.w1(32'hbbafc1c9),
	.w2(32'hbb451f7f),
	.w3(32'h3aad613b),
	.w4(32'hbb661f1f),
	.w5(32'hba67bb2d),
	.w6(32'hbb1a5b32),
	.w7(32'hba84fef0),
	.w8(32'hba4e31c7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b334b),
	.w1(32'h39cb6484),
	.w2(32'h3a5e31ff),
	.w3(32'hba8bbde8),
	.w4(32'h399e6b4c),
	.w5(32'h3a4c0853),
	.w6(32'h39b5d077),
	.w7(32'h3ab2d561),
	.w8(32'h3a81b6af),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab470d9),
	.w1(32'h39055282),
	.w2(32'h399687d2),
	.w3(32'h3a85002c),
	.w4(32'hbafe5e5f),
	.w5(32'hba39e757),
	.w6(32'h36130c3a),
	.w7(32'h3a7bee72),
	.w8(32'h3a8b8bc4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed7789),
	.w1(32'hba2063a8),
	.w2(32'h3ab7cb2d),
	.w3(32'h3b005d50),
	.w4(32'h3ab6bfc6),
	.w5(32'h3b2c42d8),
	.w6(32'hbaeb2a18),
	.w7(32'hba83a1f3),
	.w8(32'hbb16a363),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a43016),
	.w1(32'h38203498),
	.w2(32'h3a5eb8cb),
	.w3(32'h3acf6200),
	.w4(32'hb9e8ff93),
	.w5(32'h3a4be9c4),
	.w6(32'hbb047666),
	.w7(32'hba46b2d2),
	.w8(32'hba11fb8b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28dcc2),
	.w1(32'h3b0eec4d),
	.w2(32'h3a20cab8),
	.w3(32'h39a29d9c),
	.w4(32'h3a8673f3),
	.w5(32'h39d7ef4f),
	.w6(32'h3a818e72),
	.w7(32'h3b01a4ef),
	.w8(32'hb9fc7fc7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa2631),
	.w1(32'h3b6b07ba),
	.w2(32'h39d2831a),
	.w3(32'h3ba142b1),
	.w4(32'h3b35a3f1),
	.w5(32'hbaf02fe3),
	.w6(32'h3ba33f81),
	.w7(32'h3b1bc4c9),
	.w8(32'hb9c32299),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384e7868),
	.w1(32'h398dac21),
	.w2(32'hb97ee9da),
	.w3(32'h348681cd),
	.w4(32'h39b39dd9),
	.w5(32'h3a97995d),
	.w6(32'hb8037986),
	.w7(32'h39369c97),
	.w8(32'hbabc2ff0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0d2f4),
	.w1(32'hba01d7cc),
	.w2(32'hba96dc20),
	.w3(32'hbb56d22a),
	.w4(32'hbb1e4b72),
	.w5(32'hbb01f2f7),
	.w6(32'hba120510),
	.w7(32'h3b34b5c3),
	.w8(32'h3ae093e3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba625653),
	.w1(32'h3b500339),
	.w2(32'h3ba3c0a1),
	.w3(32'hbabb03d3),
	.w4(32'hbb1d949a),
	.w5(32'hbb1b5d1a),
	.w6(32'hb82e4b06),
	.w7(32'h3a68b892),
	.w8(32'hb9afb3ea),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd78e4e),
	.w1(32'h3b820e44),
	.w2(32'h3b8b49ce),
	.w3(32'h3b2f4493),
	.w4(32'h3ba67c68),
	.w5(32'h3b8c1b79),
	.w6(32'h3affb532),
	.w7(32'h3b00ad50),
	.w8(32'h3b6fecef),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11d068),
	.w1(32'h3b1605f5),
	.w2(32'h37d92e5c),
	.w3(32'h3b77159b),
	.w4(32'hb8541051),
	.w5(32'hba981dbe),
	.w6(32'h3a0fe054),
	.w7(32'h3bb2cb8a),
	.w8(32'h3b1db383),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83b4fc8),
	.w1(32'hba46b37e),
	.w2(32'hbb3c04d0),
	.w3(32'hba3ab8a1),
	.w4(32'h397aba37),
	.w5(32'hbb1e386f),
	.w6(32'h3b364823),
	.w7(32'hba3b5e52),
	.w8(32'h3a9197b0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e4265),
	.w1(32'hbb4936a4),
	.w2(32'h3a6401e2),
	.w3(32'h39ca0ba3),
	.w4(32'hbb1d5ced),
	.w5(32'h3a4f3f38),
	.w6(32'hb94ffba6),
	.w7(32'h3a42e012),
	.w8(32'hb6c2fe5f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1abfaa),
	.w1(32'h39c9a34e),
	.w2(32'hb726137a),
	.w3(32'h3b12ad7f),
	.w4(32'h39104467),
	.w5(32'h39a7a897),
	.w6(32'h3a9e6aa1),
	.w7(32'h3b3956ea),
	.w8(32'h3a9bcd4a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3912e38c),
	.w1(32'hbb2a02aa),
	.w2(32'h3b6ab047),
	.w3(32'h3a813cd3),
	.w4(32'h38cef319),
	.w5(32'h3b83cb2f),
	.w6(32'hbbf7866f),
	.w7(32'h39368ccc),
	.w8(32'hbba4e782),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67037b),
	.w1(32'h3c623a2c),
	.w2(32'h3c3908b4),
	.w3(32'h3c43d7c8),
	.w4(32'h3c4d841f),
	.w5(32'h3a9b86c8),
	.w6(32'h3c2e587f),
	.w7(32'h3bfcb4f5),
	.w8(32'hbaae0920),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b739a9b),
	.w1(32'h3bb2b7be),
	.w2(32'h3b4fed9d),
	.w3(32'h3b419fd9),
	.w4(32'h3b823cae),
	.w5(32'h3ab40cf6),
	.w6(32'h3b7dfb9a),
	.w7(32'h3b9409f1),
	.w8(32'hba774fc0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9945ec2),
	.w1(32'hba02220b),
	.w2(32'hba21c6b9),
	.w3(32'hb9b1f77a),
	.w4(32'hb99d38d6),
	.w5(32'hba0efd8c),
	.w6(32'hb9b62b6b),
	.w7(32'h3a321d3b),
	.w8(32'hba98f75e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48a44b),
	.w1(32'h3b82bf10),
	.w2(32'hba83e5ed),
	.w3(32'hb9db2785),
	.w4(32'h3993a118),
	.w5(32'hbb0f5615),
	.w6(32'h3a891573),
	.w7(32'hb9c7d60c),
	.w8(32'hba37d428),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ab087),
	.w1(32'hbb7a551a),
	.w2(32'hba3f7e81),
	.w3(32'hbafa5167),
	.w4(32'hbb80a6b4),
	.w5(32'hbb9b71c7),
	.w6(32'hba19e000),
	.w7(32'h3b0eae22),
	.w8(32'h3b2fac25),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9eada3),
	.w1(32'h3cc9865e),
	.w2(32'h3c621582),
	.w3(32'h3c98c6ed),
	.w4(32'h3c2aabff),
	.w5(32'h3aa5900c),
	.w6(32'h3c53ed9b),
	.w7(32'h3bf5959c),
	.w8(32'hbbe16571),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becec0d),
	.w1(32'hba1bcd16),
	.w2(32'hbb7befb4),
	.w3(32'hbc14c5ba),
	.w4(32'hbb176297),
	.w5(32'hbb2f91e9),
	.w6(32'hb9da4f96),
	.w7(32'h3aa265a8),
	.w8(32'h3ad623db),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fafbe),
	.w1(32'hbb660f14),
	.w2(32'hbb2fae72),
	.w3(32'hbb960a45),
	.w4(32'hbba7ec76),
	.w5(32'hbb0875d7),
	.w6(32'hbb58026f),
	.w7(32'h3a033e30),
	.w8(32'h3a9ad4fa),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabecfd),
	.w1(32'hbb4b418c),
	.w2(32'hbae9aa6d),
	.w3(32'hbb01ce93),
	.w4(32'hbba56548),
	.w5(32'hbb70aa74),
	.w6(32'hbbc560ed),
	.w7(32'hbaac5903),
	.w8(32'hbad330df),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1582c6),
	.w1(32'hba280e4c),
	.w2(32'hba886e3c),
	.w3(32'hbba7e64b),
	.w4(32'hba7e2087),
	.w5(32'hbac648b5),
	.w6(32'hba4497ba),
	.w7(32'hb7ca2823),
	.w8(32'hbae1355c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cae2e),
	.w1(32'hba9e4004),
	.w2(32'h3b624d6e),
	.w3(32'hbb7a7fd1),
	.w4(32'hbb27bbb5),
	.w5(32'h3b255571),
	.w6(32'hbb5ea832),
	.w7(32'h38bff9d8),
	.w8(32'h3b6e8b61),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec7e9e),
	.w1(32'h3ba2e657),
	.w2(32'h3c3ad081),
	.w3(32'hbb164f5a),
	.w4(32'hbadea890),
	.w5(32'h3bc2de43),
	.w6(32'hbb8cc085),
	.w7(32'h3be88a0d),
	.w8(32'hbbd28c57),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39246dd8),
	.w1(32'hbabbc50b),
	.w2(32'hbbafa2fa),
	.w3(32'hbc330c77),
	.w4(32'h3b41ccd0),
	.w5(32'h3962e64c),
	.w6(32'hbb2d4b72),
	.w7(32'hba6975f7),
	.w8(32'hbb2fcf8e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7cec0),
	.w1(32'h3af9aa51),
	.w2(32'h38acb850),
	.w3(32'hbbad96dc),
	.w4(32'hb94c7eea),
	.w5(32'hba825b13),
	.w6(32'h39160cf6),
	.w7(32'hb91f76d5),
	.w8(32'hba8718c8),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394bb031),
	.w1(32'h3ab1a9b3),
	.w2(32'h3a78c62e),
	.w3(32'hba953e6c),
	.w4(32'hba303379),
	.w5(32'hba63e34a),
	.w6(32'hb9eba391),
	.w7(32'h3a0719f5),
	.w8(32'hba3d6c24),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dd0b1),
	.w1(32'hbabcb9a6),
	.w2(32'hba857cb6),
	.w3(32'hb7fea8c4),
	.w4(32'h3919ac2f),
	.w5(32'hb9699600),
	.w6(32'h3a9bee21),
	.w7(32'h3aeae65f),
	.w8(32'hbb029d90),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef3f91),
	.w1(32'hbc045298),
	.w2(32'h37bda24b),
	.w3(32'hba996f19),
	.w4(32'hbbf2415c),
	.w5(32'h3bdca279),
	.w6(32'hbbb42b6b),
	.w7(32'h3bbe20e8),
	.w8(32'hbc039954),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66eccc),
	.w1(32'hb9e9692c),
	.w2(32'h3b18d753),
	.w3(32'hbabce72a),
	.w4(32'hbae83c45),
	.w5(32'hb9a84e4e),
	.w6(32'hbac28311),
	.w7(32'h39bf5995),
	.w8(32'hba370aa4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f7a02),
	.w1(32'h3b84fc0a),
	.w2(32'h3a19ba45),
	.w3(32'hbac076fc),
	.w4(32'h3abaa5b8),
	.w5(32'hbaa6c9ae),
	.w6(32'h3abd46d7),
	.w7(32'h3b1fb220),
	.w8(32'hba32d716),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdac515),
	.w1(32'h3b2c3b09),
	.w2(32'h3b020a90),
	.w3(32'h3bcb3b39),
	.w4(32'h3a495e61),
	.w5(32'hba33bcf7),
	.w6(32'h3b8fbb90),
	.w7(32'h3b2d70b9),
	.w8(32'hbac5fe5b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f8c9c),
	.w1(32'hbc2b88ba),
	.w2(32'hbb892687),
	.w3(32'hbc53017a),
	.w4(32'hbc03ea9d),
	.w5(32'h3a40b5ec),
	.w6(32'hbc4efefc),
	.w7(32'hbb144202),
	.w8(32'h3a88a5b7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedb8d6),
	.w1(32'hbc034945),
	.w2(32'hbaff6241),
	.w3(32'hbc15590b),
	.w4(32'hbbdcd48b),
	.w5(32'h3b3162be),
	.w6(32'hbc10e184),
	.w7(32'hbb9671c7),
	.w8(32'h3aa73c6f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0150d),
	.w1(32'hba80032a),
	.w2(32'h390ad658),
	.w3(32'hbab30b62),
	.w4(32'hba62235e),
	.w5(32'h3a212d66),
	.w6(32'hbaf05b3f),
	.w7(32'hba0767ff),
	.w8(32'hb971c7b9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6fa20),
	.w1(32'h3b2108cb),
	.w2(32'hba86ee22),
	.w3(32'hb88cdd1e),
	.w4(32'h3b9fbbb2),
	.w5(32'hba0e1b76),
	.w6(32'h3bc456f3),
	.w7(32'h3bd9aa91),
	.w8(32'hbb19881b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3449fb),
	.w1(32'h36e391f9),
	.w2(32'h3a819bb5),
	.w3(32'hbc46971f),
	.w4(32'h3a0b1463),
	.w5(32'h3a4769dc),
	.w6(32'h3a2ab220),
	.w7(32'h3a70094b),
	.w8(32'h3a42f837),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0947d5),
	.w1(32'h3aaa48bf),
	.w2(32'h3a1354d0),
	.w3(32'h3a82db9d),
	.w4(32'hba4d6ad8),
	.w5(32'hbb108f91),
	.w6(32'hbaa7a140),
	.w7(32'h350a4a1e),
	.w8(32'hba967b45),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cd330),
	.w1(32'hb9846ea6),
	.w2(32'hbb1ec90b),
	.w3(32'hba689ab3),
	.w4(32'h3a9b38ad),
	.w5(32'hba5ac7ed),
	.w6(32'h3afd9609),
	.w7(32'h3b533aff),
	.w8(32'hb9442f55),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbec0c),
	.w1(32'hb9c9075a),
	.w2(32'hbb70af2f),
	.w3(32'hbb2f7b57),
	.w4(32'hb9f60492),
	.w5(32'hba88532b),
	.w6(32'hbaaaae99),
	.w7(32'h3b071202),
	.w8(32'h3b38d432),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a96f0),
	.w1(32'hba7081e2),
	.w2(32'hbbb619c0),
	.w3(32'hbb08487f),
	.w4(32'hbad40c30),
	.w5(32'hbb79dd63),
	.w6(32'hb9f4be5e),
	.w7(32'h3b26f141),
	.w8(32'h3aa5d094),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27d22f),
	.w1(32'h3a377c62),
	.w2(32'h3ac4eb04),
	.w3(32'h39c414dd),
	.w4(32'hb8a9858d),
	.w5(32'hb9dfe14d),
	.w6(32'h3b924bd4),
	.w7(32'h3ad61913),
	.w8(32'hba611375),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f42cd),
	.w1(32'h3cbc2fe8),
	.w2(32'h3cf0770d),
	.w3(32'h3c9acc48),
	.w4(32'h3c3cb9ab),
	.w5(32'h3c7c7d99),
	.w6(32'h3c184375),
	.w7(32'h3ca71360),
	.w8(32'hbbf67af0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9d0af),
	.w1(32'hb8a80ed6),
	.w2(32'hbac5dee7),
	.w3(32'hbb7dc557),
	.w4(32'hba90daa3),
	.w5(32'hbb34f469),
	.w6(32'hbaa39bb5),
	.w7(32'h39b83e01),
	.w8(32'hbae6bd14),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f19e98),
	.w1(32'hba2cac6f),
	.w2(32'hbab4ab7c),
	.w3(32'hbadb1c39),
	.w4(32'h38f3897f),
	.w5(32'hb98194fd),
	.w6(32'hb96dd9b3),
	.w7(32'hbaa7b2c1),
	.w8(32'hb8c34f7c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b37b60),
	.w1(32'hb955ec63),
	.w2(32'h3a53fdfc),
	.w3(32'h39f682e1),
	.w4(32'hba4daeb7),
	.w5(32'hb937ec9c),
	.w6(32'h3b07dc06),
	.w7(32'h3b160ec9),
	.w8(32'h3b083044),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8031d6),
	.w1(32'h3a088274),
	.w2(32'h3b95d849),
	.w3(32'h3a8cc7b5),
	.w4(32'h3a037245),
	.w5(32'h3b0ebe4d),
	.w6(32'h3af039b1),
	.w7(32'hbae6e3e2),
	.w8(32'h3b3455a5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccb6ec),
	.w1(32'h3b22bce2),
	.w2(32'h3ae976fc),
	.w3(32'h3b911634),
	.w4(32'h3a75bfaf),
	.w5(32'hb7c80257),
	.w6(32'h3b0f712d),
	.w7(32'h3b3d5717),
	.w8(32'hb9aebdc6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ff086),
	.w1(32'h3c203bf4),
	.w2(32'h3bb7399f),
	.w3(32'h3c099bd0),
	.w4(32'h3bec13a7),
	.w5(32'hba873f6d),
	.w6(32'h3bfd4954),
	.w7(32'h3ba33d2f),
	.w8(32'hbb656f0b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab10a46),
	.w1(32'hb9f40fb4),
	.w2(32'h3adfa9ea),
	.w3(32'h3b341268),
	.w4(32'hbafffb3a),
	.w5(32'hb997b467),
	.w6(32'hbb41d547),
	.w7(32'h3a82ba89),
	.w8(32'hbaa73594),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4a7c8),
	.w1(32'h3b89105d),
	.w2(32'hbbedc8b3),
	.w3(32'hbb6867f3),
	.w4(32'h3b9c49f0),
	.w5(32'hbbd68e52),
	.w6(32'h3c5bce0d),
	.w7(32'h3ad36f0f),
	.w8(32'h3a0aad76),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dd438),
	.w1(32'h3a45a8ea),
	.w2(32'h3a86a15c),
	.w3(32'hbc283677),
	.w4(32'hba2e6200),
	.w5(32'hba5a6b9b),
	.w6(32'h3a5a1165),
	.w7(32'h3b89ba17),
	.w8(32'hba97d673),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a5ea7),
	.w1(32'hbb345194),
	.w2(32'h3a4dd8a9),
	.w3(32'hbba9a462),
	.w4(32'hb829a375),
	.w5(32'h3b17e06e),
	.w6(32'hba794ac7),
	.w7(32'h39c83988),
	.w8(32'h3a499e00),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15595d),
	.w1(32'h3a14841d),
	.w2(32'h3a8604de),
	.w3(32'h3a5bf8f2),
	.w4(32'h39b06f91),
	.w5(32'h3abf2e2f),
	.w6(32'hba6d8ecb),
	.w7(32'h39ce435e),
	.w8(32'h3aa8e1c2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a000c0c),
	.w1(32'h39b768aa),
	.w2(32'hb96e6496),
	.w3(32'h37afa9f5),
	.w4(32'h39cb2306),
	.w5(32'h3983625b),
	.w6(32'h393fa821),
	.w7(32'hb935cea5),
	.w8(32'h38f287aa),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84dfb1),
	.w1(32'h3bc3c2c8),
	.w2(32'h3b736cb6),
	.w3(32'h3b8f916f),
	.w4(32'h3b81edbe),
	.w5(32'h3ac712ce),
	.w6(32'h3b14a459),
	.w7(32'h3b5a7f3d),
	.w8(32'h3a95e53e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2a85b),
	.w1(32'h3b883448),
	.w2(32'h3b258de9),
	.w3(32'h3ba3930e),
	.w4(32'h3b37a6ab),
	.w5(32'hb89c6f23),
	.w6(32'h3b5b7829),
	.w7(32'hbaa1abec),
	.w8(32'hb95777d1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a532359),
	.w1(32'hbaeef6af),
	.w2(32'hba4b205c),
	.w3(32'h3a1a6b51),
	.w4(32'hba989c84),
	.w5(32'hbb04a588),
	.w6(32'hb86caa68),
	.w7(32'h3983c830),
	.w8(32'hb7622f54),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba533e06),
	.w1(32'hb9a74c34),
	.w2(32'h3a331a88),
	.w3(32'hba77a20b),
	.w4(32'h3a9990e3),
	.w5(32'h3b0c8cd8),
	.w6(32'h39cced50),
	.w7(32'h3a52522c),
	.w8(32'h3a5f0a53),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ffb62),
	.w1(32'hb92c4b69),
	.w2(32'hb9e872e2),
	.w3(32'h39bee130),
	.w4(32'h3a004dc0),
	.w5(32'h39e9c1a3),
	.w6(32'hb98e0b51),
	.w7(32'h3a082322),
	.w8(32'hb9a8ad75),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381a6266),
	.w1(32'hbb37b4be),
	.w2(32'hba87478c),
	.w3(32'hb978bbbb),
	.w4(32'hb9d90bd6),
	.w5(32'h3b1c9688),
	.w6(32'hbae18ace),
	.w7(32'h39aaf555),
	.w8(32'h390335a9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a39fb),
	.w1(32'h3bea3944),
	.w2(32'h3972c22a),
	.w3(32'h3b20fc62),
	.w4(32'h3c2b34f8),
	.w5(32'h39daecb2),
	.w6(32'h3c584d02),
	.w7(32'h3b9ffd4b),
	.w8(32'hbb14cd96),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e7f93),
	.w1(32'h3bfb7aa0),
	.w2(32'h3c29872a),
	.w3(32'hbbf77c0a),
	.w4(32'hba50ea31),
	.w5(32'h3bd9371a),
	.w6(32'h3a6c5c76),
	.w7(32'h3c7ee109),
	.w8(32'h3ae8b948),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72b0ac),
	.w1(32'h3c05bd97),
	.w2(32'h3b960685),
	.w3(32'h3b35b4b7),
	.w4(32'h3b393933),
	.w5(32'hb888834a),
	.w6(32'h3bbe1032),
	.w7(32'h3b0f3d6b),
	.w8(32'h3a4d24e3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf65162),
	.w1(32'hbb7c0c5d),
	.w2(32'hbb9ef038),
	.w3(32'hbb92c6f2),
	.w4(32'hba63261a),
	.w5(32'h39d8b808),
	.w6(32'hb9f854c0),
	.w7(32'h3a0384dc),
	.w8(32'h3c051725),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9468a2),
	.w1(32'hba00b039),
	.w2(32'hb947fc5d),
	.w3(32'h37e8a028),
	.w4(32'hb90bb4ed),
	.w5(32'h39ad1fcd),
	.w6(32'hba49836b),
	.w7(32'h3a41aeaf),
	.w8(32'hb9a13ff5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94108bc),
	.w1(32'h3a91f6e6),
	.w2(32'h3a008a65),
	.w3(32'hba5aa84d),
	.w4(32'h3a269225),
	.w5(32'h3a05b2c8),
	.w6(32'h3a1454ac),
	.w7(32'h3a3f20f1),
	.w8(32'h388dd038),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a2b413),
	.w1(32'h39a7461a),
	.w2(32'hb96216ad),
	.w3(32'hba280fc9),
	.w4(32'h3a006135),
	.w5(32'h3a3999f5),
	.w6(32'h3986ef3b),
	.w7(32'h3945c2f8),
	.w8(32'h3752b6f7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0941ff),
	.w1(32'h3bc989f8),
	.w2(32'h3b5851f1),
	.w3(32'h3b17717e),
	.w4(32'h3aaa8730),
	.w5(32'hba03234d),
	.w6(32'h3adac695),
	.w7(32'h3b332796),
	.w8(32'hba824b59),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd805e),
	.w1(32'h398e42d7),
	.w2(32'h3af35178),
	.w3(32'hb9b8b631),
	.w4(32'h3a746150),
	.w5(32'h3ac46881),
	.w6(32'hb977f2dd),
	.w7(32'h3a3e84ad),
	.w8(32'h39ad71c4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7ebeb),
	.w1(32'h3b84adbb),
	.w2(32'h3a976a5c),
	.w3(32'h3bfe61f4),
	.w4(32'h3b988332),
	.w5(32'hbb00c8ee),
	.w6(32'h3c0e60ba),
	.w7(32'h3b822153),
	.w8(32'hba3ad8f2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f0769),
	.w1(32'h3c2703cd),
	.w2(32'h3bc7cc95),
	.w3(32'h3c58c374),
	.w4(32'h3c4fcc3e),
	.w5(32'h3b57fb02),
	.w6(32'h3c300b66),
	.w7(32'h3c04eabe),
	.w8(32'h3acd922d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb919af8),
	.w1(32'hbb10f95d),
	.w2(32'h3a4fc35a),
	.w3(32'hbbb750ea),
	.w4(32'hbadac4dc),
	.w5(32'h3b316de0),
	.w6(32'hbb8dc5de),
	.w7(32'h3b0478eb),
	.w8(32'h3b31b20a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd9114),
	.w1(32'hb6b993b8),
	.w2(32'h3ab6644c),
	.w3(32'h3aabd9d9),
	.w4(32'hbb0b84fe),
	.w5(32'hbb10d941),
	.w6(32'hbb99439d),
	.w7(32'h3ac50038),
	.w8(32'hbb631196),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24995d),
	.w1(32'h3b839f3f),
	.w2(32'hb9d488e5),
	.w3(32'hbb229738),
	.w4(32'h3a32d6b4),
	.w5(32'hbacc9a92),
	.w6(32'h3a9d2e85),
	.w7(32'h3acfd511),
	.w8(32'hbacc962a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c1b36),
	.w1(32'h3c3fee1b),
	.w2(32'h3c698352),
	.w3(32'hbaf1b52c),
	.w4(32'hb9e3df47),
	.w5(32'h3bccb1aa),
	.w6(32'h3b9e48c1),
	.w7(32'h3c644a12),
	.w8(32'hba9c9807),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c147eaf),
	.w1(32'h3bfeb9cc),
	.w2(32'h3baa45b0),
	.w3(32'hbb67f87a),
	.w4(32'h3baf9016),
	.w5(32'h3a3e4b8e),
	.w6(32'h3b73e436),
	.w7(32'h3b767fc5),
	.w8(32'hba806eee),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38486f71),
	.w1(32'h3b25e24f),
	.w2(32'h3b128c29),
	.w3(32'hb9c88507),
	.w4(32'h39b22ae1),
	.w5(32'h38ce1e32),
	.w6(32'h3a16e3a8),
	.w7(32'h3a87b94b),
	.w8(32'hbaaaf4ad),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d43af),
	.w1(32'hb9dd6d35),
	.w2(32'hba23d155),
	.w3(32'hbae7dc9d),
	.w4(32'hb920ea5e),
	.w5(32'hb7f03f9f),
	.w6(32'hba7f23cf),
	.w7(32'h390fef77),
	.w8(32'hb93d9b53),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbf476),
	.w1(32'h3c2b13bb),
	.w2(32'h3cd0028e),
	.w3(32'hba649116),
	.w4(32'hbc2a10aa),
	.w5(32'h3c731a16),
	.w6(32'hbc035aff),
	.w7(32'h3c8ce41e),
	.w8(32'hbc1dd3c4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7bacd8),
	.w1(32'hba366f52),
	.w2(32'hba5c5d75),
	.w3(32'hbb42e139),
	.w4(32'h3a65ad6b),
	.w5(32'hb94bb707),
	.w6(32'hb9d7c47b),
	.w7(32'hb62c8dbf),
	.w8(32'hba0c8ca5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8860ac),
	.w1(32'hbb9a1449),
	.w2(32'hbb72d0d9),
	.w3(32'hbbd0a28b),
	.w4(32'hbb5416d6),
	.w5(32'hba368f3b),
	.w6(32'hbaede120),
	.w7(32'hba51ad28),
	.w8(32'h3af05f7d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07a6b9),
	.w1(32'h3b098b83),
	.w2(32'h3a126856),
	.w3(32'h3b2328d9),
	.w4(32'h37344ecb),
	.w5(32'hba4824a2),
	.w6(32'h38762e11),
	.w7(32'h3832aa71),
	.w8(32'hba54dfd8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b469319),
	.w1(32'hba187a15),
	.w2(32'hbaf59d61),
	.w3(32'hbacf6bf2),
	.w4(32'hbb44fef3),
	.w5(32'hbb43ae50),
	.w6(32'h385f82b2),
	.w7(32'h3b32bbd0),
	.w8(32'hbafaa089),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd8e5e),
	.w1(32'h3c0a2487),
	.w2(32'h3a996f73),
	.w3(32'h3c1a4919),
	.w4(32'h3b9d5a72),
	.w5(32'hbc0032e4),
	.w6(32'h3c447782),
	.w7(32'h3b01fe65),
	.w8(32'hbbf50f79),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb055563),
	.w1(32'h3b0a007c),
	.w2(32'h3b96baa9),
	.w3(32'hbb739ffc),
	.w4(32'hba77e93e),
	.w5(32'h396b2c31),
	.w6(32'hba7de2a3),
	.w7(32'hba5bdd1c),
	.w8(32'hb95e6cdf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfec29),
	.w1(32'h3b417c7e),
	.w2(32'h3ae8d518),
	.w3(32'h3b829841),
	.w4(32'h3b4982ba),
	.w5(32'hb860114e),
	.w6(32'h3b2ff171),
	.w7(32'h3b564e98),
	.w8(32'h3a8b72e8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393827b5),
	.w1(32'hba176268),
	.w2(32'hbafaeae3),
	.w3(32'hbadf7fee),
	.w4(32'hbab7dc63),
	.w5(32'hbae68f29),
	.w6(32'hbb05be4d),
	.w7(32'h3a06b2cf),
	.w8(32'hbb06d500),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a959d1f),
	.w1(32'h3c23e3c8),
	.w2(32'h3c2eb6a6),
	.w3(32'hbb0de71a),
	.w4(32'hba8331d8),
	.w5(32'h3a458a1d),
	.w6(32'h3beb5f20),
	.w7(32'h3c389c0b),
	.w8(32'hbb56cfb2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32cbb2),
	.w1(32'hba9d1486),
	.w2(32'hba4cd293),
	.w3(32'hbc3be1fb),
	.w4(32'hbb7482b4),
	.w5(32'hbb65956d),
	.w6(32'hba100a52),
	.w7(32'h3a705c9b),
	.w8(32'hba8660b3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba497448),
	.w1(32'hbb09ca58),
	.w2(32'hbb104b8b),
	.w3(32'hbb4a3f09),
	.w4(32'hbb2a7e51),
	.w5(32'h39ffc25e),
	.w6(32'hbb85ba7c),
	.w7(32'hbb30b453),
	.w8(32'hbaf498fd),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39924703),
	.w1(32'hbb88d24b),
	.w2(32'hbada67d5),
	.w3(32'hba02ecb4),
	.w4(32'hba769977),
	.w5(32'h3b283d48),
	.w6(32'hbb4a713d),
	.w7(32'h3b5c5e11),
	.w8(32'hbb4354a1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5b17f),
	.w1(32'hba89e4ed),
	.w2(32'hbb72c275),
	.w3(32'hbb5bed2b),
	.w4(32'h38db1c2b),
	.w5(32'hbb4c606a),
	.w6(32'hb9fbaaba),
	.w7(32'h3a0ba0b7),
	.w8(32'hbb29031f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f5948),
	.w1(32'h3a8a64a5),
	.w2(32'h3b37ee3e),
	.w3(32'h3b5ebfd8),
	.w4(32'hba158a54),
	.w5(32'h39ce7d55),
	.w6(32'h3aa4b1ba),
	.w7(32'h3a851241),
	.w8(32'hb8a02104),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2aedc3),
	.w1(32'h3c4182b3),
	.w2(32'h3c24631c),
	.w3(32'h3c7411ee),
	.w4(32'h3c39530f),
	.w5(32'h3a7e16ff),
	.w6(32'h3c6de93b),
	.w7(32'h3c315942),
	.w8(32'hba97e666),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef4b50),
	.w1(32'hbb8fa3d4),
	.w2(32'hbbb649f7),
	.w3(32'hbc3a914b),
	.w4(32'hbbb01bee),
	.w5(32'hba90d6e6),
	.w6(32'hbc422db9),
	.w7(32'hbbc266dc),
	.w8(32'hbb60ed60),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a38a1),
	.w1(32'hbb4c9685),
	.w2(32'hbb4c90c3),
	.w3(32'hbbaf311c),
	.w4(32'hbb066e6e),
	.w5(32'hbb3fe52e),
	.w6(32'hbbae4038),
	.w7(32'hb8fe8cf8),
	.w8(32'h3afaf038),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdae8dc),
	.w1(32'h3bbe52a4),
	.w2(32'h3a826eb9),
	.w3(32'h3bb737c1),
	.w4(32'h3b7a76dd),
	.w5(32'hb9fa5cdc),
	.w6(32'h3ba12faf),
	.w7(32'h3a5f131e),
	.w8(32'hbb0307f4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00d457),
	.w1(32'h38447176),
	.w2(32'hb9ad9446),
	.w3(32'hba068184),
	.w4(32'h378fcf4e),
	.w5(32'h3928e5eb),
	.w6(32'hb99f86d5),
	.w7(32'h3913f71c),
	.w8(32'hba592486),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c593d29),
	.w1(32'h3cbba76d),
	.w2(32'h3c6373f9),
	.w3(32'h3c67e0db),
	.w4(32'h3c902ef2),
	.w5(32'h3c079f74),
	.w6(32'h3c8a273e),
	.w7(32'h3c203669),
	.w8(32'h3a90b043),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46b0ff),
	.w1(32'hb9bbccfc),
	.w2(32'h3b6f2e98),
	.w3(32'hbb1af245),
	.w4(32'hba147428),
	.w5(32'h3bd23651),
	.w6(32'hba852658),
	.w7(32'h3a9e5ff1),
	.w8(32'h3bb85dbc),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba823c33),
	.w1(32'h3a426498),
	.w2(32'h3b1afa92),
	.w3(32'hba746a75),
	.w4(32'hb9938ce6),
	.w5(32'h3a359521),
	.w6(32'hba09aeaa),
	.w7(32'h3ab7aa14),
	.w8(32'h3a57d55e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14ef8b),
	.w1(32'h3b82f81a),
	.w2(32'h393dadfc),
	.w3(32'h3a79446c),
	.w4(32'hba60a5e1),
	.w5(32'hbb49a4d0),
	.w6(32'h399c54c2),
	.w7(32'hba532534),
	.w8(32'hbb269bd4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32e362),
	.w1(32'hbb6b591a),
	.w2(32'hbb89810c),
	.w3(32'hbb9ba385),
	.w4(32'hbb494472),
	.w5(32'hbb2936f4),
	.w6(32'hbb28db8a),
	.w7(32'hbb20e9ce),
	.w8(32'hba9ca180),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3f3c1),
	.w1(32'hbb18d421),
	.w2(32'hbb0cc9c0),
	.w3(32'hbb8abd00),
	.w4(32'hbae295cd),
	.w5(32'hbaccfd14),
	.w6(32'hbb0b8056),
	.w7(32'h3b5b9a07),
	.w8(32'h3b931855),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc8582),
	.w1(32'hb9b9e5c0),
	.w2(32'hba2a75de),
	.w3(32'h3a4a940b),
	.w4(32'hbb1148d7),
	.w5(32'h38992edb),
	.w6(32'hba2bbd5e),
	.w7(32'hba885dd2),
	.w8(32'hba9c8faf),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42b1a5),
	.w1(32'hbb11976b),
	.w2(32'hbb7287e3),
	.w3(32'h3b00464d),
	.w4(32'hb92040fc),
	.w5(32'hb9a2925c),
	.w6(32'h3b0e2e24),
	.w7(32'hba0452ed),
	.w8(32'h3961edd6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbffea3),
	.w1(32'h3b096f12),
	.w2(32'h3b3d8c86),
	.w3(32'h3bc60e5d),
	.w4(32'h3acfadda),
	.w5(32'h3b16a3c6),
	.w6(32'hba10e6c9),
	.w7(32'h3ac6d910),
	.w8(32'h3a1eaa3e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a6964),
	.w1(32'h3b5a6d23),
	.w2(32'h3b13b39c),
	.w3(32'h3b3ee476),
	.w4(32'h3a7821f1),
	.w5(32'h3a119f79),
	.w6(32'h3b457ea7),
	.w7(32'h3b138eec),
	.w8(32'h3b6210e8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d1a1d),
	.w1(32'hbb24daa8),
	.w2(32'hbb0356e7),
	.w3(32'hb9945df6),
	.w4(32'hbbbe9be5),
	.w5(32'hbb66b4c2),
	.w6(32'hbae97544),
	.w7(32'h38b2a4d8),
	.w8(32'hbacc4746),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4f909),
	.w1(32'hba456c71),
	.w2(32'hbb08da6a),
	.w3(32'hbb3a0aa9),
	.w4(32'h3979cfa2),
	.w5(32'hb9ea624d),
	.w6(32'hb98f9716),
	.w7(32'hbae0fc5f),
	.w8(32'hba6d6e94),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92d01a),
	.w1(32'h39e15f28),
	.w2(32'hb95a6c12),
	.w3(32'hb87c5509),
	.w4(32'h39ca26cd),
	.w5(32'hb737897e),
	.w6(32'hb9b5edb4),
	.w7(32'hba4b3cf8),
	.w8(32'hba5fa4f5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389a2af6),
	.w1(32'h38c8885c),
	.w2(32'h37981b87),
	.w3(32'hb9c75440),
	.w4(32'h3938d9fb),
	.w5(32'hb88c8a5e),
	.w6(32'hba4ed17c),
	.w7(32'hba927152),
	.w8(32'hbab45b8a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dbdde),
	.w1(32'h3afea946),
	.w2(32'h3b385377),
	.w3(32'hb9122bf0),
	.w4(32'h3ae4ea45),
	.w5(32'hbaa2efaf),
	.w6(32'h3a41a99f),
	.w7(32'h3a6efcc0),
	.w8(32'h3b1c2ff0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5be36a),
	.w1(32'hbad227d6),
	.w2(32'hbb0e0f9a),
	.w3(32'hbabc2178),
	.w4(32'hbb65dc78),
	.w5(32'h37592d65),
	.w6(32'hbb070c07),
	.w7(32'h3af66f78),
	.w8(32'hbb1631f8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9900e),
	.w1(32'h3b18261f),
	.w2(32'h3b67d379),
	.w3(32'hbacb01ec),
	.w4(32'hbaf37656),
	.w5(32'h3a68d1e2),
	.w6(32'h3a01b89d),
	.w7(32'h3afbc3f3),
	.w8(32'hbaaf25df),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a16f5),
	.w1(32'h3b829b08),
	.w2(32'h3b79ddb5),
	.w3(32'hb877adcd),
	.w4(32'h3aa38d00),
	.w5(32'h39774fd9),
	.w6(32'h3b072a4f),
	.w7(32'h3b1a5e92),
	.w8(32'hbae32076),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4a2b6),
	.w1(32'hbbf514cd),
	.w2(32'hbb9719d2),
	.w3(32'hbbf91ec3),
	.w4(32'hbb5ebd42),
	.w5(32'h3a0cd1ef),
	.w6(32'hbb887723),
	.w7(32'hbb44d4fd),
	.w8(32'h39970209),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a125af0),
	.w1(32'hba6c123b),
	.w2(32'h3a3efa40),
	.w3(32'h3a1ee1c0),
	.w4(32'h3abbeac8),
	.w5(32'h39f0b153),
	.w6(32'hbae20c5b),
	.w7(32'hba786915),
	.w8(32'h3a99c0a0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17ca13),
	.w1(32'h3afeefec),
	.w2(32'h3b985113),
	.w3(32'h3ab14ea3),
	.w4(32'h3701f532),
	.w5(32'h3b0a3eca),
	.w6(32'hba3a7ef7),
	.w7(32'h3b6435d6),
	.w8(32'h38e8c4bf),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae46928),
	.w1(32'h3b87dddb),
	.w2(32'h3b54890d),
	.w3(32'hbb02f330),
	.w4(32'hb7cfeda8),
	.w5(32'h39c643ce),
	.w6(32'h3a0ea587),
	.w7(32'h3b0963bd),
	.w8(32'hbac73e9c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39013ab4),
	.w1(32'hbadf98c3),
	.w2(32'hba84257d),
	.w3(32'hbb368aba),
	.w4(32'hbaff697e),
	.w5(32'hb9de2ccf),
	.w6(32'hbaa3732d),
	.w7(32'hba720fbe),
	.w8(32'h39125e01),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84ca68),
	.w1(32'h3b824e9e),
	.w2(32'h39e9a4eb),
	.w3(32'h3b27a864),
	.w4(32'h3ad67c1a),
	.w5(32'hba278c01),
	.w6(32'h3b274c82),
	.w7(32'h3a9f626e),
	.w8(32'h39021afa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b526c91),
	.w1(32'h3ae978fe),
	.w2(32'hba43ff41),
	.w3(32'h39f824dd),
	.w4(32'h38fe7b7d),
	.w5(32'hbb306ba2),
	.w6(32'h3b295d4c),
	.w7(32'h3b278215),
	.w8(32'hb97b01c0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abac371),
	.w1(32'h3b1d29b5),
	.w2(32'h3af8b5f7),
	.w3(32'h3af60b5c),
	.w4(32'h3b01c2a6),
	.w5(32'h3a7bb95c),
	.w6(32'h3ad01f3e),
	.w7(32'h3a79184d),
	.w8(32'h394422ad),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe24e4),
	.w1(32'h3a572ebe),
	.w2(32'hb976e128),
	.w3(32'h3a48c872),
	.w4(32'h39239889),
	.w5(32'hba51b83a),
	.w6(32'h38a3f02e),
	.w7(32'h397e9cd7),
	.w8(32'hba254548),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a3f9d),
	.w1(32'hba050517),
	.w2(32'hba5bf93e),
	.w3(32'hba9a5ba3),
	.w4(32'hb9a61c76),
	.w5(32'hba0b776a),
	.w6(32'hba8ccc20),
	.w7(32'hba5cb3e6),
	.w8(32'h38a882ae),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3deb51),
	.w1(32'hb826dbc5),
	.w2(32'hbaa53a37),
	.w3(32'h3992e183),
	.w4(32'hb906d6e9),
	.w5(32'hbaa388f9),
	.w6(32'h3a076c46),
	.w7(32'h39d52738),
	.w8(32'hba68e0a4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11f3a9),
	.w1(32'hbbaa7312),
	.w2(32'hbbe4474a),
	.w3(32'hbb210a01),
	.w4(32'hbb8ed801),
	.w5(32'hbbc27286),
	.w6(32'hba623261),
	.w7(32'hbb2b760e),
	.w8(32'hbb8550d9),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6981a),
	.w1(32'h3c114702),
	.w2(32'h3bad7ef8),
	.w3(32'h3c250e73),
	.w4(32'h3c02fc11),
	.w5(32'h38ca2421),
	.w6(32'h3c0c792f),
	.w7(32'h3bcc3526),
	.w8(32'h3b04d6b3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad56398),
	.w1(32'hbb1e2406),
	.w2(32'hbad8d746),
	.w3(32'hbb2fe93b),
	.w4(32'hba60856a),
	.w5(32'h395d791a),
	.w6(32'hbb161b20),
	.w7(32'hba17cc79),
	.w8(32'h38312282),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48e8c8),
	.w1(32'h3a36216c),
	.w2(32'h3a94be58),
	.w3(32'hb7fce215),
	.w4(32'h3a6c96bb),
	.w5(32'hb9c43856),
	.w6(32'h3acbb576),
	.w7(32'h3ad4256c),
	.w8(32'h3b1e2cce),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf12bdb),
	.w1(32'h3be3d644),
	.w2(32'h3b255e4c),
	.w3(32'h3bf835a6),
	.w4(32'h3bc84e0b),
	.w5(32'hbaac9054),
	.w6(32'h3bc1a9e4),
	.w7(32'h3b926e36),
	.w8(32'hbb36375f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39896c24),
	.w1(32'hbaa20d10),
	.w2(32'hbb16e63c),
	.w3(32'hba124f3b),
	.w4(32'hba1cc18d),
	.w5(32'hba9c2146),
	.w6(32'h38ca1665),
	.w7(32'h39472b6d),
	.w8(32'hb982ce24),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a801129),
	.w1(32'h3965ea77),
	.w2(32'hba3d33a4),
	.w3(32'hb92f7f9d),
	.w4(32'hba1e1649),
	.w5(32'hba7cf35a),
	.w6(32'h37b1b945),
	.w7(32'h382f82d4),
	.w8(32'hb95c6708),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05ba06),
	.w1(32'h39eda8dc),
	.w2(32'h37ef3971),
	.w3(32'hb5d9db24),
	.w4(32'h38e5a6bf),
	.w5(32'hb992d834),
	.w6(32'h39fe3fde),
	.w7(32'h3a5179f8),
	.w8(32'h39c7870a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb818d1e),
	.w1(32'hbbddbf89),
	.w2(32'hbb4f8b43),
	.w3(32'hbb990703),
	.w4(32'hbbba3abc),
	.w5(32'hba2cb8b6),
	.w6(32'hbb6afc20),
	.w7(32'hba522a30),
	.w8(32'h3a6b5f4b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2381b9),
	.w1(32'h3adc3d85),
	.w2(32'h3a576a19),
	.w3(32'h3b41f71c),
	.w4(32'h3a91ab09),
	.w5(32'hba19cfd2),
	.w6(32'h3b1a9111),
	.w7(32'h39dafc6d),
	.w8(32'hba54bc70),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb733c85f),
	.w1(32'h360dbdc2),
	.w2(32'h3743dd85),
	.w3(32'hb5be23a5),
	.w4(32'h36d9b8fc),
	.w5(32'h37991835),
	.w6(32'hb68cc006),
	.w7(32'h3743f5e5),
	.w8(32'h3743e3aa),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fe4625),
	.w1(32'hb5e625a7),
	.w2(32'hb653aefb),
	.w3(32'h36934a06),
	.w4(32'hb7273b4f),
	.w5(32'hb71b6f29),
	.w6(32'hb6e59173),
	.w7(32'hb78256c1),
	.w8(32'hb78643a6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85e01d9),
	.w1(32'h3768a041),
	.w2(32'h3943d429),
	.w3(32'hba82f1d9),
	.w4(32'h3883dbba),
	.w5(32'h3b09c87d),
	.w6(32'hba170226),
	.w7(32'h396bb15a),
	.w8(32'h3b10f62d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58c574),
	.w1(32'hbb258b62),
	.w2(32'hba24b2c9),
	.w3(32'hba33fa82),
	.w4(32'hb95c97a8),
	.w5(32'h3aa6a39c),
	.w6(32'h3a1e9333),
	.w7(32'h3a1a8383),
	.w8(32'h3a575a17),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f53379),
	.w1(32'h3a939b97),
	.w2(32'h3a1d19fd),
	.w3(32'hbad2ba6f),
	.w4(32'h39a82fcf),
	.w5(32'hb8e6ee3e),
	.w6(32'h3a2f23d8),
	.w7(32'h3b636924),
	.w8(32'h3b218b0d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70d1171),
	.w1(32'hb51594ea),
	.w2(32'hb4d3f96c),
	.w3(32'hb6a42713),
	.w4(32'h370bbced),
	.w5(32'hb70f67f9),
	.w6(32'h36db0529),
	.w7(32'h375961c1),
	.w8(32'hb6ac0540),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad588e5),
	.w1(32'h3a3bd9c5),
	.w2(32'hbace0790),
	.w3(32'hbab84fa7),
	.w4(32'hbabc35fd),
	.w5(32'hbb073c68),
	.w6(32'h397d7d38),
	.w7(32'h3abbdb59),
	.w8(32'hb8ddf0b4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dae493),
	.w1(32'hbab508d9),
	.w2(32'hbb13aeb8),
	.w3(32'hbb4995c1),
	.w4(32'hbaef46ec),
	.w5(32'hbab00b91),
	.w6(32'hba7d116a),
	.w7(32'h3a31385e),
	.w8(32'h3a2331f3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb45425),
	.w1(32'h3bd8c0a4),
	.w2(32'h3b88df84),
	.w3(32'h3ba5f237),
	.w4(32'h3b9bafcd),
	.w5(32'h3aa488d3),
	.w6(32'h3b6994ef),
	.w7(32'h3b8522f8),
	.w8(32'h3a3a669f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9479c6),
	.w1(32'h3940351f),
	.w2(32'hba35426a),
	.w3(32'hb9d52d19),
	.w4(32'hba05d0ff),
	.w5(32'h39018b38),
	.w6(32'h38719f6f),
	.w7(32'h3a61a946),
	.w8(32'h3b05d589),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab774ab),
	.w1(32'hbb0cf6d8),
	.w2(32'hbad0af08),
	.w3(32'hbade55ac),
	.w4(32'hbaeba1cc),
	.w5(32'hba4b0075),
	.w6(32'hbb064539),
	.w7(32'hba5fe217),
	.w8(32'hba931490),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba900851),
	.w1(32'hba5c9b4d),
	.w2(32'hba2c0091),
	.w3(32'hba333177),
	.w4(32'hba4ba1f3),
	.w5(32'hb9cc85ea),
	.w6(32'hba674f2e),
	.w7(32'hba217389),
	.w8(32'hba57818e),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b1d7d),
	.w1(32'hbad075ee),
	.w2(32'hba5eb21a),
	.w3(32'hbb3d6693),
	.w4(32'hbae3d139),
	.w5(32'hb907c134),
	.w6(32'hbb3e1ec9),
	.w7(32'hbabce159),
	.w8(32'h39adbb81),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba955319),
	.w1(32'hbb7721a6),
	.w2(32'hbb15d41b),
	.w3(32'hba9d694a),
	.w4(32'hbb402a19),
	.w5(32'hbae7dfb9),
	.w6(32'hbb04ed00),
	.w7(32'hbb2c0529),
	.w8(32'hbaef29ac),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e044c),
	.w1(32'hba2f561d),
	.w2(32'hb8a6bb2f),
	.w3(32'hba9d1394),
	.w4(32'hba294ea1),
	.w5(32'h392d438e),
	.w6(32'hbaada06b),
	.w7(32'hba496eff),
	.w8(32'hb86d6217),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28bf5b),
	.w1(32'h3b381133),
	.w2(32'h3adb77c4),
	.w3(32'h3b508f54),
	.w4(32'h3b21a7e9),
	.w5(32'hb8a35ca8),
	.w6(32'h3b27a16d),
	.w7(32'h3a97e213),
	.w8(32'hb9d24b5f),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9b595),
	.w1(32'hba288f98),
	.w2(32'hb989eb01),
	.w3(32'hba0d8124),
	.w4(32'hba26af6d),
	.w5(32'hb8bb46ba),
	.w6(32'hba0b52be),
	.w7(32'hba0cc384),
	.w8(32'hb98ff8b7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa6b08),
	.w1(32'h3a7a7f8b),
	.w2(32'hba28bc1d),
	.w3(32'h3a3ba5f8),
	.w4(32'h382e337f),
	.w5(32'hbaa2fe78),
	.w6(32'h3a5cbdb7),
	.w7(32'h3a0e3a34),
	.w8(32'hba37d9e0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95744ab),
	.w1(32'hb8be79bd),
	.w2(32'hb84407c6),
	.w3(32'hb8b21390),
	.w4(32'h3739f170),
	.w5(32'h38a1c602),
	.w6(32'hb894eb98),
	.w7(32'hb863b55d),
	.w8(32'h37f47609),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39674c4b),
	.w1(32'hb9a820f2),
	.w2(32'hba8541f4),
	.w3(32'hbaef2860),
	.w4(32'hbab2f8cf),
	.w5(32'hba9490fd),
	.w6(32'hba8a4f5d),
	.w7(32'hb99a30c3),
	.w8(32'h39f1004f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb848be68),
	.w1(32'h381a59fb),
	.w2(32'h398ff728),
	.w3(32'hb9aafa03),
	.w4(32'hb7b6c84f),
	.w5(32'h38caeeb8),
	.w6(32'hb8752d12),
	.w7(32'h38d26d8e),
	.w8(32'h398b34dc),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0744a),
	.w1(32'h3a00b9b8),
	.w2(32'h3930f181),
	.w3(32'h3b3d1221),
	.w4(32'h3aaed0d2),
	.w5(32'h39a8828a),
	.w6(32'h3b5fdaa1),
	.w7(32'h3b1f29bd),
	.w8(32'h3aa803ba),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b45056),
	.w1(32'h37d69a5f),
	.w2(32'hb8a62690),
	.w3(32'hb847e609),
	.w4(32'hb7addafd),
	.w5(32'hb8c76c72),
	.w6(32'hb8435112),
	.w7(32'hb8507358),
	.w8(32'hb8e7301d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980f52c),
	.w1(32'h399c0247),
	.w2(32'h395e85c8),
	.w3(32'h39d93caa),
	.w4(32'h393aa4c2),
	.w5(32'h365411a2),
	.w6(32'h39e6023f),
	.w7(32'h399bd502),
	.w8(32'h38f1338f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae53da8),
	.w1(32'hbb662341),
	.w2(32'hbb194b8c),
	.w3(32'hbb3a8a4a),
	.w4(32'hbb8284b7),
	.w5(32'hbaa3f3a7),
	.w6(32'hbb32d38d),
	.w7(32'hbb3002e5),
	.w8(32'hba94790a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13326a),
	.w1(32'h3b7ce468),
	.w2(32'hbb28ab94),
	.w3(32'h3b8d1972),
	.w4(32'h3b109da7),
	.w5(32'hbb5feeee),
	.w6(32'h3ba16dad),
	.w7(32'h3a13dcae),
	.w8(32'hbb4ed3ab),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45b45f),
	.w1(32'hb8a1cc6b),
	.w2(32'h3a09763b),
	.w3(32'hba3c5a2e),
	.w4(32'h392ffb86),
	.w5(32'h3a307cc8),
	.w6(32'hba7b60ef),
	.w7(32'hb90e1891),
	.w8(32'h3a103f45),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f821f9),
	.w1(32'hbae00e39),
	.w2(32'hbb05be26),
	.w3(32'hbb4353c6),
	.w4(32'hbb26fb67),
	.w5(32'hba8ea80b),
	.w6(32'hbb09ad80),
	.w7(32'h3939b390),
	.w8(32'h3a840f88),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9761b5f),
	.w1(32'hba1d0a01),
	.w2(32'hba5ec918),
	.w3(32'hb9c100f5),
	.w4(32'hb9eb5719),
	.w5(32'hba1b146d),
	.w6(32'hb994afba),
	.w7(32'hba083dc9),
	.w8(32'hba1a4f06),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19b719),
	.w1(32'h3b15586b),
	.w2(32'h3a9ae029),
	.w3(32'h3a91d597),
	.w4(32'h3abfadfb),
	.w5(32'hb7e16fef),
	.w6(32'h3ad18920),
	.w7(32'h3ba5c340),
	.w8(32'h3b433539),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed67b6),
	.w1(32'h3abb910f),
	.w2(32'h39e420c8),
	.w3(32'h3acbc4ea),
	.w4(32'h3a894c70),
	.w5(32'hb9df82b1),
	.w6(32'h3ac8e01f),
	.w7(32'h3a82464c),
	.w8(32'h378e0624),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb95af8),
	.w1(32'h3b3fafea),
	.w2(32'hba65f020),
	.w3(32'h3b52a2ee),
	.w4(32'h3a7a59ab),
	.w5(32'hbb81f016),
	.w6(32'h3baadbfb),
	.w7(32'h3b2b1207),
	.w8(32'hbae1713e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370cc74c),
	.w1(32'hb91badfe),
	.w2(32'hb94554da),
	.w3(32'hb9ba8bd8),
	.w4(32'hb90df2cd),
	.w5(32'hb927affd),
	.w6(32'hb9b3bca4),
	.w7(32'hb9784a9c),
	.w8(32'hb909003b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10728f),
	.w1(32'h3a251eb4),
	.w2(32'hba86858e),
	.w3(32'h3a0e4c0c),
	.w4(32'h38b51df6),
	.w5(32'hbaa62b46),
	.w6(32'h3aa0dd1e),
	.w7(32'h39f7085f),
	.w8(32'hba30f685),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7aa2fd8),
	.w1(32'hb639a4af),
	.w2(32'hb7876864),
	.w3(32'hb72be158),
	.w4(32'h370fc376),
	.w5(32'hb74d83f7),
	.w6(32'hb741a12c),
	.w7(32'h3747c3e7),
	.w8(32'hb7c02ac1),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0c482),
	.w1(32'hba7e5c4e),
	.w2(32'hba81d9f1),
	.w3(32'h3aba35d1),
	.w4(32'hba565985),
	.w5(32'hba6e1321),
	.w6(32'h3af4dc9e),
	.w7(32'hb8db65d9),
	.w8(32'h387b0862),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbb6b2),
	.w1(32'hb9264688),
	.w2(32'hba032831),
	.w3(32'h3a4f7e15),
	.w4(32'h393b9739),
	.w5(32'hb9b396be),
	.w6(32'h39535b7d),
	.w7(32'hb8999ccc),
	.w8(32'hb9dae844),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd478b),
	.w1(32'hb6e1f2b4),
	.w2(32'h39c3e8e7),
	.w3(32'hba640d15),
	.w4(32'hba6aa5e8),
	.w5(32'hb949f213),
	.w6(32'hb9e82090),
	.w7(32'h39169d8e),
	.w8(32'h3a75e792),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378ef4e0),
	.w1(32'hb706e2d1),
	.w2(32'hb7a9dfec),
	.w3(32'h376d6863),
	.w4(32'hb6db0d2b),
	.w5(32'hb7bfcf11),
	.w6(32'h376a4f64),
	.w7(32'h36ae87f2),
	.w8(32'hb73ad9fc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f29225),
	.w1(32'hb8c6bfa1),
	.w2(32'hb893923b),
	.w3(32'hb930ab19),
	.w4(32'hb8e7dc48),
	.w5(32'hb8b8c58f),
	.w6(32'hb8d346f4),
	.w7(32'hb8447807),
	.w8(32'hb7d918a1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a126df0),
	.w1(32'h3a1e263d),
	.w2(32'hb8a3b95a),
	.w3(32'hba23e66e),
	.w4(32'h3906ab46),
	.w5(32'hb9edde36),
	.w6(32'hba4010a4),
	.w7(32'h383f9e29),
	.w8(32'h3a3f7a48),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2259f),
	.w1(32'h3b06d27c),
	.w2(32'h39ee9d50),
	.w3(32'hb9a383a2),
	.w4(32'h3a3cef91),
	.w5(32'h38e666f5),
	.w6(32'hb726a685),
	.w7(32'h3a135b00),
	.w8(32'h3a8d7911),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4706e8),
	.w1(32'h39f2c15b),
	.w2(32'h38fab698),
	.w3(32'h3a05b3c9),
	.w4(32'h3945748f),
	.w5(32'hb90be2a7),
	.w6(32'h39f14f88),
	.w7(32'h3960a9eb),
	.w8(32'h38aca84c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20d223),
	.w1(32'h3a80e79e),
	.w2(32'h3907e455),
	.w3(32'h3adacf4e),
	.w4(32'h392788b6),
	.w5(32'hba7db46d),
	.w6(32'h3a1e6f2f),
	.w7(32'hb9fc65df),
	.w8(32'h38c191f7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7aae4),
	.w1(32'h3c0aaa15),
	.w2(32'h3b19ddbb),
	.w3(32'h3b6836a8),
	.w4(32'h3bc34c31),
	.w5(32'h3a0adbe4),
	.w6(32'h3b909f0d),
	.w7(32'h3c3d4ee8),
	.w8(32'h3be0070e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77fc71),
	.w1(32'hbc0e1205),
	.w2(32'hbbbe2343),
	.w3(32'hbbc0c49b),
	.w4(32'hbc03f6be),
	.w5(32'hbb762bf6),
	.w6(32'hbbcafca4),
	.w7(32'hbbecbd53),
	.w8(32'hbb3ecf5a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391a2217),
	.w1(32'h39cfaff9),
	.w2(32'h39fbfdc8),
	.w3(32'h39953480),
	.w4(32'h3a09dd7c),
	.w5(32'h39be262b),
	.w6(32'h396cb7e7),
	.w7(32'h39a47a86),
	.w8(32'h38d6bc50),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a2fe73),
	.w1(32'hb805a0b0),
	.w2(32'hb7dd7ebb),
	.w3(32'hb7bcf27b),
	.w4(32'hb7e12ab3),
	.w5(32'hb797e908),
	.w6(32'hb71f2a3a),
	.w7(32'hb7a01877),
	.w8(32'hb694accb),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9da6f),
	.w1(32'hb90a75e4),
	.w2(32'hb90465a9),
	.w3(32'hb8e71a55),
	.w4(32'hb7bb3a04),
	.w5(32'hb80b04d0),
	.w6(32'hb9638f46),
	.w7(32'hb8a3d377),
	.w8(32'h388f749a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d11300),
	.w1(32'h3604744a),
	.w2(32'h36bf0759),
	.w3(32'h37863977),
	.w4(32'hb6c5e91c),
	.w5(32'hb63d8a5d),
	.w6(32'hb6fdbdc1),
	.w7(32'hb7207d66),
	.w8(32'hb6efda94),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398599f6),
	.w1(32'hb9cf1b8e),
	.w2(32'hb9a73876),
	.w3(32'h396d3a00),
	.w4(32'hb9cf1e44),
	.w5(32'hb994d6d0),
	.w6(32'h3849a874),
	.w7(32'hba08f857),
	.w8(32'hba1323d3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62fa4e),
	.w1(32'h3a58f43f),
	.w2(32'h39e8a8ee),
	.w3(32'h3b26b64a),
	.w4(32'h3a8d84be),
	.w5(32'hb9f49c00),
	.w6(32'h3b078ccc),
	.w7(32'h3ac8a1c4),
	.w8(32'h3a78e069),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafb2ff),
	.w1(32'hbacff9fe),
	.w2(32'hbb2c1fad),
	.w3(32'hbb3eb9f6),
	.w4(32'hba2560e1),
	.w5(32'hbaa14cdb),
	.w6(32'hba5ce1c8),
	.w7(32'h3b133adc),
	.w8(32'h3a25c39c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a2028),
	.w1(32'hb8ff6cb9),
	.w2(32'hba23d3a0),
	.w3(32'hb9ebfb60),
	.w4(32'hba5729f6),
	.w5(32'hba047d7d),
	.w6(32'hb99a4a2a),
	.w7(32'hb945a355),
	.w8(32'h38c3a29e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398dbf4d),
	.w1(32'h39c9cb20),
	.w2(32'hb911ac03),
	.w3(32'hba923e85),
	.w4(32'hb9b698d8),
	.w5(32'h39388a38),
	.w6(32'hb95ad244),
	.w7(32'h3b12693d),
	.w8(32'h3b013ef1),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c6954),
	.w1(32'h3aea5c9a),
	.w2(32'h3b00ae63),
	.w3(32'hbab5b459),
	.w4(32'h3ac4e52e),
	.w5(32'h3b1a2668),
	.w6(32'hb990e4ae),
	.w7(32'h3ae5c452),
	.w8(32'h3b336c15),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ab6323),
	.w1(32'hb6b5a97d),
	.w2(32'hb48950f9),
	.w3(32'hb6c72d6f),
	.w4(32'hb71ca2e5),
	.w5(32'hb6bb0842),
	.w6(32'hb72ae92f),
	.w7(32'hb746fb8c),
	.w8(32'hb75519af),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafd611),
	.w1(32'h3b083d10),
	.w2(32'h3aa4839e),
	.w3(32'h3a8bd65e),
	.w4(32'h3b0802ef),
	.w5(32'h3a195ea2),
	.w6(32'h3a60340a),
	.w7(32'h3a6ea68c),
	.w8(32'h394bab08),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb818648a),
	.w1(32'hb81c173e),
	.w2(32'hb85bae0e),
	.w3(32'hb801f3f1),
	.w4(32'hb7d7fb5c),
	.w5(32'hb7f46708),
	.w6(32'hb8635ab1),
	.w7(32'hb82f908f),
	.w8(32'hb85a116d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4227a3),
	.w1(32'h3991bdcf),
	.w2(32'h37f1476f),
	.w3(32'h3b2299ca),
	.w4(32'h3a95d539),
	.w5(32'h3a85b36b),
	.w6(32'h3b81266d),
	.w7(32'h3a9c74c7),
	.w8(32'h3b5faec3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11ee05),
	.w1(32'hbb7875a1),
	.w2(32'hbb61d25c),
	.w3(32'hbb0689a4),
	.w4(32'hbb3f6ca6),
	.w5(32'hbad5b172),
	.w6(32'hbb29fedf),
	.w7(32'hbaec9b75),
	.w8(32'hba4c6df8),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba957294),
	.w1(32'hbad401a6),
	.w2(32'hbabfb1f0),
	.w3(32'hbb462da1),
	.w4(32'hbaf806b7),
	.w5(32'hb941a8b0),
	.w6(32'hbafc372d),
	.w7(32'hba1c7b94),
	.w8(32'h3a373fd0),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e6b65),
	.w1(32'hb92487e8),
	.w2(32'h3a123031),
	.w3(32'hb9c66a75),
	.w4(32'hb8ea1635),
	.w5(32'h3a3f2cb7),
	.w6(32'hba67a012),
	.w7(32'hb9d0ec31),
	.w8(32'h39802e70),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ff6d0),
	.w1(32'hbba8bb79),
	.w2(32'hbb1d425f),
	.w3(32'hbbca4896),
	.w4(32'hbb7c2702),
	.w5(32'hba38d128),
	.w6(32'hbbc181db),
	.w7(32'hbb1a573e),
	.w8(32'h39790742),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc43a2),
	.w1(32'h3a06943f),
	.w2(32'hba824169),
	.w3(32'h3957c734),
	.w4(32'hba1545d3),
	.w5(32'hbac01d7d),
	.w6(32'h3a6b1727),
	.w7(32'h3a57a4ab),
	.w8(32'hb949556c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2362f),
	.w1(32'h3acfdd72),
	.w2(32'hb87fe4cb),
	.w3(32'hbb24c121),
	.w4(32'h3a9aac73),
	.w5(32'h3a8edd75),
	.w6(32'hb7bdbf29),
	.w7(32'h3bb5bf7a),
	.w8(32'h3ba7f610),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f6fed2),
	.w1(32'h3812f9ea),
	.w2(32'h378547e5),
	.w3(32'h3819a70c),
	.w4(32'h381c03b8),
	.w5(32'h379ff14b),
	.w6(32'h38153cd1),
	.w7(32'h383a0973),
	.w8(32'h38054ee3),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c3d314),
	.w1(32'hb819a8ba),
	.w2(32'hb858032c),
	.w3(32'hb7ea62f8),
	.w4(32'hb893f8c6),
	.w5(32'hb8bc0dd9),
	.w6(32'h37353c5a),
	.w7(32'hb75da617),
	.w8(32'hb7f55a68),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a510088),
	.w1(32'h3b07d1d8),
	.w2(32'hba95640a),
	.w3(32'hb9e36098),
	.w4(32'h3b041541),
	.w5(32'h3a9a5712),
	.w6(32'h3a99be38),
	.w7(32'h3b196281),
	.w8(32'h3b04ff72),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43bcd4),
	.w1(32'h3c0d4265),
	.w2(32'h3aaf175b),
	.w3(32'h3b9510be),
	.w4(32'h3b19c51d),
	.w5(32'hbb4a365a),
	.w6(32'h3bd85fe4),
	.w7(32'h3b2ed1e1),
	.w8(32'h3a869b14),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8b544),
	.w1(32'hba8b5097),
	.w2(32'hbb170f8d),
	.w3(32'hbb5baf09),
	.w4(32'hbb0e6de6),
	.w5(32'hbac57859),
	.w6(32'hba6d4d56),
	.w7(32'h3adb213b),
	.w8(32'h3acc0587),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a948406),
	.w1(32'h3aa4f190),
	.w2(32'h3a2e7b2d),
	.w3(32'h3aad45e8),
	.w4(32'h3a6d684b),
	.w5(32'h38e247b9),
	.w6(32'h3a4de863),
	.w7(32'h391e4905),
	.w8(32'hb928bd53),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c0ae25),
	.w1(32'hb7fc6533),
	.w2(32'hb87c0464),
	.w3(32'hb740483b),
	.w4(32'hb848524e),
	.w5(32'hb84587c1),
	.w6(32'hb6f62b0e),
	.w7(32'hb816be99),
	.w8(32'hb847d46b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb790c440),
	.w1(32'hb88f13d9),
	.w2(32'hb86bd245),
	.w3(32'hb8511cea),
	.w4(32'hb921b762),
	.w5(32'hb9330e5d),
	.w6(32'hb7ce9d7f),
	.w7(32'hb8d34718),
	.w8(32'hb8e94a13),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2201f3),
	.w1(32'h3b674911),
	.w2(32'h3b578334),
	.w3(32'h3b58b3f6),
	.w4(32'h3b91217e),
	.w5(32'h3ad51013),
	.w6(32'h3b4bb267),
	.w7(32'h3b4cfa79),
	.w8(32'h3a19b909),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb30c0),
	.w1(32'h3c1c5a7e),
	.w2(32'h3b884c55),
	.w3(32'h3bb90340),
	.w4(32'h3bf571de),
	.w5(32'h3a581f28),
	.w6(32'h3bdda377),
	.w7(32'h3c0db9bd),
	.w8(32'h3b6ac06a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92fb28),
	.w1(32'h3c0c8b0b),
	.w2(32'h3bb1638a),
	.w3(32'h3bf69ce1),
	.w4(32'h3c09a6e3),
	.w5(32'h3b130ece),
	.w6(32'h3c07d6bd),
	.w7(32'h3bcd7d88),
	.w8(32'hba5a39ea),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa1467),
	.w1(32'hbaf50a5a),
	.w2(32'hba1ca6e5),
	.w3(32'hbb07063a),
	.w4(32'hbab7d226),
	.w5(32'h396883cc),
	.w6(32'hbac9bae8),
	.w7(32'hba27bd2f),
	.w8(32'h39cd1d9b),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb190a0c),
	.w1(32'hbb9ecfcb),
	.w2(32'hbb59380a),
	.w3(32'hbb65c191),
	.w4(32'hbb9d51fa),
	.w5(32'hba83bd18),
	.w6(32'hbb4d0f3d),
	.w7(32'hbb1cbea3),
	.w8(32'h3961e13b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb730a432),
	.w1(32'hb6b6199c),
	.w2(32'hb63074b2),
	.w3(32'hb7835656),
	.w4(32'hb7006edf),
	.w5(32'hb5965e6a),
	.w6(32'hb78db8c8),
	.w7(32'hb6c58b1f),
	.w8(32'hb6694de3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7264356),
	.w1(32'h3585b091),
	.w2(32'h363d553c),
	.w3(32'hb713e32d),
	.w4(32'h3701fd85),
	.w5(32'h37059bef),
	.w6(32'hb76dd948),
	.w7(32'hb6376161),
	.w8(32'h35aeee0d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373ed0a0),
	.w1(32'h37362eae),
	.w2(32'h36e744f5),
	.w3(32'h378b3aa2),
	.w4(32'h372406d0),
	.w5(32'hb5b63598),
	.w6(32'h36f298e8),
	.w7(32'hb7414b51),
	.w8(32'hb7582bc4),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e6ae24),
	.w1(32'hb5ebffd3),
	.w2(32'hb73afacc),
	.w3(32'hb7a6b179),
	.w4(32'hb794ee81),
	.w5(32'hb7b4548b),
	.w6(32'hb7d9cca0),
	.w7(32'hb784644d),
	.w8(32'hb71aca8e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a10ba),
	.w1(32'h396ea75d),
	.w2(32'h39ea915c),
	.w3(32'hb98d2043),
	.w4(32'h39aad3b5),
	.w5(32'h39f6e04c),
	.w6(32'hb9b7f279),
	.w7(32'hb891a5ae),
	.w8(32'h3903647c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17fef8),
	.w1(32'h3add98b0),
	.w2(32'h3a9a3e60),
	.w3(32'h3a4dde17),
	.w4(32'hba0f5cc2),
	.w5(32'hba0e44ae),
	.w6(32'h3ad8e1bb),
	.w7(32'h39084b5f),
	.w8(32'h3aa264f0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7e27d),
	.w1(32'hbac9dbad),
	.w2(32'hba6b8620),
	.w3(32'hbb1e2370),
	.w4(32'hbaacd8c7),
	.w5(32'hba1d972a),
	.w6(32'hbaffe084),
	.w7(32'hba7ac22e),
	.w8(32'h3a29e627),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cf123c),
	.w1(32'hb7b53015),
	.w2(32'hb80651a9),
	.w3(32'hb7fc620a),
	.w4(32'hb79eae9b),
	.w5(32'hb807783f),
	.w6(32'hb7dad6dc),
	.w7(32'hb69d4206),
	.w8(32'hb7a9493e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c96c4),
	.w1(32'h3c36329c),
	.w2(32'h3c0fe0b9),
	.w3(32'h3c3c90ac),
	.w4(32'h3c27385f),
	.w5(32'h3b2e78c9),
	.w6(32'h3c16a5ed),
	.w7(32'h3bf72590),
	.w8(32'h3a2058be),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cadde),
	.w1(32'h3afbb69a),
	.w2(32'hb8f3491b),
	.w3(32'h3b1ac0c8),
	.w4(32'h3abba8b8),
	.w5(32'hba4e09b0),
	.w6(32'h3b3cdabe),
	.w7(32'h3b153756),
	.w8(32'hb9da0b64),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ca513),
	.w1(32'hb8a0282d),
	.w2(32'h381595ac),
	.w3(32'hb8b03012),
	.w4(32'hb8e734e3),
	.w5(32'h382fb234),
	.w6(32'hb86df59a),
	.w7(32'hb8663bf4),
	.w8(32'h38242645),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ec214),
	.w1(32'h3b63a2f2),
	.w2(32'h3acaf77f),
	.w3(32'h3b5291ab),
	.w4(32'h3b334cca),
	.w5(32'h39738b2c),
	.w6(32'h3b4039d7),
	.w7(32'h3b079a63),
	.w8(32'h39639d87),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9307636),
	.w1(32'hb8a0c0ab),
	.w2(32'hb868e51c),
	.w3(32'hb91c6f0e),
	.w4(32'hb88615ca),
	.w5(32'hb877c034),
	.w6(32'hb8ea8986),
	.w7(32'hb893d70c),
	.w8(32'hb8ac192f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9525cfe),
	.w1(32'hb83a9015),
	.w2(32'h37d24d31),
	.w3(32'hb991a7ed),
	.w4(32'hb906627c),
	.w5(32'hb79d337b),
	.w6(32'hb814f9a2),
	.w7(32'h37b0d59e),
	.w8(32'hb611bd3c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73099ae),
	.w1(32'hb7a5eea7),
	.w2(32'hb7c27f8a),
	.w3(32'hb78e7278),
	.w4(32'hb755feae),
	.w5(32'hb73e0cd7),
	.w6(32'hb599f24c),
	.w7(32'hb79020d7),
	.w8(32'hb7c2d175),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68ab1b0),
	.w1(32'hb6ae04d6),
	.w2(32'hb6104cff),
	.w3(32'hb6248254),
	.w4(32'h37a803d9),
	.w5(32'hb66f5c5d),
	.w6(32'hb78d7fbc),
	.w7(32'h36f35532),
	.w8(32'h36befa4f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5acd1e),
	.w1(32'hba87f637),
	.w2(32'hb98e9828),
	.w3(32'hbabfab5c),
	.w4(32'hba64660f),
	.w5(32'hba14e330),
	.w6(32'hbaa25ae7),
	.w7(32'hb91e74e3),
	.w8(32'h397129c9),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85f4a4),
	.w1(32'h3b071e18),
	.w2(32'hbad4f9e1),
	.w3(32'h3a831b49),
	.w4(32'h39a72f73),
	.w5(32'hbb403f43),
	.w6(32'h3b25bef6),
	.w7(32'h3b09be3d),
	.w8(32'hba7ea438),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b303a68),
	.w1(32'h3b3a4537),
	.w2(32'h3897347f),
	.w3(32'h3acc0312),
	.w4(32'h3ab51add),
	.w5(32'hbaa44f0c),
	.w6(32'h3b0310e4),
	.w7(32'h3b04b911),
	.w8(32'hb9a8899e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7f03b),
	.w1(32'h3a66c9e8),
	.w2(32'hba980dcb),
	.w3(32'h3a6f9f09),
	.w4(32'hb8bb7c46),
	.w5(32'hbb0ac357),
	.w6(32'h3a58e97c),
	.w7(32'h3b01228c),
	.w8(32'h3887b594),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b8b92),
	.w1(32'hb8fb41f3),
	.w2(32'h3875bcb7),
	.w3(32'hb9359b83),
	.w4(32'hb91a383e),
	.w5(32'h37cab573),
	.w6(32'hb8b6083f),
	.w7(32'hb895bb63),
	.w8(32'h383c9504),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37016b2d),
	.w1(32'h371162f8),
	.w2(32'h37143534),
	.w3(32'h3716daab),
	.w4(32'h36f862bf),
	.w5(32'h34aa8554),
	.w6(32'h355be0b9),
	.w7(32'h3336cec6),
	.w8(32'hb605ce6a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80b29e7),
	.w1(32'hb899159f),
	.w2(32'hb8940661),
	.w3(32'hb809fd6a),
	.w4(32'hb8a57e64),
	.w5(32'hb8838521),
	.w6(32'hb7979164),
	.w7(32'hb8a1bd52),
	.w8(32'hb825db50),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f0f1df),
	.w1(32'h376bdaeb),
	.w2(32'h37af441e),
	.w3(32'hb8062779),
	.w4(32'hb784ec94),
	.w5(32'h36232ef0),
	.w6(32'hb7622917),
	.w7(32'h368163d6),
	.w8(32'h37a938d0),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26a52b),
	.w1(32'h3af6d392),
	.w2(32'h39ef82c3),
	.w3(32'h3b1b7167),
	.w4(32'h3abc4b25),
	.w5(32'hba5bca5d),
	.w6(32'h3b1b83c1),
	.w7(32'h3ac47744),
	.w8(32'hb9c56003),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4552308),
	.w1(32'h37ce6c2b),
	.w2(32'h3799b098),
	.w3(32'h37f36c22),
	.w4(32'h389945f7),
	.w5(32'h39003067),
	.w6(32'hb6695c44),
	.w7(32'h381d1cff),
	.w8(32'h39405d30),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05ef85),
	.w1(32'hb96465bb),
	.w2(32'h39db9218),
	.w3(32'hb95c46ba),
	.w4(32'hb9705708),
	.w5(32'h3a0db923),
	.w6(32'hb92058fd),
	.w7(32'hb98ee637),
	.w8(32'h3916e8e0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d155ff),
	.w1(32'h393de0b4),
	.w2(32'h3a0a4241),
	.w3(32'hb99222eb),
	.w4(32'h38cf94ce),
	.w5(32'h39e28891),
	.w6(32'hba1e40a0),
	.w7(32'hba153df0),
	.w8(32'hb7b7da87),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92fd88a),
	.w1(32'hb84a629f),
	.w2(32'hb7b02c11),
	.w3(32'hb91cb50c),
	.w4(32'hb59d233f),
	.w5(32'h382c3022),
	.w6(32'hb90016ae),
	.w7(32'h383019cc),
	.w8(32'h38d299be),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ad3d6),
	.w1(32'h39ddf9d0),
	.w2(32'h3a6a5a4e),
	.w3(32'hb95629f9),
	.w4(32'h39fc53a4),
	.w5(32'h39e948ea),
	.w6(32'hb96838b3),
	.w7(32'h3a627fed),
	.w8(32'h3a86b5be),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88792f3),
	.w1(32'hb83ef834),
	.w2(32'hb7b993c3),
	.w3(32'hb8a5157e),
	.w4(32'hb88b5f69),
	.w5(32'hb837af10),
	.w6(32'hb7d404d0),
	.w7(32'hb814a6de),
	.w8(32'hb708b3e7),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6e799),
	.w1(32'h3bbaa2c1),
	.w2(32'h39de49f3),
	.w3(32'h3bc2e694),
	.w4(32'h3b3cbfbf),
	.w5(32'hba83f94d),
	.w6(32'h3b57d21e),
	.w7(32'h3aa8f249),
	.w8(32'hbb0675ab),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89a8c06),
	.w1(32'hb670edae),
	.w2(32'hb7d2fc57),
	.w3(32'hb866adb3),
	.w4(32'hb76460af),
	.w5(32'hb780f6a2),
	.w6(32'hb85323a6),
	.w7(32'hb5ddb806),
	.w8(32'h3788233e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb36a15),
	.w1(32'h3b7e86cf),
	.w2(32'h3a202e07),
	.w3(32'hba1b7f85),
	.w4(32'hba8080b4),
	.w5(32'hbae0e363),
	.w6(32'hb99fa654),
	.w7(32'hba760ff4),
	.w8(32'hb9a1bc7a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule