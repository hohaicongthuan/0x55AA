module layer_6_featuremap_106(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc38bca),
	.w1(32'hbbc6e09f),
	.w2(32'hbc00302b),
	.w3(32'hbb9c3f78),
	.w4(32'hbbdfa41b),
	.w5(32'hbb92b428),
	.w6(32'hbb919db0),
	.w7(32'hbbe341a9),
	.w8(32'hbb1982d5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb793f8ab),
	.w1(32'hbba1acd7),
	.w2(32'hbb3f1eea),
	.w3(32'hbaf2149d),
	.w4(32'hbad613c9),
	.w5(32'h38be6ec5),
	.w6(32'hbb686521),
	.w7(32'hbb820e36),
	.w8(32'hbb8d9134),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb003cc6),
	.w1(32'h3ba81756),
	.w2(32'hbcc01585),
	.w3(32'h3c69c57c),
	.w4(32'hbaf2d4a0),
	.w5(32'hbbee41b5),
	.w6(32'h3c62a9f0),
	.w7(32'hbcc5dffa),
	.w8(32'hbc7d9367),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c7c5d),
	.w1(32'hbb32c005),
	.w2(32'hbbd494f0),
	.w3(32'hbc24623e),
	.w4(32'hbc3ded9b),
	.w5(32'hbc0f1362),
	.w6(32'hbc2a4d55),
	.w7(32'hbc49e322),
	.w8(32'hbc0ea7cc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cbdbf0),
	.w1(32'hbc1d89d9),
	.w2(32'hbcba1ee6),
	.w3(32'h3b27b8e4),
	.w4(32'hbc482ad2),
	.w5(32'hbc705c6d),
	.w6(32'h3b52b424),
	.w7(32'hbd19f8ae),
	.w8(32'hbce7e901),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc865f6f),
	.w1(32'h3b2af09a),
	.w2(32'hbafa74f8),
	.w3(32'h3bacf5b9),
	.w4(32'hbae662c7),
	.w5(32'hbb823531),
	.w6(32'h3baff27f),
	.w7(32'hbaeb1286),
	.w8(32'hbaa56e2c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7f880),
	.w1(32'h3bbf103d),
	.w2(32'h3b9bf299),
	.w3(32'h3b0207f2),
	.w4(32'h3bafcc1a),
	.w5(32'h3bbe7fde),
	.w6(32'h3b110e56),
	.w7(32'h3b95e1c5),
	.w8(32'h3b2c3399),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2584d),
	.w1(32'h3d04a6e8),
	.w2(32'h3d213070),
	.w3(32'h3ce87a8d),
	.w4(32'h3cf246bb),
	.w5(32'h3d1232ca),
	.w6(32'h3cd45606),
	.w7(32'h3d1dc145),
	.w8(32'h3d284fbc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d313b29),
	.w1(32'hbc2d9faf),
	.w2(32'hbc432f67),
	.w3(32'hbc50c210),
	.w4(32'hbbaa8b77),
	.w5(32'hbaf58087),
	.w6(32'hbc5e2a39),
	.w7(32'hbc8972be),
	.w8(32'h3b589131),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9401d9b),
	.w1(32'hbb15d303),
	.w2(32'hbb9b8e26),
	.w3(32'h3aa64b55),
	.w4(32'hb91af272),
	.w5(32'h396ad538),
	.w6(32'h3b2d92d9),
	.w7(32'h3ab42e01),
	.w8(32'h3b97f847),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3e6f8),
	.w1(32'h3c13df4f),
	.w2(32'h3c26696a),
	.w3(32'h3af90891),
	.w4(32'h3934938b),
	.w5(32'hbbb467f7),
	.w6(32'h3a39afda),
	.w7(32'h3b6e6aa3),
	.w8(32'h3bb4b937),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc216746),
	.w1(32'hbc45eb20),
	.w2(32'hbc59a04a),
	.w3(32'h3a048e7e),
	.w4(32'hbb46b548),
	.w5(32'h3c9b504a),
	.w6(32'hbb85bcf8),
	.w7(32'hbc015694),
	.w8(32'h3c745dcc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40c519),
	.w1(32'hb8e6a820),
	.w2(32'hbb982d44),
	.w3(32'h3a98caef),
	.w4(32'hbb50bb13),
	.w5(32'hb90663f7),
	.w6(32'h3966baec),
	.w7(32'hbb75fcc9),
	.w8(32'hba187d02),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c0261),
	.w1(32'hbb15916e),
	.w2(32'hbbbf3d85),
	.w3(32'hbacc065a),
	.w4(32'h3b6e2c1c),
	.w5(32'hbb36e47d),
	.w6(32'h3c83b63a),
	.w7(32'h3ace10b3),
	.w8(32'hba5210c5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b222632),
	.w1(32'h3a295cb4),
	.w2(32'hba19edac),
	.w3(32'h3a5c093c),
	.w4(32'hbbc055ce),
	.w5(32'hba0e77bd),
	.w6(32'hbb4b38d1),
	.w7(32'hbc201af2),
	.w8(32'hbb47313b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d57dc),
	.w1(32'hb98e82ee),
	.w2(32'hbb919d5a),
	.w3(32'h38fe6347),
	.w4(32'hba8c61ce),
	.w5(32'hbb93f907),
	.w6(32'hba809b50),
	.w7(32'hbb81edc8),
	.w8(32'hbbc62ddc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46b687),
	.w1(32'hbba2c3de),
	.w2(32'hbb8eb0c5),
	.w3(32'hbbbdf44e),
	.w4(32'hbc1dd746),
	.w5(32'hbb555948),
	.w6(32'hbb7df9e4),
	.w7(32'hbc73fabf),
	.w8(32'hbc3dd345),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76322f),
	.w1(32'hbb1933e0),
	.w2(32'hbb44de52),
	.w3(32'hba1f1dc0),
	.w4(32'hbaccca39),
	.w5(32'h3a0b6d38),
	.w6(32'h3ab3ac5b),
	.w7(32'h3a57460e),
	.w8(32'h3bc166ef),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e5983),
	.w1(32'h3b1d8aa3),
	.w2(32'hbb4841af),
	.w3(32'h3b2ed272),
	.w4(32'hbb337123),
	.w5(32'hbba1c36c),
	.w6(32'h3b0f3457),
	.w7(32'hbb7b77ed),
	.w8(32'hbbc932fe),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ff589),
	.w1(32'h3bfae482),
	.w2(32'hbc1070aa),
	.w3(32'h3c47f58d),
	.w4(32'hbb2cf2f6),
	.w5(32'h3b9be1bf),
	.w6(32'h3c05e4b8),
	.w7(32'hbb78b7d8),
	.w8(32'hbbb658d7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcea99),
	.w1(32'hba762618),
	.w2(32'h3a4bf932),
	.w3(32'hbaf8df67),
	.w4(32'hba34dc50),
	.w5(32'hbb0d39cc),
	.w6(32'hbb06ddcb),
	.w7(32'hbacc4dc8),
	.w8(32'hbac20073),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2633ef),
	.w1(32'hbbc7a315),
	.w2(32'hbc135b9b),
	.w3(32'hbc143368),
	.w4(32'hbbd5c56a),
	.w5(32'hbb3e2711),
	.w6(32'hbc7ddb91),
	.w7(32'hbc2821c3),
	.w8(32'hb916ab89),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83df82),
	.w1(32'hbc1ac8db),
	.w2(32'hbc1009e4),
	.w3(32'hbc53777c),
	.w4(32'hbb9d4729),
	.w5(32'h3c814068),
	.w6(32'hbcaf883f),
	.w7(32'hbc037894),
	.w8(32'h3d1727ba),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d20f9c8),
	.w1(32'hbc2c30c7),
	.w2(32'hbbc0ae02),
	.w3(32'h3be120dd),
	.w4(32'h3b83285a),
	.w5(32'h3c66ede4),
	.w6(32'hbbdfc0d1),
	.w7(32'h3c4b5bb4),
	.w8(32'h3cc0e883),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0a84e),
	.w1(32'hbc813cef),
	.w2(32'hbc88e4a8),
	.w3(32'hbc2eef8b),
	.w4(32'hbcc61e92),
	.w5(32'hbc45dfb3),
	.w6(32'hbc27cc01),
	.w7(32'hbcb946f6),
	.w8(32'hbc3388ca),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af96090),
	.w1(32'h3b6a96d7),
	.w2(32'hbc44cac4),
	.w3(32'h3bb89b51),
	.w4(32'h38963b6e),
	.w5(32'hbb922b01),
	.w6(32'h3c02d833),
	.w7(32'hbb909808),
	.w8(32'hbbc2c331),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5937f9),
	.w1(32'hbc9444de),
	.w2(32'hbcb06ec5),
	.w3(32'hbc331d86),
	.w4(32'hbc928919),
	.w5(32'hbbd9a987),
	.w6(32'hbc4a651f),
	.w7(32'hbc837126),
	.w8(32'hbc261cfa),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1928a2),
	.w1(32'h3b59058e),
	.w2(32'h3ab5e1ff),
	.w3(32'hb9c246dd),
	.w4(32'hbad5b6a9),
	.w5(32'hba2c3098),
	.w6(32'h3ad659ed),
	.w7(32'hb9469020),
	.w8(32'hbbaf7997),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc08944),
	.w1(32'h3b06717d),
	.w2(32'hb9259f2f),
	.w3(32'h3ac6d2a4),
	.w4(32'h3a9938e7),
	.w5(32'h3aff84c5),
	.w6(32'hb92f5fd8),
	.w7(32'hbab7859d),
	.w8(32'hbaec0fcd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d1180),
	.w1(32'hbc3ecb33),
	.w2(32'hbcbdd433),
	.w3(32'hbb968723),
	.w4(32'hbc2e56ca),
	.w5(32'hbccf65f2),
	.w6(32'hbc1496b1),
	.w7(32'hbce46995),
	.w8(32'hbc1fcdd4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05d553),
	.w1(32'h3cb49f5d),
	.w2(32'h3a838f5c),
	.w3(32'h3b2cd2ea),
	.w4(32'hbc8ca0fc),
	.w5(32'hbd17679e),
	.w6(32'h3c940261),
	.w7(32'hbbf498e7),
	.w8(32'hbcc8065f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb871a2a),
	.w1(32'h3bfc2a47),
	.w2(32'hbcbbc613),
	.w3(32'h3bec260b),
	.w4(32'hbcd10cde),
	.w5(32'hbd6a67e7),
	.w6(32'h3bb68a60),
	.w7(32'hbd0454eb),
	.w8(32'hbd729eee),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3a2069),
	.w1(32'h3ad2d129),
	.w2(32'h3aceaa22),
	.w3(32'h3c5579f7),
	.w4(32'h3b905562),
	.w5(32'h3cb9e673),
	.w6(32'h3b33ded0),
	.w7(32'h3bc10fdc),
	.w8(32'h3d1a2edf),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c885e74),
	.w1(32'hbb20c68b),
	.w2(32'hbc9589c0),
	.w3(32'hbc35c6e9),
	.w4(32'hbcbcc03f),
	.w5(32'hbb6d5060),
	.w6(32'hba8cc68d),
	.w7(32'hbce65326),
	.w8(32'h3a8f98ad),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a574209),
	.w1(32'hba87048e),
	.w2(32'hbb06c3c3),
	.w3(32'hba476426),
	.w4(32'hbb3b2570),
	.w5(32'hbac50d42),
	.w6(32'hb9ba2fa4),
	.w7(32'hbb2b0a7a),
	.w8(32'h38433d57),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393eeb3f),
	.w1(32'h3b46cbb1),
	.w2(32'hbc1e4e35),
	.w3(32'hbb33b151),
	.w4(32'hbc3c2085),
	.w5(32'hbc35e9c0),
	.w6(32'h3b3aa1f5),
	.w7(32'hbc548f6c),
	.w8(32'hbc4834d1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe06046),
	.w1(32'hb9b6c3cd),
	.w2(32'hbb66adc7),
	.w3(32'hbb9c2da0),
	.w4(32'hbbe2eb4e),
	.w5(32'hbbc5079f),
	.w6(32'h3aa9f406),
	.w7(32'hbb95cbeb),
	.w8(32'hbb921578),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48a30c),
	.w1(32'h37dabf23),
	.w2(32'hb7648a1b),
	.w3(32'hbb0f11cb),
	.w4(32'hba1c7877),
	.w5(32'h3ad2de3d),
	.w6(32'hbb24bda0),
	.w7(32'hbb15da08),
	.w8(32'hbad62637),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f56530),
	.w1(32'h3a143976),
	.w2(32'h3bf9d1a4),
	.w3(32'h3ac5ceb2),
	.w4(32'h3ba04403),
	.w5(32'h3c85b072),
	.w6(32'h3b61767d),
	.w7(32'h3c3fbab8),
	.w8(32'h3bd75bb2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f2f37),
	.w1(32'h3c1b73b1),
	.w2(32'h3c0327a7),
	.w3(32'h3aaa1325),
	.w4(32'hbb904211),
	.w5(32'hbcd516c7),
	.w6(32'h3c784e08),
	.w7(32'h3bf9bccc),
	.w8(32'hbd255ba9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba309a7),
	.w1(32'hbc954c48),
	.w2(32'hbc641245),
	.w3(32'hbc80435b),
	.w4(32'h3b8913af),
	.w5(32'h3cabe307),
	.w6(32'hbc4d051a),
	.w7(32'hba3479a1),
	.w8(32'h3bc7aa27),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ac1d0),
	.w1(32'h3b3f423b),
	.w2(32'h3b2c23bc),
	.w3(32'hbb1104f3),
	.w4(32'hba20dee6),
	.w5(32'h3a62bbe9),
	.w6(32'hbb61fcf3),
	.w7(32'hbb0aa026),
	.w8(32'hbb33b2ff),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84a43a),
	.w1(32'hbbd21576),
	.w2(32'h3b83089c),
	.w3(32'hba7b48c1),
	.w4(32'h3b2f9b55),
	.w5(32'h3c81b62f),
	.w6(32'hbb2490d3),
	.w7(32'h3af60214),
	.w8(32'h3ca96a7c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca79f16),
	.w1(32'hbae6a5f0),
	.w2(32'hbb45c55d),
	.w3(32'hbba82957),
	.w4(32'hbacb2698),
	.w5(32'hbbad4a3d),
	.w6(32'hbbaa3059),
	.w7(32'hbc1157eb),
	.w8(32'hbc3c5415),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4421b),
	.w1(32'hbba65739),
	.w2(32'hbbf26cb0),
	.w3(32'hbb011e66),
	.w4(32'hbb25defa),
	.w5(32'hbbb2bb13),
	.w6(32'hbba46711),
	.w7(32'hbb4ed16c),
	.w8(32'hbbae130d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f38fb),
	.w1(32'hbc279750),
	.w2(32'hbc3d03c1),
	.w3(32'h3c3489ac),
	.w4(32'hb9645f33),
	.w5(32'hba6416b2),
	.w6(32'hbb612692),
	.w7(32'hbc72bd67),
	.w8(32'h3c61e14f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83423e),
	.w1(32'h3c0f5ce1),
	.w2(32'h3c3bc22c),
	.w3(32'h3b736471),
	.w4(32'hbaceb77c),
	.w5(32'hbbce0dc3),
	.w6(32'h3b8cec8a),
	.w7(32'h3ac47a4b),
	.w8(32'hbbf24fb8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc905195),
	.w1(32'hbb5e6fc5),
	.w2(32'hbba84b70),
	.w3(32'h3b7408dd),
	.w4(32'hbc48d377),
	.w5(32'h3b9fa21f),
	.w6(32'hbae9aaa5),
	.w7(32'hbc52fcbd),
	.w8(32'h3c19cd17),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6ebaf),
	.w1(32'hbb38c152),
	.w2(32'hbbb021ea),
	.w3(32'hbb1ee338),
	.w4(32'hbc1db3b0),
	.w5(32'hbc32cb33),
	.w6(32'hbb8bf126),
	.w7(32'hbc2eb9c0),
	.w8(32'hbc4c87e9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb8993),
	.w1(32'h3c9bb437),
	.w2(32'hbbd68ecd),
	.w3(32'hbb452028),
	.w4(32'hbc2b7158),
	.w5(32'hbc6b987d),
	.w6(32'h3c7f8d16),
	.w7(32'h3b0333f3),
	.w8(32'hbbf23d31),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abccaf8),
	.w1(32'hbb9a1305),
	.w2(32'hbc1caae7),
	.w3(32'hb9d3f23d),
	.w4(32'hbb82ce6e),
	.w5(32'hbb04841b),
	.w6(32'hbb30919e),
	.w7(32'hbbb44347),
	.w8(32'hbb273843),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcb283),
	.w1(32'h3a97f3db),
	.w2(32'h3baccbe3),
	.w3(32'h3a50eafa),
	.w4(32'h3bf3eed3),
	.w5(32'h3c661b26),
	.w6(32'h39a9b34f),
	.w7(32'h3bee684c),
	.w8(32'h3c74176f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c135248),
	.w1(32'hbb3e8d91),
	.w2(32'hbc061e88),
	.w3(32'hba96a638),
	.w4(32'hbbdbf420),
	.w5(32'hbb8fd85e),
	.w6(32'hbb2f092c),
	.w7(32'hbbab5072),
	.w8(32'hbba8ea7d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3100ca),
	.w1(32'hbada547f),
	.w2(32'hbb0b4add),
	.w3(32'hbaa13ac3),
	.w4(32'hbb4be108),
	.w5(32'hb84d2433),
	.w6(32'hbc3a5417),
	.w7(32'hbc3ff466),
	.w8(32'hbc49b016),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7113b),
	.w1(32'hbc0ac410),
	.w2(32'hbc00ddb4),
	.w3(32'hba635000),
	.w4(32'hbb60bdc4),
	.w5(32'hb98d04b0),
	.w6(32'hbbb2fc34),
	.w7(32'hbc092a69),
	.w8(32'hbbe6b590),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaafb2f),
	.w1(32'h3b76c2a1),
	.w2(32'h3bc4f768),
	.w3(32'h3a5e660c),
	.w4(32'h394e8fb3),
	.w5(32'h3b5f40b0),
	.w6(32'hbc0929c5),
	.w7(32'hbc39334d),
	.w8(32'hbb8a8fa3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c94e8),
	.w1(32'h3c1bc12f),
	.w2(32'h3b9fb4e1),
	.w3(32'h3c0c2277),
	.w4(32'h3bd294a7),
	.w5(32'hba0bcef6),
	.w6(32'h3b9e29af),
	.w7(32'h3b9a0e71),
	.w8(32'h3a557d8a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbde1e),
	.w1(32'h39cc17fb),
	.w2(32'hbb68810e),
	.w3(32'hba378039),
	.w4(32'hbb4aa0dc),
	.w5(32'hbb79f943),
	.w6(32'hbc0ed871),
	.w7(32'hbb8aaf0f),
	.w8(32'hbc6894e9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8c946),
	.w1(32'h3b8ce122),
	.w2(32'h3a9d2868),
	.w3(32'h3b19c8d6),
	.w4(32'h3b1e1066),
	.w5(32'hba705144),
	.w6(32'hbb977e17),
	.w7(32'hbbafa135),
	.w8(32'hbc35f632),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b2120),
	.w1(32'h3c2cb956),
	.w2(32'h3c3c9429),
	.w3(32'hbca22a0e),
	.w4(32'hbcfaad98),
	.w5(32'hbb86d4b8),
	.w6(32'hbc5bc62e),
	.w7(32'hbcfc45c1),
	.w8(32'hbb94a353),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96cf47),
	.w1(32'h3b5441d3),
	.w2(32'h3b1dae27),
	.w3(32'h3bf6a63b),
	.w4(32'h3c9ca00d),
	.w5(32'h3c0f9531),
	.w6(32'h3bdee6f1),
	.w7(32'h3c9f296f),
	.w8(32'h3be2d4b9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7475b0),
	.w1(32'hbb8c00d8),
	.w2(32'hbc477e26),
	.w3(32'hbb1e495c),
	.w4(32'hbc49a230),
	.w5(32'hbc83b1b6),
	.w6(32'hbb558855),
	.w7(32'hbc6361e6),
	.w8(32'hbc9a6590),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb37bb),
	.w1(32'hba8b4feb),
	.w2(32'hbc413e6c),
	.w3(32'hbc38f913),
	.w4(32'hbc992562),
	.w5(32'h39a00e7d),
	.w6(32'h3bcb4f37),
	.w7(32'hbc2c3028),
	.w8(32'h3bbdb6cc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1db64e),
	.w1(32'h3c3990c9),
	.w2(32'hbaa2c5a7),
	.w3(32'h3b8e9e98),
	.w4(32'hba6816cc),
	.w5(32'hbbb45590),
	.w6(32'h3aebb99c),
	.w7(32'hbc11963c),
	.w8(32'hbc8b43ba),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule