module layer_10_featuremap_333(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7b523),
	.w1(32'hbbd52e7c),
	.w2(32'h392822e4),
	.w3(32'hbbd62b56),
	.w4(32'hbbe1a9d2),
	.w5(32'h3a579870),
	.w6(32'hbb78e790),
	.w7(32'hbaf8ae51),
	.w8(32'hbb9cb822),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee1257),
	.w1(32'hbb894012),
	.w2(32'hbbc99092),
	.w3(32'hba87e2f5),
	.w4(32'hbb9646d2),
	.w5(32'h3a3ae482),
	.w6(32'h3a716f9e),
	.w7(32'hbbae0f0d),
	.w8(32'hb94aae13),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cb042),
	.w1(32'hbadc29da),
	.w2(32'h3a8cb102),
	.w3(32'hb86fc4c5),
	.w4(32'hbb68fac8),
	.w5(32'h3baa2e8a),
	.w6(32'h39cd102b),
	.w7(32'h3b077465),
	.w8(32'h3b8afde5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc32cf6),
	.w1(32'h3bd3a31c),
	.w2(32'h3b894b49),
	.w3(32'h3b6ddde1),
	.w4(32'h3b77f809),
	.w5(32'hb8eb9d12),
	.w6(32'h3b0e5695),
	.w7(32'h3ac4f3aa),
	.w8(32'h3b1b7dff),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad73001),
	.w1(32'hbb9e5d95),
	.w2(32'hba57bdc7),
	.w3(32'hbba45943),
	.w4(32'hbb84fcad),
	.w5(32'hb914ccdc),
	.w6(32'hbb83554c),
	.w7(32'hba8cb54d),
	.w8(32'h3b521ca1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb44480),
	.w1(32'h3b938a11),
	.w2(32'h3b9ef758),
	.w3(32'hb96fd570),
	.w4(32'hbab91906),
	.w5(32'h3a89ffe7),
	.w6(32'h3b20f14f),
	.w7(32'h3aed1151),
	.w8(32'hbb1a4e25),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5095a2),
	.w1(32'h3af57dc6),
	.w2(32'hbbe7ded1),
	.w3(32'h39747046),
	.w4(32'h3b5bb29f),
	.w5(32'hbc1202c7),
	.w6(32'hbb357b5d),
	.w7(32'hba142197),
	.w8(32'hbba09765),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec6b4f),
	.w1(32'hbb99de1b),
	.w2(32'hbbd1951d),
	.w3(32'h3b4041b2),
	.w4(32'h3bdf43d2),
	.w5(32'h3b3b1640),
	.w6(32'hbb94d949),
	.w7(32'hbc1833d8),
	.w8(32'hba594c51),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e3666),
	.w1(32'h3b0a6836),
	.w2(32'h3b2a75f3),
	.w3(32'hba4c9b64),
	.w4(32'hb87a19bd),
	.w5(32'hb9bd7a3e),
	.w6(32'h3b3af1bd),
	.w7(32'h3b0be9fe),
	.w8(32'h3b656f0f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd20a18),
	.w1(32'h3b28b116),
	.w2(32'h3ad77d02),
	.w3(32'h397b66c2),
	.w4(32'hba92de8e),
	.w5(32'hbb638849),
	.w6(32'h3adce02a),
	.w7(32'h3b2bf574),
	.w8(32'h3b2f3200),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf74421),
	.w1(32'h3c06eb4f),
	.w2(32'h3c035027),
	.w3(32'h3a917f81),
	.w4(32'h39298003),
	.w5(32'hbb5209c3),
	.w6(32'h3b59302b),
	.w7(32'h3b1a703d),
	.w8(32'h3ab6de88),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5e4ae),
	.w1(32'h39ec53e5),
	.w2(32'hbc182fc5),
	.w3(32'hbbbd8aca),
	.w4(32'h3a0cc4f7),
	.w5(32'hbbd4c784),
	.w6(32'hb9698658),
	.w7(32'h39230fda),
	.w8(32'h3b8b5a3e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1915a),
	.w1(32'hbabbe58c),
	.w2(32'hbbbf3508),
	.w3(32'hba3cb180),
	.w4(32'hbb07a06e),
	.w5(32'hbbae6b6b),
	.w6(32'h3b9ab122),
	.w7(32'h3bc68c49),
	.w8(32'hbb91b516),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d49b1),
	.w1(32'hbb83af72),
	.w2(32'hbb80e9c4),
	.w3(32'h3b0fe3d1),
	.w4(32'hba1fab50),
	.w5(32'h3aa0f204),
	.w6(32'hb9e1bebd),
	.w7(32'hbaa286ae),
	.w8(32'hbaee4d52),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8faa2c),
	.w1(32'h3b9bb78d),
	.w2(32'h3b6c3778),
	.w3(32'h3b2a3088),
	.w4(32'h39c4dbf9),
	.w5(32'hbb26d8f4),
	.w6(32'h3a43afa0),
	.w7(32'hbadebdb9),
	.w8(32'hbb7c7f81),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65f58b),
	.w1(32'hbbd212ad),
	.w2(32'hbb296cc6),
	.w3(32'h3bc518de),
	.w4(32'hbbc638c4),
	.w5(32'hbb4d8dfb),
	.w6(32'h3b7a148a),
	.w7(32'h3b896cf9),
	.w8(32'h3b1a5868),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2a3bc),
	.w1(32'h3c1e8455),
	.w2(32'h3bef6e02),
	.w3(32'hb9d980c9),
	.w4(32'h3abb3c47),
	.w5(32'h3a881bcd),
	.w6(32'h3bb4d896),
	.w7(32'h3b545254),
	.w8(32'h3a2ad035),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace6806),
	.w1(32'hbb28f93a),
	.w2(32'hbc1a7546),
	.w3(32'h3ba33159),
	.w4(32'h3b97b89a),
	.w5(32'hbbb93529),
	.w6(32'hbad98e9b),
	.w7(32'h3b6cc4ad),
	.w8(32'hbb7d659e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2afd1c),
	.w1(32'hb8578d31),
	.w2(32'hbb8c35bb),
	.w3(32'h3a4358f9),
	.w4(32'h3abe521f),
	.w5(32'hbba0c9a2),
	.w6(32'hbab0fb96),
	.w7(32'h3b6fb038),
	.w8(32'hbacdf864),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8a5b3),
	.w1(32'hba53d7aa),
	.w2(32'hb9850bf9),
	.w3(32'h3a8a8ee7),
	.w4(32'h3b299a1d),
	.w5(32'hba9e2f6b),
	.w6(32'hbabbb9b0),
	.w7(32'h3a8c8cee),
	.w8(32'h3a6dc029),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c9a5b),
	.w1(32'hbb12d544),
	.w2(32'h3b1f5d6f),
	.w3(32'h3b00818d),
	.w4(32'h3a0285a8),
	.w5(32'h3ba361df),
	.w6(32'h38de2b93),
	.w7(32'h3b9693fd),
	.w8(32'h3b6e124a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe6a9b),
	.w1(32'h3c04af1d),
	.w2(32'h3c08a432),
	.w3(32'h3b7b0d1e),
	.w4(32'h3bee5088),
	.w5(32'hbacc4609),
	.w6(32'h3a5996e0),
	.w7(32'h3aaed258),
	.w8(32'hbb0938d8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d6742),
	.w1(32'h3bcba337),
	.w2(32'hbbc5d728),
	.w3(32'h3b029575),
	.w4(32'h3afd6777),
	.w5(32'hbbc1c473),
	.w6(32'h3b330c40),
	.w7(32'h3b560a04),
	.w8(32'hbbbf8431),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab7ab0),
	.w1(32'hbb116cb8),
	.w2(32'hbb9b946e),
	.w3(32'h3acbaa30),
	.w4(32'hbc0d9fd1),
	.w5(32'h3a54073b),
	.w6(32'h39e98092),
	.w7(32'hbb7ca210),
	.w8(32'hbb3ff6ab),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc6444),
	.w1(32'h399bffc2),
	.w2(32'h3b4ff8b6),
	.w3(32'hbb092e87),
	.w4(32'hba9abc44),
	.w5(32'h3c07dcda),
	.w6(32'hbb79e04a),
	.w7(32'hbb22575a),
	.w8(32'h3a5dcfdb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89c88a),
	.w1(32'h3b7eccd7),
	.w2(32'h3bbfdd71),
	.w3(32'h3a04ab98),
	.w4(32'h3b20f0ea),
	.w5(32'h3a81c2e6),
	.w6(32'hbb6dde8d),
	.w7(32'hb9eb0f53),
	.w8(32'h3aac286c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab37fe),
	.w1(32'h3b0dad0d),
	.w2(32'h3b92bfc3),
	.w3(32'hb9a45cb7),
	.w4(32'h3b8ce9d5),
	.w5(32'hbad8cac3),
	.w6(32'hbaf470c5),
	.w7(32'h3b3b599d),
	.w8(32'h3b54907a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca37f),
	.w1(32'hbade604c),
	.w2(32'h3bc92509),
	.w3(32'hbc414c19),
	.w4(32'hba220aa0),
	.w5(32'hbb8bdec5),
	.w6(32'hbb4ceac3),
	.w7(32'h3c0da1cf),
	.w8(32'hbaba40a2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb976026),
	.w1(32'hbb68db4b),
	.w2(32'hbb519961),
	.w3(32'h3af473d8),
	.w4(32'h3ace8b4a),
	.w5(32'hba288402),
	.w6(32'hbb92ae75),
	.w7(32'hbb0088c3),
	.w8(32'hb9f8e292),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20ad0e),
	.w1(32'hbb2be7e4),
	.w2(32'hb9fa98f9),
	.w3(32'hba89b5aa),
	.w4(32'hbaa65f68),
	.w5(32'h3a4f219f),
	.w6(32'hbaf1df98),
	.w7(32'hbb1668c5),
	.w8(32'hbb951010),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21132c),
	.w1(32'hbc584e27),
	.w2(32'hbc399da6),
	.w3(32'h3b228524),
	.w4(32'h3ab27ac8),
	.w5(32'hbb70c542),
	.w6(32'hbbaf3315),
	.w7(32'hbbb7c094),
	.w8(32'h3b5711a3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80c21a),
	.w1(32'h3ae37d9c),
	.w2(32'h3b4efb71),
	.w3(32'hbbaee4db),
	.w4(32'hbbd10a78),
	.w5(32'hb987f6ad),
	.w6(32'h399b43bd),
	.w7(32'hbb37732b),
	.w8(32'hba8ce98a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f892e),
	.w1(32'hbb80b58d),
	.w2(32'hbb5ada63),
	.w3(32'h3a287b5f),
	.w4(32'h3bd687ad),
	.w5(32'h39797741),
	.w6(32'hbb8b91b3),
	.w7(32'hbb6eecab),
	.w8(32'hbaaa94a0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13b3dd),
	.w1(32'h3a34a684),
	.w2(32'hba30aa3c),
	.w3(32'h3ab01add),
	.w4(32'hb94bf2ba),
	.w5(32'h393d70c0),
	.w6(32'h3b0915ec),
	.w7(32'hbae878cc),
	.w8(32'hbb49afb9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c32caa),
	.w1(32'hbb21ca85),
	.w2(32'hba0266e2),
	.w3(32'h393e8b8b),
	.w4(32'h3ba6fbd6),
	.w5(32'hba590d91),
	.w6(32'hbacdd90c),
	.w7(32'h3ac3f0df),
	.w8(32'hba44428c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5a5bc),
	.w1(32'hba112a77),
	.w2(32'hbb87bf49),
	.w3(32'h39bf7abc),
	.w4(32'h3abdbc69),
	.w5(32'h3ba916d6),
	.w6(32'hbabd5be3),
	.w7(32'h3b7a491f),
	.w8(32'hbbded0a4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc787d08),
	.w1(32'h3be44fb6),
	.w2(32'hbc765ea2),
	.w3(32'hbbbadea8),
	.w4(32'h3c9e6bb2),
	.w5(32'hbb3f88c1),
	.w6(32'hbc2fcc8d),
	.w7(32'hbc42f23a),
	.w8(32'h3b8af14f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde4c6c),
	.w1(32'h3b23b74e),
	.w2(32'h3ca6315e),
	.w3(32'hbbbdf5d3),
	.w4(32'h3a43f589),
	.w5(32'h39e57181),
	.w6(32'hbb791f51),
	.w7(32'h3c0f5585),
	.w8(32'h3a00b7c6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0666ac),
	.w1(32'hbba7d328),
	.w2(32'h3a756328),
	.w3(32'hbc59eed5),
	.w4(32'hbc36f7cd),
	.w5(32'h3b9a78c3),
	.w6(32'hbb9200df),
	.w7(32'hba168cf8),
	.w8(32'h3ae303ae),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8b835),
	.w1(32'h3bc58e4e),
	.w2(32'h3c0a833a),
	.w3(32'hbae56fa4),
	.w4(32'h3aa840cb),
	.w5(32'hbb27e051),
	.w6(32'hbaf8a1aa),
	.w7(32'h3a833dc0),
	.w8(32'hbb89094e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5f939),
	.w1(32'hbb583abe),
	.w2(32'hbb6bb4cb),
	.w3(32'hbb31abfb),
	.w4(32'hbb3f2c55),
	.w5(32'h3a882023),
	.w6(32'hbaa8f2b3),
	.w7(32'hbb247226),
	.w8(32'hba011dd0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b982909),
	.w1(32'h3bab5cf7),
	.w2(32'h3bc77f5c),
	.w3(32'hbb071088),
	.w4(32'h3b36031b),
	.w5(32'hbb1c05e4),
	.w6(32'hbbbe7ed9),
	.w7(32'hba421703),
	.w8(32'hba9e2f8b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7519b9),
	.w1(32'hbbee6b7c),
	.w2(32'hbb109db7),
	.w3(32'hbb137dff),
	.w4(32'hbb0f6afb),
	.w5(32'hbab31df5),
	.w6(32'hbb31376b),
	.w7(32'h3b60ba60),
	.w8(32'h3af0623d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72a946),
	.w1(32'hbbc8ed07),
	.w2(32'hbc2c1d72),
	.w3(32'hba074b11),
	.w4(32'hbb15379f),
	.w5(32'hbbb6b885),
	.w6(32'h3b5592f3),
	.w7(32'h3c040bfa),
	.w8(32'hbaa7d695),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8d6a8),
	.w1(32'h3b3a4793),
	.w2(32'h3b5f29dd),
	.w3(32'hbb93c802),
	.w4(32'hb943c5ac),
	.w5(32'h3b04b218),
	.w6(32'hbbf2522c),
	.w7(32'hbb8f34f7),
	.w8(32'hbb05b868),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb39b1),
	.w1(32'h3c3a8dd9),
	.w2(32'h3b405e2c),
	.w3(32'h398e5aeb),
	.w4(32'h3a848401),
	.w5(32'h3ad88f98),
	.w6(32'h3b6d46d8),
	.w7(32'hbaffb7fc),
	.w8(32'hbbd61245),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b242524),
	.w1(32'h3b198d74),
	.w2(32'h3b5de39f),
	.w3(32'hb988931e),
	.w4(32'hbacd0603),
	.w5(32'h3b3fb107),
	.w6(32'h39c5b942),
	.w7(32'h3a7f353d),
	.w8(32'h3b97bdec),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93543c),
	.w1(32'h3bbe9cd0),
	.w2(32'hbb4c676f),
	.w3(32'h3c0c6050),
	.w4(32'h3c4e3415),
	.w5(32'hbba92649),
	.w6(32'h3b99bfaa),
	.w7(32'h3c02276e),
	.w8(32'hba053e8e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8057d8),
	.w1(32'hbbb5a437),
	.w2(32'hbbc3e5c9),
	.w3(32'h3a4769ba),
	.w4(32'hbb3cc72e),
	.w5(32'h3b20e5ac),
	.w6(32'hb9f052a2),
	.w7(32'hba8f60d5),
	.w8(32'h3a138ede),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13ae58),
	.w1(32'h3bdbfeb4),
	.w2(32'h3c08e88b),
	.w3(32'h3b2a8a77),
	.w4(32'h3c0c5bcd),
	.w5(32'h3b789272),
	.w6(32'hbb9b4248),
	.w7(32'h39bdcbd8),
	.w8(32'h3be532ea),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922492f),
	.w1(32'hbbb4be28),
	.w2(32'hbbaf0a9f),
	.w3(32'hbb0d6c61),
	.w4(32'hbb5fb076),
	.w5(32'hb9832701),
	.w6(32'h3a837e29),
	.w7(32'hbab68482),
	.w8(32'h3b7aa7bd),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18990b),
	.w1(32'hbabe9226),
	.w2(32'hbb8036e3),
	.w3(32'hbb4f168f),
	.w4(32'hbafa4ea4),
	.w5(32'hbac5e933),
	.w6(32'hb9a81454),
	.w7(32'h3a7e1ad0),
	.w8(32'hbb157a2c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42eed0),
	.w1(32'h39bd5e5a),
	.w2(32'h3ac3cd9f),
	.w3(32'hba3fde70),
	.w4(32'hba36eedd),
	.w5(32'hba1d9644),
	.w6(32'h3ab9c499),
	.w7(32'h3b06d299),
	.w8(32'hbbbb8392),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4002cc),
	.w1(32'hbba54001),
	.w2(32'hbc2b95e4),
	.w3(32'h3c1196b0),
	.w4(32'h3bf67c5d),
	.w5(32'hbc317035),
	.w6(32'hbae25f66),
	.w7(32'h3b9f72f4),
	.w8(32'h390b3a30),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad677b4),
	.w1(32'hba765b19),
	.w2(32'hbb21b666),
	.w3(32'hbb58f854),
	.w4(32'hba5471dc),
	.w5(32'hba7e7dbf),
	.w6(32'hba250aff),
	.w7(32'h3acbae28),
	.w8(32'hb91c7df6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01dd17),
	.w1(32'h38f26ea0),
	.w2(32'h3afa23a7),
	.w3(32'h3aadfb26),
	.w4(32'h3ad2d3e2),
	.w5(32'hb9cac47a),
	.w6(32'h38aa9e0d),
	.w7(32'h3a43cd3b),
	.w8(32'hbad220f3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba643665),
	.w1(32'h3a812da8),
	.w2(32'hb615a05e),
	.w3(32'h3a2f496f),
	.w4(32'h38a8055f),
	.w5(32'hbb8c8012),
	.w6(32'h3aea37a5),
	.w7(32'h3a2e1c6a),
	.w8(32'hbbb32448),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfb7fd),
	.w1(32'hbb84893f),
	.w2(32'hbaa7681c),
	.w3(32'h3a50e891),
	.w4(32'h3b1b3ba4),
	.w5(32'h3b2eae07),
	.w6(32'hbb2c068e),
	.w7(32'h3ae75982),
	.w8(32'h3a875bb7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf029f),
	.w1(32'h3ba06c24),
	.w2(32'h3c00f83b),
	.w3(32'hba456821),
	.w4(32'h3badd57c),
	.w5(32'h3a83e686),
	.w6(32'hbbc57b55),
	.w7(32'h39a11bf8),
	.w8(32'h3b456243),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7f4d3),
	.w1(32'h3c61a3c7),
	.w2(32'h3c35b586),
	.w3(32'h3ac17b02),
	.w4(32'h3c007752),
	.w5(32'hbb858f59),
	.w6(32'h3b14ca68),
	.w7(32'h3bbfc6fa),
	.w8(32'hba9df89b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadeb5d8),
	.w1(32'hbb3633f4),
	.w2(32'hbb930429),
	.w3(32'hbad5636c),
	.w4(32'hbb167d60),
	.w5(32'hbb70dbfb),
	.w6(32'h39478946),
	.w7(32'h3afca7d7),
	.w8(32'hbad7a86c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9333cd),
	.w1(32'h3b7b7b01),
	.w2(32'hbb25af0c),
	.w3(32'h391d3f83),
	.w4(32'hbb8a4bee),
	.w5(32'hbb45af0f),
	.w6(32'hbaaa912e),
	.w7(32'hbb50159b),
	.w8(32'h3b253446),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb249777),
	.w1(32'hbb94ca20),
	.w2(32'hbb6aa3d6),
	.w3(32'hbad46b49),
	.w4(32'hbad538ca),
	.w5(32'hbac4701a),
	.w6(32'h3afed2d3),
	.w7(32'h3b62c8ad),
	.w8(32'hbb510d29),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08e50e),
	.w1(32'hbb61a354),
	.w2(32'hba48597e),
	.w3(32'h3a496858),
	.w4(32'h3b196e99),
	.w5(32'hbaecfc23),
	.w6(32'hbb325c9e),
	.w7(32'h39db9409),
	.w8(32'h391bd6ef),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb843473a),
	.w1(32'hbb8ae1b7),
	.w2(32'hbb96eb96),
	.w3(32'hb8d2686d),
	.w4(32'hba8cdc24),
	.w5(32'hbbbecdaa),
	.w6(32'hbaf9eae3),
	.w7(32'hbaf3d892),
	.w8(32'h3ba63977),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28ba43),
	.w1(32'hbad30df2),
	.w2(32'h3a3d72cc),
	.w3(32'hbbad91b9),
	.w4(32'hbbd46e0b),
	.w5(32'hbb607d7e),
	.w6(32'h3b836963),
	.w7(32'h3b808263),
	.w8(32'hbba85475),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a4b0b),
	.w1(32'hbc2a2cbf),
	.w2(32'hbc72981f),
	.w3(32'h3a8664f1),
	.w4(32'hbb1b8d31),
	.w5(32'hbb573d47),
	.w6(32'h3b7b85c6),
	.w7(32'hb9f65078),
	.w8(32'h3b6874a2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28bde6),
	.w1(32'h3a97da53),
	.w2(32'hbbb91ca2),
	.w3(32'h3c06f7e0),
	.w4(32'h3c3a734b),
	.w5(32'h3bbf1638),
	.w6(32'h3c18411d),
	.w7(32'h3ba61d87),
	.w8(32'hbb1759a0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb41d6e),
	.w1(32'hbb1c851a),
	.w2(32'hbb6f079b),
	.w3(32'hbab8df9b),
	.w4(32'hbb674f70),
	.w5(32'hbb16f98f),
	.w6(32'hbb9ce174),
	.w7(32'hbadaa8b3),
	.w8(32'hbb699093),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b170a53),
	.w1(32'h3b854f2c),
	.w2(32'h3b9ac338),
	.w3(32'hbbbf05d6),
	.w4(32'hbb9a5d3d),
	.w5(32'h3ba9f167),
	.w6(32'hbb6b3ce2),
	.w7(32'hba9c4dd4),
	.w8(32'hbb937de1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bd4ae),
	.w1(32'hbb6f439e),
	.w2(32'h3a5109c6),
	.w3(32'h3a6ca3e2),
	.w4(32'h3b98fba4),
	.w5(32'hbb44b0ec),
	.w6(32'hbba8238e),
	.w7(32'hba0c3a99),
	.w8(32'hbb40e984),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbcbf6),
	.w1(32'hbb7b3859),
	.w2(32'h3985f965),
	.w3(32'hbb040ce5),
	.w4(32'hbba6f4ae),
	.w5(32'hb7d25e78),
	.w6(32'h38117c41),
	.w7(32'h3a24de5d),
	.w8(32'h3b9c9964),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39933dfc),
	.w1(32'h3b829e18),
	.w2(32'h3b986992),
	.w3(32'hb99b9f43),
	.w4(32'hbb6bf4a1),
	.w5(32'h3a3147c6),
	.w6(32'h3b5269bb),
	.w7(32'h3b55f25c),
	.w8(32'hbb4cf05c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e5515),
	.w1(32'hbb94b6d5),
	.w2(32'hbbf6446a),
	.w3(32'h3b2a2913),
	.w4(32'h3b0e3c23),
	.w5(32'hbbd2f465),
	.w6(32'hbaa2b843),
	.w7(32'hb9c86375),
	.w8(32'h3b43382c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39dd4c),
	.w1(32'h3b25986a),
	.w2(32'h3b49c08b),
	.w3(32'hb7efee12),
	.w4(32'hba31b91b),
	.w5(32'hba206685),
	.w6(32'h3c107e6c),
	.w7(32'h3ba4fee8),
	.w8(32'h3a5637d9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb61945),
	.w1(32'hbbb34dd4),
	.w2(32'hbc228af4),
	.w3(32'h3a664b49),
	.w4(32'hba85f086),
	.w5(32'hbbb6a37a),
	.w6(32'h3b86709e),
	.w7(32'h3aec5e3a),
	.w8(32'hbac58a0f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdd3bc),
	.w1(32'h3921403b),
	.w2(32'hbba55142),
	.w3(32'h3b002d80),
	.w4(32'h3bc257dc),
	.w5(32'hbbb71fcd),
	.w6(32'h3b3db825),
	.w7(32'h3aa37ae7),
	.w8(32'hbb1bc353),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ed4e1a),
	.w1(32'hba25f582),
	.w2(32'hb979fdd7),
	.w3(32'hbbe3db9c),
	.w4(32'hbbb2165e),
	.w5(32'h3add4f80),
	.w6(32'hbbb342e9),
	.w7(32'hbb87d9d6),
	.w8(32'h37adf644),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba23e52),
	.w1(32'h3b79bfd7),
	.w2(32'h3a3062ef),
	.w3(32'h3b69f61e),
	.w4(32'h398ecbbe),
	.w5(32'h39fa5653),
	.w6(32'h3bdd1538),
	.w7(32'h3b787afa),
	.w8(32'h3a990b26),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dc06a),
	.w1(32'h3b5064f6),
	.w2(32'hbb99507f),
	.w3(32'h3b0204c0),
	.w4(32'hb9d0c9bb),
	.w5(32'hbc1fc784),
	.w6(32'h3be1d490),
	.w7(32'h39dcf624),
	.w8(32'hbc08bb0c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd60656),
	.w1(32'hbc12c4be),
	.w2(32'hbbec936d),
	.w3(32'hbb01f003),
	.w4(32'hbb4d7d00),
	.w5(32'hb94a8b1e),
	.w6(32'hbb5fae10),
	.w7(32'hbb472460),
	.w8(32'hbb3e6679),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb030c30),
	.w1(32'hbaafe2f0),
	.w2(32'hbb9286a0),
	.w3(32'h3adfdd17),
	.w4(32'h3adeb624),
	.w5(32'hbb2e39c1),
	.w6(32'hbb17daf8),
	.w7(32'h39fb606b),
	.w8(32'hba12b8bb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c153c),
	.w1(32'hbb2e4967),
	.w2(32'hbae4eab9),
	.w3(32'hba771a25),
	.w4(32'hbb49caaa),
	.w5(32'h3be1f04a),
	.w6(32'hbb147ec6),
	.w7(32'hbb285874),
	.w8(32'h3c4d9293),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c587dc9),
	.w1(32'h3c1b595d),
	.w2(32'h3c363b60),
	.w3(32'h3b82ceb1),
	.w4(32'h3b14f320),
	.w5(32'hbac58e8b),
	.w6(32'h3c46f4be),
	.w7(32'h3c2fdf18),
	.w8(32'hbb117cdb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a001a33),
	.w1(32'hbaa3b55a),
	.w2(32'hba19011c),
	.w3(32'hbb14edf1),
	.w4(32'hbb093030),
	.w5(32'hbb4f9d86),
	.w6(32'hbb67eb6e),
	.w7(32'hbb3467ea),
	.w8(32'h3afb794b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c1d68),
	.w1(32'h3bc0bb79),
	.w2(32'h3bbcd81f),
	.w3(32'hba768466),
	.w4(32'hbc01a843),
	.w5(32'hbaef915b),
	.w6(32'h3b8fd112),
	.w7(32'h3a5ee95b),
	.w8(32'hbb622030),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7aa8d),
	.w1(32'h3b7120e0),
	.w2(32'h3b79dff4),
	.w3(32'hbb648177),
	.w4(32'hbb8fff55),
	.w5(32'hba8ad21e),
	.w6(32'hbbeb80b4),
	.w7(32'hbb11cb91),
	.w8(32'hb999b240),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a57d69),
	.w1(32'hb9c107ce),
	.w2(32'h3a9b0a32),
	.w3(32'hbb211292),
	.w4(32'hba047729),
	.w5(32'h3adae950),
	.w6(32'h3ac3fa90),
	.w7(32'h3b32bb56),
	.w8(32'h3ac3bd14),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba046fc),
	.w1(32'h3bd7d2fd),
	.w2(32'h3b397f74),
	.w3(32'hb9284cc6),
	.w4(32'h3b1a7315),
	.w5(32'h3ba2ed7e),
	.w6(32'hb9c6740c),
	.w7(32'hbade88cd),
	.w8(32'hbacb0479),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f05721),
	.w1(32'hbb33e168),
	.w2(32'hbbc2f2b8),
	.w3(32'h3b96d8d0),
	.w4(32'h3b18dd71),
	.w5(32'h39a7e09a),
	.w6(32'h3a7952d8),
	.w7(32'hba9130fc),
	.w8(32'h3a7eb43f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e85e6),
	.w1(32'h398a525f),
	.w2(32'h37f6e93f),
	.w3(32'hbb5e591f),
	.w4(32'hbb8a74cd),
	.w5(32'h3b4e0426),
	.w6(32'h3b01b4b0),
	.w7(32'hbb8347a6),
	.w8(32'h3b597f54),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca990e),
	.w1(32'h38100968),
	.w2(32'hbc525c81),
	.w3(32'h3c07acf6),
	.w4(32'h3b03a7f0),
	.w5(32'hbc5890f1),
	.w6(32'h3b9152d2),
	.w7(32'hbb652279),
	.w8(32'hbbeeba73),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11de9d),
	.w1(32'h3b58653f),
	.w2(32'h3ba35361),
	.w3(32'hbc03971c),
	.w4(32'h39a16376),
	.w5(32'h3b2a5785),
	.w6(32'hbc45dc56),
	.w7(32'hbbbd575a),
	.w8(32'h3ba191b1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55a4f1),
	.w1(32'hbb6e37d2),
	.w2(32'hbbbb3038),
	.w3(32'h3bd9baa8),
	.w4(32'h3a0c1fe9),
	.w5(32'hbb9a5b4c),
	.w6(32'h3ba147fd),
	.w7(32'h3b7b9f08),
	.w8(32'hbacea64a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17699c),
	.w1(32'hbbcc3a47),
	.w2(32'h3b1b67c5),
	.w3(32'hbb15e415),
	.w4(32'hbb719349),
	.w5(32'hbc38be01),
	.w6(32'hbb75995b),
	.w7(32'h3a7bbcc5),
	.w8(32'h3bc8cdfe),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf18cf9),
	.w1(32'hbbcd5cec),
	.w2(32'h3bf6d6d3),
	.w3(32'hbc0dd508),
	.w4(32'hbbcbe1a8),
	.w5(32'h3b890dfb),
	.w6(32'h3b405db1),
	.w7(32'h3c0d282f),
	.w8(32'h3b78554f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48065f),
	.w1(32'h3b468cea),
	.w2(32'hbaf34c7a),
	.w3(32'h39ee2f05),
	.w4(32'hbb4f26bd),
	.w5(32'h3b830945),
	.w6(32'h3bca123f),
	.w7(32'h3ad12b4a),
	.w8(32'h3b087b0c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16f753),
	.w1(32'hbaa5c30e),
	.w2(32'hbb8980b8),
	.w3(32'h3bef6699),
	.w4(32'h3c008276),
	.w5(32'hbaf36958),
	.w6(32'h3a7cbcaf),
	.w7(32'h3a9727d1),
	.w8(32'hb9a5c270),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab069cb),
	.w1(32'h39bf000d),
	.w2(32'hbbf5ca6e),
	.w3(32'h3afc4e63),
	.w4(32'h3af25566),
	.w5(32'hbb9b148f),
	.w6(32'h3a8e1533),
	.w7(32'hb9be8f12),
	.w8(32'h3a184635),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eb329),
	.w1(32'h3c5d82b4),
	.w2(32'hb9f9c374),
	.w3(32'hbb7085fe),
	.w4(32'h3c071dbc),
	.w5(32'h3b825cbb),
	.w6(32'h3aae465f),
	.w7(32'hbb826fc8),
	.w8(32'h3a195d2d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdb61d),
	.w1(32'h3bf49e61),
	.w2(32'h3c0eb6ce),
	.w3(32'hbace1da3),
	.w4(32'h3a30d20d),
	.w5(32'h3ba1df45),
	.w6(32'hbae28d93),
	.w7(32'h3b10776c),
	.w8(32'h3bbb7f2e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b543874),
	.w1(32'h3b5a198d),
	.w2(32'h3b8e3837),
	.w3(32'hbb20595b),
	.w4(32'hba70a5ea),
	.w5(32'h3b131173),
	.w6(32'h3a1a092f),
	.w7(32'h38fadc9d),
	.w8(32'hbb5f6102),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba163628),
	.w1(32'h3b69e413),
	.w2(32'hbc21e02d),
	.w3(32'hbb311272),
	.w4(32'h3aa4978c),
	.w5(32'hbb90f36a),
	.w6(32'hb9539581),
	.w7(32'hbb9ae270),
	.w8(32'h3b244a0e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6020c),
	.w1(32'hb511738b),
	.w2(32'hba507e22),
	.w3(32'hb935aeb1),
	.w4(32'hbaeccd21),
	.w5(32'hbb119e49),
	.w6(32'h38f037a0),
	.w7(32'hbaa2b971),
	.w8(32'hbb358aea),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf04160),
	.w1(32'h3c0977ac),
	.w2(32'hbc2c8350),
	.w3(32'hbbc8fb19),
	.w4(32'h3a7faa8e),
	.w5(32'hbb7047ad),
	.w6(32'hbba1d962),
	.w7(32'hbbd144d5),
	.w8(32'hbb45f9a6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86bd4f),
	.w1(32'h39bb8b9d),
	.w2(32'hbb67f870),
	.w3(32'hbb2c34fb),
	.w4(32'h3afd905c),
	.w5(32'h3a5b2a57),
	.w6(32'hbabe25b6),
	.w7(32'hb9c03705),
	.w8(32'h3a93a968),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375efc58),
	.w1(32'hb98dee32),
	.w2(32'h39b7cfab),
	.w3(32'hb9a138e0),
	.w4(32'hb941a786),
	.w5(32'h3905085a),
	.w6(32'h37673392),
	.w7(32'hb95a43f4),
	.w8(32'h38078b0a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904a521),
	.w1(32'h38f05340),
	.w2(32'hba32f37f),
	.w3(32'h39c91b79),
	.w4(32'hbacc26a1),
	.w5(32'h3a070eb8),
	.w6(32'h3a227aa4),
	.w7(32'hba15ec5c),
	.w8(32'hbb0017bc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ada0a1),
	.w1(32'hba017421),
	.w2(32'hbb701968),
	.w3(32'h3a9d5339),
	.w4(32'h3ac445b2),
	.w5(32'hbb3c7908),
	.w6(32'hb9d07e9e),
	.w7(32'h3ac91f37),
	.w8(32'hbada2a48),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cdacdb),
	.w1(32'h3a9be9c8),
	.w2(32'h3b0b092c),
	.w3(32'hbb0fdc30),
	.w4(32'hbaa0ca79),
	.w5(32'h3ae779c0),
	.w6(32'hbac78037),
	.w7(32'hba1dbbbd),
	.w8(32'h39c834cb),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d4042),
	.w1(32'hba6fbc60),
	.w2(32'h3b050464),
	.w3(32'hbb1ef50b),
	.w4(32'hbb2cbed6),
	.w5(32'h3b497f92),
	.w6(32'hbb17fa48),
	.w7(32'hb9e937a3),
	.w8(32'h3b430234),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b584e6f),
	.w1(32'h3b18d1ce),
	.w2(32'h3b17f1d6),
	.w3(32'h3b3c8e22),
	.w4(32'h39cb3914),
	.w5(32'h39becf20),
	.w6(32'h3b6dffad),
	.w7(32'hb8f8c8e5),
	.w8(32'hbad5e3ff),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64c703),
	.w1(32'h3b528ff7),
	.w2(32'hbac964fb),
	.w3(32'h3bb98e9c),
	.w4(32'h3bad9f3e),
	.w5(32'h3b377d63),
	.w6(32'hb9e5c8cc),
	.w7(32'h391a928e),
	.w8(32'hbb8dcf62),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a236a67),
	.w1(32'hbb41a27b),
	.w2(32'hbb892dea),
	.w3(32'h3b64a00f),
	.w4(32'hbb3a3ccc),
	.w5(32'hbbaf2a66),
	.w6(32'h3b57ee56),
	.w7(32'h3a89c208),
	.w8(32'hbb88e7ca),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a315a),
	.w1(32'h3a8a517b),
	.w2(32'h396ca68b),
	.w3(32'h39905bd5),
	.w4(32'h39c0a132),
	.w5(32'h3a0cff10),
	.w6(32'h3a0c50c5),
	.w7(32'hb8e038bf),
	.w8(32'h3a7f440a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af34951),
	.w1(32'h3aeb0fd4),
	.w2(32'h3acaa0e0),
	.w3(32'h3b207947),
	.w4(32'h3ab0638a),
	.w5(32'hb93fc89b),
	.w6(32'h3b85062a),
	.w7(32'h3a9d1d65),
	.w8(32'hb93626b7),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1f334),
	.w1(32'hb8dbd792),
	.w2(32'hba2829de),
	.w3(32'h39e0874f),
	.w4(32'hb9904692),
	.w5(32'hbb10f408),
	.w6(32'h3983a1bf),
	.w7(32'hba202a70),
	.w8(32'hbaf1e966),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba678bdf),
	.w1(32'hbaaa57e5),
	.w2(32'hba89a12f),
	.w3(32'hba8697b5),
	.w4(32'hbaa84702),
	.w5(32'hb9f0b051),
	.w6(32'hba20009e),
	.w7(32'hba801100),
	.w8(32'hba06bd8d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba512783),
	.w1(32'hba9bb034),
	.w2(32'hbaa00d6f),
	.w3(32'hba6bb909),
	.w4(32'hba6a3e4d),
	.w5(32'hb9ed5490),
	.w6(32'hba916e99),
	.w7(32'hba6ca169),
	.w8(32'h38c53642),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a4a27),
	.w1(32'hba1e0181),
	.w2(32'h39b82b00),
	.w3(32'hbaa1d3a3),
	.w4(32'hba4b3115),
	.w5(32'hba2f3fe5),
	.w6(32'hbacd0b1d),
	.w7(32'hb93c8ab3),
	.w8(32'hbb04d788),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a704586),
	.w1(32'h3ab231e1),
	.w2(32'h39ad7d4a),
	.w3(32'h3a4fe7a4),
	.w4(32'h3a8ba219),
	.w5(32'hb9db6b0b),
	.w6(32'h3b04bcdf),
	.w7(32'h3a0a10c5),
	.w8(32'hb9b89e8c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00d4c5),
	.w1(32'h3a01ad13),
	.w2(32'hbb34fb3b),
	.w3(32'h3ae70c1d),
	.w4(32'h3b007b86),
	.w5(32'hbafcddd1),
	.w6(32'h3b04706d),
	.w7(32'h3acddfc7),
	.w8(32'h3a9d2a1d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985dacf),
	.w1(32'hbb0619f7),
	.w2(32'h3b093eab),
	.w3(32'hbadf6a27),
	.w4(32'hbba027f2),
	.w5(32'h3851032f),
	.w6(32'hb822a763),
	.w7(32'hbb4a3573),
	.w8(32'hbb154498),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba509c76),
	.w1(32'hba2fd5f0),
	.w2(32'hba5c302f),
	.w3(32'hba2422ec),
	.w4(32'hb936f169),
	.w5(32'hb97f0f60),
	.w6(32'hba63a056),
	.w7(32'hba056d2d),
	.w8(32'h39027d0b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b537f),
	.w1(32'hb99c7066),
	.w2(32'hba5a6efd),
	.w3(32'hba3150ee),
	.w4(32'hba3fc763),
	.w5(32'h38770575),
	.w6(32'hba037f4a),
	.w7(32'hba75d040),
	.w8(32'hba6e3de3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba278fd8),
	.w1(32'hba2afe91),
	.w2(32'hb9a86dab),
	.w3(32'hba49f1e1),
	.w4(32'hba79b448),
	.w5(32'h390299e9),
	.w6(32'hba9df292),
	.w7(32'hb9a357e6),
	.w8(32'h3901cdff),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dc2c2),
	.w1(32'hb9fb67a3),
	.w2(32'hba2bd6fd),
	.w3(32'hb990f13a),
	.w4(32'hba397217),
	.w5(32'h3a83d36f),
	.w6(32'h38859769),
	.w7(32'hb87347db),
	.w8(32'h3a445af6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4552cf),
	.w1(32'h3b7f29af),
	.w2(32'hbc14a149),
	.w3(32'h3baf5f4e),
	.w4(32'h3bb8d907),
	.w5(32'h3b866c96),
	.w6(32'h3a1bb8d9),
	.w7(32'hb9df9e23),
	.w8(32'hbad408b2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d657be),
	.w1(32'hbb7f0a1a),
	.w2(32'hbbb83301),
	.w3(32'h3b302025),
	.w4(32'h3a9ec5e5),
	.w5(32'hbbc8ab04),
	.w6(32'h3a2822a9),
	.w7(32'h3b067352),
	.w8(32'hbb065d95),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c14f7),
	.w1(32'hbaaaf667),
	.w2(32'hbb67833b),
	.w3(32'hb9ee7f50),
	.w4(32'hba2ee25b),
	.w5(32'hba94f45a),
	.w6(32'h3a198e77),
	.w7(32'hbaa864f8),
	.w8(32'h390624c7),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14106f),
	.w1(32'h3a83f7ee),
	.w2(32'hbac00722),
	.w3(32'h39b3651c),
	.w4(32'h3ae8f361),
	.w5(32'h39c43b71),
	.w6(32'h3ab75840),
	.w7(32'hbab7b221),
	.w8(32'hba4ad192),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03b1dc),
	.w1(32'h3a5f7d64),
	.w2(32'h3a30da15),
	.w3(32'hb943ccd4),
	.w4(32'h39b465dc),
	.w5(32'hb9e825de),
	.w6(32'hb929e563),
	.w7(32'h39615171),
	.w8(32'hb9c9c523),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b19b7),
	.w1(32'hba24bce2),
	.w2(32'hbaea9e27),
	.w3(32'hba51947d),
	.w4(32'hba06ce33),
	.w5(32'hbb0eb8b4),
	.w6(32'hb9f5e6aa),
	.w7(32'hba15c649),
	.w8(32'hbafbc171),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5443be),
	.w1(32'hbab4d720),
	.w2(32'hb627d862),
	.w3(32'hba1b4f08),
	.w4(32'hbaf67c26),
	.w5(32'hbb02d13d),
	.w6(32'h3a4de330),
	.w7(32'hb8e0f89f),
	.w8(32'hbb2388a0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba616785),
	.w1(32'hbb17da2d),
	.w2(32'hbc0841e3),
	.w3(32'h3b4e1bf0),
	.w4(32'h3b26f695),
	.w5(32'hbbc30d87),
	.w6(32'h3b30ac6e),
	.w7(32'h3b04ab5d),
	.w8(32'h39ca0dd3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a5a57),
	.w1(32'h3b062adf),
	.w2(32'h3b54c482),
	.w3(32'hb95b7317),
	.w4(32'hb988dad4),
	.w5(32'h3a77699b),
	.w6(32'h3999e852),
	.w7(32'h39560442),
	.w8(32'hb9d840bb),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabb98d),
	.w1(32'h39054ee0),
	.w2(32'hbb7d60e0),
	.w3(32'h3b18f54c),
	.w4(32'hba87a502),
	.w5(32'hbb40f00a),
	.w6(32'h3afd9734),
	.w7(32'hba25feee),
	.w8(32'hbb049db8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a509643),
	.w1(32'h3a6cc323),
	.w2(32'hbbd0fc49),
	.w3(32'h3b2fcd5f),
	.w4(32'h3b223dd6),
	.w5(32'hbb428325),
	.w6(32'h3ad99509),
	.w7(32'h3ae561b6),
	.w8(32'hba330283),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ff8e8),
	.w1(32'h3b2de04a),
	.w2(32'h3a38859d),
	.w3(32'hbad35e2b),
	.w4(32'h3a5d9557),
	.w5(32'h3b6920d3),
	.w6(32'hba42e3e3),
	.w7(32'hbac255a9),
	.w8(32'hbaf69949),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac77c09),
	.w1(32'hba498d6e),
	.w2(32'hbb67e95a),
	.w3(32'h3af20595),
	.w4(32'h39419679),
	.w5(32'hbb8db930),
	.w6(32'h3b0376f4),
	.w7(32'h39b42d94),
	.w8(32'hbb022e83),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b2fe96),
	.w1(32'h38ab3a18),
	.w2(32'hba9da05d),
	.w3(32'h38899a97),
	.w4(32'hb998e47e),
	.w5(32'h384f121a),
	.w6(32'hba185ae8),
	.w7(32'hba161c85),
	.w8(32'hb9143d04),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87a1050),
	.w1(32'h3af5fad0),
	.w2(32'h3b1c63e1),
	.w3(32'h3a8cc6b4),
	.w4(32'hb86f1548),
	.w5(32'h3b217465),
	.w6(32'hba43dbb4),
	.w7(32'hb9a56bec),
	.w8(32'h3af40862),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b062909),
	.w1(32'h3a479519),
	.w2(32'hb9e43ccd),
	.w3(32'h39dce44e),
	.w4(32'hb9b587e7),
	.w5(32'hba0b7281),
	.w6(32'hba57a101),
	.w7(32'hb9ef596b),
	.w8(32'hb96c7d44),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87b70ce),
	.w1(32'hba381d79),
	.w2(32'hba337537),
	.w3(32'hb9f2af62),
	.w4(32'hb8e562d1),
	.w5(32'hb847c248),
	.w6(32'h396c43b6),
	.w7(32'h397d90a9),
	.w8(32'hb967d9be),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb763a),
	.w1(32'hb91fe6bd),
	.w2(32'hb9b5918b),
	.w3(32'hb61407f6),
	.w4(32'hb952451e),
	.w5(32'hb8c18f4e),
	.w6(32'h3959d2ce),
	.w7(32'h389b3945),
	.w8(32'h38e37240),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a0ec4e),
	.w1(32'h3a8fddcb),
	.w2(32'hb9997977),
	.w3(32'hb9b164a6),
	.w4(32'h3a08435f),
	.w5(32'h3a8ed3be),
	.w6(32'hb95a10a4),
	.w7(32'hb9e8e970),
	.w8(32'h3b0cfea5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b081ff3),
	.w1(32'h3aea1667),
	.w2(32'h3b3c62ba),
	.w3(32'hba961729),
	.w4(32'hb9cf9703),
	.w5(32'h3b21cdad),
	.w6(32'h39cfc473),
	.w7(32'h39e9b428),
	.w8(32'hba6efbf3),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a49faf),
	.w1(32'hb9a33d00),
	.w2(32'hbb1c1afc),
	.w3(32'h3a167d5e),
	.w4(32'h3a191e77),
	.w5(32'hba93be6c),
	.w6(32'hb9d7e5ba),
	.w7(32'h3a5fe29b),
	.w8(32'hb8c27cfd),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394100d7),
	.w1(32'hb86ad74d),
	.w2(32'hb9193be0),
	.w3(32'hb9e9f7cc),
	.w4(32'h391994b7),
	.w5(32'h3a1b8487),
	.w6(32'h3a1a85ac),
	.w7(32'h3a1d0b75),
	.w8(32'h3a111179),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a904e92),
	.w1(32'hb9987e27),
	.w2(32'hbb420447),
	.w3(32'h3ab36285),
	.w4(32'h3b00571e),
	.w5(32'hbb589694),
	.w6(32'h3a5f0dc0),
	.w7(32'h3b281d4e),
	.w8(32'hbac17844),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97b359),
	.w1(32'hba877fa6),
	.w2(32'hb99fdfea),
	.w3(32'hba1086da),
	.w4(32'hb6ad061e),
	.w5(32'hb9e5deb0),
	.w6(32'h3a10b453),
	.w7(32'hb9993604),
	.w8(32'h3a54812a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b83495),
	.w1(32'h38cdddcc),
	.w2(32'hbbca943d),
	.w3(32'h3a9d9c5f),
	.w4(32'h3a26db6f),
	.w5(32'hbb9362d5),
	.w6(32'h3b011e83),
	.w7(32'h39c595ca),
	.w8(32'h3aa20d3d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39802d00),
	.w1(32'h39728f2e),
	.w2(32'h3ba8849a),
	.w3(32'hbb1a3c57),
	.w4(32'hba4632ac),
	.w5(32'h3b315770),
	.w6(32'hbb1c4c0e),
	.w7(32'h3b720e99),
	.w8(32'h3803dbcf),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd0431),
	.w1(32'h39fd8de3),
	.w2(32'h3964d5a0),
	.w3(32'hb6507c24),
	.w4(32'hba85f536),
	.w5(32'h39c0fc1e),
	.w6(32'h3aea9231),
	.w7(32'h3a13aa1b),
	.w8(32'hba441232),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b3bcf8),
	.w1(32'hb8fc64d6),
	.w2(32'hba5f5fe6),
	.w3(32'hba633772),
	.w4(32'hbac0ecf5),
	.w5(32'hbb3614ca),
	.w6(32'hba98f4c8),
	.w7(32'hbabc73f8),
	.w8(32'hbb220bba),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b9ab63),
	.w1(32'hba230637),
	.w2(32'h3924ffa8),
	.w3(32'hbace3c82),
	.w4(32'hba482850),
	.w5(32'h39f5baa6),
	.w6(32'hbb2042ec),
	.w7(32'hbaf78219),
	.w8(32'hbae05422),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd1797),
	.w1(32'h3a70f81e),
	.w2(32'h38938a54),
	.w3(32'hba7b798f),
	.w4(32'hba858aee),
	.w5(32'h3a4ad277),
	.w6(32'hbab7c625),
	.w7(32'h39a0eeec),
	.w8(32'h3a3f12eb),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955ce3b),
	.w1(32'h3a1f9103),
	.w2(32'h3b0717f6),
	.w3(32'hba38f860),
	.w4(32'hba25abf7),
	.w5(32'h390f1df6),
	.w6(32'h3a0a4a74),
	.w7(32'h39339daa),
	.w8(32'h3a7e7de1),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93afe00),
	.w1(32'hba002010),
	.w2(32'hbb1ac08a),
	.w3(32'h3a4e80ae),
	.w4(32'hb96e9a5b),
	.w5(32'hba57e735),
	.w6(32'h3ac5cb3d),
	.w7(32'hba88410a),
	.w8(32'h3a9f1fb4),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399be1bc),
	.w1(32'h3a20f527),
	.w2(32'h3a62abd9),
	.w3(32'h3a1fe3e5),
	.w4(32'h39ee82df),
	.w5(32'h3af6a3f6),
	.w6(32'h39de43d2),
	.w7(32'h3a2b6943),
	.w8(32'h3b244961),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fe341),
	.w1(32'h3b04509e),
	.w2(32'hbb175ca0),
	.w3(32'h3b93a333),
	.w4(32'h3b31103a),
	.w5(32'hbb45d89b),
	.w6(32'h3ba33b49),
	.w7(32'h3b451fd2),
	.w8(32'hba889ed4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3d151),
	.w1(32'h38bd0a3f),
	.w2(32'hbaf08096),
	.w3(32'hb937ee53),
	.w4(32'h3a3f8809),
	.w5(32'hbaecb02d),
	.w6(32'hb91444d1),
	.w7(32'h3a1e8a61),
	.w8(32'h39194f66),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89c219),
	.w1(32'hba4bea5d),
	.w2(32'h3ae8de47),
	.w3(32'hbb1584b7),
	.w4(32'hbacc0f11),
	.w5(32'h3ab3c4be),
	.w6(32'hbb51b4e8),
	.w7(32'hbae7c149),
	.w8(32'hba402aee),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d9fec),
	.w1(32'h39ef9f37),
	.w2(32'hb9a43e30),
	.w3(32'h39e7f76b),
	.w4(32'h397189b1),
	.w5(32'hb9e6eb73),
	.w6(32'h3a860e89),
	.w7(32'hb8de281c),
	.w8(32'h392b4969),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb357988),
	.w1(32'hbb8455f3),
	.w2(32'hbb6ce324),
	.w3(32'hba8e510e),
	.w4(32'hb8dface3),
	.w5(32'hba6df51b),
	.w6(32'hba8611c9),
	.w7(32'h3937e52e),
	.w8(32'h399e8452),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394bdb4c),
	.w1(32'h3a1cea86),
	.w2(32'hb7330f69),
	.w3(32'h395ff22f),
	.w4(32'hba2deacb),
	.w5(32'hb95885e5),
	.w6(32'h3a1516f3),
	.w7(32'hb9d5c079),
	.w8(32'hba96435d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e8fe6),
	.w1(32'hb9227536),
	.w2(32'hba1decb8),
	.w3(32'hb9919545),
	.w4(32'hb9854c03),
	.w5(32'h3b085353),
	.w6(32'hba7d2d9a),
	.w7(32'hb9e1bf0e),
	.w8(32'h3b5b470e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cebcd),
	.w1(32'h3b5a1e9b),
	.w2(32'h3b8ae6c1),
	.w3(32'h3b126886),
	.w4(32'h3a5e77cb),
	.w5(32'h3ab868ce),
	.w6(32'h3af946bd),
	.w7(32'h3acca851),
	.w8(32'hba050f0b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fbcc9),
	.w1(32'h3b20e9e8),
	.w2(32'hbb655dff),
	.w3(32'h3b3cbe21),
	.w4(32'h3bd3d853),
	.w5(32'h3b0bd568),
	.w6(32'h3ae88c85),
	.w7(32'h3b06d871),
	.w8(32'h3a3afa72),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0f934),
	.w1(32'hba600b12),
	.w2(32'hba561fba),
	.w3(32'hba65d32f),
	.w4(32'hba5141b1),
	.w5(32'hba479a87),
	.w6(32'hb9cc1023),
	.w7(32'hba0c626b),
	.w8(32'h39493ee8),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad39e8b),
	.w1(32'h3a351864),
	.w2(32'h3b0bd6b8),
	.w3(32'hbaa2b867),
	.w4(32'hbabe0d2c),
	.w5(32'h398754fb),
	.w6(32'hba1638ea),
	.w7(32'hb9b0c616),
	.w8(32'hbabf0fbc),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb086a04),
	.w1(32'hbb00b4d3),
	.w2(32'hbafb79aa),
	.w3(32'hbb3cbfeb),
	.w4(32'hbaa10a4b),
	.w5(32'h3a2b5729),
	.w6(32'hbb1b524c),
	.w7(32'hb8b98d98),
	.w8(32'h3ac9b0cd),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c272a4),
	.w1(32'hbb270e3f),
	.w2(32'hbb64f965),
	.w3(32'hbabd4dee),
	.w4(32'hba925647),
	.w5(32'hbb31fd86),
	.w6(32'hbaebdcfe),
	.w7(32'h3b03c186),
	.w8(32'h3a34b21a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b106dfc),
	.w1(32'h3a92967b),
	.w2(32'h38805301),
	.w3(32'h3b0b5a3a),
	.w4(32'h3a3bd22d),
	.w5(32'h39dc0401),
	.w6(32'h3b5e6a17),
	.w7(32'h3b1a2df1),
	.w8(32'h3a03ecbf),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b117fe9),
	.w1(32'hb8c5c144),
	.w2(32'hbb4bea43),
	.w3(32'h3b6f9b18),
	.w4(32'h3b1e81c5),
	.w5(32'hbb652898),
	.w6(32'h3ad44222),
	.w7(32'h3b36a590),
	.w8(32'hbaae45e9),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94c6c4f),
	.w1(32'h38c0ee08),
	.w2(32'h3991c7f8),
	.w3(32'h39305dc4),
	.w4(32'h39e701e2),
	.w5(32'hba641499),
	.w6(32'hb8e00122),
	.w7(32'hb91698c6),
	.w8(32'hba85bcdd),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f446a),
	.w1(32'hbac7ab8a),
	.w2(32'hbb10a361),
	.w3(32'h3b00ba73),
	.w4(32'hb9dc5441),
	.w5(32'hbb173282),
	.w6(32'h3ac96740),
	.w7(32'h3a9f3a6f),
	.w8(32'hba086256),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5eb067),
	.w1(32'h3a4c8911),
	.w2(32'h39d48a27),
	.w3(32'h3a320192),
	.w4(32'h3a42c4a0),
	.w5(32'hba5667fe),
	.w6(32'h39dc0c54),
	.w7(32'h3a12f785),
	.w8(32'hba1aaa5a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32be34),
	.w1(32'h3aa72314),
	.w2(32'h3ac7c329),
	.w3(32'h3a00df9f),
	.w4(32'h3a2fd66c),
	.w5(32'hb98b0abf),
	.w6(32'h3ac104b0),
	.w7(32'h3aeb8f66),
	.w8(32'hb8f014cd),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3812b636),
	.w1(32'hb911db97),
	.w2(32'hb98a35a1),
	.w3(32'hb9d7a6d2),
	.w4(32'hba612a66),
	.w5(32'h3a18b91b),
	.w6(32'hb95db6cb),
	.w7(32'hbacbd281),
	.w8(32'h3a132a9e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae652d7),
	.w1(32'hbb25a1b6),
	.w2(32'hbaf5bb53),
	.w3(32'h3aff4fd3),
	.w4(32'hbb26458c),
	.w5(32'hbb884958),
	.w6(32'h3ba8b74c),
	.w7(32'h3a9909d6),
	.w8(32'hbb2400d9),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad0cce),
	.w1(32'hba0fa9d1),
	.w2(32'hba0fd08e),
	.w3(32'hb98f84b1),
	.w4(32'hba0fe6f0),
	.w5(32'h3a272a50),
	.w6(32'hb9a5dbcf),
	.w7(32'hb98bbe15),
	.w8(32'h38cda2d7),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b0910e),
	.w1(32'h3921db12),
	.w2(32'h3789b1fa),
	.w3(32'h39ca2e1e),
	.w4(32'h3a1d8201),
	.w5(32'hba8afe67),
	.w6(32'hb9a23750),
	.w7(32'h3934f3d9),
	.w8(32'hba407752),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a372855),
	.w1(32'hb9ee7568),
	.w2(32'h39ad224c),
	.w3(32'hbb330739),
	.w4(32'hbb2c1e7f),
	.w5(32'hb99501af),
	.w6(32'hbad32559),
	.w7(32'hbb0211b2),
	.w8(32'hbb2a8fb7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb399c40),
	.w1(32'h3b041fb0),
	.w2(32'hbb0dad27),
	.w3(32'hbb72d744),
	.w4(32'hb85651c0),
	.w5(32'hbb84a74d),
	.w6(32'hbab253e2),
	.w7(32'hbbb32d1c),
	.w8(32'hbb85af83),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac5a4e),
	.w1(32'h3b263e99),
	.w2(32'hbb8f2354),
	.w3(32'hbb83d5df),
	.w4(32'h3aecb422),
	.w5(32'hba8b1118),
	.w6(32'hba23fb2d),
	.w7(32'hbb127675),
	.w8(32'h3a9afe97),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8756398),
	.w1(32'h39c300a4),
	.w2(32'h39b882be),
	.w3(32'h39036365),
	.w4(32'h398a3a5f),
	.w5(32'h3adbbed0),
	.w6(32'hb8ea812b),
	.w7(32'h38922b3d),
	.w8(32'h3aaae40a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b742c1c),
	.w1(32'h3a5dbc86),
	.w2(32'hbbab7ab2),
	.w3(32'h3b885b5a),
	.w4(32'h3b5169f9),
	.w5(32'hbb47aece),
	.w6(32'h3a2a893d),
	.w7(32'h3b5f7717),
	.w8(32'hbad6b2e2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a715006),
	.w1(32'hbb7262b9),
	.w2(32'h3aee0a87),
	.w3(32'hbb2e7853),
	.w4(32'hbb8044b2),
	.w5(32'hba68d86d),
	.w6(32'hbb70c2c6),
	.w7(32'h39a41f70),
	.w8(32'hbb32b390),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f627b5),
	.w1(32'h3918d2ef),
	.w2(32'hbb116a7b),
	.w3(32'h3a86a666),
	.w4(32'h3af92bec),
	.w5(32'hbb18e3d6),
	.w6(32'h3ac9f169),
	.w7(32'h3abc1610),
	.w8(32'h397368be),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927bd00),
	.w1(32'hb963e7aa),
	.w2(32'h3863a342),
	.w3(32'hba22924a),
	.w4(32'hb9b687a4),
	.w5(32'hba2f7eb5),
	.w6(32'h39590d35),
	.w7(32'h39c0bce3),
	.w8(32'hba92e33c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4c623),
	.w1(32'h3906521c),
	.w2(32'h3a1049ed),
	.w3(32'hba3255cd),
	.w4(32'h384d386d),
	.w5(32'hba24f8b4),
	.w6(32'hba3ea930),
	.w7(32'hb99fa3f5),
	.w8(32'hbaa23c5f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac041af),
	.w1(32'hba8b5098),
	.w2(32'hba2102b2),
	.w3(32'hba8a4ee4),
	.w4(32'h37fd805b),
	.w5(32'h39f5f046),
	.w6(32'hbacc717c),
	.w7(32'hba0db279),
	.w8(32'h3962a412),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b57a64),
	.w1(32'h3997cdbe),
	.w2(32'hbb73bebf),
	.w3(32'h3a1ef93f),
	.w4(32'h3b4672c4),
	.w5(32'hba380fbc),
	.w6(32'h3a6f148d),
	.w7(32'h3a6e8d3d),
	.w8(32'h3b023e93),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aded057),
	.w1(32'h3aa60c60),
	.w2(32'hba492e32),
	.w3(32'h3a79cfcc),
	.w4(32'h3a855f26),
	.w5(32'h3948b8a0),
	.w6(32'h39e43c96),
	.w7(32'h3a46476c),
	.w8(32'hba3bb291),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36f84b),
	.w1(32'h3b266a3e),
	.w2(32'h3ae234c5),
	.w3(32'hbae87c65),
	.w4(32'hba7f344e),
	.w5(32'h39bcb959),
	.w6(32'hba8a34bc),
	.w7(32'hbb2e3b8f),
	.w8(32'hbb1a8aea),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96441fe),
	.w1(32'h39d98735),
	.w2(32'h39c56a26),
	.w3(32'h393548c4),
	.w4(32'h39e13c03),
	.w5(32'h39aadb04),
	.w6(32'hb89358a0),
	.w7(32'hba443a98),
	.w8(32'hba20b6f3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9ef09),
	.w1(32'hb9ef867d),
	.w2(32'hbb7d3ea9),
	.w3(32'h3aec60c9),
	.w4(32'h3abef096),
	.w5(32'hba35e78b),
	.w6(32'hbab7582e),
	.w7(32'h3a32cd6e),
	.w8(32'h39d65030),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc6bd6),
	.w1(32'h3a8bd6bb),
	.w2(32'hba107860),
	.w3(32'hbaf190f2),
	.w4(32'h3a447b08),
	.w5(32'h3b131715),
	.w6(32'hba7eacf7),
	.w7(32'hbae6d992),
	.w8(32'hba3fc5bd),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f35799),
	.w1(32'hba37b1ba),
	.w2(32'h39ed2b8f),
	.w3(32'h39a8e72c),
	.w4(32'hb9549ec3),
	.w5(32'h39acd607),
	.w6(32'h38eedc12),
	.w7(32'hb9486580),
	.w8(32'h38814000),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3bda0),
	.w1(32'hb9811880),
	.w2(32'hbb42d2c6),
	.w3(32'h3a58bf61),
	.w4(32'h3a118505),
	.w5(32'hbb31d701),
	.w6(32'hba4473e5),
	.w7(32'hbb795189),
	.w8(32'hbb522dad),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83ab25),
	.w1(32'hba5dd2f7),
	.w2(32'hbaaf0800),
	.w3(32'hba0503bb),
	.w4(32'h38223edb),
	.w5(32'h39e091d2),
	.w6(32'hb9f1b900),
	.w7(32'hb9b24ccc),
	.w8(32'h3928c195),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f7135),
	.w1(32'hb9b16a6a),
	.w2(32'hbb2ab471),
	.w3(32'hba09a5ce),
	.w4(32'h3784dcf8),
	.w5(32'hbaec2b5e),
	.w6(32'h36a6a364),
	.w7(32'h3948e63f),
	.w8(32'hbad4261a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a2b930),
	.w1(32'h39baa190),
	.w2(32'h3a79d8c4),
	.w3(32'hbb1e5c48),
	.w4(32'hbb6b608d),
	.w5(32'hb957a73c),
	.w6(32'hbb211e16),
	.w7(32'hbb0f5971),
	.w8(32'hbb8dc2b5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33b0d7),
	.w1(32'hb9370031),
	.w2(32'h3a14c4dd),
	.w3(32'hbb12c098),
	.w4(32'hba54881f),
	.w5(32'h3a8caf98),
	.w6(32'hba331854),
	.w7(32'hba58ad85),
	.w8(32'hb9ab3abd),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92910be),
	.w1(32'hb7a0ee8b),
	.w2(32'hb869c64a),
	.w3(32'hb964081f),
	.w4(32'hb98e6e8c),
	.w5(32'h39020ee0),
	.w6(32'hb8f67d40),
	.w7(32'hb5689431),
	.w8(32'h39bae23c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa039f4),
	.w1(32'hba1ab0ef),
	.w2(32'h3afdc83c),
	.w3(32'hbb163aba),
	.w4(32'hbace5dbe),
	.w5(32'h3a0cc28b),
	.w6(32'hbab4d1fa),
	.w7(32'hbaab3c0c),
	.w8(32'hbb2c6ced),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4725d8),
	.w1(32'hba51c3d9),
	.w2(32'hbb02a99a),
	.w3(32'h3a951ca7),
	.w4(32'h3a60dcfa),
	.w5(32'hb9f00c4b),
	.w6(32'h3a3b9e48),
	.w7(32'h388a363c),
	.w8(32'h389893b4),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6aaebd),
	.w1(32'h3a062a25),
	.w2(32'hba900523),
	.w3(32'h3ac81f46),
	.w4(32'h3a8ac75b),
	.w5(32'hbacbf88b),
	.w6(32'h3a3f971c),
	.w7(32'h3ace276a),
	.w8(32'hba28b90d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a8f7ad),
	.w1(32'hb994c529),
	.w2(32'hba55c3b6),
	.w3(32'hb9a7e645),
	.w4(32'hba30feb1),
	.w5(32'hb8d7af69),
	.w6(32'hb923bbd6),
	.w7(32'hba227bc8),
	.w8(32'hba45a4e1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dde2dd),
	.w1(32'hba3bdbb9),
	.w2(32'hba55768b),
	.w3(32'hb9e6e221),
	.w4(32'hb9832ff8),
	.w5(32'h38d1ab61),
	.w6(32'h3a89dec8),
	.w7(32'hb999c8db),
	.w8(32'h3909ba11),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba8bc1),
	.w1(32'h3b48333c),
	.w2(32'hbb39ddcf),
	.w3(32'hb99fb670),
	.w4(32'h3b8e4917),
	.w5(32'h3b607d7b),
	.w6(32'h3aa9784a),
	.w7(32'hbb09b471),
	.w8(32'hbb91865d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82cd6a),
	.w1(32'h3ac68384),
	.w2(32'hbb506894),
	.w3(32'h3ae05f63),
	.w4(32'h3a66b97f),
	.w5(32'h3a86cda8),
	.w6(32'h3af89dd0),
	.w7(32'hba341cf1),
	.w8(32'hbb146d54),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7edd59),
	.w1(32'h3a881752),
	.w2(32'h3aad48a7),
	.w3(32'hba52a483),
	.w4(32'h3a0af1d7),
	.w5(32'h38bb8c02),
	.w6(32'h398bd5aa),
	.w7(32'hb84dd7ff),
	.w8(32'hbb3db665),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390588c9),
	.w1(32'hba9b2b4e),
	.w2(32'hbc1e3ae2),
	.w3(32'h3a0bdbff),
	.w4(32'h3a6f2415),
	.w5(32'hbc2a13f7),
	.w6(32'h3b5ec175),
	.w7(32'hbb31c3f6),
	.w8(32'hbba16146),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba876db5),
	.w1(32'hbaecac2c),
	.w2(32'hbadb9b2f),
	.w3(32'hb9c32f06),
	.w4(32'hbaab68cc),
	.w5(32'hba04851b),
	.w6(32'hbacd2a28),
	.w7(32'hba68c962),
	.w8(32'hb9c80d66),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace29fd),
	.w1(32'h39d00920),
	.w2(32'hbacbd8f6),
	.w3(32'h3ac0f92c),
	.w4(32'h39a3bc1a),
	.w5(32'h3a194857),
	.w6(32'h3a970962),
	.w7(32'hba317ba3),
	.w8(32'h39efd2a7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d9bc2),
	.w1(32'h3be2d1a7),
	.w2(32'hbb8f6773),
	.w3(32'hbb602ac8),
	.w4(32'h3c58562e),
	.w5(32'h3afe8ec4),
	.w6(32'h393d1d85),
	.w7(32'h3baca719),
	.w8(32'h3b03585f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93244c),
	.w1(32'h3afcc3b6),
	.w2(32'hbbe1c50c),
	.w3(32'h3b8eb5ac),
	.w4(32'h3b9532b9),
	.w5(32'hbad40c92),
	.w6(32'h3a066ae7),
	.w7(32'h3b6c88c3),
	.w8(32'h39f5384d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb150d08),
	.w1(32'h3add8193),
	.w2(32'hbb60b867),
	.w3(32'h3a9847ac),
	.w4(32'h3b2a9811),
	.w5(32'hba19d95f),
	.w6(32'h3aceb1eb),
	.w7(32'hba513d98),
	.w8(32'h3a556c33),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58b1b7),
	.w1(32'h3a30306c),
	.w2(32'h3b0afcba),
	.w3(32'hbb140bd6),
	.w4(32'hbb293703),
	.w5(32'h3a8f4e03),
	.w6(32'hbaf53cf5),
	.w7(32'hba80f493),
	.w8(32'h394bad77),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64e5a8),
	.w1(32'h390729b0),
	.w2(32'h3b5b96b7),
	.w3(32'hba54fdba),
	.w4(32'hbb2fcaa8),
	.w5(32'h39fe90e0),
	.w6(32'hb964eb2d),
	.w7(32'hba5ebbbc),
	.w8(32'hbaaf9bb2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394667bd),
	.w1(32'h380ef74e),
	.w2(32'hb91af5f6),
	.w3(32'h37f444f6),
	.w4(32'hb9c588d3),
	.w5(32'h3a6abfe6),
	.w6(32'h3a26ad4d),
	.w7(32'hb8563596),
	.w8(32'h3a866682),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff9962),
	.w1(32'h39ae09e2),
	.w2(32'h3989f676),
	.w3(32'h38595c6e),
	.w4(32'hba03512c),
	.w5(32'hba3da17c),
	.w6(32'h3a175ba4),
	.w7(32'h394c4d53),
	.w8(32'hb8b4ff68),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e430c2),
	.w1(32'hba5e525f),
	.w2(32'hbab6abdf),
	.w3(32'h3ab07e13),
	.w4(32'h3a085c30),
	.w5(32'h3985a93c),
	.w6(32'h3862ce2e),
	.w7(32'h399c3038),
	.w8(32'hb87b89f7),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99979ff),
	.w1(32'h39c4ef66),
	.w2(32'hb92038b6),
	.w3(32'h38b49801),
	.w4(32'h3987f9a7),
	.w5(32'h3b16e3b9),
	.w6(32'h3b109fbe),
	.w7(32'h399ef9fe),
	.w8(32'h3a4fbc6b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab30efb),
	.w1(32'h3aaf8644),
	.w2(32'hbb9def69),
	.w3(32'hba1144d8),
	.w4(32'hbb2e1227),
	.w5(32'hbbac08ae),
	.w6(32'hba26ebe7),
	.w7(32'hbb933956),
	.w8(32'h3c1ef102),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badb6c5),
	.w1(32'h3c340bf6),
	.w2(32'hbb973c21),
	.w3(32'hba8913b2),
	.w4(32'h3b384451),
	.w5(32'h3a820406),
	.w6(32'h3c0e630b),
	.w7(32'hbc00be1c),
	.w8(32'h3bc4cdd0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aead600),
	.w1(32'h3c7ab60a),
	.w2(32'h3c48d801),
	.w3(32'h3c213ec6),
	.w4(32'h3c01dcfd),
	.w5(32'hbb02d819),
	.w6(32'hbc190008),
	.w7(32'h3c1d905a),
	.w8(32'hbbb7df64),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3715ac8d),
	.w1(32'h3bc02bfb),
	.w2(32'h3aaa6d0f),
	.w3(32'h3b85f0cb),
	.w4(32'hbb367c3e),
	.w5(32'hb9a6a3ef),
	.w6(32'hbbabab45),
	.w7(32'hbb320206),
	.w8(32'hba33b18e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab168c),
	.w1(32'hb9bf3a93),
	.w2(32'hbbfa9c98),
	.w3(32'h3b27871f),
	.w4(32'h3ba82bee),
	.w5(32'hbbc2e442),
	.w6(32'h3aa70040),
	.w7(32'hbb8dd0b2),
	.w8(32'h3c194840),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba875e69),
	.w1(32'h3b382afd),
	.w2(32'hbae7d1b5),
	.w3(32'hbaf15c22),
	.w4(32'h3a203799),
	.w5(32'h3b573de8),
	.w6(32'hbbefedd6),
	.w7(32'h3b613760),
	.w8(32'hbc0765aa),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5489f),
	.w1(32'h3b8e0a71),
	.w2(32'h3b831de9),
	.w3(32'h3bdef679),
	.w4(32'h3c7cdb6e),
	.w5(32'h3c070546),
	.w6(32'hbb586b4f),
	.w7(32'hbb134b5e),
	.w8(32'hbb71db82),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0b587),
	.w1(32'h3bdff806),
	.w2(32'hb9422a42),
	.w3(32'h3b68b386),
	.w4(32'h3bf33b61),
	.w5(32'h3bb33c50),
	.w6(32'h3b025243),
	.w7(32'hb901f08e),
	.w8(32'hbbf8fc93),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ccadc),
	.w1(32'hbb889993),
	.w2(32'h3aa94d03),
	.w3(32'h3b30c28e),
	.w4(32'h3b80c650),
	.w5(32'h3b864d8b),
	.w6(32'h3c57b0ef),
	.w7(32'hbb1f5b7f),
	.w8(32'hb8e0a648),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf06b62),
	.w1(32'h3b8b4b52),
	.w2(32'h3b6807fb),
	.w3(32'h3bb6c3b0),
	.w4(32'h3b2c5a95),
	.w5(32'hba69ad57),
	.w6(32'h3ac79eb3),
	.w7(32'h3b0f4e75),
	.w8(32'h3b04b3b3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b37b0),
	.w1(32'h3b161d8e),
	.w2(32'hbb6aa7c0),
	.w3(32'hbae578fb),
	.w4(32'hbb6620ee),
	.w5(32'h3bf2b0ff),
	.w6(32'hbbcbe186),
	.w7(32'hbb9dcee1),
	.w8(32'h3a1212c5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98c359),
	.w1(32'hbac6abf8),
	.w2(32'hbac7e802),
	.w3(32'h3b007c21),
	.w4(32'h3b6a6102),
	.w5(32'hbc1118f9),
	.w6(32'hbb934fed),
	.w7(32'hbb0902b4),
	.w8(32'hbbbcea72),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fd662),
	.w1(32'hbb86f490),
	.w2(32'hbb2f934f),
	.w3(32'hbc288c23),
	.w4(32'hbc403dae),
	.w5(32'hbb629030),
	.w6(32'h3a320f6c),
	.w7(32'hbb598849),
	.w8(32'hbb1102c9),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f4a52),
	.w1(32'hbbb0539e),
	.w2(32'hbc163a90),
	.w3(32'hbb940f0d),
	.w4(32'hbbb66ad7),
	.w5(32'hbc314516),
	.w6(32'hbb4da33a),
	.w7(32'h3a11e78e),
	.w8(32'hbc13cc1a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5803d),
	.w1(32'hbb8e84d5),
	.w2(32'hbbd6ba57),
	.w3(32'hbade1c5f),
	.w4(32'hb93b9d4d),
	.w5(32'hba6a6919),
	.w6(32'hbbd3eaa1),
	.w7(32'hbb223cb0),
	.w8(32'h3a1fb50f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37cb2c),
	.w1(32'h3b1f59ab),
	.w2(32'h39bfe3da),
	.w3(32'h3a9f24ec),
	.w4(32'hbae585a9),
	.w5(32'h39b31eb2),
	.w6(32'hbab5cdd0),
	.w7(32'h3b86ab23),
	.w8(32'hbc2457af),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a335e),
	.w1(32'hbc3e79bb),
	.w2(32'hbb3b9af4),
	.w3(32'hbbc56a55),
	.w4(32'h3b0f9e90),
	.w5(32'hbbaf16f1),
	.w6(32'h3c33834f),
	.w7(32'hbc46f84f),
	.w8(32'hba6caa25),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a43dd),
	.w1(32'h3a450de6),
	.w2(32'hbb7f9159),
	.w3(32'hbb20e183),
	.w4(32'hbc00d34f),
	.w5(32'hbb764f35),
	.w6(32'hbbb4b099),
	.w7(32'hbc038174),
	.w8(32'hbba85198),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d0bca),
	.w1(32'hbb3503aa),
	.w2(32'hba6c0a6c),
	.w3(32'hbaa83d7f),
	.w4(32'hbab72603),
	.w5(32'h3c208b3a),
	.w6(32'hbb9745b4),
	.w7(32'hbb89cfce),
	.w8(32'h3aa7629e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b355bc2),
	.w1(32'h3bbbc100),
	.w2(32'h3821ffeb),
	.w3(32'h3c07d699),
	.w4(32'h3bacbd9a),
	.w5(32'h3c6eb1e3),
	.w6(32'h3bf8b68a),
	.w7(32'h3ca2cc2b),
	.w8(32'h3be94f4b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abec5c4),
	.w1(32'hb961fe33),
	.w2(32'hbc004c83),
	.w3(32'h3c2c6950),
	.w4(32'h3b8a032a),
	.w5(32'hbb2c74d3),
	.w6(32'h3b8f7361),
	.w7(32'h3a838c2e),
	.w8(32'hbb81a1bc),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8309ae),
	.w1(32'h3b9695cd),
	.w2(32'hbae4353a),
	.w3(32'h3bd86408),
	.w4(32'hba2641a5),
	.w5(32'h3a90c0ac),
	.w6(32'h3ad89cad),
	.w7(32'hbc7d48f8),
	.w8(32'hbb6fff5b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a843fc),
	.w1(32'h3bf31734),
	.w2(32'h3af3f71e),
	.w3(32'hba80bb1e),
	.w4(32'h376bc952),
	.w5(32'hbb37bbb8),
	.w6(32'hba85996b),
	.w7(32'h3bb25dcc),
	.w8(32'hbb9cbf37),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e251a),
	.w1(32'hbad29664),
	.w2(32'hbbcd7c3e),
	.w3(32'hbb660cd9),
	.w4(32'hbbd144ae),
	.w5(32'hbb5c05e4),
	.w6(32'hbb6351d9),
	.w7(32'hbb9bc3d3),
	.w8(32'hbb722c72),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f5109),
	.w1(32'h3b4d0381),
	.w2(32'h3a1df4b8),
	.w3(32'hbba92a50),
	.w4(32'hbac026c3),
	.w5(32'hb97586f9),
	.w6(32'h3b5a082a),
	.w7(32'hbb9e0c8b),
	.w8(32'h3accd5eb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2d390),
	.w1(32'h3999b6f9),
	.w2(32'hbb3a6a55),
	.w3(32'hbbb74ae3),
	.w4(32'hbbde1bfd),
	.w5(32'hbbd7ec4e),
	.w6(32'h3c107e00),
	.w7(32'hbb54e17b),
	.w8(32'h3bdd5f63),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93d1d1),
	.w1(32'hbb72d6fd),
	.w2(32'hbb599df6),
	.w3(32'h3a79ec01),
	.w4(32'hbbcbb893),
	.w5(32'h3ba36cb1),
	.w6(32'h3c32a2ce),
	.w7(32'h3b497e2c),
	.w8(32'hbb04c693),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab983a2),
	.w1(32'hbba9ea3e),
	.w2(32'hbb904c3a),
	.w3(32'h3bcaafb5),
	.w4(32'hbb5c3c0f),
	.w5(32'hbb9c1a28),
	.w6(32'h3b7a875a),
	.w7(32'h3c30fdd0),
	.w8(32'hbb8d1711),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba409205),
	.w1(32'hba2c6bc9),
	.w2(32'hbb5da40b),
	.w3(32'h3b147f74),
	.w4(32'hb9639cc9),
	.w5(32'hbba17996),
	.w6(32'h3b7ce1b3),
	.w7(32'h39ff17c2),
	.w8(32'h3955ba51),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc84776),
	.w1(32'h3c511e31),
	.w2(32'h3c5b8b09),
	.w3(32'hba3f4349),
	.w4(32'h3ba0fcdc),
	.w5(32'h3b49e40c),
	.w6(32'hbc2db96d),
	.w7(32'hbb1ab026),
	.w8(32'hbc3e80df),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule