module layer_10_featuremap_473(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ffbef),
	.w1(32'hbc450ab1),
	.w2(32'h3bebeb2a),
	.w3(32'hbc0ef159),
	.w4(32'hbd10a8dd),
	.w5(32'hbc93b632),
	.w6(32'h39d75f3c),
	.w7(32'hbc2ca58b),
	.w8(32'hbbb0ab98),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce29e81),
	.w1(32'hbc33aa8f),
	.w2(32'hbc1c7f26),
	.w3(32'h3d2983cb),
	.w4(32'hbc45db41),
	.w5(32'h3a49dc02),
	.w6(32'h3c9dd231),
	.w7(32'hbc3f0f98),
	.w8(32'hbc339945),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b359b),
	.w1(32'hbc124043),
	.w2(32'hbc0beb52),
	.w3(32'hbc1ba954),
	.w4(32'hbbe9eae1),
	.w5(32'h3ac321ef),
	.w6(32'hbb3fff5e),
	.w7(32'hbc17fb11),
	.w8(32'hbc3682b1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13e487),
	.w1(32'h3a8db84d),
	.w2(32'h3ac0e76e),
	.w3(32'h3bb61289),
	.w4(32'h3c025d6f),
	.w5(32'hbc1e28b7),
	.w6(32'hbb8281ab),
	.w7(32'hbb646912),
	.w8(32'h3b83d0ed),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc211dce),
	.w1(32'h39805702),
	.w2(32'hbbcbe742),
	.w3(32'hbbf89a6f),
	.w4(32'h3bc83e8b),
	.w5(32'hbb9b904f),
	.w6(32'hbc315220),
	.w7(32'hbba5af17),
	.w8(32'hbb888d05),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934b0a6),
	.w1(32'hba24aac0),
	.w2(32'hbb18c955),
	.w3(32'hb8f047ec),
	.w4(32'hb74d0fcf),
	.w5(32'h3b7201cb),
	.w6(32'hbb222c80),
	.w7(32'h3c47b059),
	.w8(32'hb9fa7f5f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb017b9c),
	.w1(32'h3bf9f720),
	.w2(32'h3adab707),
	.w3(32'hbc5c4fae),
	.w4(32'h3a0a23c7),
	.w5(32'hbc6f4ce2),
	.w6(32'h3c02e9db),
	.w7(32'h3bc9b6b1),
	.w8(32'h3b45cbab),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3e9a9),
	.w1(32'hbb86e0cd),
	.w2(32'hba6e921f),
	.w3(32'hbb5208ed),
	.w4(32'hbb40ac6e),
	.w5(32'hbba238d9),
	.w6(32'hbb40369c),
	.w7(32'hbba69149),
	.w8(32'hbbbf02f0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eec683),
	.w1(32'hbbe4e206),
	.w2(32'hbc8f41fa),
	.w3(32'h3b0faef7),
	.w4(32'hbc0d9250),
	.w5(32'hbc480db4),
	.w6(32'hbb6aab3a),
	.w7(32'hbbd35a66),
	.w8(32'hbc1bfa5f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32050a),
	.w1(32'h3ba008e8),
	.w2(32'h3abaec1f),
	.w3(32'hbc2d7eb7),
	.w4(32'h3b89f11b),
	.w5(32'hbb42214c),
	.w6(32'hbb740c18),
	.w7(32'hbb584715),
	.w8(32'hbbd1e761),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a675aeb),
	.w1(32'h3af29e85),
	.w2(32'h3b31fb04),
	.w3(32'h3c11317c),
	.w4(32'hbbc720c9),
	.w5(32'hbba6cd02),
	.w6(32'hbac615d2),
	.w7(32'hbad5bc94),
	.w8(32'hbb6cabc0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd7943),
	.w1(32'h3b9b6ab3),
	.w2(32'h39169246),
	.w3(32'hbc12a81c),
	.w4(32'h3c533c55),
	.w5(32'h3c6d4d86),
	.w6(32'hbb94f2fb),
	.w7(32'h3ba31b37),
	.w8(32'hbb5ded5d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38de6a),
	.w1(32'hbc245e1c),
	.w2(32'hbc85dd63),
	.w3(32'hbcbe4998),
	.w4(32'h3c341242),
	.w5(32'h3c2144dc),
	.w6(32'hbc68e32e),
	.w7(32'h3b7549d4),
	.w8(32'hbbcd88ef),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65d5e1),
	.w1(32'hbc344b5d),
	.w2(32'hbc14b42c),
	.w3(32'hbca7a790),
	.w4(32'hbc02c0cc),
	.w5(32'hbaa73ae1),
	.w6(32'hbb4e74c1),
	.w7(32'hbc336470),
	.w8(32'hbba13daf),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81934c),
	.w1(32'hbbe66321),
	.w2(32'hbc5040a5),
	.w3(32'hbbb9a947),
	.w4(32'hbbd78812),
	.w5(32'h39e1b04a),
	.w6(32'hbbfb8829),
	.w7(32'hbbcd372b),
	.w8(32'hbc13c217),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11317d),
	.w1(32'hbc652243),
	.w2(32'hbb7be2c4),
	.w3(32'hbc86a357),
	.w4(32'hbb9238a9),
	.w5(32'hb9387346),
	.w6(32'hbc689776),
	.w7(32'hbbacd6d3),
	.w8(32'h3a24eefc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf4bc2),
	.w1(32'h3a10f66f),
	.w2(32'h3c1606c8),
	.w3(32'hbbb8f53e),
	.w4(32'h3b2f9888),
	.w5(32'h3c1c2566),
	.w6(32'hbbfa6325),
	.w7(32'h39f4702d),
	.w8(32'h3c672a98),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71b5dd),
	.w1(32'hbc76c4b7),
	.w2(32'hba940c40),
	.w3(32'h3bac2be7),
	.w4(32'hbd1e82a1),
	.w5(32'hbb490bed),
	.w6(32'hbb3f26ee),
	.w7(32'hbcc1bec2),
	.w8(32'hbc5c4e33),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47b73c),
	.w1(32'hbbe904d8),
	.w2(32'hbc01e2ca),
	.w3(32'h3cfd60d1),
	.w4(32'h3ba72014),
	.w5(32'h3c1a4dd0),
	.w6(32'h3c9be3fc),
	.w7(32'hba7d313d),
	.w8(32'hbb311bf8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1602d6),
	.w1(32'hbc7469bb),
	.w2(32'hbc0dc3c0),
	.w3(32'hbc92d1d8),
	.w4(32'hbc887ba3),
	.w5(32'hbbae13f5),
	.w6(32'hbc291c55),
	.w7(32'hbc10d5f3),
	.w8(32'hbc69ee33),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18d9e6),
	.w1(32'h3c550eb7),
	.w2(32'h3bc435c2),
	.w3(32'hbb8e52e7),
	.w4(32'h3c9ad81a),
	.w5(32'h3ca8757d),
	.w6(32'hbb644ae1),
	.w7(32'h3c802bbd),
	.w8(32'h3c06e6d9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fee51),
	.w1(32'hbc0adf5f),
	.w2(32'hbca07954),
	.w3(32'hbc8bcfca),
	.w4(32'hbbba2e4a),
	.w5(32'hbbc3e411),
	.w6(32'hbc0bf7cc),
	.w7(32'hbbccab14),
	.w8(32'hbc687285),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c66d1),
	.w1(32'hba85f296),
	.w2(32'hbc1f3ea2),
	.w3(32'hbc1b0da1),
	.w4(32'h3bba1ea3),
	.w5(32'hba648a62),
	.w6(32'hbbd97d71),
	.w7(32'h3afeb9e7),
	.w8(32'hbc16fda3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c947e),
	.w1(32'hbb38aed4),
	.w2(32'hbc526504),
	.w3(32'h3ad853e1),
	.w4(32'h3c372919),
	.w5(32'h39f2c5ca),
	.w6(32'hba480157),
	.w7(32'hba2467f3),
	.w8(32'hbbb4b2a6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c045a),
	.w1(32'hbc705f8c),
	.w2(32'hbcccb020),
	.w3(32'h3c2d77a3),
	.w4(32'hbbf3c4bf),
	.w5(32'hbbd89a31),
	.w6(32'hbb308794),
	.w7(32'hbc02ec15),
	.w8(32'hbcb06480),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca32bc8),
	.w1(32'h3c90577b),
	.w2(32'h3a300b9a),
	.w3(32'hbc3536cf),
	.w4(32'h3c9ef5d5),
	.w5(32'hbbf97387),
	.w6(32'hbcadec7b),
	.w7(32'h3c26870a),
	.w8(32'h3c244390),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87f74d),
	.w1(32'h3be2d263),
	.w2(32'hbafedaf5),
	.w3(32'h3c90d833),
	.w4(32'hb8c0fdc6),
	.w5(32'hbbba250b),
	.w6(32'h3c9a5c4c),
	.w7(32'h3b9ed083),
	.w8(32'h3bd4454b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf320b),
	.w1(32'h3b70d735),
	.w2(32'hbb279ea0),
	.w3(32'h3c1c429d),
	.w4(32'hb891b18f),
	.w5(32'hbb978f43),
	.w6(32'h3b1b2291),
	.w7(32'hbad4c971),
	.w8(32'hbb11267d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa1d02),
	.w1(32'h3ba87d70),
	.w2(32'hbb900f61),
	.w3(32'hb9d78dfb),
	.w4(32'hba8b4453),
	.w5(32'h3b664a03),
	.w6(32'hbc1ea767),
	.w7(32'h3bb29061),
	.w8(32'hba60c7cb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d10f1),
	.w1(32'h3c5f082d),
	.w2(32'hbb9b360c),
	.w3(32'hbc12c8b3),
	.w4(32'h3ce3158e),
	.w5(32'hbb6cec06),
	.w6(32'h3af36c98),
	.w7(32'h3ca1a546),
	.w8(32'h3abd9af1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc45c3d),
	.w1(32'h3b0b773a),
	.w2(32'h3c48bc23),
	.w3(32'hbd1e7d86),
	.w4(32'h3be14bed),
	.w5(32'h3b80b853),
	.w6(32'hbc525c23),
	.w7(32'hbad9ab63),
	.w8(32'h3b454a52),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcca0f3),
	.w1(32'h3a65a868),
	.w2(32'hbb761f80),
	.w3(32'h3c626e37),
	.w4(32'hbb43a026),
	.w5(32'hbc18118a),
	.w6(32'h3c03816c),
	.w7(32'hb9091c5a),
	.w8(32'hbbfd3697),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb256e1c),
	.w1(32'hbb2f056b),
	.w2(32'hba9e0bb4),
	.w3(32'hbbbc2ef6),
	.w4(32'h3b65ab56),
	.w5(32'hbb22f8b0),
	.w6(32'hbb0d449b),
	.w7(32'hb92521eb),
	.w8(32'hbab721d4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde5894),
	.w1(32'h3bce8a91),
	.w2(32'h3b094e80),
	.w3(32'hbb8bca12),
	.w4(32'h3b0749ac),
	.w5(32'hbbb92525),
	.w6(32'hbc1f27e8),
	.w7(32'h3bc37690),
	.w8(32'h3b911489),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf834f5),
	.w1(32'h39088b94),
	.w2(32'h3b647ee2),
	.w3(32'h3c04aa3d),
	.w4(32'h3b54e2e6),
	.w5(32'h3acd0421),
	.w6(32'hba16b309),
	.w7(32'hbbb4f07f),
	.w8(32'h39bce5c4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f0390),
	.w1(32'hbb380c79),
	.w2(32'hbaf5ebc1),
	.w3(32'h3b4dd413),
	.w4(32'hbc4f20ee),
	.w5(32'h39ddad94),
	.w6(32'hbc228b1e),
	.w7(32'hbb70109b),
	.w8(32'h3ab3519f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a047c),
	.w1(32'hbc2f12cf),
	.w2(32'hbc3938c5),
	.w3(32'h3b877922),
	.w4(32'hbc6eed32),
	.w5(32'hbc23cae5),
	.w6(32'hba5a196c),
	.w7(32'hbc23b331),
	.w8(32'hbc5101ac),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86edeb),
	.w1(32'hbbb646a2),
	.w2(32'hbb095a2a),
	.w3(32'hbbcdf886),
	.w4(32'hbc14a9cf),
	.w5(32'h3b5fda65),
	.w6(32'hbbf06d9a),
	.w7(32'hbb69b0e1),
	.w8(32'hbbd23356),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb3f0b),
	.w1(32'hba9a986f),
	.w2(32'h3a883390),
	.w3(32'hbbb65fd2),
	.w4(32'hbcfe44fb),
	.w5(32'hbb3342fe),
	.w6(32'h3b8802e0),
	.w7(32'hbc812744),
	.w8(32'hbc09d3ca),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c672b11),
	.w1(32'hbb72284c),
	.w2(32'h38860218),
	.w3(32'h3ca617e8),
	.w4(32'hbc242e2c),
	.w5(32'hbc490ec1),
	.w6(32'h3bb23d3d),
	.w7(32'hbc1a305b),
	.w8(32'hb9d9cfa3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88fc0a1),
	.w1(32'hb9d4458e),
	.w2(32'hbc186bef),
	.w3(32'h3c0e2194),
	.w4(32'h3ba54d3e),
	.w5(32'hbc207196),
	.w6(32'hb9f432de),
	.w7(32'hbbc13459),
	.w8(32'hbab5df93),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb576576),
	.w1(32'hbbf87983),
	.w2(32'hbc68d354),
	.w3(32'h38637e1d),
	.w4(32'hbba9f1e5),
	.w5(32'hbb3a9ac1),
	.w6(32'hbbb04560),
	.w7(32'hbbd8785a),
	.w8(32'hbc313a03),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4db7e4),
	.w1(32'hb9de0e77),
	.w2(32'hbba1ec50),
	.w3(32'hbc4679ae),
	.w4(32'h3c5975ec),
	.w5(32'hbc8adae7),
	.w6(32'hbc4cf623),
	.w7(32'h3b2a7198),
	.w8(32'hbb2e44ec),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3ca4e),
	.w1(32'hbba6d75c),
	.w2(32'h3b70a27c),
	.w3(32'hba666968),
	.w4(32'hbc00d581),
	.w5(32'hbb5d7522),
	.w6(32'h3b51fc03),
	.w7(32'hbbfbbfc3),
	.w8(32'hbb617b57),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc134574),
	.w1(32'hbabd4134),
	.w2(32'hbba99830),
	.w3(32'h3c2a3f7c),
	.w4(32'h3c1b0e54),
	.w5(32'hbb44cb5b),
	.w6(32'hbb2ae3ed),
	.w7(32'hb9d6778e),
	.w8(32'hbbc6ced8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc67bcd),
	.w1(32'hba023475),
	.w2(32'hbb32df2d),
	.w3(32'hbbb0e371),
	.w4(32'hbbb5c7ff),
	.w5(32'hbc4038e8),
	.w6(32'hbb81f227),
	.w7(32'hbc2d8f60),
	.w8(32'hbbe24c8b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03c295),
	.w1(32'hbabeec50),
	.w2(32'hbba486cd),
	.w3(32'hbc14a2c9),
	.w4(32'h3b7ddb1b),
	.w5(32'h3bd898eb),
	.w6(32'hbc3bb7a1),
	.w7(32'hb9c8e7da),
	.w8(32'hbbd61f0f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dbf7b),
	.w1(32'hbbfe1ffa),
	.w2(32'hbbe75840),
	.w3(32'hbb1f4ca7),
	.w4(32'hbc6ae1ff),
	.w5(32'hbc0fc891),
	.w6(32'hbb8e6944),
	.w7(32'hbc090476),
	.w8(32'hbc20cbd9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11df54),
	.w1(32'h3a05bf83),
	.w2(32'h3bc665d6),
	.w3(32'hbb6987e5),
	.w4(32'h3bda0355),
	.w5(32'h3c28fc0a),
	.w6(32'hbab7e8eb),
	.w7(32'hbb1af472),
	.w8(32'h3ac350d2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c033f8f),
	.w1(32'h3ae17a3e),
	.w2(32'h3bdea907),
	.w3(32'h3b99fbd8),
	.w4(32'h3b95502d),
	.w5(32'h3b9cd1e8),
	.w6(32'hbb539ed4),
	.w7(32'h3b871f25),
	.w8(32'h3a4e94d0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c053819),
	.w1(32'hbc5c93fc),
	.w2(32'hbbfb8581),
	.w3(32'h3c4d3d28),
	.w4(32'hbba7ccf3),
	.w5(32'h3d11f414),
	.w6(32'h397bbb1b),
	.w7(32'hba1eabc6),
	.w8(32'h3ad28495),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21f397),
	.w1(32'hbb943976),
	.w2(32'hbc22f533),
	.w3(32'hbc17daed),
	.w4(32'hbc072ae5),
	.w5(32'hbc6457ac),
	.w6(32'hbbf08a9a),
	.w7(32'hbc357990),
	.w8(32'hbc448969),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04ae09),
	.w1(32'h3b2b7132),
	.w2(32'h3baf0990),
	.w3(32'hbc385194),
	.w4(32'h3ae90927),
	.w5(32'hbb79a68a),
	.w6(32'hbc3e5e2e),
	.w7(32'h3b090646),
	.w8(32'hbb582385),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a2f45),
	.w1(32'hbb3c540f),
	.w2(32'hbbe955f1),
	.w3(32'h3baca7ac),
	.w4(32'hbc0063d1),
	.w5(32'hbbc773ab),
	.w6(32'h3b55b23d),
	.w7(32'h3b1c4e16),
	.w8(32'hbbbc881f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa28b4b),
	.w1(32'hbb596f36),
	.w2(32'hbaa31a8a),
	.w3(32'hba8a30ec),
	.w4(32'hbb5a794b),
	.w5(32'hbbda4f78),
	.w6(32'h3b52ad60),
	.w7(32'h3ade1188),
	.w8(32'hbbb3d21c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99b66b),
	.w1(32'hbb71e9ef),
	.w2(32'hbb4e7afb),
	.w3(32'hb924eb1a),
	.w4(32'hbb999674),
	.w5(32'hbbe56733),
	.w6(32'hbb6156f8),
	.w7(32'h3b0fe68a),
	.w8(32'hbbdb0ebb),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f207c),
	.w1(32'h3bb05494),
	.w2(32'h399380ff),
	.w3(32'h3b110545),
	.w4(32'h3cf88eea),
	.w5(32'h3b4871a2),
	.w6(32'h3b0d8584),
	.w7(32'h3c9ecf17),
	.w8(32'h3c04fcef),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca82f6),
	.w1(32'hbc35452b),
	.w2(32'hbc59b268),
	.w3(32'hbd022ae3),
	.w4(32'hbc64641e),
	.w5(32'h3b3f9d31),
	.w6(32'hbbad861a),
	.w7(32'hbcd3e361),
	.w8(32'h3be41579),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc105dc1),
	.w1(32'hbb3c5073),
	.w2(32'hbbd02df6),
	.w3(32'hbbdeaefa),
	.w4(32'hbbb5dc1c),
	.w5(32'hbc449852),
	.w6(32'hbc205189),
	.w7(32'hbbe9e5bb),
	.w8(32'hbc058e82),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8bcd4),
	.w1(32'hbc5bba6a),
	.w2(32'hbc8e054e),
	.w3(32'hbbcc4581),
	.w4(32'hbc2a6263),
	.w5(32'h3bf21ce3),
	.w6(32'hbbb17e13),
	.w7(32'h3b271b41),
	.w8(32'hbbc0dcc7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5d055),
	.w1(32'h3a6497fa),
	.w2(32'h3ba349aa),
	.w3(32'h3927c27c),
	.w4(32'h3ba00678),
	.w5(32'h3ad640e1),
	.w6(32'hbb14369e),
	.w7(32'h3c50b254),
	.w8(32'hbb1f3dc6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8904e7),
	.w1(32'h3b67087b),
	.w2(32'hbbc7e425),
	.w3(32'h3c18ab3a),
	.w4(32'hba9903e8),
	.w5(32'hbabef45b),
	.w6(32'hbacbe2a2),
	.w7(32'h3b4b0b90),
	.w8(32'hbc065b79),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03ea68),
	.w1(32'hbb9be63e),
	.w2(32'hbc19ae12),
	.w3(32'hba3c68bc),
	.w4(32'hbc1ead32),
	.w5(32'hbab98b22),
	.w6(32'h3a47ac85),
	.w7(32'hbc07f873),
	.w8(32'hbbfcd6fd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc105623),
	.w1(32'h3c44e87c),
	.w2(32'h3b985acc),
	.w3(32'h3c6b944f),
	.w4(32'h3caebc90),
	.w5(32'h3c5c92b6),
	.w6(32'hbc23f61a),
	.w7(32'h3c40f07d),
	.w8(32'hba86cb2c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce0efe),
	.w1(32'h3b13bb1c),
	.w2(32'h3bc4bdc4),
	.w3(32'hbc5eb7b5),
	.w4(32'h3baca552),
	.w5(32'hbb2880b0),
	.w6(32'h3b94dc9e),
	.w7(32'hb9d09ba1),
	.w8(32'h3bbcfa5b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c033cef),
	.w1(32'h394d5e06),
	.w2(32'h38980ff0),
	.w3(32'h3c301678),
	.w4(32'hbc905b72),
	.w5(32'hbb354c50),
	.w6(32'h3bcfb0f1),
	.w7(32'hbbbce2d1),
	.w8(32'h39715ca3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7665a6),
	.w1(32'hbb8d25c3),
	.w2(32'h39fcb98a),
	.w3(32'h3cbe19e0),
	.w4(32'hba3791fb),
	.w5(32'h3c1895bb),
	.w6(32'h3c22b8b8),
	.w7(32'hb713be41),
	.w8(32'hbc02a162),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b654992),
	.w1(32'h3c05f4eb),
	.w2(32'hba9e4002),
	.w3(32'hbbd1609f),
	.w4(32'hbaa30ecf),
	.w5(32'hb96a045d),
	.w6(32'h3b479d69),
	.w7(32'h3a821a96),
	.w8(32'hbb5cad54),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8700bd),
	.w1(32'hba6efaa5),
	.w2(32'hbc2095e1),
	.w3(32'hbaabfda7),
	.w4(32'hbbb6ffb7),
	.w5(32'hbb931d98),
	.w6(32'hba986ea1),
	.w7(32'hbbbcaa34),
	.w8(32'hbc83ca4f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc805b6e),
	.w1(32'h3bf5beb8),
	.w2(32'h3a85cb07),
	.w3(32'hbc6c2187),
	.w4(32'h3bb1064c),
	.w5(32'hbbf1bb95),
	.w6(32'hbcb8e546),
	.w7(32'h3ac5cd2b),
	.w8(32'hbbecb816),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dc184),
	.w1(32'h3bb156a5),
	.w2(32'h3bc1fc9a),
	.w3(32'hbb9d2978),
	.w4(32'h3b1952fb),
	.w5(32'h3c272dbf),
	.w6(32'hbb7e884a),
	.w7(32'h3ab6258e),
	.w8(32'hbaf850e6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bede8b2),
	.w1(32'hba59d86a),
	.w2(32'hbb839ce5),
	.w3(32'h3c037417),
	.w4(32'hbb7534f2),
	.w5(32'h3b5c7d19),
	.w6(32'hbac840e5),
	.w7(32'h3c049b57),
	.w8(32'h3bcf88d7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab97d98),
	.w1(32'hba5115be),
	.w2(32'h39a785a2),
	.w3(32'h3b969d98),
	.w4(32'hbb1f4226),
	.w5(32'hbbe4d894),
	.w6(32'h3b73a8ab),
	.w7(32'hba8c99d1),
	.w8(32'hbae59af4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64f1fe),
	.w1(32'h39d99ee7),
	.w2(32'hbb0afbb2),
	.w3(32'hbbfd6791),
	.w4(32'h3af2a9b3),
	.w5(32'h3b1c495a),
	.w6(32'hbb92f964),
	.w7(32'hba29393b),
	.w8(32'h39877498),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e8a6f5),
	.w1(32'hbad9426e),
	.w2(32'hbb3a51ac),
	.w3(32'hbb1b2a94),
	.w4(32'hbc115593),
	.w5(32'hbbbaf1b5),
	.w6(32'hbb4fc0c5),
	.w7(32'hba971315),
	.w8(32'hba5c4cbc),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9b006),
	.w1(32'hbb8d6186),
	.w2(32'hbbe7858a),
	.w3(32'hbc1aec15),
	.w4(32'hbb62da8c),
	.w5(32'h3b036ee6),
	.w6(32'hbb25dbbd),
	.w7(32'hbbeb02d6),
	.w8(32'hbbf44e79),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc007a09),
	.w1(32'h3be6a323),
	.w2(32'h3b3df1e7),
	.w3(32'hbbb41efa),
	.w4(32'h3bbf2e68),
	.w5(32'h3b53c0d8),
	.w6(32'hbbfcd017),
	.w7(32'hbb4786b8),
	.w8(32'h3a0f1b15),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be91fc5),
	.w1(32'h3acb7312),
	.w2(32'hbbe135a6),
	.w3(32'h3c252a01),
	.w4(32'hba48a261),
	.w5(32'hbb0f5add),
	.w6(32'hba95e8b9),
	.w7(32'hbb44ea98),
	.w8(32'h3848800d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1e215),
	.w1(32'h3a95a29b),
	.w2(32'hbb786728),
	.w3(32'hbba5383d),
	.w4(32'h3ad78904),
	.w5(32'h3af4863c),
	.w6(32'hba8ebd7b),
	.w7(32'h3b352e8e),
	.w8(32'h3b14bdd1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b910369),
	.w1(32'h3b41777d),
	.w2(32'hbb65223e),
	.w3(32'h3b77006d),
	.w4(32'hbb8bb6b8),
	.w5(32'hbb814779),
	.w6(32'h3ad90724),
	.w7(32'hbb2bc6be),
	.w8(32'hbbe1501e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b2799),
	.w1(32'hb9788bd9),
	.w2(32'hbbcd4f90),
	.w3(32'h3b19e4dc),
	.w4(32'h3a80e370),
	.w5(32'hbbb1cf60),
	.w6(32'hbb0f5570),
	.w7(32'h3b1a988a),
	.w8(32'hbb6e8579),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4a3ab),
	.w1(32'h3b0ad7ff),
	.w2(32'hb9e1e006),
	.w3(32'hbacb1181),
	.w4(32'hbb8d693a),
	.w5(32'hbb9e2416),
	.w6(32'hbb62448e),
	.w7(32'hba8aae12),
	.w8(32'hbb6f31db),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acc065),
	.w1(32'hbbb73992),
	.w2(32'hbba5a0b1),
	.w3(32'hbb8bd556),
	.w4(32'hb97190f4),
	.w5(32'hbb34bcca),
	.w6(32'hbaf83e3e),
	.w7(32'h3ba0185a),
	.w8(32'h3b269dfa),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a994d),
	.w1(32'hbae45687),
	.w2(32'h3b58a552),
	.w3(32'hbab7bca0),
	.w4(32'h3c176dab),
	.w5(32'h3c5865bf),
	.w6(32'h3ab95f0e),
	.w7(32'h3b87d3a3),
	.w8(32'hbc2f644a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bdda3),
	.w1(32'hbaf859be),
	.w2(32'h39fd2169),
	.w3(32'h3b0e0ee2),
	.w4(32'hbb442fd6),
	.w5(32'hbaa16554),
	.w6(32'hb8f2eb76),
	.w7(32'h3b0842e1),
	.w8(32'hbadc3501),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfdcfc),
	.w1(32'h3aca5bc7),
	.w2(32'hbaff5de1),
	.w3(32'hbb98db26),
	.w4(32'h3c0d918a),
	.w5(32'h388be4c0),
	.w6(32'h3a6d6421),
	.w7(32'hbbca6d3c),
	.w8(32'hbb74f5d4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33a7cc),
	.w1(32'h3b23b1c9),
	.w2(32'hba101232),
	.w3(32'hbba2155f),
	.w4(32'h3b097c44),
	.w5(32'h3b9a40ae),
	.w6(32'hb98f4ed9),
	.w7(32'hbb528403),
	.w8(32'hb994217d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad20be),
	.w1(32'hbadb5905),
	.w2(32'hbbbd03b8),
	.w3(32'h3b231402),
	.w4(32'hbae6f5b1),
	.w5(32'h3b89b1ed),
	.w6(32'hb9831716),
	.w7(32'hba82d630),
	.w8(32'h3b3b62cc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b571d),
	.w1(32'h3b42c3c2),
	.w2(32'hb9c096e3),
	.w3(32'hbb83f44b),
	.w4(32'h3c27d7a5),
	.w5(32'h3c854d9c),
	.w6(32'hbb023795),
	.w7(32'h3a58a06f),
	.w8(32'hbb1ce38e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace127e),
	.w1(32'hbb713efb),
	.w2(32'h3a10c0bd),
	.w3(32'h3c28c666),
	.w4(32'hbac07357),
	.w5(32'h3a6aa6ca),
	.w6(32'hbc3422fd),
	.w7(32'hbc0ec631),
	.w8(32'hbb900ff1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7acdc1),
	.w1(32'h3a1a7a8f),
	.w2(32'hba5472c6),
	.w3(32'h3b19c3b3),
	.w4(32'h3a1a9b51),
	.w5(32'h38047826),
	.w6(32'h3991cd72),
	.w7(32'hb9f07834),
	.w8(32'hba0d4e66),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbece216),
	.w1(32'h3adc88ad),
	.w2(32'h3c0b9e3a),
	.w3(32'hbb7a3210),
	.w4(32'h3bf95ef2),
	.w5(32'h3b983e3b),
	.w6(32'hbbb6798f),
	.w7(32'hbba122fd),
	.w8(32'hbc1f5a8d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f3f8b),
	.w1(32'hbaf49b1c),
	.w2(32'h3b05e728),
	.w3(32'h3a72ab8e),
	.w4(32'h3a5a3753),
	.w5(32'h3aa685c7),
	.w6(32'h3b239d88),
	.w7(32'h3ab052bd),
	.w8(32'hbbf62e62),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65d423),
	.w1(32'h37c8696d),
	.w2(32'hba0032e5),
	.w3(32'hbb4226a4),
	.w4(32'h3b814a78),
	.w5(32'h3c13a18f),
	.w6(32'hbc0e70b9),
	.w7(32'h39ab68a4),
	.w8(32'hbb791be8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eb71e),
	.w1(32'h3aa6a2eb),
	.w2(32'hbb8a2531),
	.w3(32'h3b81b8aa),
	.w4(32'h3c64591d),
	.w5(32'h3cea68e7),
	.w6(32'hbb540453),
	.w7(32'hbc09b93d),
	.w8(32'hbc629a3f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9db3c5),
	.w1(32'hba6cad67),
	.w2(32'hbc1e35dc),
	.w3(32'h3c68051d),
	.w4(32'hbb00bb23),
	.w5(32'hbb3ab09b),
	.w6(32'hbbec551b),
	.w7(32'h3ba8134a),
	.w8(32'h3aedf45f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb833eb91),
	.w1(32'hbbb7bea8),
	.w2(32'hbc1a37a7),
	.w3(32'h38e991ff),
	.w4(32'hbb21124d),
	.w5(32'h3ba03fe0),
	.w6(32'h3b8bd211),
	.w7(32'hbba72f82),
	.w8(32'hbb67a088),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadde660),
	.w1(32'h3b02b1fe),
	.w2(32'hbb764029),
	.w3(32'h3b3ad0ac),
	.w4(32'hba62bbd0),
	.w5(32'hbb8f37d4),
	.w6(32'h3ac29501),
	.w7(32'hbbfa605e),
	.w8(32'hbbe2f0cc),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eae7e),
	.w1(32'h3a9b5b2c),
	.w2(32'hbb7e9e4d),
	.w3(32'hbb8dfd38),
	.w4(32'h3afc67e5),
	.w5(32'hbb8ba510),
	.w6(32'hbbe95871),
	.w7(32'hbc088bf3),
	.w8(32'hbbd35dd7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fef9f),
	.w1(32'hbc1479d9),
	.w2(32'hbb0787a0),
	.w3(32'hbc01025c),
	.w4(32'hbba23b40),
	.w5(32'h3a81797e),
	.w6(32'hbc0d62a8),
	.w7(32'h3b40a7c1),
	.w8(32'h3c297ec5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0b2ba),
	.w1(32'h3b64bdc3),
	.w2(32'hbba1fad4),
	.w3(32'h3a580b66),
	.w4(32'h3c383095),
	.w5(32'h3c9ca6f6),
	.w6(32'h3b667ca1),
	.w7(32'h3abfbf1e),
	.w8(32'h3a7a4ff3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fcc4c8),
	.w1(32'hbb6bf959),
	.w2(32'hbafcc708),
	.w3(32'h3bb50e85),
	.w4(32'hbb0e4734),
	.w5(32'hbb50dc25),
	.w6(32'hbb7ae882),
	.w7(32'hbbc680d7),
	.w8(32'hbc142f17),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba67351),
	.w1(32'hbb94ba6d),
	.w2(32'hbbb78444),
	.w3(32'hba8e3c90),
	.w4(32'hbaeac5b8),
	.w5(32'h3aea8415),
	.w6(32'h39c17b5b),
	.w7(32'h3acae284),
	.w8(32'h3b5d0d09),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59c5c6),
	.w1(32'hb953a8d6),
	.w2(32'hbace5bdb),
	.w3(32'hbad99e36),
	.w4(32'h39b0a817),
	.w5(32'hbba9b69e),
	.w6(32'h3c109cde),
	.w7(32'h3a83ffc8),
	.w8(32'hb9949e06),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb342d6b),
	.w1(32'hbbc7e2d5),
	.w2(32'hbbf002b8),
	.w3(32'hbbadfd35),
	.w4(32'h3aaad75e),
	.w5(32'h3c37ef1e),
	.w6(32'hbab99871),
	.w7(32'hbb315544),
	.w8(32'hbb24728f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c76fd),
	.w1(32'hbacf4e41),
	.w2(32'hbbd423a0),
	.w3(32'h3bc2cf67),
	.w4(32'hbacd1ac0),
	.w5(32'hbada5104),
	.w6(32'hbb66ba4f),
	.w7(32'hbb9fbd96),
	.w8(32'hbbbb15ef),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cb372),
	.w1(32'h3ad57825),
	.w2(32'h3aaa53f3),
	.w3(32'hbb07f679),
	.w4(32'hb9185bff),
	.w5(32'hb9daae71),
	.w6(32'hbb474572),
	.w7(32'hb9985aa1),
	.w8(32'hba934781),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07e378),
	.w1(32'hbba15ed9),
	.w2(32'h3be29b03),
	.w3(32'hba97cfe4),
	.w4(32'hbad423b8),
	.w5(32'hbafc17de),
	.w6(32'hbb2c4d8b),
	.w7(32'h3b3f6830),
	.w8(32'hbb0456af),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dc77c),
	.w1(32'hba87ddc7),
	.w2(32'hba083dcf),
	.w3(32'hbc259ae1),
	.w4(32'h3a6d5f79),
	.w5(32'h3ba246d3),
	.w6(32'hbab93ef5),
	.w7(32'hbb6852c6),
	.w8(32'hbb6aee58),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9ffe4),
	.w1(32'hbb558a38),
	.w2(32'hbaacc44d),
	.w3(32'h3ad1a6dc),
	.w4(32'h3ba23060),
	.w5(32'h3bd90cf4),
	.w6(32'hbb1ab740),
	.w7(32'hba4b99be),
	.w8(32'hbb30cbd7),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ab41eb),
	.w1(32'h3bf5a007),
	.w2(32'h3b36cb36),
	.w3(32'h3c09ef05),
	.w4(32'hbbfd3c8e),
	.w5(32'hbbaf03bf),
	.w6(32'hbb686230),
	.w7(32'hbb8842a3),
	.w8(32'h39c54dd8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d1f11),
	.w1(32'hb9f59230),
	.w2(32'hbb5abf01),
	.w3(32'hbb90e9f5),
	.w4(32'hba646511),
	.w5(32'hbb9de885),
	.w6(32'h3a544412),
	.w7(32'hbaa11a1f),
	.w8(32'hbb69e711),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6e97e),
	.w1(32'hbb1fc358),
	.w2(32'hbad75546),
	.w3(32'hbadf6297),
	.w4(32'h3a0a36dc),
	.w5(32'hb9d7edc6),
	.w6(32'h3a8515bc),
	.w7(32'hb9fa9644),
	.w8(32'h39a916e2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ad192),
	.w1(32'hbc24ba7c),
	.w2(32'hbb9121e3),
	.w3(32'hbbbe4aa9),
	.w4(32'hbac05245),
	.w5(32'h3c653414),
	.w6(32'hbae8bc35),
	.w7(32'hbacc2f5e),
	.w8(32'hbb91414a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c5dce),
	.w1(32'hbaecd8ab),
	.w2(32'hbb4a2606),
	.w3(32'h3a11bb1f),
	.w4(32'h3a82ac49),
	.w5(32'hbb8ac5e8),
	.w6(32'hbb1f1c79),
	.w7(32'h3b193e02),
	.w8(32'hba6b9012),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba995857),
	.w1(32'h3b9b7201),
	.w2(32'h3b8bf920),
	.w3(32'h3aadd367),
	.w4(32'h3ba72890),
	.w5(32'h3b00a95f),
	.w6(32'hbb8ef208),
	.w7(32'h3c0c6965),
	.w8(32'h3beadadc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b470b75),
	.w1(32'h3b932eb0),
	.w2(32'h3b67c73c),
	.w3(32'h3a20138e),
	.w4(32'hb8dc7594),
	.w5(32'h3b1a28b1),
	.w6(32'h3bb0fcab),
	.w7(32'h3bce363d),
	.w8(32'h3ab31816),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b955a3),
	.w1(32'h398b1cca),
	.w2(32'h3a9dbc82),
	.w3(32'h3b977e0e),
	.w4(32'hbb61390d),
	.w5(32'hb9d85463),
	.w6(32'hba78586a),
	.w7(32'hba31fee8),
	.w8(32'hbb9103a1),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15d038),
	.w1(32'h3a041c4c),
	.w2(32'hbb920849),
	.w3(32'hbb235da8),
	.w4(32'hbbb0995e),
	.w5(32'hbb7aed63),
	.w6(32'hbbd38a0c),
	.w7(32'hbb627ebe),
	.w8(32'hbaa0700b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb230302),
	.w1(32'h3b2e8ffd),
	.w2(32'h39a3bb3e),
	.w3(32'hb9ac6bee),
	.w4(32'hbb10c649),
	.w5(32'hbbf92d21),
	.w6(32'hbbf43464),
	.w7(32'h3b1ba845),
	.w8(32'h3b48aeed),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad76a00),
	.w1(32'hbab524da),
	.w2(32'h3a5d84e2),
	.w3(32'h3a7eae9e),
	.w4(32'h3b80cfaf),
	.w5(32'hbb35c313),
	.w6(32'h3bb0f035),
	.w7(32'hbb2fc86f),
	.w8(32'h38ece340),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e22f5),
	.w1(32'hbac59f62),
	.w2(32'h3b72f6a7),
	.w3(32'hbb68e68c),
	.w4(32'hba3f3037),
	.w5(32'hbb01f650),
	.w6(32'hbba22101),
	.w7(32'hbb8ab4b7),
	.w8(32'hbad5944b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6709c8),
	.w1(32'hbb4b2071),
	.w2(32'hbb6036f0),
	.w3(32'hbb2e1f8e),
	.w4(32'h3ad80b21),
	.w5(32'h3c091fee),
	.w6(32'hbb4af5a5),
	.w7(32'hbb32ab12),
	.w8(32'hbbbec497),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61a59c),
	.w1(32'h3a9600fd),
	.w2(32'h3a3e7ef3),
	.w3(32'h3b4be6e6),
	.w4(32'h3a0e56e4),
	.w5(32'hba76508c),
	.w6(32'h3b42378b),
	.w7(32'h3b34040f),
	.w8(32'hb8431472),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c89dd3),
	.w1(32'hbb922333),
	.w2(32'hbb8a8c41),
	.w3(32'h3b50a247),
	.w4(32'hbb47f8c5),
	.w5(32'h3bcef714),
	.w6(32'h3b9ec34f),
	.w7(32'hba3ba7da),
	.w8(32'hbb83bcef),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2343b),
	.w1(32'hbab5b5db),
	.w2(32'h3b2a62a9),
	.w3(32'hba1eafb7),
	.w4(32'h3b30adf5),
	.w5(32'h3c227eb3),
	.w6(32'hbb582bba),
	.w7(32'h3b297593),
	.w8(32'h39bc73e9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeaed45),
	.w1(32'hbbce4902),
	.w2(32'hbb87b234),
	.w3(32'h3b961b70),
	.w4(32'hbc4d093e),
	.w5(32'h39a4112f),
	.w6(32'h3b06011b),
	.w7(32'hbba03f6d),
	.w8(32'hbba4d3ed),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85bf02),
	.w1(32'h3aa8e9c8),
	.w2(32'h3ba140df),
	.w3(32'hbb11223d),
	.w4(32'h3c0c30e7),
	.w5(32'h3a2ec8dd),
	.w6(32'hbb4bc978),
	.w7(32'hbb4784b4),
	.w8(32'hbbf7f6e3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7d279),
	.w1(32'h3aef00c2),
	.w2(32'h3a0f5b4d),
	.w3(32'h398a47bb),
	.w4(32'h3c0d85e7),
	.w5(32'h3c421843),
	.w6(32'hba0584c1),
	.w7(32'hbbd9ddf8),
	.w8(32'hbb205599),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06b715),
	.w1(32'h3ade8e0b),
	.w2(32'hbb008a1c),
	.w3(32'h3c338fae),
	.w4(32'hbb5122f2),
	.w5(32'h3abd64e1),
	.w6(32'hbb50e297),
	.w7(32'hbaad9713),
	.w8(32'hb9dce354),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64a375),
	.w1(32'hbb0d9594),
	.w2(32'hbbd37d07),
	.w3(32'hbb3ff28f),
	.w4(32'h3b5ba508),
	.w5(32'h3c338712),
	.w6(32'hba5634fe),
	.w7(32'hbad8f835),
	.w8(32'hbbc02c27),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7252cd),
	.w1(32'h399bb97c),
	.w2(32'h3a26b47c),
	.w3(32'h3c1cc3f9),
	.w4(32'hbb84260a),
	.w5(32'h3b80c6f2),
	.w6(32'hbb466ecf),
	.w7(32'h39929b15),
	.w8(32'h3a5de79a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cf831),
	.w1(32'h3acb9efe),
	.w2(32'h3a0d8344),
	.w3(32'h3bcef199),
	.w4(32'hb8317d17),
	.w5(32'hba5b7ec1),
	.w6(32'h3b043d2c),
	.w7(32'hbb62e1b5),
	.w8(32'hb9e00c7d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0947),
	.w1(32'hbbd012d9),
	.w2(32'hbbc7cbd9),
	.w3(32'hba3284b7),
	.w4(32'hbafaf735),
	.w5(32'hbb5919ab),
	.w6(32'h39a2c26c),
	.w7(32'h3a474f94),
	.w8(32'hbb665144),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92bf91),
	.w1(32'hba1d893e),
	.w2(32'hbc62cc47),
	.w3(32'hbb91ef98),
	.w4(32'hbba1f32d),
	.w5(32'hbae89385),
	.w6(32'hbacbbd77),
	.w7(32'h3994339e),
	.w8(32'hbb752449),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d9b00),
	.w1(32'h3b1cb82b),
	.w2(32'h3b12dcdf),
	.w3(32'h3a3f8658),
	.w4(32'h3a048efc),
	.w5(32'hb9da98a6),
	.w6(32'h38d2970c),
	.w7(32'h3b29fbdd),
	.w8(32'h3b414367),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c73bb),
	.w1(32'hbafe9738),
	.w2(32'hba9a8be2),
	.w3(32'h3b277679),
	.w4(32'hba99f7fb),
	.w5(32'h3a84cc30),
	.w6(32'h3aaf5da3),
	.w7(32'hbadd13c9),
	.w8(32'hbbba3e82),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bbf3c),
	.w1(32'hba87ba68),
	.w2(32'hbad835ab),
	.w3(32'hbc2f2b47),
	.w4(32'h3b19c574),
	.w5(32'h3bc9cf95),
	.w6(32'hbc05e4a9),
	.w7(32'hbb1f5ba2),
	.w8(32'hbaed15fe),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa670b),
	.w1(32'h3bb4a25c),
	.w2(32'h3c0e321e),
	.w3(32'h3c1469e4),
	.w4(32'hbb42df66),
	.w5(32'h3af6632e),
	.w6(32'hbabd1b5a),
	.w7(32'hbac41ef5),
	.w8(32'hbb4039d1),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b882e12),
	.w1(32'h3b5acf63),
	.w2(32'hbbca2df0),
	.w3(32'hba328dad),
	.w4(32'hb9cd24b0),
	.w5(32'hbc077cbb),
	.w6(32'hbb78f9dc),
	.w7(32'hbb556879),
	.w8(32'hbbbeaa42),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fbbc0),
	.w1(32'hbbc9f14f),
	.w2(32'hbb95492d),
	.w3(32'hbb0ef50c),
	.w4(32'hbaff49b0),
	.w5(32'hbac75a1b),
	.w6(32'hbb3c85e9),
	.w7(32'h36a01511),
	.w8(32'hba94d0ed),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6be1c3),
	.w1(32'h3bb06c88),
	.w2(32'h3a39bc22),
	.w3(32'hbbb6a6ad),
	.w4(32'h3a019522),
	.w5(32'hbb8c7edb),
	.w6(32'hbb560422),
	.w7(32'h3b5b411e),
	.w8(32'hbada0aed),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b147cad),
	.w1(32'h3ab93a1b),
	.w2(32'h3abc6b6a),
	.w3(32'h3a2f1a39),
	.w4(32'hbb8df4c1),
	.w5(32'hbb3eeeca),
	.w6(32'h3b9bd53b),
	.w7(32'hb9e5bf94),
	.w8(32'hbba1b2c5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95c62f),
	.w1(32'hbaef5760),
	.w2(32'hbbace2b5),
	.w3(32'hba502c52),
	.w4(32'hbabfaca0),
	.w5(32'hbb6a741e),
	.w6(32'h3b3c7238),
	.w7(32'hba3c64ca),
	.w8(32'hbb21c97d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87485d),
	.w1(32'hba73d2dd),
	.w2(32'hbb9333f9),
	.w3(32'hbb4a3547),
	.w4(32'hbae4e13d),
	.w5(32'hbb3d9836),
	.w6(32'h3bb06923),
	.w7(32'hba580c45),
	.w8(32'h3b582d4b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bf51e),
	.w1(32'h3ad44dd0),
	.w2(32'h3a398a87),
	.w3(32'hbb07e8fb),
	.w4(32'h3b9b60d8),
	.w5(32'h3b5dbecc),
	.w6(32'h3a22268e),
	.w7(32'hbb6edd72),
	.w8(32'h3a4e0dab),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dff60d),
	.w1(32'hb9d13a45),
	.w2(32'hbb5470f0),
	.w3(32'h3b605789),
	.w4(32'h3a20666c),
	.w5(32'hbb08416e),
	.w6(32'hbb7089eb),
	.w7(32'h3a87237f),
	.w8(32'hbba5d37b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d2746),
	.w1(32'hbb8bdf3d),
	.w2(32'h3a9e57db),
	.w3(32'hb9ec0257),
	.w4(32'hbb80f0d6),
	.w5(32'hbb3000dd),
	.w6(32'hbaa3f5c9),
	.w7(32'h3a9fdb1c),
	.w8(32'h3bb42079),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be42da8),
	.w1(32'hb89443db),
	.w2(32'hbbd67000),
	.w3(32'hbbc49c4a),
	.w4(32'hb9c61637),
	.w5(32'hbb8d9fb8),
	.w6(32'hba6fe74c),
	.w7(32'hba012f35),
	.w8(32'hbb7afd95),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fa09b),
	.w1(32'hbbbaf506),
	.w2(32'hbc21b7f4),
	.w3(32'hba35a177),
	.w4(32'hbb769fa8),
	.w5(32'hb995f87e),
	.w6(32'hbb9bbe21),
	.w7(32'hba984abf),
	.w8(32'hbc15781c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae4401),
	.w1(32'h3b81c3f3),
	.w2(32'hbb0fd4a5),
	.w3(32'hbb8f4580),
	.w4(32'hba07f9e0),
	.w5(32'hbba77ddd),
	.w6(32'hbbb09544),
	.w7(32'h3b1d2c0f),
	.w8(32'h3b45a8d3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37821c61),
	.w1(32'hbc12d62f),
	.w2(32'hbc46de1e),
	.w3(32'hbbc87661),
	.w4(32'hbaa74b03),
	.w5(32'h3acac81c),
	.w6(32'hbb821cb1),
	.w7(32'h3a0f3402),
	.w8(32'hbb6ea0d5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb490895),
	.w1(32'hba9e04be),
	.w2(32'hbb192f1b),
	.w3(32'h3b142648),
	.w4(32'hbb99bb1a),
	.w5(32'hbbd51a48),
	.w6(32'h39f8a3f9),
	.w7(32'hbb4caf9e),
	.w8(32'hbb457dba),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977d5c1),
	.w1(32'hb9685841),
	.w2(32'hb9a82fc1),
	.w3(32'hb82d7dd8),
	.w4(32'h3b1382e2),
	.w5(32'h3abe6375),
	.w6(32'hbb104c25),
	.w7(32'h3aa91e37),
	.w8(32'hb9cd2af3),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4853b),
	.w1(32'h3bce9e72),
	.w2(32'h3b2bab64),
	.w3(32'hbba1e5ec),
	.w4(32'h3a68a36f),
	.w5(32'hbb5f79b6),
	.w6(32'hbb4b1508),
	.w7(32'h3b244f6f),
	.w8(32'h3b128297),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7db4a4),
	.w1(32'hbaa34377),
	.w2(32'hb9a3723a),
	.w3(32'hbbb121bf),
	.w4(32'h3b3a0814),
	.w5(32'h3a9edc9c),
	.w6(32'h3b0237bb),
	.w7(32'hba741cfc),
	.w8(32'hb859d637),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984dd0f),
	.w1(32'h3bfc2461),
	.w2(32'hba9e6cf2),
	.w3(32'hba0a221e),
	.w4(32'hbb14ee65),
	.w5(32'hbab42fbf),
	.w6(32'h3a3029bd),
	.w7(32'h3bc3c9a3),
	.w8(32'h3c04db75),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ea0f5),
	.w1(32'h3b544355),
	.w2(32'hb9051b55),
	.w3(32'h3c31a30b),
	.w4(32'hbb298ca3),
	.w5(32'hbb82a602),
	.w6(32'h3bc5d2d6),
	.w7(32'hbb562725),
	.w8(32'hbad99803),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47c2ce),
	.w1(32'hbaedb66a),
	.w2(32'hbc0da80c),
	.w3(32'hbb7d51a3),
	.w4(32'h3bcdd8b7),
	.w5(32'h3bbd7883),
	.w6(32'hbb52870f),
	.w7(32'h3b78ce68),
	.w8(32'h3bdf7806),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc43412),
	.w1(32'hb9adb9d2),
	.w2(32'h3a08bbe3),
	.w3(32'h3c0a9fad),
	.w4(32'hbbb6ccd0),
	.w5(32'hbbda3afd),
	.w6(32'h3b08d23d),
	.w7(32'hbb1233c3),
	.w8(32'hba6e2b00),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0badac),
	.w1(32'h3c0081d5),
	.w2(32'h3aeca6f2),
	.w3(32'hbb44b323),
	.w4(32'h3baf7a94),
	.w5(32'h3b4bcfad),
	.w6(32'hba84d9dd),
	.w7(32'hbb05803c),
	.w8(32'hba4f3ef7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad6ac2),
	.w1(32'h3988a81a),
	.w2(32'hbac02df6),
	.w3(32'h3b7a5568),
	.w4(32'h3a4c8d71),
	.w5(32'h3b64522d),
	.w6(32'hbb88169e),
	.w7(32'hba928502),
	.w8(32'h3ba47b01),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcd410),
	.w1(32'hba89e38d),
	.w2(32'hb9bc0ee7),
	.w3(32'hbae0fe48),
	.w4(32'hbb4696f1),
	.w5(32'hbb96062e),
	.w6(32'h39a84b4e),
	.w7(32'h3b8fb738),
	.w8(32'hba95a7ad),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6066b3),
	.w1(32'h3bae959b),
	.w2(32'h3af57e61),
	.w3(32'hba93585d),
	.w4(32'h3b9f9548),
	.w5(32'h3ab17e9b),
	.w6(32'h3b96a9a8),
	.w7(32'h3b272304),
	.w8(32'h385f7490),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70a0a3),
	.w1(32'hbaf26f3c),
	.w2(32'hbb99d99a),
	.w3(32'h3b829a76),
	.w4(32'hbb84f8bf),
	.w5(32'hbb9c0f85),
	.w6(32'hbb32827f),
	.w7(32'hbbc05828),
	.w8(32'hbbb76864),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3971c97b),
	.w1(32'h3b811e6b),
	.w2(32'h38612b08),
	.w3(32'h3b77576a),
	.w4(32'hbb6b4cd0),
	.w5(32'hbb4635ef),
	.w6(32'h3b024981),
	.w7(32'hbb822f2a),
	.w8(32'h3a61423a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff589b),
	.w1(32'hb9f5013a),
	.w2(32'h3967ae54),
	.w3(32'hbb2866dc),
	.w4(32'h3a949b69),
	.w5(32'h3b08a80e),
	.w6(32'hbb12b9a1),
	.w7(32'hbab13411),
	.w8(32'h3a46114a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0bf23),
	.w1(32'hbb357828),
	.w2(32'h3b961275),
	.w3(32'h3b27a4e5),
	.w4(32'hbb36c086),
	.w5(32'hba23a008),
	.w6(32'h397729de),
	.w7(32'h393ee0ab),
	.w8(32'h3b517b7e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad709f2),
	.w1(32'h3b97af9e),
	.w2(32'h3c070764),
	.w3(32'hbaddca98),
	.w4(32'hbb85ed59),
	.w5(32'hbbddae15),
	.w6(32'hba4e28cb),
	.w7(32'h3a9452a0),
	.w8(32'h3b59c6f5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c0323),
	.w1(32'hbadf3df0),
	.w2(32'hba9c0f6b),
	.w3(32'h3b8febe4),
	.w4(32'hbadcb0f6),
	.w5(32'hbbc18d81),
	.w6(32'h3c2fc115),
	.w7(32'hbb1f83e5),
	.w8(32'hbad780a4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2b1e8),
	.w1(32'hbb4da84e),
	.w2(32'h3a81e6c1),
	.w3(32'hbb3463c5),
	.w4(32'hbb84427f),
	.w5(32'h3797020c),
	.w6(32'h3a6c595f),
	.w7(32'hba3291d4),
	.w8(32'h3ad9d07d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h32ddc800),
	.w1(32'hbb9af030),
	.w2(32'hbb79fe53),
	.w3(32'h3a444a06),
	.w4(32'hbbaf8dee),
	.w5(32'hbbcfbea2),
	.w6(32'hbb0c81c4),
	.w7(32'hbb0d446a),
	.w8(32'hba02fff4),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f2057),
	.w1(32'h3af6db3a),
	.w2(32'h3af3d54e),
	.w3(32'hbaf93eb6),
	.w4(32'h3bf74713),
	.w5(32'h3b4d2e99),
	.w6(32'h3b0c9b7a),
	.w7(32'h3a66b4ac),
	.w8(32'hbbbe239d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0a386),
	.w1(32'h3b8068fb),
	.w2(32'h39211832),
	.w3(32'hba816b16),
	.w4(32'h3a5db081),
	.w5(32'hbbb5769e),
	.w6(32'hbac048fe),
	.w7(32'h3ae37f65),
	.w8(32'h395621cf),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b934840),
	.w1(32'hb895476a),
	.w2(32'h3b1e3133),
	.w3(32'hbb2f5f88),
	.w4(32'h3a6bc890),
	.w5(32'h3aea8998),
	.w6(32'h3bd48071),
	.w7(32'hbb6983a3),
	.w8(32'hbbc5f83e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ebfcb),
	.w1(32'h3bb448db),
	.w2(32'h3b9fcbeb),
	.w3(32'h3abbf594),
	.w4(32'h3a5f6abc),
	.w5(32'hb88ea9ff),
	.w6(32'hbbe80906),
	.w7(32'h3b724da6),
	.w8(32'h3b559c66),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba432b79),
	.w1(32'h3b4f888e),
	.w2(32'hbaa14aad),
	.w3(32'hb99fcadb),
	.w4(32'hb90985e9),
	.w5(32'h3b5c42a7),
	.w6(32'h3a1917de),
	.w7(32'h3bf3b7df),
	.w8(32'h3b7fbd85),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b256a43),
	.w1(32'hbac90d28),
	.w2(32'hbb94a216),
	.w3(32'h38e7c2b7),
	.w4(32'hbb4a42b1),
	.w5(32'h39fc8e9b),
	.w6(32'h3a5393b5),
	.w7(32'h3b64f7ee),
	.w8(32'h3ba3b481),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e04d9),
	.w1(32'h390dce36),
	.w2(32'hbbd16cf8),
	.w3(32'h3c0a0c10),
	.w4(32'h3b2acbfb),
	.w5(32'hbbc51246),
	.w6(32'h3bbb3ad6),
	.w7(32'h3b14e62c),
	.w8(32'h3a6a5750),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca3887),
	.w1(32'h3aaa754c),
	.w2(32'hba8d8672),
	.w3(32'hba993493),
	.w4(32'hbbc25fcd),
	.w5(32'hbc0e50c6),
	.w6(32'h3ba39e16),
	.w7(32'h3b816dc1),
	.w8(32'hbbbc38e2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b0248),
	.w1(32'h393d6b41),
	.w2(32'h3aa0907d),
	.w3(32'hbad89b8a),
	.w4(32'h3a477257),
	.w5(32'h3a0a712b),
	.w6(32'hbbaf7991),
	.w7(32'hbaa97c68),
	.w8(32'h3b347f06),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b016891),
	.w1(32'h3a5fe931),
	.w2(32'hbb70c658),
	.w3(32'hbb0523dc),
	.w4(32'h3b893a2e),
	.w5(32'h3a8cc4af),
	.w6(32'hbb552e2f),
	.w7(32'h3b3b953a),
	.w8(32'h3ba4f959),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4894c2),
	.w1(32'hbb8e0107),
	.w2(32'hba81b418),
	.w3(32'h3a75abbe),
	.w4(32'hbbfba1fd),
	.w5(32'hb992dc95),
	.w6(32'h3b9de248),
	.w7(32'h3ac32856),
	.w8(32'h3bb15005),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfa138),
	.w1(32'h3b398713),
	.w2(32'h3a6861d7),
	.w3(32'hbb869ee7),
	.w4(32'h3b8f5118),
	.w5(32'h3b2ee514),
	.w6(32'h39061ebd),
	.w7(32'hbb1cbf3f),
	.w8(32'h39b46d9f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13840b),
	.w1(32'h3b37babd),
	.w2(32'hba4ff1ae),
	.w3(32'hbadd7241),
	.w4(32'h3a0c0ebf),
	.w5(32'hbbfe7dd4),
	.w6(32'hba0e086f),
	.w7(32'hba9eee7c),
	.w8(32'hbb087b1d),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0493e),
	.w1(32'hbb4c9afc),
	.w2(32'hbb5932d8),
	.w3(32'h3b270a9b),
	.w4(32'h3b8acfdd),
	.w5(32'hbb9850cb),
	.w6(32'h3be3a7e0),
	.w7(32'hbb295841),
	.w8(32'hba10608e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395c114a),
	.w1(32'hbbfd303e),
	.w2(32'hbb9f0f25),
	.w3(32'hbb820766),
	.w4(32'hba2235a1),
	.w5(32'hbb83cc83),
	.w6(32'hbb970bc4),
	.w7(32'hbace1afe),
	.w8(32'hbae8c260),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc202742),
	.w1(32'hbb749ba7),
	.w2(32'h3a8eade6),
	.w3(32'hbb27c1df),
	.w4(32'hbba1f25e),
	.w5(32'hbba95cd3),
	.w6(32'h39b39edf),
	.w7(32'h3a572fd4),
	.w8(32'hbbb36ccd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc322b44),
	.w1(32'h3bc90acf),
	.w2(32'h3c08baee),
	.w3(32'h3aa591d4),
	.w4(32'h3b8db4c8),
	.w5(32'hbbe59cf8),
	.w6(32'hbbada36f),
	.w7(32'h3af6d152),
	.w8(32'hbb9b0651),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba33fb0),
	.w1(32'hbb1434a0),
	.w2(32'hba9798dc),
	.w3(32'hbbe429e5),
	.w4(32'h3712fcc0),
	.w5(32'hbb2505e1),
	.w6(32'hbb8332c1),
	.w7(32'h3ad747bb),
	.w8(32'h3b08acc1),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99719c6),
	.w1(32'hbbc658bd),
	.w2(32'hba645a37),
	.w3(32'hbb216c4b),
	.w4(32'hbb6e1d9b),
	.w5(32'hbb5d2e91),
	.w6(32'hb9fc7dd3),
	.w7(32'hbaee6c28),
	.w8(32'hbb6901af),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a82fc),
	.w1(32'h3b16e5ee),
	.w2(32'h38871921),
	.w3(32'h3bd7e756),
	.w4(32'h3a060020),
	.w5(32'hba922e4b),
	.w6(32'hba0512da),
	.w7(32'hbb82cb75),
	.w8(32'h39d22603),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeccc57),
	.w1(32'h3a168f10),
	.w2(32'hba6e2f60),
	.w3(32'h3b9f405d),
	.w4(32'h3b835a9e),
	.w5(32'h3b11c442),
	.w6(32'h3afcf039),
	.w7(32'h3b38cb48),
	.w8(32'h3a80dcff),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aeaae),
	.w1(32'hbaff4267),
	.w2(32'hbba3f120),
	.w3(32'h3b374a6d),
	.w4(32'h3b4a542a),
	.w5(32'h3b32632f),
	.w6(32'h3a8eb833),
	.w7(32'h3b1087fb),
	.w8(32'hbb07e757),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa214d),
	.w1(32'h3a2c3d0f),
	.w2(32'h3b0c5ae1),
	.w3(32'h3aa71d8c),
	.w4(32'hbae044c1),
	.w5(32'h3b21a371),
	.w6(32'h3a9c5720),
	.w7(32'hbb0ff571),
	.w8(32'hbaa545cb),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4771e4),
	.w1(32'hbbddfcfa),
	.w2(32'hbbcff6d1),
	.w3(32'hba4a09ca),
	.w4(32'h3a8c26b6),
	.w5(32'h3b0210f3),
	.w6(32'hbb3bddef),
	.w7(32'hbb8e5f17),
	.w8(32'hbad022e9),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36e217),
	.w1(32'hbb40e8f1),
	.w2(32'hbb9b644e),
	.w3(32'hbb258eeb),
	.w4(32'hbbcbc1c0),
	.w5(32'hba90e89a),
	.w6(32'h37aa4085),
	.w7(32'hbbb272dd),
	.w8(32'h3977f0b4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb097441),
	.w1(32'hb9956cf0),
	.w2(32'hbba2c252),
	.w3(32'h3bfe4dc6),
	.w4(32'hbba27c10),
	.w5(32'hbc88ad34),
	.w6(32'h3ba5c222),
	.w7(32'hbba1048d),
	.w8(32'hbc1a93fa),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe37d54),
	.w1(32'h3b15d6ef),
	.w2(32'h39fed5ad),
	.w3(32'hbba795df),
	.w4(32'h3b4270b6),
	.w5(32'h3bed6687),
	.w6(32'h3aed61c3),
	.w7(32'hbb1f76e0),
	.w8(32'hbbb4f37c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cc60f),
	.w1(32'h3bd6e942),
	.w2(32'h3c206702),
	.w3(32'hbad41cef),
	.w4(32'h3aee3859),
	.w5(32'hbbbaa376),
	.w6(32'hbb373829),
	.w7(32'hbbe09063),
	.w8(32'h3983d240),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0e295),
	.w1(32'hbaf9a434),
	.w2(32'hbb788f23),
	.w3(32'hbc04371a),
	.w4(32'hbb92364c),
	.w5(32'hbc0b67a6),
	.w6(32'h3b005d50),
	.w7(32'hba99f20d),
	.w8(32'hbb57980d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe5fc0),
	.w1(32'hba790b90),
	.w2(32'h3a8bd670),
	.w3(32'h3a2e0cb1),
	.w4(32'hbaef8285),
	.w5(32'h3a74de71),
	.w6(32'hba65d9e0),
	.w7(32'h3a3fd101),
	.w8(32'h3a3217e3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4117b),
	.w1(32'hbc028e2d),
	.w2(32'hbc10f38b),
	.w3(32'h3bb87492),
	.w4(32'hbbea32e1),
	.w5(32'hbc0cfcbf),
	.w6(32'hbb60f402),
	.w7(32'hbc2cfbe7),
	.w8(32'hbb81f2e0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb596043),
	.w1(32'h3b252131),
	.w2(32'h39d8b097),
	.w3(32'hbc528256),
	.w4(32'h390c7196),
	.w5(32'hbab15747),
	.w6(32'h3aecf1e1),
	.w7(32'hba7b3031),
	.w8(32'h3b135833),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399281a8),
	.w1(32'h3bbe2ac6),
	.w2(32'h3beac742),
	.w3(32'hb923e197),
	.w4(32'h3b6c390b),
	.w5(32'hbc5bded0),
	.w6(32'h3b404956),
	.w7(32'hba643c18),
	.w8(32'hbbf56057),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c200d10),
	.w1(32'h39fa08ca),
	.w2(32'h3bf2d50d),
	.w3(32'hba1ae480),
	.w4(32'hbc2f9ba7),
	.w5(32'hbc824d65),
	.w6(32'hb9965534),
	.w7(32'h3b3440a8),
	.w8(32'h3c7c5a97),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba721412),
	.w1(32'h3b9b694e),
	.w2(32'hba9ac29a),
	.w3(32'h3acaca01),
	.w4(32'h3be8770f),
	.w5(32'hba863422),
	.w6(32'h3877d013),
	.w7(32'h39c0642e),
	.w8(32'hba0ec410),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad26a07),
	.w1(32'h3b7fee52),
	.w2(32'h3ad302c7),
	.w3(32'hbb8bd866),
	.w4(32'h3ba9d4ad),
	.w5(32'h3b364221),
	.w6(32'h3ae574c5),
	.w7(32'hbbc7ecea),
	.w8(32'hbc4df164),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0aa09),
	.w1(32'h3ba2247f),
	.w2(32'h3ad76bb6),
	.w3(32'hbb9371ff),
	.w4(32'h3ba6956a),
	.w5(32'hbbba9655),
	.w6(32'hbb9dce81),
	.w7(32'h3af819f0),
	.w8(32'h3b1eb4d3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beeb5b7),
	.w1(32'hba73a880),
	.w2(32'h3ad04eed),
	.w3(32'hbb1887d0),
	.w4(32'hba66bd72),
	.w5(32'h3aa14984),
	.w6(32'hbafc80f2),
	.w7(32'h3ba4d414),
	.w8(32'h39d59df0),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84c56c),
	.w1(32'hbb87cb73),
	.w2(32'hbb0feca0),
	.w3(32'h3b820d90),
	.w4(32'h3ab015bb),
	.w5(32'h3c17fa59),
	.w6(32'hbab88cf1),
	.w7(32'h3ad495c8),
	.w8(32'h39974aab),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba921939),
	.w1(32'h3ad71f8b),
	.w2(32'hbbba4c81),
	.w3(32'h3b69ad59),
	.w4(32'hbb0f6f20),
	.w5(32'h3d1b3569),
	.w6(32'hba844725),
	.w7(32'h3c055cce),
	.w8(32'h3a10d734),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5018fd),
	.w1(32'h3af72995),
	.w2(32'h3b232f2d),
	.w3(32'h3cc3174d),
	.w4(32'hbbd8c055),
	.w5(32'hbc402c3e),
	.w6(32'hbc717828),
	.w7(32'h3b379630),
	.w8(32'hba58d8f0),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1037c6),
	.w1(32'hbb6bb08d),
	.w2(32'hbc1e9d67),
	.w3(32'hbc1842d2),
	.w4(32'h3c892175),
	.w5(32'h3cc6bbaf),
	.w6(32'hbc4b5f37),
	.w7(32'hbc3260c6),
	.w8(32'hbc1ebaa7),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82159b),
	.w1(32'h3c028190),
	.w2(32'h3abb9b98),
	.w3(32'hba7a1fc5),
	.w4(32'h3bdb1095),
	.w5(32'h3bcadd4e),
	.w6(32'h3aaace70),
	.w7(32'hbb8e759c),
	.w8(32'hbbad4012),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b376a7c),
	.w1(32'h3a63a3f0),
	.w2(32'h3a3bcc61),
	.w3(32'h3b85e0bf),
	.w4(32'hbaaaa47b),
	.w5(32'h3c603e7e),
	.w6(32'hbbb2a2b9),
	.w7(32'hba1a55e3),
	.w8(32'hbc31a2c4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6d88c),
	.w1(32'h3b9fb0a8),
	.w2(32'hba2ae502),
	.w3(32'hbb69fb58),
	.w4(32'hbba403a4),
	.w5(32'hbaf10ae5),
	.w6(32'hbbc80401),
	.w7(32'h3c4d9603),
	.w8(32'h3d02b578),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfda31),
	.w1(32'hbbe2a1d7),
	.w2(32'hbbbf59bf),
	.w3(32'h3c8496ad),
	.w4(32'hbb1b973a),
	.w5(32'hbb1050c1),
	.w6(32'hbbc0a684),
	.w7(32'hbb652bb0),
	.w8(32'hba1447c2),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dc0ed),
	.w1(32'hbc0b1274),
	.w2(32'hbb5e28b1),
	.w3(32'hbadc2d7c),
	.w4(32'hbbb8bcac),
	.w5(32'hbc1476d6),
	.w6(32'h38b1e5de),
	.w7(32'h391e3713),
	.w8(32'hbb65b8c4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a696448),
	.w1(32'hbc2dfea7),
	.w2(32'hba24ea59),
	.w3(32'hbb0759cf),
	.w4(32'h3bc99b8a),
	.w5(32'h3d81a92f),
	.w6(32'hbc6091f2),
	.w7(32'hbbcd475c),
	.w8(32'hbbf4a4d9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec101d),
	.w1(32'h3a92ce02),
	.w2(32'hbb0dddfe),
	.w3(32'h3cab7610),
	.w4(32'h3b80ada3),
	.w5(32'h3c6f097b),
	.w6(32'h3a69d3f7),
	.w7(32'hbbc80b42),
	.w8(32'hbc592c89),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb514617),
	.w1(32'hba45bdec),
	.w2(32'hbbb5f935),
	.w3(32'h3bd6da9c),
	.w4(32'h3c2663ed),
	.w5(32'h3c80b29a),
	.w6(32'hbc0565d1),
	.w7(32'hbb557934),
	.w8(32'hbc19d064),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb35b4),
	.w1(32'hbb36e13c),
	.w2(32'hbb09d420),
	.w3(32'h3c2fb20d),
	.w4(32'h3c7f3324),
	.w5(32'h3d69a1da),
	.w6(32'hbbb1f919),
	.w7(32'hbb57225d),
	.w8(32'hbc4e46f3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d145a),
	.w1(32'hb9f75d6b),
	.w2(32'h3b85bc5e),
	.w3(32'h3bb73c19),
	.w4(32'hbbeb380b),
	.w5(32'hbc33fb6e),
	.w6(32'hbc4f40ec),
	.w7(32'hba5f7011),
	.w8(32'h3b7cd00a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdbf1d),
	.w1(32'h3c1085bb),
	.w2(32'h3ac78466),
	.w3(32'hbb2e7b5e),
	.w4(32'h3b5e1301),
	.w5(32'h3c258f6d),
	.w6(32'h3b78078d),
	.w7(32'hbbab7a7c),
	.w8(32'hbc49d9cb),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e679c),
	.w1(32'h3ac1fc56),
	.w2(32'hbbc5d945),
	.w3(32'h3874375d),
	.w4(32'hbaf14dc9),
	.w5(32'hbbb8081f),
	.w6(32'hbbfff604),
	.w7(32'hbb5ab026),
	.w8(32'h3a3dabe1),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44c530),
	.w1(32'hbc96c409),
	.w2(32'hbc648bae),
	.w3(32'hbbc691ab),
	.w4(32'hbc2cb055),
	.w5(32'hbc44c7a2),
	.w6(32'hb9d26f41),
	.w7(32'hbb0bf084),
	.w8(32'hbc1173cd),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb368fa9),
	.w1(32'hba8ffb3e),
	.w2(32'h3bdc56b7),
	.w3(32'hbb3f7e29),
	.w4(32'hbbb5a8e7),
	.w5(32'hbc5b5190),
	.w6(32'hbb863a09),
	.w7(32'hbb0ce90a),
	.w8(32'h3c522428),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fdffa),
	.w1(32'h3b3dba30),
	.w2(32'hbbe59c5a),
	.w3(32'hbbeff90a),
	.w4(32'h3b01bcc1),
	.w5(32'h3c57131d),
	.w6(32'h3adbc7b4),
	.w7(32'hbb73fb42),
	.w8(32'hbc061366),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba643e1),
	.w1(32'hbb453b16),
	.w2(32'hbb66cab5),
	.w3(32'h3ad0e63d),
	.w4(32'hbb61a763),
	.w5(32'hbc1403ad),
	.w6(32'hbc307c4d),
	.w7(32'h3a4570cb),
	.w8(32'hbb3e910f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6103d),
	.w1(32'hbc3604e8),
	.w2(32'hbb418f7c),
	.w3(32'hbbc3dfd4),
	.w4(32'hbb2e2f3c),
	.w5(32'hba819c39),
	.w6(32'hbb18d845),
	.w7(32'hbb7e2bf9),
	.w8(32'hbb984fe7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b250f3a),
	.w1(32'hbac3c836),
	.w2(32'hbb994f31),
	.w3(32'h3a94af0c),
	.w4(32'hbbbdfa22),
	.w5(32'hbb81d22c),
	.w6(32'h3b9b8db2),
	.w7(32'hbb3d2af4),
	.w8(32'hbb15881a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab16894),
	.w1(32'hbb23ec3e),
	.w2(32'hbc15a49b),
	.w3(32'hbb736b2f),
	.w4(32'h3bb5d1d0),
	.w5(32'h3cabb4dd),
	.w6(32'hbabf477d),
	.w7(32'h3b77afb2),
	.w8(32'h3a0eedbd),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9feb793),
	.w1(32'h38f19774),
	.w2(32'hbbd3809f),
	.w3(32'h3bf56b34),
	.w4(32'h3b851ee6),
	.w5(32'h3bf774ff),
	.w6(32'h3888e9a2),
	.w7(32'hbb74037c),
	.w8(32'hbbccf8a7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e2462),
	.w1(32'hbb831832),
	.w2(32'h3b435067),
	.w3(32'h3ad56153),
	.w4(32'h3aef9de6),
	.w5(32'h3babca99),
	.w6(32'hbbe35931),
	.w7(32'h3acc90f9),
	.w8(32'hbb52e380),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe842d),
	.w1(32'hbc3dba52),
	.w2(32'hbc14c140),
	.w3(32'h3baa6079),
	.w4(32'hbbab22a1),
	.w5(32'hbc289d74),
	.w6(32'h3889688f),
	.w7(32'hbbb8106d),
	.w8(32'hbbf75c63),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff1d34),
	.w1(32'h3a8ec3ad),
	.w2(32'hbb90f230),
	.w3(32'hbbf03bd3),
	.w4(32'hbba652a5),
	.w5(32'hbb4f9680),
	.w6(32'hbb3b7375),
	.w7(32'hbb823684),
	.w8(32'hbb9ea4d7),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22781a),
	.w1(32'h3b10ac92),
	.w2(32'hb9c0233c),
	.w3(32'hba9e7b45),
	.w4(32'hb904b978),
	.w5(32'h3bf3ba5e),
	.w6(32'h3b9003f2),
	.w7(32'h3bae663f),
	.w8(32'hbb59bd39),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e2f5b),
	.w1(32'hbc79bb86),
	.w2(32'hbcbd044d),
	.w3(32'h3b737d4d),
	.w4(32'hbc8fdd4a),
	.w5(32'h3b982c2f),
	.w6(32'h3ac0316f),
	.w7(32'hbaa97eff),
	.w8(32'h3b022b57),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4adc41),
	.w1(32'h3a9dfe3e),
	.w2(32'hbc3448d3),
	.w3(32'hb9b7324d),
	.w4(32'hbb12a792),
	.w5(32'hba9b664b),
	.w6(32'hbb123a16),
	.w7(32'h3a131558),
	.w8(32'h38c6f6f0),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91f518),
	.w1(32'h3b567214),
	.w2(32'h3b458d67),
	.w3(32'h3acc927a),
	.w4(32'h3ba09529),
	.w5(32'h3b2e753c),
	.w6(32'h3bc88646),
	.w7(32'h3b3134e8),
	.w8(32'hbb897327),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d6e82),
	.w1(32'h3a4b569b),
	.w2(32'h3ab3d0c2),
	.w3(32'h39dd9cfc),
	.w4(32'hbc03e9da),
	.w5(32'hbb9fc6e2),
	.w6(32'h3b2681c4),
	.w7(32'h3b660b72),
	.w8(32'h3c3dca7b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02aaf0),
	.w1(32'hbaf7f334),
	.w2(32'hbbf17b1d),
	.w3(32'h3bd87d0f),
	.w4(32'h3929d035),
	.w5(32'h3aa60f3e),
	.w6(32'h3b8f0e01),
	.w7(32'h3a828166),
	.w8(32'hbb8b7dd1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b4ae1),
	.w1(32'h3bb2851b),
	.w2(32'h3bd5deef),
	.w3(32'h37456078),
	.w4(32'hba7541a7),
	.w5(32'hbc5459fb),
	.w6(32'hbaa1fd83),
	.w7(32'hbc07e7ae),
	.w8(32'hbae14f45),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc161202),
	.w1(32'h3b877dc5),
	.w2(32'h3b6b0acc),
	.w3(32'hbbbba385),
	.w4(32'h3ba5db15),
	.w5(32'hbb2903aa),
	.w6(32'h3b85aea0),
	.w7(32'h3ba9c60c),
	.w8(32'h3b61efb1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56e8d4),
	.w1(32'h3b066536),
	.w2(32'h3bbfab0c),
	.w3(32'hba497d48),
	.w4(32'h3b87dc26),
	.w5(32'hbb56433e),
	.w6(32'h3b8226cf),
	.w7(32'hbb6bc302),
	.w8(32'hba317c80),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66468a),
	.w1(32'h39b2308b),
	.w2(32'h3ab3913a),
	.w3(32'h3bd6d904),
	.w4(32'h390b5072),
	.w5(32'hba324cbf),
	.w6(32'hbbaa933f),
	.w7(32'hbb999897),
	.w8(32'hbb7e54e8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f9a2b),
	.w1(32'hb938fa14),
	.w2(32'hba851ad0),
	.w3(32'hbb98db45),
	.w4(32'h392fdbbf),
	.w5(32'hbb9790ce),
	.w6(32'hbb8034ea),
	.w7(32'hbc0025d5),
	.w8(32'h39c0b5ec),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba0a1b),
	.w1(32'h3bd01ffc),
	.w2(32'hba1ff660),
	.w3(32'hbb783d93),
	.w4(32'h392cae01),
	.w5(32'hbc69e98a),
	.w6(32'h3bdc2065),
	.w7(32'h3b7eb5e5),
	.w8(32'h39ea3245),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b91a6),
	.w1(32'hbb4bdd85),
	.w2(32'h3b3a5be0),
	.w3(32'h3b386c89),
	.w4(32'hbbbf0ab5),
	.w5(32'hbc4007ea),
	.w6(32'h3ab1ce69),
	.w7(32'hbc1f1a6f),
	.w8(32'hbbf9bed0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9a547),
	.w1(32'hbae714e6),
	.w2(32'hba365a87),
	.w3(32'hbc16bc8f),
	.w4(32'h3beff2c3),
	.w5(32'h3ca61e32),
	.w6(32'h3bc23e60),
	.w7(32'hbb4bfeae),
	.w8(32'hbc74f70e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56cbe6),
	.w1(32'hbb947257),
	.w2(32'hba36fd5e),
	.w3(32'h3a4ce49d),
	.w4(32'h3b7090a5),
	.w5(32'h3b7b2dd7),
	.w6(32'hbbd2da10),
	.w7(32'hbb9c8b5b),
	.w8(32'hbb079a93),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12fd1c),
	.w1(32'h3b581a61),
	.w2(32'h3b8265b2),
	.w3(32'h3b828fd5),
	.w4(32'h39a0055c),
	.w5(32'hbb2cc5a0),
	.w6(32'h3beefc05),
	.w7(32'hbb181d9f),
	.w8(32'h3babd2ad),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80103b),
	.w1(32'hbb2c669c),
	.w2(32'hba2a481f),
	.w3(32'hbb8155b5),
	.w4(32'hb9aeef25),
	.w5(32'h3c52a69e),
	.w6(32'h3b53e6bd),
	.w7(32'hb826d0d7),
	.w8(32'hbc184430),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39284a3a),
	.w1(32'hbc932770),
	.w2(32'hbc874faf),
	.w3(32'hbbc2b923),
	.w4(32'hbb6c5502),
	.w5(32'h3c572b4d),
	.w6(32'hbae20934),
	.w7(32'hbb1ac90a),
	.w8(32'hbadde387),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb910c55),
	.w1(32'h3b380578),
	.w2(32'hbba1264a),
	.w3(32'h3c07ecd3),
	.w4(32'hbb27daf3),
	.w5(32'h3c5a6806),
	.w6(32'hbb7f3d05),
	.w7(32'hbbc6d940),
	.w8(32'hbc5808ed),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule