module layer_10_featuremap_71(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59e1a8),
	.w1(32'h3aab5000),
	.w2(32'h3c009885),
	.w3(32'h3c853283),
	.w4(32'h3aa88e66),
	.w5(32'h3b54fce8),
	.w6(32'h3b0bafae),
	.w7(32'hbc4f358e),
	.w8(32'h3b9c95d9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b1f71),
	.w1(32'h3b5fbecc),
	.w2(32'hbc924e2e),
	.w3(32'h3c39d9fe),
	.w4(32'h3c1fb848),
	.w5(32'hbca7058d),
	.w6(32'hbb6a6657),
	.w7(32'h3b4c8f0a),
	.w8(32'hbc2a823c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8dca5f),
	.w1(32'hbbd3b389),
	.w2(32'hbb04b9e3),
	.w3(32'hbcd8a90b),
	.w4(32'hbbb09ca7),
	.w5(32'hbb3df4ad),
	.w6(32'hbc1aa5fb),
	.w7(32'h3c1be4ed),
	.w8(32'h3b878d67),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a228ae1),
	.w1(32'hbb91f831),
	.w2(32'h3bb97da7),
	.w3(32'h3c2d441b),
	.w4(32'h3b8c080a),
	.w5(32'h3af49649),
	.w6(32'h3c3c1f3a),
	.w7(32'h3b6d96aa),
	.w8(32'hbaa96148),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b965203),
	.w1(32'hba33e2bd),
	.w2(32'hba832d64),
	.w3(32'hb8300dde),
	.w4(32'h3a58ba02),
	.w5(32'hbba96222),
	.w6(32'h3beec03b),
	.w7(32'h3c17b8d1),
	.w8(32'hba03de49),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f0f44),
	.w1(32'hbacbfeef),
	.w2(32'hbb8a806f),
	.w3(32'hbc87db9b),
	.w4(32'hbb69e0ce),
	.w5(32'hbc4ebe70),
	.w6(32'hbc7e7aab),
	.w7(32'h3b737142),
	.w8(32'hbbe90841),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd48c65),
	.w1(32'hbac7cc94),
	.w2(32'hbba5891f),
	.w3(32'hbd11cd1c),
	.w4(32'hbbbba3ed),
	.w5(32'h3c0c4881),
	.w6(32'hbce66d3d),
	.w7(32'hbacc4850),
	.w8(32'hbbccd3d3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65fd69),
	.w1(32'hbb88de84),
	.w2(32'hbba8cd42),
	.w3(32'h3d007e71),
	.w4(32'h3c4119f4),
	.w5(32'h3b15de5f),
	.w6(32'hb9d8985a),
	.w7(32'hbc50dc05),
	.w8(32'h3c29729e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4c650),
	.w1(32'hbc2d90f8),
	.w2(32'h388e15f9),
	.w3(32'h3a7b4329),
	.w4(32'hbc069084),
	.w5(32'h3bb417fb),
	.w6(32'h3c5c9296),
	.w7(32'hbbc43750),
	.w8(32'hbb888db8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48a19b),
	.w1(32'h39874492),
	.w2(32'h3b3d3446),
	.w3(32'h3c17740d),
	.w4(32'h3bcc9b47),
	.w5(32'h3a8b8e01),
	.w6(32'hbb420678),
	.w7(32'h3b422baa),
	.w8(32'h3af611cb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b687c19),
	.w1(32'h3b6050eb),
	.w2(32'hbaa0591b),
	.w3(32'h3b95579c),
	.w4(32'h3b9db456),
	.w5(32'hbb1c7b82),
	.w6(32'h3b20b23a),
	.w7(32'h3b239cda),
	.w8(32'h3b125dd1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a2a0a3),
	.w1(32'hbb01b147),
	.w2(32'h3ba6a42e),
	.w3(32'h3b3e6f80),
	.w4(32'h3b81fbc2),
	.w5(32'h3c39e554),
	.w6(32'h3b3a9b64),
	.w7(32'hbb9e203a),
	.w8(32'h3c48ff8e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7b890),
	.w1(32'h3b5057d7),
	.w2(32'h3c142420),
	.w3(32'h3c8ad841),
	.w4(32'h3c1fb383),
	.w5(32'h3c1c5f8a),
	.w6(32'h3c76bfde),
	.w7(32'h3c235935),
	.w8(32'h3c5929d7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba55ee),
	.w1(32'hb9550e4b),
	.w2(32'hbbc0ec0e),
	.w3(32'h3ce3490f),
	.w4(32'h3c2c4d0f),
	.w5(32'h3bc65553),
	.w6(32'h3ce0480a),
	.w7(32'h3c0a1fd3),
	.w8(32'h3ad4fe8a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc004ff5),
	.w1(32'hbac14aa4),
	.w2(32'hbbdba142),
	.w3(32'h3be5ed9d),
	.w4(32'h37621d79),
	.w5(32'hbc3d6312),
	.w6(32'h3bf72441),
	.w7(32'h3ba0af7b),
	.w8(32'hbc7acaf5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b974198),
	.w1(32'h3b3b5ba3),
	.w2(32'h3bec3a22),
	.w3(32'h3b5ba9cd),
	.w4(32'h3b4c2f4d),
	.w5(32'h3bb2aca1),
	.w6(32'hbaa9e4d6),
	.w7(32'hbb83088a),
	.w8(32'h3bca1e18),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14b2ab),
	.w1(32'h3be3f028),
	.w2(32'hba114046),
	.w3(32'h3c1fab35),
	.w4(32'h3bebb8be),
	.w5(32'hba86b8f5),
	.w6(32'h3c07fb8a),
	.w7(32'h3bb2c9ee),
	.w8(32'hbb89542a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05cb8a),
	.w1(32'hbb6328db),
	.w2(32'h3b9f152a),
	.w3(32'hbb71217b),
	.w4(32'hbaa712b4),
	.w5(32'h3c0a404c),
	.w6(32'hbc0d478d),
	.w7(32'hbb6b635c),
	.w8(32'h3ba828d7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d7a14),
	.w1(32'h3bcd4c3c),
	.w2(32'hbc4090ae),
	.w3(32'h3ca0b906),
	.w4(32'h3c226474),
	.w5(32'hbbe26c84),
	.w6(32'h3c9b1898),
	.w7(32'h3bbeed5b),
	.w8(32'h3b2042b5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c8d95),
	.w1(32'h3b2f1541),
	.w2(32'hbab7de00),
	.w3(32'h3baafd37),
	.w4(32'hbb8d2029),
	.w5(32'hbbc441d8),
	.w6(32'h3bd8728d),
	.w7(32'hbb975f62),
	.w8(32'hb739e4d4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d3731),
	.w1(32'h395898ba),
	.w2(32'hbbf926eb),
	.w3(32'hbb80b4d4),
	.w4(32'h3a86a7ca),
	.w5(32'hbc12b953),
	.w6(32'hbb9a228b),
	.w7(32'h3b91547e),
	.w8(32'hb94b96ad),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef3709),
	.w1(32'h3ac89a69),
	.w2(32'hbc511b44),
	.w3(32'h38db6e6b),
	.w4(32'hbae87dea),
	.w5(32'hbc2b2cbe),
	.w6(32'h3ad74d6b),
	.w7(32'hbb52712c),
	.w8(32'hbc432494),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0186d),
	.w1(32'hbba3bbfd),
	.w2(32'hbb8d9c7e),
	.w3(32'h3bebc74f),
	.w4(32'hbb751388),
	.w5(32'hbbd45e00),
	.w6(32'hba7876bb),
	.w7(32'hba90a72e),
	.w8(32'hbba66362),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaa007),
	.w1(32'hbbda4b71),
	.w2(32'h3b72af7d),
	.w3(32'hbb6d0df4),
	.w4(32'hbc10e0f0),
	.w5(32'h3bdee3b6),
	.w6(32'hbbd51e7c),
	.w7(32'hbc1093f8),
	.w8(32'h3bd08b64),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4abd92),
	.w1(32'h3b805126),
	.w2(32'hba873cc5),
	.w3(32'h3c8cd628),
	.w4(32'h3be9d797),
	.w5(32'h3bfd0469),
	.w6(32'h3c631a48),
	.w7(32'h3a89c830),
	.w8(32'h3c37d4ac),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22f296),
	.w1(32'h3bfb3e9f),
	.w2(32'hb9b87fa5),
	.w3(32'h3c111079),
	.w4(32'h3b295459),
	.w5(32'h3b5a5681),
	.w6(32'h3b9a4e0d),
	.w7(32'h3a12fabb),
	.w8(32'h38a27a43),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c77b7f),
	.w1(32'h3b12798a),
	.w2(32'hba2ab304),
	.w3(32'h3ba5f33a),
	.w4(32'h3bc5d0db),
	.w5(32'hba03faea),
	.w6(32'hb99cec3d),
	.w7(32'h3bdb67be),
	.w8(32'hb9f8f52b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb148b3c),
	.w1(32'hba0f45bd),
	.w2(32'h3c85a798),
	.w3(32'hbb0d5995),
	.w4(32'hba716990),
	.w5(32'h3c08a545),
	.w6(32'hba9de1ff),
	.w7(32'hba98472d),
	.w8(32'h3b129e9d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ba588),
	.w1(32'hbcaab7e5),
	.w2(32'hbc7bc71f),
	.w3(32'hbc65c0ae),
	.w4(32'hbc3ef431),
	.w5(32'hbc86fd01),
	.w6(32'hbbdbdcd6),
	.w7(32'h3c4e2821),
	.w8(32'hbca40b53),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc889377),
	.w1(32'hbb2c9055),
	.w2(32'hbaa57e51),
	.w3(32'hbd0ef9ef),
	.w4(32'hbcc0ee09),
	.w5(32'hbb52673d),
	.w6(32'hbc88f37b),
	.w7(32'hbc2e2f32),
	.w8(32'hb914427a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb08ab),
	.w1(32'h3b82d74e),
	.w2(32'hbb4c92ff),
	.w3(32'hbbb6baca),
	.w4(32'hba9d7b6f),
	.w5(32'hbbadd9c5),
	.w6(32'hbb986e84),
	.w7(32'hbb1ddcc8),
	.w8(32'hbbc5299d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be08d9b),
	.w1(32'h3a3f8148),
	.w2(32'hbb9ed8c9),
	.w3(32'h3be8c5e0),
	.w4(32'h3c10fb59),
	.w5(32'hbb1f3338),
	.w6(32'h3a894e49),
	.w7(32'hbbb4b21e),
	.w8(32'hbc01fb75),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaacff),
	.w1(32'hbaa1b2c7),
	.w2(32'h3b6e2356),
	.w3(32'h3bc55f69),
	.w4(32'h3c0436b2),
	.w5(32'hba182aa5),
	.w6(32'h3b0fcec4),
	.w7(32'hba0ebd65),
	.w8(32'h3a9d0d39),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33d98f),
	.w1(32'h3b6c6d17),
	.w2(32'hbbd2194e),
	.w3(32'hba88d2a4),
	.w4(32'h3b157f1e),
	.w5(32'hbb986f74),
	.w6(32'h3b4c1662),
	.w7(32'h3c08d468),
	.w8(32'h3ae051f8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be23298),
	.w1(32'h3b02a22b),
	.w2(32'h3b8ecf3f),
	.w3(32'hbb8e1bb7),
	.w4(32'hba9c4106),
	.w5(32'h3b93c249),
	.w6(32'hbb9f4254),
	.w7(32'hbc02fff9),
	.w8(32'hbb176927),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fc39e),
	.w1(32'h3b9fd3cc),
	.w2(32'h3c5a5c4f),
	.w3(32'h3bb5ec84),
	.w4(32'h3bbee463),
	.w5(32'h3bd095a5),
	.w6(32'h3b0c2427),
	.w7(32'h3b6678e4),
	.w8(32'h3bde90ed),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0de9d),
	.w1(32'hbbf2b84c),
	.w2(32'hbbb026de),
	.w3(32'hbc41a4b9),
	.w4(32'hbc5c6f95),
	.w5(32'hbb15a7e1),
	.w6(32'hbba2232b),
	.w7(32'hbc00bcc8),
	.w8(32'h3bbd600a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4d78e),
	.w1(32'hbc3ba92d),
	.w2(32'hbc60affb),
	.w3(32'hbc1eee78),
	.w4(32'hbbb06672),
	.w5(32'hbc5024dc),
	.w6(32'h3bb454a0),
	.w7(32'h3bd6de45),
	.w8(32'hbc629078),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf660c),
	.w1(32'hbc4d834b),
	.w2(32'h3c6c1e33),
	.w3(32'hbc9c700e),
	.w4(32'hbc744add),
	.w5(32'h3ba9d696),
	.w6(32'hbc8dacce),
	.w7(32'hbbaf5e09),
	.w8(32'h3b487204),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd6276c),
	.w1(32'h3c45153c),
	.w2(32'hbb17e789),
	.w3(32'h3c306b7b),
	.w4(32'h3b5cd4a9),
	.w5(32'hbb3ea3b3),
	.w6(32'h3ab00ef3),
	.w7(32'hbbcb26a9),
	.w8(32'hb9cad1f1),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39124829),
	.w1(32'hbbcc5862),
	.w2(32'hbc020dbf),
	.w3(32'hbbb57321),
	.w4(32'hbbfe810b),
	.w5(32'hbbff7c12),
	.w6(32'hbba71dfa),
	.w7(32'hbc4eacc1),
	.w8(32'h3b6cdc75),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d7408),
	.w1(32'hbc1cca1c),
	.w2(32'hbb6bbb3f),
	.w3(32'hbcc87694),
	.w4(32'hbcabd701),
	.w5(32'h3ba21a04),
	.w6(32'hbc29d4b6),
	.w7(32'h3b9b3d05),
	.w8(32'hbc24a6fa),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a7a38),
	.w1(32'h3c3e6c97),
	.w2(32'hba002e31),
	.w3(32'h3b1fb620),
	.w4(32'h3bd14564),
	.w5(32'h38f49c1b),
	.w6(32'hbb76e1fc),
	.w7(32'hbb67425b),
	.w8(32'hbabf78ce),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf7abe),
	.w1(32'hbc01d509),
	.w2(32'hbbea2466),
	.w3(32'hba04f003),
	.w4(32'hbb74cb9e),
	.w5(32'hbc25222a),
	.w6(32'hb9a86e7d),
	.w7(32'hbb8e7d27),
	.w8(32'hbc1d1547),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbdd9a),
	.w1(32'h3c270f9e),
	.w2(32'h3995f13a),
	.w3(32'hbc36803e),
	.w4(32'h3be52e4f),
	.w5(32'h3b025941),
	.w6(32'hbb770270),
	.w7(32'h3c3223e7),
	.w8(32'h3ad3957b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0870c),
	.w1(32'h3b8e2e55),
	.w2(32'h3b77f40e),
	.w3(32'h3a2f5b99),
	.w4(32'h3bcd9f95),
	.w5(32'h3be76e2c),
	.w6(32'h3c15a02a),
	.w7(32'h3b0d3a12),
	.w8(32'hb8ffe23f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c310148),
	.w1(32'h3c9f7e5d),
	.w2(32'hbbf67b8f),
	.w3(32'h3c53b727),
	.w4(32'h3c3fe4c8),
	.w5(32'hbc7ad121),
	.w6(32'h3c0f2b8c),
	.w7(32'h3ba655f4),
	.w8(32'hbb972012),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c303c8f),
	.w1(32'h3c8c7509),
	.w2(32'h3ae6e5c5),
	.w3(32'hbc21c34e),
	.w4(32'h37bb2cf9),
	.w5(32'h3b4a9c81),
	.w6(32'hbc88dce7),
	.w7(32'hbc258a41),
	.w8(32'h3ad1afbd),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95dab27),
	.w1(32'hbb68fa88),
	.w2(32'h3c5db93d),
	.w3(32'h3b5f53b6),
	.w4(32'h3a8e3d9f),
	.w5(32'h3c874b4d),
	.w6(32'h3b5b28ea),
	.w7(32'h3a8bbe10),
	.w8(32'h3b981eda),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a83a7),
	.w1(32'h3b980a5f),
	.w2(32'h397d6ae5),
	.w3(32'h3cc06188),
	.w4(32'h3c2790f4),
	.w5(32'hbbe80930),
	.w6(32'hb9169662),
	.w7(32'hbac2cd0f),
	.w8(32'hbb0b98f5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b468f46),
	.w1(32'h3c90982a),
	.w2(32'h3b8b09bd),
	.w3(32'h3b463689),
	.w4(32'h3c24b438),
	.w5(32'h381c6808),
	.w6(32'hbab7a8b4),
	.w7(32'h3b9a488d),
	.w8(32'hbc729b9d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32e774),
	.w1(32'h3c38cbad),
	.w2(32'hbbb5a25c),
	.w3(32'h3b057a56),
	.w4(32'hbc1d6f65),
	.w5(32'h3b91d1ad),
	.w6(32'hbc82fbb6),
	.w7(32'hbc3f37ff),
	.w8(32'hbb448815),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e89fd),
	.w1(32'h3c156500),
	.w2(32'hbbba89ec),
	.w3(32'h3bab3ecb),
	.w4(32'h3c832ff7),
	.w5(32'hbbbcafb7),
	.w6(32'h3b85d3e5),
	.w7(32'h3bafaa96),
	.w8(32'hbbc8ebd2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d2f7a),
	.w1(32'h3c480953),
	.w2(32'h3bb9ad40),
	.w3(32'h3c4e97e0),
	.w4(32'h3c2bab6b),
	.w5(32'hbc799ebc),
	.w6(32'hbbe1c6f8),
	.w7(32'hbc36f91d),
	.w8(32'hbc705ec7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d40fb),
	.w1(32'hbb20b07d),
	.w2(32'hbb57dddf),
	.w3(32'hbc507713),
	.w4(32'hbbcadf93),
	.w5(32'hbc4fbe99),
	.w6(32'hbcbd7eee),
	.w7(32'hbc6fe035),
	.w8(32'hbc388f5d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c708ec9),
	.w1(32'h3ca788e0),
	.w2(32'h3c9ed5a4),
	.w3(32'hbbcb4f46),
	.w4(32'h3c4229df),
	.w5(32'h3c6076ce),
	.w6(32'hbbb51856),
	.w7(32'hbb82d637),
	.w8(32'h3c6c77cf),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4d2e0),
	.w1(32'h3b2e1b6a),
	.w2(32'h3a4f2e0d),
	.w3(32'h3c3d7642),
	.w4(32'hbad59511),
	.w5(32'hbb092c1f),
	.w6(32'h3c14cfac),
	.w7(32'h3a765729),
	.w8(32'hbbb280e1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c512b26),
	.w1(32'h39dca52c),
	.w2(32'hb864c4c0),
	.w3(32'h3b2ba3e6),
	.w4(32'hbbdd7f93),
	.w5(32'hba8a99ab),
	.w6(32'hbb586714),
	.w7(32'hbb595f71),
	.w8(32'h3c5ebb9b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5a31c),
	.w1(32'h3bb622f7),
	.w2(32'h3c109e2e),
	.w3(32'hbaa57079),
	.w4(32'h3aa8b3c5),
	.w5(32'hb7097457),
	.w6(32'h3c39194d),
	.w7(32'h3c3e16ec),
	.w8(32'h3b90e040),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89407c),
	.w1(32'h3c5f6b2c),
	.w2(32'hbc013442),
	.w3(32'hbc11d565),
	.w4(32'h3b14f545),
	.w5(32'hbbcd4f34),
	.w6(32'h3a82e49a),
	.w7(32'h3b751fdf),
	.w8(32'h3ab28b8f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0623c1),
	.w1(32'h3b8aa4c3),
	.w2(32'hbb0b652d),
	.w3(32'hbb77fb0c),
	.w4(32'hbb27d933),
	.w5(32'h3b177f19),
	.w6(32'hb8aa451a),
	.w7(32'h3a71efa1),
	.w8(32'h3a538fe9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1701f),
	.w1(32'hbbb732e0),
	.w2(32'hbbaaacfb),
	.w3(32'h3b84b240),
	.w4(32'hbbc451ca),
	.w5(32'hbbb22cee),
	.w6(32'hbb8d315c),
	.w7(32'hbbe9264b),
	.w8(32'hbc176e16),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52e3b0),
	.w1(32'hbba03942),
	.w2(32'hbbc31924),
	.w3(32'hbb83242a),
	.w4(32'hba6ca63d),
	.w5(32'hbb1a90dc),
	.w6(32'h36951425),
	.w7(32'hbb538c6e),
	.w8(32'h3bfae969),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a0698),
	.w1(32'hbc25aef5),
	.w2(32'h3c224e4e),
	.w3(32'hbc7c9d1b),
	.w4(32'hbc700450),
	.w5(32'h3bdf2440),
	.w6(32'h3ba767aa),
	.w7(32'h3b096884),
	.w8(32'h3b4c5434),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba387fb),
	.w1(32'h3b4ca09f),
	.w2(32'h3bd106db),
	.w3(32'hbb4d64fc),
	.w4(32'hbb487bda),
	.w5(32'h3c5d3edc),
	.w6(32'h3affaf67),
	.w7(32'hbbed0d2f),
	.w8(32'h3bfc2bdc),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be784f9),
	.w1(32'h3a24420c),
	.w2(32'hbb067c07),
	.w3(32'h3c63794f),
	.w4(32'h3bbc477e),
	.w5(32'h3b0a1ced),
	.w6(32'h3be8490e),
	.w7(32'h3bbc09f3),
	.w8(32'h3be1977a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fa5c0),
	.w1(32'hbc48ce3a),
	.w2(32'hb9816a35),
	.w3(32'h3a39967e),
	.w4(32'hbb07cad5),
	.w5(32'hbb504c5d),
	.w6(32'h3c12791b),
	.w7(32'h3b85a33c),
	.w8(32'hbc22f87d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30516b),
	.w1(32'h3b2ad672),
	.w2(32'hbad015f8),
	.w3(32'hbb8567b6),
	.w4(32'h3ba8d117),
	.w5(32'hbb414050),
	.w6(32'hbc86812b),
	.w7(32'h3a8747ca),
	.w8(32'hbb71d07a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b12af),
	.w1(32'h3aae0c2c),
	.w2(32'hbc154fdf),
	.w3(32'h3a26a9f0),
	.w4(32'h3bd0f03f),
	.w5(32'hbb9c186a),
	.w6(32'hba81f3c6),
	.w7(32'hbaa070d0),
	.w8(32'h3b16bb4e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8117c5),
	.w1(32'hbc86e963),
	.w2(32'h3b6f6d82),
	.w3(32'hbc4a6cb9),
	.w4(32'hbc41fc44),
	.w5(32'hba7aabaf),
	.w6(32'hbbf1123e),
	.w7(32'hbbab5fbc),
	.w8(32'h3b875527),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65b6b9),
	.w1(32'h3c76668c),
	.w2(32'h3c083cf7),
	.w3(32'hb94038da),
	.w4(32'h3c35e14f),
	.w5(32'h3c10e3b6),
	.w6(32'hbba2a009),
	.w7(32'h3a863425),
	.w8(32'h3b81be60),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3703e),
	.w1(32'h3a809dbf),
	.w2(32'h3b5709a1),
	.w3(32'h3c509e04),
	.w4(32'hbbeda9a7),
	.w5(32'h3b217d68),
	.w6(32'hbab47a36),
	.w7(32'hbbc157e4),
	.w8(32'h3a052db9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20c222),
	.w1(32'h3c98a17b),
	.w2(32'hba619c44),
	.w3(32'h3b31745b),
	.w4(32'h3b94cde8),
	.w5(32'h3afcc5ae),
	.w6(32'h3ba10d29),
	.w7(32'hbaa5ebe0),
	.w8(32'h3b3d570b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a47cd),
	.w1(32'hba6a5ae2),
	.w2(32'h3b8418de),
	.w3(32'hbbb5f0c9),
	.w4(32'hbab6eb1e),
	.w5(32'h3afe6c28),
	.w6(32'hbc06ede4),
	.w7(32'hbc026b32),
	.w8(32'hba8c650e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86a8fb1),
	.w1(32'hba8a2ea3),
	.w2(32'h3b87b444),
	.w3(32'hbb25be46),
	.w4(32'hbb149bed),
	.w5(32'hbc511ce7),
	.w6(32'hbb6a3ba1),
	.w7(32'hbb666d98),
	.w8(32'hbcccf910),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca726b4),
	.w1(32'h3caaa807),
	.w2(32'h3b67ab20),
	.w3(32'hbae4d019),
	.w4(32'h3b5dd056),
	.w5(32'h3b21a3a2),
	.w6(32'hbcec7259),
	.w7(32'hbca8139f),
	.w8(32'h3c10b005),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17b7f4),
	.w1(32'h3bf83129),
	.w2(32'h3ba15caa),
	.w3(32'h3c1fe9ef),
	.w4(32'h3c1cce7e),
	.w5(32'hbb065fbe),
	.w6(32'h3bcab91f),
	.w7(32'h3b27666a),
	.w8(32'h39868dff),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2420d6),
	.w1(32'h3bb103aa),
	.w2(32'h3a695942),
	.w3(32'hba457020),
	.w4(32'hba565e03),
	.w5(32'hbb0798cf),
	.w6(32'hba5afea4),
	.w7(32'hbc28e056),
	.w8(32'h3b8a92de),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c928c22),
	.w1(32'h3c83e60e),
	.w2(32'hbb0c59d9),
	.w3(32'h3c1f60d0),
	.w4(32'h3c042b10),
	.w5(32'h396e39ed),
	.w6(32'h3b5e7459),
	.w7(32'hbb875d9e),
	.w8(32'hba0395d7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11e81b),
	.w1(32'hbaf2662e),
	.w2(32'hbae183d9),
	.w3(32'hbb71c4ef),
	.w4(32'h3b09eb21),
	.w5(32'hbb122a25),
	.w6(32'hbc001c76),
	.w7(32'hb9f0a526),
	.w8(32'h3c25ba09),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a1d7d),
	.w1(32'h3c25f00c),
	.w2(32'h3b69458d),
	.w3(32'h3b24b883),
	.w4(32'h3b2de1f0),
	.w5(32'h3a93a27b),
	.w6(32'h3b575e3f),
	.w7(32'h3b259343),
	.w8(32'h3b8345ed),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19fab8),
	.w1(32'h39e72735),
	.w2(32'h3c023102),
	.w3(32'hbac662be),
	.w4(32'h3a85ce63),
	.w5(32'h3c262115),
	.w6(32'h3b136010),
	.w7(32'h3b98012f),
	.w8(32'h3b815ec2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81e319),
	.w1(32'hbc560c7e),
	.w2(32'hbbf1d014),
	.w3(32'h3983d70d),
	.w4(32'hbc0f89c2),
	.w5(32'hbbc7861c),
	.w6(32'hba878868),
	.w7(32'h3a8889bc),
	.w8(32'hb9895afd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbe105),
	.w1(32'h39cb905d),
	.w2(32'hbbc0e359),
	.w3(32'hbc058376),
	.w4(32'hbc1c8703),
	.w5(32'h3b93ab96),
	.w6(32'hbc4a78ca),
	.w7(32'hbc3714ec),
	.w8(32'hbb902ba0),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cdd30),
	.w1(32'h3b3ad5b0),
	.w2(32'h3ba196ac),
	.w3(32'h3c0037ac),
	.w4(32'h3bfe90dc),
	.w5(32'hbc9007ec),
	.w6(32'h3a4570c9),
	.w7(32'h3ba87087),
	.w8(32'hbc117bc9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96fd9f),
	.w1(32'h3aa8c103),
	.w2(32'h3c054f59),
	.w3(32'hbc587ada),
	.w4(32'hbc0dfb59),
	.w5(32'h3c156438),
	.w6(32'hbc7a7e32),
	.w7(32'hbb624027),
	.w8(32'h3b7a84a8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27cf90),
	.w1(32'hb89d7b63),
	.w2(32'hbab6f427),
	.w3(32'h3b9ee414),
	.w4(32'hbb887c61),
	.w5(32'hbb73e58b),
	.w6(32'h3aba63d7),
	.w7(32'hbb73a198),
	.w8(32'hbbdae1a4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adee0db),
	.w1(32'h3a1f40a0),
	.w2(32'h3bd3cdd6),
	.w3(32'hbb991ac2),
	.w4(32'hbb5223c1),
	.w5(32'hb7d57057),
	.w6(32'hbbc1d07a),
	.w7(32'hbc097232),
	.w8(32'hba13be8c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c869754),
	.w1(32'h3bd907aa),
	.w2(32'hbb497a5b),
	.w3(32'h3c1fb0ef),
	.w4(32'h3c74b1e6),
	.w5(32'hbc05cdec),
	.w6(32'h3b5deffc),
	.w7(32'h3c16d35a),
	.w8(32'hbc4954f8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a8206),
	.w1(32'h3c22adf8),
	.w2(32'hbb1e6d26),
	.w3(32'h3c2da13f),
	.w4(32'h3c4717ce),
	.w5(32'h3c4b1c18),
	.w6(32'hbc32df5c),
	.w7(32'hbbaccd4c),
	.w8(32'h3c7d3bee),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94fec5),
	.w1(32'h3aa5cac3),
	.w2(32'h3a488cb2),
	.w3(32'h3d0dff77),
	.w4(32'h3cd484cd),
	.w5(32'h3c877965),
	.w6(32'h3cd50f1e),
	.w7(32'h3c57acd8),
	.w8(32'h3cc95886),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc603810),
	.w1(32'hbc7dfd7f),
	.w2(32'hbb8ed8c1),
	.w3(32'h3c062dcb),
	.w4(32'h3afe45a9),
	.w5(32'hbbabe852),
	.w6(32'h3cf62cda),
	.w7(32'h3cb7d56e),
	.w8(32'hbc0f7d33),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b6694),
	.w1(32'hbbfc96ed),
	.w2(32'h3b8b9186),
	.w3(32'hbc1bfde0),
	.w4(32'hbc45a3e8),
	.w5(32'h3b014701),
	.w6(32'hbc698725),
	.w7(32'hbc8d4693),
	.w8(32'hbab6584d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40b1c1),
	.w1(32'h3c153e37),
	.w2(32'h3aded73f),
	.w3(32'h3b5bf057),
	.w4(32'h3b616245),
	.w5(32'hbb3e83be),
	.w6(32'hbb33850b),
	.w7(32'hbbb97f3b),
	.w8(32'hbafcdff7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d8c1f),
	.w1(32'h3a38dc8f),
	.w2(32'hbc38b8ff),
	.w3(32'h3b7e96a7),
	.w4(32'h3b9bfa45),
	.w5(32'hbbc9c21b),
	.w6(32'hbb4dc62f),
	.w7(32'hbbc697eb),
	.w8(32'hbc4650ea),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c1032),
	.w1(32'hbc2343e1),
	.w2(32'h3c4a382e),
	.w3(32'hbcb13aae),
	.w4(32'hbc9972dc),
	.w5(32'h3b63def3),
	.w6(32'hbc6bc3ec),
	.w7(32'hbb98d1e9),
	.w8(32'hbb8bdb61),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a6a9f),
	.w1(32'h3bbef52e),
	.w2(32'hbb9a5916),
	.w3(32'h3b684026),
	.w4(32'hbb9ba360),
	.w5(32'hbbdc78bf),
	.w6(32'hbc3adefd),
	.w7(32'hbc44a3f6),
	.w8(32'hbc20ab24),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b668406),
	.w1(32'h3c3c7eea),
	.w2(32'hbaee61e6),
	.w3(32'hbb430a19),
	.w4(32'h3bd2609c),
	.w5(32'hbb38fa59),
	.w6(32'hbba43938),
	.w7(32'h3b22cb48),
	.w8(32'hbbe22603),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8daed),
	.w1(32'h3c2a5694),
	.w2(32'hbcb0fcae),
	.w3(32'h3c039ea7),
	.w4(32'h3c12b1e2),
	.w5(32'hbc5314ba),
	.w6(32'hbbd3b8b9),
	.w7(32'h392366f8),
	.w8(32'h3aad2716),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce706b),
	.w1(32'hbbb0bfbb),
	.w2(32'hb90cbbab),
	.w3(32'hbc6ed722),
	.w4(32'hbbf5d3e8),
	.w5(32'hbc0ec2b3),
	.w6(32'hbb062a7c),
	.w7(32'hbc499a1c),
	.w8(32'hbb9916c5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c2dcb),
	.w1(32'h3ae80940),
	.w2(32'hbb3d6f47),
	.w3(32'hbc5b9275),
	.w4(32'hbbf11f1a),
	.w5(32'hbc015c7d),
	.w6(32'hbc1d0278),
	.w7(32'hbc48e475),
	.w8(32'hbc181863),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77e14e),
	.w1(32'h3a6deb7d),
	.w2(32'hb8849b09),
	.w3(32'hbc55aca1),
	.w4(32'hbbaa8349),
	.w5(32'h3acd549d),
	.w6(32'hbc957a5f),
	.w7(32'hbc2f63e3),
	.w8(32'h3bdf9f00),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf72928),
	.w1(32'hbb064510),
	.w2(32'hbc0c9545),
	.w3(32'h3b6fc29a),
	.w4(32'h3beb98e5),
	.w5(32'hbc0e32b8),
	.w6(32'h3c04885b),
	.w7(32'h3ba90616),
	.w8(32'hbad324fe),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c541774),
	.w1(32'h3c74f0a0),
	.w2(32'h3c1c3208),
	.w3(32'h3c6216bb),
	.w4(32'h3c75475a),
	.w5(32'h3b8290c7),
	.w6(32'h3ba8fde7),
	.w7(32'hbb41631a),
	.w8(32'hbbb36e0d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac1580),
	.w1(32'hba4d6c47),
	.w2(32'h3bf9002a),
	.w3(32'h3bd06009),
	.w4(32'hba14c628),
	.w5(32'h3b29411f),
	.w6(32'h3bb290db),
	.w7(32'hbb3bd0c7),
	.w8(32'hbb032b8f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cec0d),
	.w1(32'hbb30e98a),
	.w2(32'h3c74b345),
	.w3(32'h3b6feb9e),
	.w4(32'hbb7a5568),
	.w5(32'h3bf195d8),
	.w6(32'hbbce4d15),
	.w7(32'hbc02fd0d),
	.w8(32'hbb5cb386),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c917bd8),
	.w1(32'h3a46e658),
	.w2(32'hbc394024),
	.w3(32'h3bc4ebee),
	.w4(32'hbb33f7c7),
	.w5(32'hbc40768e),
	.w6(32'hbc395979),
	.w7(32'hbb5cbdd8),
	.w8(32'hbbed4c40),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93b338),
	.w1(32'hbb9bed33),
	.w2(32'h38b9dd46),
	.w3(32'hbc8cc37f),
	.w4(32'hbc5093c6),
	.w5(32'h3c0a259d),
	.w6(32'hbc82514a),
	.w7(32'hbc1e743d),
	.w8(32'h3c092433),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67c80d),
	.w1(32'h3c783ed4),
	.w2(32'h3ab94e6b),
	.w3(32'h3ba0f83f),
	.w4(32'h3bf504a6),
	.w5(32'hbb2c3ee8),
	.w6(32'h3ba7d8da),
	.w7(32'h3c07a783),
	.w8(32'hbb0ae3d0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba11967),
	.w1(32'h3a73b1c5),
	.w2(32'hbbbedfa7),
	.w3(32'h3b5ae43e),
	.w4(32'h3bb3ee77),
	.w5(32'hbb5f3611),
	.w6(32'hbb3ef012),
	.w7(32'hbbf6d368),
	.w8(32'h3b3efe5b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb602d5),
	.w1(32'h3c0a59f4),
	.w2(32'hbb3de86c),
	.w3(32'h3c1f66a3),
	.w4(32'h3bbfc396),
	.w5(32'hbb624f34),
	.w6(32'h39fd3359),
	.w7(32'h3a45862a),
	.w8(32'h3be648ba),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b177f46),
	.w1(32'h3ba2ed99),
	.w2(32'hbb97b760),
	.w3(32'h3b53a3a4),
	.w4(32'h3b9b1063),
	.w5(32'hbafebd7b),
	.w6(32'h3bd828d3),
	.w7(32'hba9b2b0f),
	.w8(32'h3b1b79ad),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf70b9b),
	.w1(32'h3c7402e0),
	.w2(32'hbba0f6d9),
	.w3(32'hbb315096),
	.w4(32'h3bc77622),
	.w5(32'hbc01fead),
	.w6(32'hbba40bb2),
	.w7(32'hbbdd27c9),
	.w8(32'hbc1b12c3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0a8ad),
	.w1(32'h3c273956),
	.w2(32'h3c0bba9f),
	.w3(32'h3c28aa24),
	.w4(32'h3b7218eb),
	.w5(32'h3bf512b8),
	.w6(32'hba311c1e),
	.w7(32'hbb06c5fe),
	.w8(32'h3b84de7c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a5969),
	.w1(32'h3c283d01),
	.w2(32'hbc8d8205),
	.w3(32'hbbb2406e),
	.w4(32'hbae057df),
	.w5(32'hbc81fe65),
	.w6(32'h39d39dab),
	.w7(32'h3ab8bf9c),
	.w8(32'h3b624800),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf990a6),
	.w1(32'hbc98dd60),
	.w2(32'hbc304277),
	.w3(32'hbd044747),
	.w4(32'hbcaeb3e5),
	.w5(32'hbc21cad0),
	.w6(32'hbb90a264),
	.w7(32'hba1400ae),
	.w8(32'hbc7a879b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39272425),
	.w1(32'hbbe779b9),
	.w2(32'hbc35effc),
	.w3(32'h3b91f49b),
	.w4(32'hbb597383),
	.w5(32'hbc6c1499),
	.w6(32'hbc47f80b),
	.w7(32'hbc82dca7),
	.w8(32'hbb040c83),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc992fdd),
	.w1(32'hbc2b062d),
	.w2(32'hbc0648a1),
	.w3(32'hbce7f6f9),
	.w4(32'hbc9cd879),
	.w5(32'hbc30b0c5),
	.w6(32'hbc2ec54b),
	.w7(32'hbbceae63),
	.w8(32'hbc25a7a7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0202b),
	.w1(32'h3b9ea2df),
	.w2(32'h3ba577e9),
	.w3(32'hbbec2969),
	.w4(32'hba89ff25),
	.w5(32'h39ef106c),
	.w6(32'hbc3a8ba0),
	.w7(32'hbb9a6071),
	.w8(32'hbb6c008c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c64e9),
	.w1(32'h3b5fae05),
	.w2(32'hbba17f1d),
	.w3(32'hbb66e147),
	.w4(32'hbbf489e8),
	.w5(32'hbb871a6e),
	.w6(32'hbc060f59),
	.w7(32'hbbde1200),
	.w8(32'hbba30eec),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab9c9d),
	.w1(32'h3a435bec),
	.w2(32'hbaef446c),
	.w3(32'h3a76cf26),
	.w4(32'h3b3fea6e),
	.w5(32'hb8b27e2a),
	.w6(32'h399a5750),
	.w7(32'hbb9fddda),
	.w8(32'hbb0d74d3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a1fa1),
	.w1(32'hbb2d9022),
	.w2(32'h3956fc95),
	.w3(32'hbb1f329b),
	.w4(32'hbacd7cbb),
	.w5(32'hbb9841f1),
	.w6(32'h39710cbc),
	.w7(32'hba33351b),
	.w8(32'hbbdbc96a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f8bb5),
	.w1(32'h3c305317),
	.w2(32'h3b9f7bf1),
	.w3(32'hbb3e024a),
	.w4(32'h3a93265e),
	.w5(32'h3ac58d31),
	.w6(32'hbc109146),
	.w7(32'hbba2057d),
	.w8(32'hbb920195),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c485564),
	.w1(32'hb9d412eb),
	.w2(32'h3b3de11c),
	.w3(32'h3b32260f),
	.w4(32'hbb5cb53a),
	.w5(32'hbb117a5f),
	.w6(32'hbbac1de1),
	.w7(32'hbbc6c721),
	.w8(32'h3aa88e02),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc86809),
	.w1(32'hbc224416),
	.w2(32'h3b553762),
	.w3(32'hbc5e48e8),
	.w4(32'hbc55da31),
	.w5(32'h3b55017d),
	.w6(32'hbbc223f4),
	.w7(32'hbadca46d),
	.w8(32'h374e8432),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80484a),
	.w1(32'h3c440459),
	.w2(32'h3ba53013),
	.w3(32'h3c0023e3),
	.w4(32'h3bef0bbf),
	.w5(32'h3aaf85e6),
	.w6(32'h3b274fcd),
	.w7(32'h3ab80640),
	.w8(32'hbb91a2fd),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2fe1f),
	.w1(32'h3b7dd5fa),
	.w2(32'hba54368c),
	.w3(32'hbb93fbfc),
	.w4(32'hbb263303),
	.w5(32'hbb711fd4),
	.w6(32'hbbcb421a),
	.w7(32'h3a21bc33),
	.w8(32'hbc093d9b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf6e24),
	.w1(32'h3bfd0a36),
	.w2(32'h3ca09154),
	.w3(32'hbad2f248),
	.w4(32'h3bdc2715),
	.w5(32'h3b619e69),
	.w6(32'hbc1af8c4),
	.w7(32'h3ad54fb8),
	.w8(32'hbbe533ae),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1bd5fa),
	.w1(32'h3c90ce29),
	.w2(32'h3c224500),
	.w3(32'h3ae3b523),
	.w4(32'hbb46389e),
	.w5(32'h3c331a38),
	.w6(32'hbc785081),
	.w7(32'hbc7b548f),
	.w8(32'h3bbf1b29),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88c128),
	.w1(32'h3bceb84e),
	.w2(32'hbc19e20e),
	.w3(32'h3caa3398),
	.w4(32'h3bb6e21f),
	.w5(32'hbc39ce19),
	.w6(32'h3c1e75f8),
	.w7(32'hba72296f),
	.w8(32'hbbfe9cea),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94cf53),
	.w1(32'hbc5f926c),
	.w2(32'h3a4dcc65),
	.w3(32'hbcd43191),
	.w4(32'hbcba761d),
	.w5(32'h3bfde964),
	.w6(32'hbce3348b),
	.w7(32'hbc9a2e24),
	.w8(32'h3a99ef03),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51c59e),
	.w1(32'h3b83a010),
	.w2(32'h3946ff8a),
	.w3(32'h3c205636),
	.w4(32'h3c158df0),
	.w5(32'hbb3c6c23),
	.w6(32'h3bc0a2e2),
	.w7(32'h3b9bc5b5),
	.w8(32'hbbf755b2),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2984a6),
	.w1(32'hbc0488f5),
	.w2(32'h3c3c9c48),
	.w3(32'hba2c3c91),
	.w4(32'hbb3401e6),
	.w5(32'h3bd37be7),
	.w6(32'hbb9fed98),
	.w7(32'hbb0f2931),
	.w8(32'h3c26e62c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb912e3),
	.w1(32'h3c1fc174),
	.w2(32'h38d55d1b),
	.w3(32'hbb87ab31),
	.w4(32'h3bb2265f),
	.w5(32'hb8f1045b),
	.w6(32'hba414e4f),
	.w7(32'h3c4a4b39),
	.w8(32'hbb7b41fe),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896a8a8),
	.w1(32'hb97c4a71),
	.w2(32'hbc38d962),
	.w3(32'hbb19d8e1),
	.w4(32'hba6a3c50),
	.w5(32'hbc9f3b5c),
	.w6(32'hbbb008cf),
	.w7(32'hbbe0ce7f),
	.w8(32'hbc7cd083),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ed060),
	.w1(32'hbb83896b),
	.w2(32'h3a5c8839),
	.w3(32'hbcd36cc4),
	.w4(32'hbc62475d),
	.w5(32'h3c350396),
	.w6(32'hbcb8e22d),
	.w7(32'hbc155985),
	.w8(32'h3b2f828c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4e719),
	.w1(32'h3b0dc05f),
	.w2(32'h3c3d4569),
	.w3(32'h3c899f05),
	.w4(32'h3b5d3431),
	.w5(32'h3c46c526),
	.w6(32'h3b69c820),
	.w7(32'hbb7e91b7),
	.w8(32'h3bf78927),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb835c8ee),
	.w1(32'hbb86c64d),
	.w2(32'h39039623),
	.w3(32'h3bd9cd5b),
	.w4(32'h3b0a7c3f),
	.w5(32'hba8d9797),
	.w6(32'h3c2aa68a),
	.w7(32'h3bba9c76),
	.w8(32'h3a821714),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11ec40),
	.w1(32'h3b8aac7f),
	.w2(32'h3c06cd7d),
	.w3(32'hbaae8481),
	.w4(32'h3a3b25a1),
	.w5(32'h3b9d72f6),
	.w6(32'hb96c051b),
	.w7(32'h3a362d68),
	.w8(32'hbb0b743c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1644da),
	.w1(32'h3c3d1521),
	.w2(32'h3bd07271),
	.w3(32'h3c3fe8bd),
	.w4(32'h3c285042),
	.w5(32'hba7b613b),
	.w6(32'h3bb60c0a),
	.w7(32'h399df6b8),
	.w8(32'hbbed5672),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6356ee),
	.w1(32'h3c610a88),
	.w2(32'hbbfd8905),
	.w3(32'h3af03736),
	.w4(32'h3b720fd0),
	.w5(32'h3936e9c9),
	.w6(32'hbbff185b),
	.w7(32'hbbabfbe5),
	.w8(32'h3b4d6710),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f7094),
	.w1(32'h39e7154f),
	.w2(32'hbc302766),
	.w3(32'hba06447a),
	.w4(32'h3a8fda52),
	.w5(32'hbc4cd8b8),
	.w6(32'h3a867560),
	.w7(32'h3bb0682b),
	.w8(32'hbc549d48),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73850d),
	.w1(32'hbabd1fad),
	.w2(32'hbc01e2c1),
	.w3(32'hbccfb800),
	.w4(32'hbcf01888),
	.w5(32'hbbe7e6e7),
	.w6(32'hbcd1a1a8),
	.w7(32'hbc6a5d64),
	.w8(32'h3befc173),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc507e0c),
	.w1(32'hbafc1d19),
	.w2(32'h3a989e51),
	.w3(32'hbc8e415a),
	.w4(32'hbb8493bb),
	.w5(32'hba5929c0),
	.w6(32'hbb4c66df),
	.w7(32'h3b9c47b7),
	.w8(32'h3a1ea331),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a2762),
	.w1(32'h3b2f4f81),
	.w2(32'hbb918c53),
	.w3(32'hba3629bc),
	.w4(32'hbae025ee),
	.w5(32'hbb8777d3),
	.w6(32'hbb0b6a1a),
	.w7(32'hbb1257e1),
	.w8(32'h3ac45423),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdc327),
	.w1(32'h3b5739ca),
	.w2(32'hbb0a3392),
	.w3(32'h3ba94579),
	.w4(32'h3c4bc6de),
	.w5(32'hbb45d083),
	.w6(32'h3b8039bc),
	.w7(32'h3c17dce0),
	.w8(32'hbb99767b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ff089),
	.w1(32'hbb54891e),
	.w2(32'hbc845554),
	.w3(32'hba28d6eb),
	.w4(32'h3ab91e41),
	.w5(32'hbc995933),
	.w6(32'hbb15168a),
	.w7(32'hbb53c8c1),
	.w8(32'hbca72e62),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fc405),
	.w1(32'hbaf989f7),
	.w2(32'hbb094a5e),
	.w3(32'hbc8fbe78),
	.w4(32'hbc5cdc97),
	.w5(32'hbbf2d957),
	.w6(32'hbc990062),
	.w7(32'hbc552e79),
	.w8(32'h3b1bd99d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2efe36),
	.w1(32'h3c11dfb8),
	.w2(32'hbb17788e),
	.w3(32'h3b0ffea1),
	.w4(32'h3bd70184),
	.w5(32'hbbce0a97),
	.w6(32'h3b8acfc3),
	.w7(32'h3b0384ca),
	.w8(32'hbc495cfa),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b374a42),
	.w1(32'h3c31ed3c),
	.w2(32'hbc638964),
	.w3(32'hbb7bb1d9),
	.w4(32'hbb881c24),
	.w5(32'hbc44932f),
	.w6(32'h3bda6d12),
	.w7(32'hbb23baf0),
	.w8(32'hbc370402),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb735fda),
	.w1(32'h3b444460),
	.w2(32'h39c17526),
	.w3(32'hbc82503b),
	.w4(32'hbc41b219),
	.w5(32'hbb45ce7f),
	.w6(32'hbc87c60f),
	.w7(32'hbbb42f78),
	.w8(32'hbb81d9b2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefc48a),
	.w1(32'h3b732403),
	.w2(32'h3b191934),
	.w3(32'hbbba46a4),
	.w4(32'hbb63b8ce),
	.w5(32'h3ba7926a),
	.w6(32'hbc04edef),
	.w7(32'hbb8cea09),
	.w8(32'h3b838751),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89b1e3),
	.w1(32'h39a34104),
	.w2(32'hbc3ec0e9),
	.w3(32'hba7f2ef8),
	.w4(32'h3b4dd983),
	.w5(32'hbc71fa85),
	.w6(32'h3b0e1f3b),
	.w7(32'h3b5e5c13),
	.w8(32'hbc2e1893),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9777f5),
	.w1(32'hbade4a77),
	.w2(32'hbb9ff259),
	.w3(32'hbc9a1a73),
	.w4(32'h39822781),
	.w5(32'hba3e0e08),
	.w6(32'hbb96d814),
	.w7(32'hbc2abc81),
	.w8(32'h3bc7b3f1),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfa061),
	.w1(32'h3c0e2768),
	.w2(32'hba86012f),
	.w3(32'h3bfefa8e),
	.w4(32'h3c808d3f),
	.w5(32'hb9b08218),
	.w6(32'h3c06fd9a),
	.w7(32'hbb1f5bec),
	.w8(32'hba1d9922),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c1a61),
	.w1(32'hba7c26c2),
	.w2(32'h3b87c554),
	.w3(32'h3afa4f69),
	.w4(32'h37b32210),
	.w5(32'h3b5c803b),
	.w6(32'h3a98e8fe),
	.w7(32'hb9aa3f2c),
	.w8(32'h3b70866d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb0fa8),
	.w1(32'h3be20cd2),
	.w2(32'h3b923c6d),
	.w3(32'h3ba6ed35),
	.w4(32'h3ba4ed08),
	.w5(32'h3bc5e918),
	.w6(32'h3bbd21d4),
	.w7(32'h3b8f70bc),
	.w8(32'h3b9568fc),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dce8f),
	.w1(32'h3b9d2999),
	.w2(32'h3b21f52e),
	.w3(32'h3abca7d8),
	.w4(32'hbabc8148),
	.w5(32'h3c28b85f),
	.w6(32'h3a0a117c),
	.w7(32'hbabe82b5),
	.w8(32'h3b948caf),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15d4ce),
	.w1(32'h3bb95a89),
	.w2(32'h3b9a63fc),
	.w3(32'h3caf50ce),
	.w4(32'h3c7be6be),
	.w5(32'h3b06568e),
	.w6(32'h3c6d34c0),
	.w7(32'h3c162bba),
	.w8(32'h3bec2972),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b844481),
	.w1(32'h3b4677e5),
	.w2(32'hb8fc9e2a),
	.w3(32'h3a9612c3),
	.w4(32'h3a98f920),
	.w5(32'hba7b3bef),
	.w6(32'h3bc45ee8),
	.w7(32'h3bc1bef1),
	.w8(32'h3bc10ef8),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacedcc8),
	.w1(32'hbab314d0),
	.w2(32'h3b70d402),
	.w3(32'hbae88a6f),
	.w4(32'hba9cbf8d),
	.w5(32'h3c8163f2),
	.w6(32'h3b4fd6a6),
	.w7(32'h3b0484a5),
	.w8(32'h3c050020),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c571413),
	.w1(32'h3bdfbab3),
	.w2(32'h3a3704c8),
	.w3(32'h3cf096da),
	.w4(32'h3ca4669b),
	.w5(32'h3aae4b92),
	.w6(32'h3ca6ea20),
	.w7(32'h3c3aa948),
	.w8(32'h3b2116a5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c28b5),
	.w1(32'h3b180c66),
	.w2(32'hbba69d33),
	.w3(32'h3ba12c91),
	.w4(32'h3b326cd9),
	.w5(32'hbc26984b),
	.w6(32'h3b39f96c),
	.w7(32'h3b9828a1),
	.w8(32'hbbe360c1),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a9898),
	.w1(32'hbbe08608),
	.w2(32'h3a7c446c),
	.w3(32'hbc90aac2),
	.w4(32'hbc5ee214),
	.w5(32'hbac7f7a5),
	.w6(32'hbc62241a),
	.w7(32'hbc2ac95b),
	.w8(32'hbb4162f3),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fee63),
	.w1(32'h3b4e9e88),
	.w2(32'hbbdf0e21),
	.w3(32'hbb0cc760),
	.w4(32'hbb0b70b7),
	.w5(32'h3af7ab13),
	.w6(32'hbb51db90),
	.w7(32'hbb8349d7),
	.w8(32'hbb9dec9c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add9d9c),
	.w1(32'hbb9e99e9),
	.w2(32'h3bb2a010),
	.w3(32'h3c58c332),
	.w4(32'h3b3d56da),
	.w5(32'h3bd3a3c1),
	.w6(32'h3b9284d5),
	.w7(32'hbb9f48fc),
	.w8(32'hb8ecf5fd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95b5be),
	.w1(32'h3b9d03d8),
	.w2(32'h3b955170),
	.w3(32'h3bb85425),
	.w4(32'h3bed71b4),
	.w5(32'h3b0a0c39),
	.w6(32'hba883dfe),
	.w7(32'hbb0b76dd),
	.w8(32'h3bb8ddd4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc950d7),
	.w1(32'hb9bfc5db),
	.w2(32'h3b641805),
	.w3(32'h3b9caa6a),
	.w4(32'hbb630259),
	.w5(32'h3b26a630),
	.w6(32'h3ba341b4),
	.w7(32'hbb9a83fd),
	.w8(32'h3939bda9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67bc68),
	.w1(32'h3b7ab74e),
	.w2(32'h3b27e827),
	.w3(32'h3a3b760d),
	.w4(32'h3b2a213d),
	.w5(32'h39e932f0),
	.w6(32'hba3d9d0c),
	.w7(32'hba5846c5),
	.w8(32'h386a473d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b139bf9),
	.w1(32'h3aabe452),
	.w2(32'h3aeca9cb),
	.w3(32'h3aba0357),
	.w4(32'hba981cd9),
	.w5(32'hbb48637f),
	.w6(32'h3aaa282a),
	.w7(32'hba8329c0),
	.w8(32'hbadf2044),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fdcf79),
	.w1(32'h3ad95f8f),
	.w2(32'h3b7cbe4e),
	.w3(32'hb96e5c2d),
	.w4(32'hbbc201e6),
	.w5(32'hbb891738),
	.w6(32'hbb17171d),
	.w7(32'hbb1a576c),
	.w8(32'h3b674be3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a6548),
	.w1(32'h3b9028ac),
	.w2(32'h3b94161e),
	.w3(32'hbc3f600a),
	.w4(32'hbb83da72),
	.w5(32'h3b3af3b7),
	.w6(32'hbb630bcc),
	.w7(32'h3b5a6016),
	.w8(32'h3b177c02),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a954441),
	.w1(32'h3aa01d8c),
	.w2(32'h3be2e95f),
	.w3(32'h3b509b9f),
	.w4(32'hb792dbb1),
	.w5(32'h3b2cf4b5),
	.w6(32'h3b416486),
	.w7(32'h3b0cbeff),
	.w8(32'h3b9682a2),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29d48d),
	.w1(32'h3be0453a),
	.w2(32'hba909164),
	.w3(32'hba7e2bb2),
	.w4(32'h3860487f),
	.w5(32'hbbaaba32),
	.w6(32'h3a055b6b),
	.w7(32'h3a050f4c),
	.w8(32'hbb68e865),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f7c5a),
	.w1(32'hbb1eb137),
	.w2(32'h3add523e),
	.w3(32'hba84db6f),
	.w4(32'hbb96a8f0),
	.w5(32'hbaa07154),
	.w6(32'hbb37d74f),
	.w7(32'hba040fe4),
	.w8(32'h3b81acf4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fa868),
	.w1(32'h3c08d771),
	.w2(32'h3aa127ef),
	.w3(32'h3a2b21db),
	.w4(32'h3bd5a3ea),
	.w5(32'hbc2984c1),
	.w6(32'h3b8e76ef),
	.w7(32'h3bc03aa7),
	.w8(32'hbb48b292),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01c2fe),
	.w1(32'hbb733d48),
	.w2(32'h3bab39f2),
	.w3(32'hbcbea305),
	.w4(32'hbc8eb3e7),
	.w5(32'h3b7481fd),
	.w6(32'hbc7f4d51),
	.w7(32'hbc245ba0),
	.w8(32'h3b3a188d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8ef75),
	.w1(32'h3b22b798),
	.w2(32'h39e1114e),
	.w3(32'h3bcced49),
	.w4(32'h3c0c07f4),
	.w5(32'h39a44b93),
	.w6(32'h3b84846f),
	.w7(32'h3b1e861d),
	.w8(32'hbaddda4f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaadcbb),
	.w1(32'h39123fa9),
	.w2(32'h3bf03792),
	.w3(32'hba59769e),
	.w4(32'hbaa61bf5),
	.w5(32'h3b8c4f99),
	.w6(32'hba824f82),
	.w7(32'hbab1a624),
	.w8(32'h3b19c6cb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0cec0),
	.w1(32'h3b739356),
	.w2(32'h3b208d57),
	.w3(32'h3a5f830f),
	.w4(32'h39059ae3),
	.w5(32'h37a76b85),
	.w6(32'hba410f11),
	.w7(32'h3a4e1534),
	.w8(32'hba8298e7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f7620),
	.w1(32'h3b8d7cce),
	.w2(32'h3b977156),
	.w3(32'hbb2b89a6),
	.w4(32'hbb7138ca),
	.w5(32'h3ba5c713),
	.w6(32'hba83d6d0),
	.w7(32'hbafef9f4),
	.w8(32'h3bc88647),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba74772),
	.w1(32'h3b88e59e),
	.w2(32'h3bd35a6b),
	.w3(32'h3b9365c3),
	.w4(32'h3b6e24ef),
	.w5(32'h3babb4cc),
	.w6(32'h3be34e70),
	.w7(32'h3bc54ed0),
	.w8(32'h39a21995),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cd0af),
	.w1(32'h3be6c32d),
	.w2(32'h3b4fbd05),
	.w3(32'h3ba73cd1),
	.w4(32'h3b0b11aa),
	.w5(32'hb9fd9bfc),
	.w6(32'h3b4c48f5),
	.w7(32'hba0af9c3),
	.w8(32'h3bc39533),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b420d2f),
	.w1(32'h3bb4b3d4),
	.w2(32'hbade5298),
	.w3(32'h3a37880a),
	.w4(32'h3ab35456),
	.w5(32'hb9a32839),
	.w6(32'h3b7a8abe),
	.w7(32'h3c1667ea),
	.w8(32'h3b316c62),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc159acf),
	.w1(32'hbc0b1150),
	.w2(32'h3b96c298),
	.w3(32'hbbf78777),
	.w4(32'hbc01c9c4),
	.w5(32'h3b66b98e),
	.w6(32'hbb865dee),
	.w7(32'hbbb10b35),
	.w8(32'h3b0a05ff),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d21a8),
	.w1(32'h3b70d69d),
	.w2(32'h3836e4f3),
	.w3(32'h3a8096b2),
	.w4(32'h3b00c9e1),
	.w5(32'h3ac1eb4f),
	.w6(32'h3abda68f),
	.w7(32'h3b4620be),
	.w8(32'h3aa9d9a1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e8471),
	.w1(32'h3b1e3f13),
	.w2(32'h3b6890a3),
	.w3(32'h3baa9b3e),
	.w4(32'h3b4e5c10),
	.w5(32'h3a934e6a),
	.w6(32'h3b67475e),
	.w7(32'h3a9c75c4),
	.w8(32'h3a28397f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1cccf),
	.w1(32'h3bc343b4),
	.w2(32'hbafcc5b7),
	.w3(32'h3b5eade3),
	.w4(32'h3bb85b17),
	.w5(32'hbb42dd76),
	.w6(32'h3b778c2c),
	.w7(32'h3bb2a188),
	.w8(32'hbb5ebf42),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b7b6e),
	.w1(32'h3b1b3b0b),
	.w2(32'h3b7078b8),
	.w3(32'hba29761e),
	.w4(32'h3a2c29f2),
	.w5(32'h39afa083),
	.w6(32'hbaa51391),
	.w7(32'hba10ba77),
	.w8(32'h3b3b9fda),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82d135),
	.w1(32'h3b776d82),
	.w2(32'h38598d84),
	.w3(32'h3be0ea31),
	.w4(32'h3bb2d9ba),
	.w5(32'h3af18992),
	.w6(32'h3b3588fe),
	.w7(32'h3ba9df1f),
	.w8(32'hbb018b18),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6cee9),
	.w1(32'h3aec3591),
	.w2(32'h3b06db80),
	.w3(32'h3b00fb15),
	.w4(32'h3a92239d),
	.w5(32'hbac9c49a),
	.w6(32'hba482bcf),
	.w7(32'h3b0d5a19),
	.w8(32'hba98c07a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cff9e3),
	.w1(32'hba47c10d),
	.w2(32'hbb784c16),
	.w3(32'hbba24b32),
	.w4(32'hbb6f4d42),
	.w5(32'hb9e45e71),
	.w6(32'hba8b6969),
	.w7(32'hba2e52ee),
	.w8(32'hb9dd6579),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb515444),
	.w1(32'hbb32192b),
	.w2(32'h3b1f436d),
	.w3(32'hba0ae656),
	.w4(32'h3af08db9),
	.w5(32'h3b096c4b),
	.w6(32'h3adf5ed6),
	.w7(32'hb918c6f6),
	.w8(32'h3ae93377),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe32d7),
	.w1(32'h3b09d295),
	.w2(32'h3ad385a9),
	.w3(32'h3b05fb69),
	.w4(32'h3aa78be7),
	.w5(32'h3b9d429b),
	.w6(32'h3a9cce96),
	.w7(32'h3ac19535),
	.w8(32'h3b9c8f8d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beefd2a),
	.w1(32'h3bf17fab),
	.w2(32'h3a0ce957),
	.w3(32'h3c58a6ac),
	.w4(32'h3c4c24dd),
	.w5(32'hbac8e394),
	.w6(32'h3c3d29d4),
	.w7(32'h3c3cec7c),
	.w8(32'hbabf8ddc),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfc0c2),
	.w1(32'hb8d5c34c),
	.w2(32'hba1b1cb0),
	.w3(32'hbad55a4e),
	.w4(32'hba81a446),
	.w5(32'h3bb507a8),
	.w6(32'hbaffc1ad),
	.w7(32'hbabe2106),
	.w8(32'h3b34a0f4),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7aa3a),
	.w1(32'hb9ce3259),
	.w2(32'h3bb42312),
	.w3(32'h3b0cbdd2),
	.w4(32'h3ae6bae1),
	.w5(32'h3b9bb40b),
	.w6(32'hb98b93c8),
	.w7(32'hbae9ca2f),
	.w8(32'h3b87ac47),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6b56c),
	.w1(32'h3bcf776f),
	.w2(32'h3a876801),
	.w3(32'h3b9a68a5),
	.w4(32'h3bbcfa91),
	.w5(32'hba3bfc5c),
	.w6(32'h3b8c3ad6),
	.w7(32'h3bb5684a),
	.w8(32'hb9f9c9ca),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bf3a9),
	.w1(32'h3b2b5dae),
	.w2(32'h3af3b367),
	.w3(32'h3b8c6762),
	.w4(32'h3ae2f7de),
	.w5(32'hb8eeb6e0),
	.w6(32'h3ab32047),
	.w7(32'h3998abf9),
	.w8(32'h3aca74ab),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a020d04),
	.w1(32'h3a9eb70a),
	.w2(32'h3a7071c2),
	.w3(32'h3ac8c6ff),
	.w4(32'h3b18f992),
	.w5(32'h3a80c4a0),
	.w6(32'h3a6f3e1b),
	.w7(32'h3aba8f56),
	.w8(32'h3a70a920),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b024b27),
	.w1(32'h39b0d612),
	.w2(32'hbab000ed),
	.w3(32'h3b675108),
	.w4(32'h3b82c97b),
	.w5(32'hba3ade2d),
	.w6(32'h3b0af114),
	.w7(32'h3b069702),
	.w8(32'hb9a4b433),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e605c),
	.w1(32'hbbd61496),
	.w2(32'hbc85a904),
	.w3(32'hbb732769),
	.w4(32'hbb591d75),
	.w5(32'hbcccc8f7),
	.w6(32'hbb90a352),
	.w7(32'hbbae8a33),
	.w8(32'hbc9efd61),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd1c67d),
	.w1(32'hbcaa74f6),
	.w2(32'h3b33fbf3),
	.w3(32'hbd178d2c),
	.w4(32'hbcff2e73),
	.w5(32'h3b8932a5),
	.w6(32'hbcfb4591),
	.w7(32'hbcd1d124),
	.w8(32'h3bae4e59),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2028ae),
	.w1(32'h3aa317b1),
	.w2(32'hbb6d697a),
	.w3(32'h3a4356ba),
	.w4(32'h3b29f69f),
	.w5(32'h3adc8309),
	.w6(32'h3b1dc218),
	.w7(32'h3b0fc048),
	.w8(32'h3b29eb65),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb443f37),
	.w1(32'hba6145d5),
	.w2(32'hb9f05d05),
	.w3(32'hbb4f0638),
	.w4(32'h37a3f6c4),
	.w5(32'hb891e3c9),
	.w6(32'hb9d7f628),
	.w7(32'h3b0db459),
	.w8(32'h3a88b244),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fc115),
	.w1(32'hbb03361b),
	.w2(32'hbb44f60f),
	.w3(32'hbb81db37),
	.w4(32'hba2b23f9),
	.w5(32'hbadfa1b3),
	.w6(32'h39e4abf9),
	.w7(32'h3ab523ec),
	.w8(32'hbb641c6b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf476d),
	.w1(32'hbb8b3cc6),
	.w2(32'h3a447cd8),
	.w3(32'hba78c257),
	.w4(32'hbbb80d5b),
	.w5(32'h3a291537),
	.w6(32'hbb10c8e0),
	.w7(32'hbbccbf59),
	.w8(32'h3a956f40),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c252f),
	.w1(32'h3a93451e),
	.w2(32'hb9b7ae1b),
	.w3(32'hb9273154),
	.w4(32'h3ac2b282),
	.w5(32'hb9f44559),
	.w6(32'h3a21d42c),
	.w7(32'h3b1ea8b2),
	.w8(32'hba46808b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0307b9),
	.w1(32'hba193f95),
	.w2(32'hbbca2f07),
	.w3(32'h3b1641e7),
	.w4(32'hb98caab1),
	.w5(32'hb82f3869),
	.w6(32'h3b0400d5),
	.w7(32'hbb050446),
	.w8(32'hbb10aa4b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9619c53),
	.w1(32'hbb6730a2),
	.w2(32'h3ad10716),
	.w3(32'h3c297b8f),
	.w4(32'h3ba25026),
	.w5(32'h3aca7d7c),
	.w6(32'h3bbb02bc),
	.w7(32'h3af104c6),
	.w8(32'hba8c63df),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49b831),
	.w1(32'h3b34f3d2),
	.w2(32'hba984faa),
	.w3(32'hbad5b898),
	.w4(32'h3b8c5378),
	.w5(32'hbb2c9183),
	.w6(32'hbb8d48b9),
	.w7(32'hb9193399),
	.w8(32'hbb5ff211),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba84988),
	.w1(32'h3b749d1a),
	.w2(32'hbb4769db),
	.w3(32'hb99eec0d),
	.w4(32'h3b462396),
	.w5(32'hb83d844d),
	.w6(32'h3a9c4d07),
	.w7(32'hbb7660cb),
	.w8(32'hb9f13f92),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1d853),
	.w1(32'hb990a813),
	.w2(32'h3b8c062b),
	.w3(32'h3a560fe6),
	.w4(32'hba12cb1e),
	.w5(32'h3ae5a809),
	.w6(32'hb92a376f),
	.w7(32'h3aa25a55),
	.w8(32'hb9c27440),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afaeb40),
	.w1(32'h3a25a5b4),
	.w2(32'h3b3f59bf),
	.w3(32'h3b1d0a1d),
	.w4(32'h37fd8dee),
	.w5(32'h3b7f26a2),
	.w6(32'h3ab15f67),
	.w7(32'hbb0728f0),
	.w8(32'h3b76bf55),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16c771),
	.w1(32'h391bc2fe),
	.w2(32'hbb503e9e),
	.w3(32'h3b638500),
	.w4(32'h39ef65c1),
	.w5(32'hbb707640),
	.w6(32'h3b54e9e2),
	.w7(32'h3a5a186b),
	.w8(32'hbb82c58c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8955a1),
	.w1(32'hbb426e36),
	.w2(32'hbae0004a),
	.w3(32'hbba5446c),
	.w4(32'hbb856de0),
	.w5(32'h39019966),
	.w6(32'hbba1e8f5),
	.w7(32'hbb87b97a),
	.w8(32'h3a06ceea),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ff5ea),
	.w1(32'hb9984fa4),
	.w2(32'h3a9e8d6e),
	.w3(32'hbb9e034d),
	.w4(32'hba0881a2),
	.w5(32'h3b920ce6),
	.w6(32'hbb8a0b62),
	.w7(32'hbb7e1e46),
	.w8(32'h3b4444ac),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83235f),
	.w1(32'h3b1a0194),
	.w2(32'hbb798d33),
	.w3(32'h3ba812a3),
	.w4(32'h3b84dd5e),
	.w5(32'hbb4d84ac),
	.w6(32'h3a7500f1),
	.w7(32'h3a5fe980),
	.w8(32'hba6cf484),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3511a),
	.w1(32'h3a41e96f),
	.w2(32'h3c06e586),
	.w3(32'hbac3a125),
	.w4(32'hba3d4a3c),
	.w5(32'h3bfe8120),
	.w6(32'hba39455d),
	.w7(32'h3a3af577),
	.w8(32'h3ba15120),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ae415),
	.w1(32'h3c4d99bc),
	.w2(32'h3b0c46c4),
	.w3(32'h3c5547d3),
	.w4(32'h3c422ef4),
	.w5(32'h3b288ded),
	.w6(32'h3c1b197d),
	.w7(32'h3c2175cf),
	.w8(32'h3a97030e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b192398),
	.w1(32'h3b1ed10a),
	.w2(32'hbbacbc23),
	.w3(32'h3b2f413b),
	.w4(32'h3b3d2308),
	.w5(32'hbbe6d66e),
	.w6(32'h3adcf7af),
	.w7(32'h3ad5f57e),
	.w8(32'hbba80353),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba302eb),
	.w1(32'hbb006b65),
	.w2(32'h3b6d2fe1),
	.w3(32'hbbd5c132),
	.w4(32'hbb458f00),
	.w5(32'h3b803612),
	.w6(32'hbb8ab398),
	.w7(32'hba97828c),
	.w8(32'h3b42a429),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90b113),
	.w1(32'h3b25e968),
	.w2(32'h39c996df),
	.w3(32'h3ad6e33b),
	.w4(32'h3a46137c),
	.w5(32'h3b24977a),
	.w6(32'h3b431bf4),
	.w7(32'h3abea772),
	.w8(32'h3b965486),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac5ea6),
	.w1(32'hbac37947),
	.w2(32'h3bef988c),
	.w3(32'hbb9d1670),
	.w4(32'h39a3f35e),
	.w5(32'h3bbf3424),
	.w6(32'h3908119a),
	.w7(32'h3b23f5d9),
	.w8(32'h3b95cc37),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86778b),
	.w1(32'h3b8ce14e),
	.w2(32'hbb7f1eaa),
	.w3(32'h3ba1a801),
	.w4(32'h3b75c350),
	.w5(32'hbb8f3635),
	.w6(32'h3a774d94),
	.w7(32'h3a835517),
	.w8(32'hbbac98d9),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3255b8),
	.w1(32'hbbe6ef03),
	.w2(32'h3aa6d8dc),
	.w3(32'hbb637b13),
	.w4(32'hbba77815),
	.w5(32'h3a707ad7),
	.w6(32'hbbb27d08),
	.w7(32'hbab08092),
	.w8(32'h3adf50cc),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b268a25),
	.w1(32'h3aaa3487),
	.w2(32'hbbb195fd),
	.w3(32'hb7437246),
	.w4(32'h3b71970e),
	.w5(32'hbb8493b8),
	.w6(32'hb95dfb4f),
	.w7(32'h3b066bae),
	.w8(32'hbb2d5c2f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a1886),
	.w1(32'h3ad171f9),
	.w2(32'hb7043002),
	.w3(32'hbb1a2b7d),
	.w4(32'h39963c8b),
	.w5(32'h3ae69234),
	.w6(32'hba96d1a9),
	.w7(32'h3b1d90db),
	.w8(32'h3acaac83),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a17cee),
	.w1(32'hbb0beb33),
	.w2(32'hba9da94b),
	.w3(32'h3b29f1c5),
	.w4(32'h3b41bb71),
	.w5(32'h3b13c64a),
	.w6(32'h3b562099),
	.w7(32'h3aa52d52),
	.w8(32'h3b580e6e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d4e9f),
	.w1(32'hb9ea46f2),
	.w2(32'h3a8bb204),
	.w3(32'h395d5574),
	.w4(32'h3aaeaee4),
	.w5(32'h3ada28db),
	.w6(32'hba8b5043),
	.w7(32'h3a936b44),
	.w8(32'h3aa50e57),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5d0c3),
	.w1(32'hb90998f2),
	.w2(32'hb9d7f02c),
	.w3(32'h3a755591),
	.w4(32'hba13f4a5),
	.w5(32'hbaca9999),
	.w6(32'h3b6949ca),
	.w7(32'hba395a5c),
	.w8(32'hbb314a2d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac805de),
	.w1(32'h3a8cab0e),
	.w2(32'hbaab9998),
	.w3(32'hbabbe01d),
	.w4(32'hbaea0490),
	.w5(32'hba8e59e9),
	.w6(32'hb9d28adc),
	.w7(32'hbaef1322),
	.w8(32'hbb173057),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89e496),
	.w1(32'hbb48913b),
	.w2(32'h3ac82a9f),
	.w3(32'hbbd88bdb),
	.w4(32'hbbef0946),
	.w5(32'h3b6a8de1),
	.w6(32'hbbe42fc2),
	.w7(32'hbbcc9827),
	.w8(32'h3ab333da),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ce7b0),
	.w1(32'h3a82a668),
	.w2(32'h3ab34c15),
	.w3(32'h3b005d21),
	.w4(32'h3b30e81f),
	.w5(32'h3aef182f),
	.w6(32'h3b42b088),
	.w7(32'h3a6b8b70),
	.w8(32'h3abed1fe),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fd6d0),
	.w1(32'h3a31c7b3),
	.w2(32'hbacac478),
	.w3(32'h39dfda55),
	.w4(32'h3a994640),
	.w5(32'hbaf39314),
	.w6(32'h3a96dff3),
	.w7(32'h399803e3),
	.w8(32'h3b4eca42),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f5ea3),
	.w1(32'hb80a7c1e),
	.w2(32'hbb199f24),
	.w3(32'hba8811c0),
	.w4(32'h396e4dea),
	.w5(32'hba2a1dbb),
	.w6(32'h3b86a714),
	.w7(32'h3b602b63),
	.w8(32'hbaba17b8),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb019113),
	.w1(32'hb91efe49),
	.w2(32'h3ba5f602),
	.w3(32'h3904eec7),
	.w4(32'hba862851),
	.w5(32'h3b6964af),
	.w6(32'hba2e09e4),
	.w7(32'h3b08793a),
	.w8(32'h3bd1d0be),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f80d2),
	.w1(32'h3ba930f7),
	.w2(32'h3a8754ec),
	.w3(32'h3bd8dcf8),
	.w4(32'h3b9a93d9),
	.w5(32'hb9af53e4),
	.w6(32'h3bb1677e),
	.w7(32'h3bc1c97b),
	.w8(32'hbb3d5625),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1457b6),
	.w1(32'h3995fd43),
	.w2(32'hba7cae87),
	.w3(32'hbb8a2c63),
	.w4(32'hbb09f2d3),
	.w5(32'hb79bb093),
	.w6(32'hbba3f424),
	.w7(32'hbb2dfc8a),
	.w8(32'h3a94c40e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8327e8),
	.w1(32'hbab13c6a),
	.w2(32'hba926093),
	.w3(32'h3b40287a),
	.w4(32'hbb0b62f2),
	.w5(32'hba7035b0),
	.w6(32'h3b639d30),
	.w7(32'hba16af08),
	.w8(32'h3b78f2f3),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9511af),
	.w1(32'h3b07c737),
	.w2(32'h3ba0de54),
	.w3(32'h3af3f812),
	.w4(32'h3bad9bce),
	.w5(32'h3b74f884),
	.w6(32'h3bb188d0),
	.w7(32'h3c0df84a),
	.w8(32'h3b2de9d1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae42ca4),
	.w1(32'h3b19f5d7),
	.w2(32'h3a08d0b3),
	.w3(32'h3b1a9081),
	.w4(32'h3b37c547),
	.w5(32'hbb94bddf),
	.w6(32'h3ac9542a),
	.w7(32'hbaa001fe),
	.w8(32'h3a381c18),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39899c4e),
	.w1(32'hbb056f35),
	.w2(32'hbb2c1116),
	.w3(32'hbbd3ce7e),
	.w4(32'hbb9b5f54),
	.w5(32'hbb1c9166),
	.w6(32'h3ab9e475),
	.w7(32'h3990508f),
	.w8(32'hbaa30215),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5886d2),
	.w1(32'hbaa4c708),
	.w2(32'h39d53178),
	.w3(32'hbb455ada),
	.w4(32'hba7b7685),
	.w5(32'h3b60d70c),
	.w6(32'hbaae318f),
	.w7(32'hb92fddb4),
	.w8(32'h3b3239e9),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b120eb7),
	.w1(32'h3b332083),
	.w2(32'h3b234f3a),
	.w3(32'h3b86f708),
	.w4(32'h3b2f8db6),
	.w5(32'h3ab37371),
	.w6(32'h3ba52a20),
	.w7(32'h3b17c24a),
	.w8(32'h39137acb),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c6ce2),
	.w1(32'h3b0f991f),
	.w2(32'h3b005574),
	.w3(32'h3a8b4249),
	.w4(32'h3aa3f51a),
	.w5(32'h3bc0226b),
	.w6(32'h39c21610),
	.w7(32'hb74905b2),
	.w8(32'h3b8b07a6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19f18d),
	.w1(32'h3b51e5c4),
	.w2(32'hbb98d658),
	.w3(32'h3bcd60ac),
	.w4(32'h3c1329de),
	.w5(32'hbaa7fa10),
	.w6(32'h3b444450),
	.w7(32'h3b5b7ff1),
	.w8(32'hb937bb91),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6897e2),
	.w1(32'hb9c66ebf),
	.w2(32'h3968c416),
	.w3(32'hbb11c3d6),
	.w4(32'hba2baf6a),
	.w5(32'h3abb431b),
	.w6(32'h3ab52299),
	.w7(32'h3964bac8),
	.w8(32'h3b1df955),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b18b2),
	.w1(32'hbab2ea3b),
	.w2(32'hbb8dd9fc),
	.w3(32'h3b1a44f7),
	.w4(32'h3ad1d9ad),
	.w5(32'hbb974c92),
	.w6(32'h3b5d87cf),
	.w7(32'h3b50fb53),
	.w8(32'hbbb9b7e4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b82aa),
	.w1(32'hbbaf2942),
	.w2(32'hbbae5d7f),
	.w3(32'hbb6815cc),
	.w4(32'hbbb62ace),
	.w5(32'hbb19afe1),
	.w6(32'hbbc98abe),
	.w7(32'hbbfbf244),
	.w8(32'hbb9c427e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb134ca7),
	.w1(32'hbb8c5392),
	.w2(32'hbb6f5158),
	.w3(32'h3ab41888),
	.w4(32'hba69c94b),
	.w5(32'hbb2b89ed),
	.w6(32'hba92df63),
	.w7(32'hbb79905e),
	.w8(32'hbb365bc4),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f8ff9),
	.w1(32'hbb4a0e61),
	.w2(32'h3accb344),
	.w3(32'hbaa00031),
	.w4(32'hbb82698c),
	.w5(32'h3ad520fb),
	.w6(32'hbad2547f),
	.w7(32'hbbf28b17),
	.w8(32'h3b1c4b0f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2577e9),
	.w1(32'h3a0f0561),
	.w2(32'hbb26d8a4),
	.w3(32'h39862ae5),
	.w4(32'h38b08f31),
	.w5(32'hba864eff),
	.w6(32'h3aa91656),
	.w7(32'h3a5ea6e5),
	.w8(32'hba386314),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6e649),
	.w1(32'h3a24cb8c),
	.w2(32'hb9ab9235),
	.w3(32'h3af91746),
	.w4(32'h3b5af6c2),
	.w5(32'h3a0bf7ea),
	.w6(32'h397ae3a1),
	.w7(32'h3b2b8e94),
	.w8(32'h3b42f28f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f35a9),
	.w1(32'h3a32be53),
	.w2(32'hbb50b2e1),
	.w3(32'hbb2fc8ec),
	.w4(32'h3b7f2123),
	.w5(32'hbb474c39),
	.w6(32'hba70d893),
	.w7(32'h39c1a386),
	.w8(32'hbb37c969),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59d3d5),
	.w1(32'hba8abec4),
	.w2(32'h3b7e0a6e),
	.w3(32'hbbaf320f),
	.w4(32'hbb886dfd),
	.w5(32'h3b347161),
	.w6(32'hbb9df819),
	.w7(32'hbafbcc99),
	.w8(32'h3bcabdea),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule