module layer_10_featuremap_114(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93446b4),
	.w1(32'hb939d394),
	.w2(32'h38616f30),
	.w3(32'hb9426d4c),
	.w4(32'h38b38ffb),
	.w5(32'h39f84248),
	.w6(32'hb9904784),
	.w7(32'h39425ba5),
	.w8(32'h394df4fe),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbbcac),
	.w1(32'h38f25f41),
	.w2(32'hb8e67f91),
	.w3(32'h3862e3ad),
	.w4(32'h3908381e),
	.w5(32'hb92a08be),
	.w6(32'h39fdaa01),
	.w7(32'h398bc97a),
	.w8(32'hb9179ac8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d113c),
	.w1(32'hba4300d0),
	.w2(32'hba287edd),
	.w3(32'hb9c90041),
	.w4(32'hb9f2e7aa),
	.w5(32'hba13e569),
	.w6(32'hba259360),
	.w7(32'hba2a1d4d),
	.w8(32'hba17a75f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b065e),
	.w1(32'hba3e4a0c),
	.w2(32'hba3d5f66),
	.w3(32'hba02e975),
	.w4(32'hb9e056fe),
	.w5(32'hb99c6db8),
	.w6(32'h3816809d),
	.w7(32'hb866f754),
	.w8(32'hb8a55f02),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2818d),
	.w1(32'h39ea8cd8),
	.w2(32'h388a03f7),
	.w3(32'hb8a040da),
	.w4(32'h3a32a9a9),
	.w5(32'hb82c36e0),
	.w6(32'h3a43c2c9),
	.w7(32'hb9d3b940),
	.w8(32'h39d2fbc1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b0b60),
	.w1(32'hb9d3d199),
	.w2(32'hb987f201),
	.w3(32'h380a552a),
	.w4(32'hb9fb9a86),
	.w5(32'hba08d162),
	.w6(32'hb96eff2d),
	.w7(32'hb9e8dd8e),
	.w8(32'hb9535416),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f4ff4d),
	.w1(32'h39170f77),
	.w2(32'hb75c8728),
	.w3(32'hb9d09f48),
	.w4(32'h399c07c9),
	.w5(32'hb7341363),
	.w6(32'hb82d499e),
	.w7(32'hb9089373),
	.w8(32'hb99e65ed),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a153111),
	.w1(32'h37c8650f),
	.w2(32'hb9895cd0),
	.w3(32'h39fd78f9),
	.w4(32'h39841a65),
	.w5(32'h38d75fb8),
	.w6(32'hb7eee521),
	.w7(32'hb9aebe9f),
	.w8(32'hb99f969f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38901a6c),
	.w1(32'hb9684acf),
	.w2(32'hb9f9f09b),
	.w3(32'h38c552d1),
	.w4(32'hb7ea9fbc),
	.w5(32'hb9ca5678),
	.w6(32'hb91ebcbd),
	.w7(32'hb9cd23d3),
	.w8(32'hb97be194),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7e80e),
	.w1(32'h3ac6b1fa),
	.w2(32'hb9dc5491),
	.w3(32'h3af4fcf1),
	.w4(32'h3af6d732),
	.w5(32'h38f8c094),
	.w6(32'h3b1473ee),
	.w7(32'h3a86b322),
	.w8(32'hb9265778),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a357cc),
	.w1(32'hb9031874),
	.w2(32'hb88819ce),
	.w3(32'h39a54897),
	.w4(32'hb91005d6),
	.w5(32'hb716a6ce),
	.w6(32'h394701e5),
	.w7(32'h39352d79),
	.w8(32'h390814a6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967bb77),
	.w1(32'hb96bde68),
	.w2(32'h392b8675),
	.w3(32'hba59eaa4),
	.w4(32'hba944a8d),
	.w5(32'hb9a3a055),
	.w6(32'hb9edfec9),
	.w7(32'h37aae3bc),
	.w8(32'h3941463d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a52ad),
	.w1(32'h393d38e8),
	.w2(32'hba2c19fd),
	.w3(32'h3acb3d52),
	.w4(32'h3a616222),
	.w5(32'hb9fd4758),
	.w6(32'h3a1aafc2),
	.w7(32'h39b2842b),
	.w8(32'hba5698bc),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea7472),
	.w1(32'hb848d43a),
	.w2(32'hba46feb8),
	.w3(32'h39d9c1d0),
	.w4(32'h38f07839),
	.w5(32'hba3fe6ef),
	.w6(32'h3a330c55),
	.w7(32'hb9a66880),
	.w8(32'hba3a4e76),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e1433),
	.w1(32'hba80760d),
	.w2(32'hbaba9a6c),
	.w3(32'h3a345925),
	.w4(32'hb968bb75),
	.w5(32'hbabebbb3),
	.w6(32'h3a7bb6ab),
	.w7(32'h3a585c72),
	.w8(32'h39a59848),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a286009),
	.w1(32'h391c9151),
	.w2(32'hba701e9b),
	.w3(32'h39d7cb45),
	.w4(32'h3a31f6db),
	.w5(32'hb991b593),
	.w6(32'h3ac76911),
	.w7(32'h3a429fcd),
	.w8(32'h3822bb87),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9081e37),
	.w1(32'h39c2dd5d),
	.w2(32'h39ae2d1e),
	.w3(32'h392f0da8),
	.w4(32'h39d53138),
	.w5(32'hb97cb85d),
	.w6(32'h39f0dfc3),
	.w7(32'h3982b391),
	.w8(32'h3997101d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00c1ad),
	.w1(32'h3acfbb1e),
	.w2(32'h3a0498a5),
	.w3(32'h3a8a3adc),
	.w4(32'h3a829158),
	.w5(32'hb8648c0f),
	.w6(32'h3a33a0f8),
	.w7(32'hb958e6c1),
	.w8(32'hba7c6905),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a873c30),
	.w1(32'h39c95301),
	.w2(32'hba37d8ff),
	.w3(32'h3aa28f4b),
	.w4(32'h3a25343c),
	.w5(32'hb9a8caa9),
	.w6(32'h3a40b20f),
	.w7(32'h386a93ef),
	.w8(32'hb9a39594),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc4ce4),
	.w1(32'h3754948e),
	.w2(32'h3817cd3f),
	.w3(32'hb9cf2a1d),
	.w4(32'h3802446f),
	.w5(32'hb8ca20c7),
	.w6(32'hb80b36ec),
	.w7(32'hb91c22f6),
	.w8(32'hb6848709),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d2ec34),
	.w1(32'hba107d2a),
	.w2(32'hb9f1f9af),
	.w3(32'hb7a3cf67),
	.w4(32'hba1ac697),
	.w5(32'hba0dccd4),
	.w6(32'hb9c0244c),
	.w7(32'hb9bea983),
	.w8(32'h37dcf804),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38adfdef),
	.w1(32'hb96a7143),
	.w2(32'hb9c82868),
	.w3(32'hb91a182d),
	.w4(32'h3a39862f),
	.w5(32'h3a0f52a5),
	.w6(32'hb8b07339),
	.w7(32'h399b05cf),
	.w8(32'hb9be7a0a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd620b),
	.w1(32'h39de69a5),
	.w2(32'hba2d2a68),
	.w3(32'h3ae1323d),
	.w4(32'h3a00e01f),
	.w5(32'hbaa1c302),
	.w6(32'h3b063f17),
	.w7(32'h3ae25de2),
	.w8(32'h397e7d79),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac96c65),
	.w1(32'h386fe77e),
	.w2(32'hba9a0fe0),
	.w3(32'h3accbd5e),
	.w4(32'h39b6f7e6),
	.w5(32'hba550536),
	.w6(32'h3acc45f0),
	.w7(32'h3a213c61),
	.w8(32'hb96798aa),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a105ccc),
	.w1(32'hb990a890),
	.w2(32'hb9f99c5a),
	.w3(32'h3a0986aa),
	.w4(32'hb702a4dd),
	.w5(32'hb993c8a2),
	.w6(32'h3ab2c56c),
	.w7(32'h3a2685a6),
	.w8(32'h39bd7e25),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a2581),
	.w1(32'hb9682144),
	.w2(32'hb9c9be0d),
	.w3(32'h37d533a0),
	.w4(32'hb8e9e433),
	.w5(32'hb969ea53),
	.w6(32'h39388dd2),
	.w7(32'h39b253a4),
	.w8(32'hb7defa71),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc643a),
	.w1(32'h385f18fb),
	.w2(32'h39413a80),
	.w3(32'hb940d6b3),
	.w4(32'h38b3e25f),
	.w5(32'h390c94d7),
	.w6(32'hb7804b34),
	.w7(32'h390753a8),
	.w8(32'h3899b3fc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883b975),
	.w1(32'hba8f66f3),
	.w2(32'hb9f553bb),
	.w3(32'h3904f302),
	.w4(32'hba07aad4),
	.w5(32'hb9ee4eaa),
	.w6(32'hba3ce9aa),
	.w7(32'hba218464),
	.w8(32'hba0fd12a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1a649),
	.w1(32'hba0c8254),
	.w2(32'hba2e3f98),
	.w3(32'h3784ed0c),
	.w4(32'hba002aba),
	.w5(32'hbaaa4724),
	.w6(32'hb830ec1c),
	.w7(32'hba34f931),
	.w8(32'hb94af38a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a801c2d),
	.w1(32'hb8c8b547),
	.w2(32'hba8433b3),
	.w3(32'h3ab4d1e0),
	.w4(32'h39620218),
	.w5(32'hba499ed3),
	.w6(32'h3ab83ceb),
	.w7(32'h39d077ba),
	.w8(32'h388f5fbe),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab2c76),
	.w1(32'hb976fb6a),
	.w2(32'hb7a83003),
	.w3(32'h395bc796),
	.w4(32'hb97a75ae),
	.w5(32'hb8c6213a),
	.w6(32'hb8ca0b93),
	.w7(32'hb88447eb),
	.w8(32'h38cb8e45),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ea497),
	.w1(32'hb905a1ca),
	.w2(32'h38905db1),
	.w3(32'h393ee804),
	.w4(32'hb918729b),
	.w5(32'hb87b2e1e),
	.w6(32'hb9639774),
	.w7(32'hb8a943ad),
	.w8(32'hb8de6c52),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0820c6),
	.w1(32'h3a40c0fe),
	.w2(32'h39e741ab),
	.w3(32'h3a1d01e8),
	.w4(32'h3a330430),
	.w5(32'hb8bc1890),
	.w6(32'h3a623e4c),
	.w7(32'h39222f3d),
	.w8(32'h39b9a11b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a9f8c),
	.w1(32'hb9826df3),
	.w2(32'h3abf6f22),
	.w3(32'hb76bc7d5),
	.w4(32'hba474529),
	.w5(32'h3a8395e1),
	.w6(32'hba088130),
	.w7(32'h3a455e0f),
	.w8(32'hb9860a05),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996ca0f),
	.w1(32'hb94bcac0),
	.w2(32'h37d4fcad),
	.w3(32'hb96814d4),
	.w4(32'hb82b2b55),
	.w5(32'hb7cf7f59),
	.w6(32'hb8822b4b),
	.w7(32'hb953641f),
	.w8(32'hb992def4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0718bf),
	.w1(32'h3922e288),
	.w2(32'h39eccbe3),
	.w3(32'hb9c1d6d0),
	.w4(32'h372da807),
	.w5(32'h39222113),
	.w6(32'h38439a74),
	.w7(32'h394971d0),
	.w8(32'h391c67e5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a986605),
	.w1(32'h3a799262),
	.w2(32'hb8291c4e),
	.w3(32'h3abc154c),
	.w4(32'h3a98c218),
	.w5(32'hb90e2d48),
	.w6(32'h3aa68a0f),
	.w7(32'h3a6f428e),
	.w8(32'h3960a9b7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a01746),
	.w1(32'h39ff8eb3),
	.w2(32'h3a47baef),
	.w3(32'hbae2efad),
	.w4(32'hb9fc911b),
	.w5(32'h36f0560c),
	.w6(32'hba0abd41),
	.w7(32'hb8f84ce9),
	.w8(32'hb84f16ae),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cf598),
	.w1(32'hba90bfce),
	.w2(32'hb95e60ac),
	.w3(32'hba61c971),
	.w4(32'hba85c12a),
	.w5(32'hba639477),
	.w6(32'h39834f90),
	.w7(32'h3a310eb3),
	.w8(32'h398b770e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9209d2b),
	.w1(32'hb9473c55),
	.w2(32'hb95a8de8),
	.w3(32'hb931ed53),
	.w4(32'hb915c749),
	.w5(32'hb925d45e),
	.w6(32'h37de8637),
	.w7(32'hb9607adc),
	.w8(32'hb93993e0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb910c390),
	.w1(32'hb79ac240),
	.w2(32'hb886b29b),
	.w3(32'hb9a12351),
	.w4(32'hb7e965b3),
	.w5(32'hb90f654e),
	.w6(32'hb916214b),
	.w7(32'hb80fc3c9),
	.w8(32'h398ab863),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38191dac),
	.w1(32'hba00470e),
	.w2(32'hb8f0104f),
	.w3(32'hb7b1f73e),
	.w4(32'hb9fc04f5),
	.w5(32'hb919f2a7),
	.w6(32'hb9d4135c),
	.w7(32'hb98a5d36),
	.w8(32'hb98fe40b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8250d9a),
	.w1(32'hb8929111),
	.w2(32'hb9982fd7),
	.w3(32'h38ff8029),
	.w4(32'hb8f0bc3a),
	.w5(32'hb9aaf742),
	.w6(32'hb8841ab2),
	.w7(32'h3798a4d5),
	.w8(32'hb99da1ac),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33a216),
	.w1(32'h3aead78f),
	.w2(32'hb93fbd40),
	.w3(32'h3b0b1193),
	.w4(32'h3b1d5924),
	.w5(32'h397d4c8d),
	.w6(32'h3b85b7db),
	.w7(32'h3aecdc5e),
	.w8(32'hb9bdfceb),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2ce72),
	.w1(32'h39c1db41),
	.w2(32'hba963388),
	.w3(32'h3aed3012),
	.w4(32'h3a9e7179),
	.w5(32'hb997fdf8),
	.w6(32'h3aee4498),
	.w7(32'h3a1fa309),
	.w8(32'hb9c25dc3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a910c27),
	.w1(32'hb85e5b63),
	.w2(32'hba990f71),
	.w3(32'h3ac2927d),
	.w4(32'h39c0640f),
	.w5(32'hba37d79e),
	.w6(32'h3aade482),
	.w7(32'h39ae0618),
	.w8(32'hba4f57d5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26d352),
	.w1(32'hb9d34e01),
	.w2(32'hbad8f9a0),
	.w3(32'h3a91f4e0),
	.w4(32'hb99cae20),
	.w5(32'hba340e94),
	.w6(32'h3a9de50e),
	.w7(32'h39a5d395),
	.w8(32'hb9daa98f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad41d8c),
	.w1(32'h3a68eb7f),
	.w2(32'hba4fa990),
	.w3(32'h3b280aeb),
	.w4(32'h3aac3546),
	.w5(32'hb9ed3dae),
	.w6(32'h3b101068),
	.w7(32'h3a5adc29),
	.w8(32'h35e8595d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a901c0),
	.w1(32'hb90380fd),
	.w2(32'h390af71a),
	.w3(32'h38ceb8bd),
	.w4(32'hb867eda3),
	.w5(32'h37b9f6d6),
	.w6(32'h37dd3163),
	.w7(32'h38806cc5),
	.w8(32'hb89a384a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e7e3f),
	.w1(32'hb9925fec),
	.w2(32'hb9f3b5a7),
	.w3(32'hb984556d),
	.w4(32'h368b9707),
	.w5(32'hb923bd3d),
	.w6(32'hb9b1caa5),
	.w7(32'hb9268447),
	.w8(32'h39156a6c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb851d369),
	.w1(32'hb990c34b),
	.w2(32'hb995950e),
	.w3(32'hb9140540),
	.w4(32'h3718ee29),
	.w5(32'hb92f5fbe),
	.w6(32'h3728ad88),
	.w7(32'h378daab3),
	.w8(32'hb8aa6bb1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d73ebc),
	.w1(32'h38c6388e),
	.w2(32'h3a9d9e53),
	.w3(32'h3998b011),
	.w4(32'h398aacaa),
	.w5(32'h3a3377bd),
	.w6(32'h39d63945),
	.w7(32'h3a073d2c),
	.w8(32'h36c71eb6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a089db8),
	.w1(32'hb6a7cd11),
	.w2(32'hb952ae9a),
	.w3(32'h39b1c62c),
	.w4(32'hb894861d),
	.w5(32'hb931fe2a),
	.w6(32'h39292732),
	.w7(32'hb9707b57),
	.w8(32'hb8cb257f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a839fe8),
	.w1(32'h3a94c007),
	.w2(32'hb82640e9),
	.w3(32'h3a9d66a4),
	.w4(32'h3a5df7f8),
	.w5(32'hb9320aa3),
	.w6(32'h3aaf9ba9),
	.w7(32'hb9abc360),
	.w8(32'h3951b6e2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399df2b9),
	.w1(32'hb85731c8),
	.w2(32'h37e68ac8),
	.w3(32'hb7e5336d),
	.w4(32'hb8002264),
	.w5(32'h37edb2a8),
	.w6(32'h386b9ac4),
	.w7(32'h3867ea43),
	.w8(32'h3939f0d0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387205bf),
	.w1(32'hb8822ad4),
	.w2(32'hb9768c4d),
	.w3(32'h37d3985b),
	.w4(32'h391bef3e),
	.w5(32'hb9d184e7),
	.w6(32'h37c7a87a),
	.w7(32'hb8cbb2f1),
	.w8(32'h39a0e527),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16ada7),
	.w1(32'hb94a0037),
	.w2(32'hb93fd6fe),
	.w3(32'h39b2d094),
	.w4(32'hb9931049),
	.w5(32'hb9aa415e),
	.w6(32'hb9d67b00),
	.w7(32'hb9667781),
	.w8(32'hb99063d7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5bc6b),
	.w1(32'hb980d413),
	.w2(32'h3a413b8a),
	.w3(32'hb9856aec),
	.w4(32'hb85f073d),
	.w5(32'hb95c4ca0),
	.w6(32'h399dd9d6),
	.w7(32'h37b72bf3),
	.w8(32'h3a2f1408),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab2182),
	.w1(32'hb949ad6b),
	.w2(32'h3843e53b),
	.w3(32'hb944f93e),
	.w4(32'hb8e4d01c),
	.w5(32'h390ae248),
	.w6(32'h390bd04e),
	.w7(32'h39c3974f),
	.w8(32'h37f27640),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eb0045),
	.w1(32'hba10c3b0),
	.w2(32'hba144a5f),
	.w3(32'h394f49a9),
	.w4(32'hb98934c1),
	.w5(32'hb9d296c5),
	.w6(32'hb92d44ee),
	.w7(32'hb94c36de),
	.w8(32'hb9b167ed),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f10d0c),
	.w1(32'hb99afac3),
	.w2(32'hb97495e3),
	.w3(32'h39b63d08),
	.w4(32'h38e7121a),
	.w5(32'hb97d29fc),
	.w6(32'h39c56d87),
	.w7(32'hb8afd3ce),
	.w8(32'hb9feeec8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd1e76),
	.w1(32'h389d450a),
	.w2(32'hb99d97ab),
	.w3(32'hb96e8ce3),
	.w4(32'h3992674d),
	.w5(32'h38714069),
	.w6(32'h38fa0736),
	.w7(32'hb9f02b13),
	.w8(32'hb93ec1bd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a5cd1),
	.w1(32'h3a59b96f),
	.w2(32'h3aa50ec4),
	.w3(32'hb872bb3e),
	.w4(32'h3a4c6800),
	.w5(32'h3a387da3),
	.w6(32'h39a4cdc9),
	.w7(32'h39c4d602),
	.w8(32'h3a398562),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a296452),
	.w1(32'h3a693f4d),
	.w2(32'h39d94310),
	.w3(32'h38d1086a),
	.w4(32'h3a91e5ce),
	.w5(32'h3a2c4a9d),
	.w6(32'h3a7ee428),
	.w7(32'h3a15c2a6),
	.w8(32'h39b12b41),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387412f5),
	.w1(32'hb9ba9b82),
	.w2(32'hb98067ff),
	.w3(32'h3986e7f3),
	.w4(32'hb99fb2a8),
	.w5(32'hba194895),
	.w6(32'hb9cb0b81),
	.w7(32'hba032901),
	.w8(32'hb99d2ed5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990772b),
	.w1(32'hb8b9315f),
	.w2(32'h3a4e929f),
	.w3(32'hb9d4d426),
	.w4(32'hb847a064),
	.w5(32'h397d89b8),
	.w6(32'hb7104dad),
	.w7(32'hb9206dea),
	.w8(32'hb766fd6c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393460fd),
	.w1(32'h39daea12),
	.w2(32'h395db218),
	.w3(32'h3a7041c3),
	.w4(32'h3a40eeed),
	.w5(32'h3a0eb385),
	.w6(32'h3a6171ac),
	.w7(32'h39d0eea4),
	.w8(32'h3a205592),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad27d7a),
	.w1(32'h393f794c),
	.w2(32'hba15e3fa),
	.w3(32'h3ac02a17),
	.w4(32'h37907e31),
	.w5(32'hba023011),
	.w6(32'h3ac1bd41),
	.w7(32'h3a924cb9),
	.w8(32'h3984b4a8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a736908),
	.w1(32'h38158246),
	.w2(32'hb950b420),
	.w3(32'h39f37af2),
	.w4(32'hb93445e0),
	.w5(32'hb9923f73),
	.w6(32'h3a42e602),
	.w7(32'h39e77385),
	.w8(32'h391fba54),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a834968),
	.w1(32'hb885b860),
	.w2(32'hba0dad39),
	.w3(32'h3aac12fb),
	.w4(32'h39b79649),
	.w5(32'hba18ab74),
	.w6(32'h3af4df73),
	.w7(32'h3a4afb0c),
	.w8(32'h389472b7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39886061),
	.w1(32'h38b76768),
	.w2(32'h39a54583),
	.w3(32'h39e81d65),
	.w4(32'h38c125c8),
	.w5(32'h395744e7),
	.w6(32'h38edc231),
	.w7(32'h3976021c),
	.w8(32'hb897480a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f1992),
	.w1(32'hb9c8edd0),
	.w2(32'h37dcb173),
	.w3(32'hb95722fe),
	.w4(32'hb9b67bb4),
	.w5(32'hb7e0449a),
	.w6(32'hb9a91619),
	.w7(32'hb9329b4e),
	.w8(32'hb91184ba),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ea415c),
	.w1(32'hb9cce21b),
	.w2(32'hb997729a),
	.w3(32'hb6d4d7ae),
	.w4(32'hb996dfd5),
	.w5(32'hb969e267),
	.w6(32'hb9afd0d0),
	.w7(32'hb9929971),
	.w8(32'hb98f36ba),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9468ba6),
	.w1(32'hb9854260),
	.w2(32'h3929c34b),
	.w3(32'hb94cadf7),
	.w4(32'hb9cfc78d),
	.w5(32'hb8cd88eb),
	.w6(32'hb97e20f9),
	.w7(32'hb953f266),
	.w8(32'hb93568b7),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb861c081),
	.w1(32'hb9ba3081),
	.w2(32'h3880ae05),
	.w3(32'hb9003281),
	.w4(32'hb950dd53),
	.w5(32'hb899429c),
	.w6(32'hb69caca7),
	.w7(32'hb8ac2adf),
	.w8(32'hb89e0d4a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb872a444),
	.w1(32'h39b55950),
	.w2(32'h37a5cca2),
	.w3(32'h381f9380),
	.w4(32'hb976f3fa),
	.w5(32'h39a156ee),
	.w6(32'h3a92e36e),
	.w7(32'h3a52c46a),
	.w8(32'hb8aa271b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a906eec),
	.w1(32'hb87253ed),
	.w2(32'hba3b82b0),
	.w3(32'h3a843e46),
	.w4(32'h39a638d8),
	.w5(32'hb9390d08),
	.w6(32'h3ab5763c),
	.w7(32'hb92deebb),
	.w8(32'hb913c180),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a530ae0),
	.w1(32'h369ece28),
	.w2(32'hb943f1fa),
	.w3(32'h3ac458c3),
	.w4(32'h3a15ee17),
	.w5(32'hb98c4180),
	.w6(32'h3a924b4c),
	.w7(32'h3a0062a2),
	.w8(32'hb9d3a87b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44f968),
	.w1(32'h39fa3a45),
	.w2(32'h359fe7a4),
	.w3(32'h3a4623ba),
	.w4(32'h39f54561),
	.w5(32'hb94dd593),
	.w6(32'h3a70cabd),
	.w7(32'h39c100ed),
	.w8(32'h388b4bf9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9574537),
	.w1(32'hb987405a),
	.w2(32'hb9e7a984),
	.w3(32'h3a0deb3d),
	.w4(32'h38bacacc),
	.w5(32'hb8e8d16d),
	.w6(32'h3965db1e),
	.w7(32'hb89786d0),
	.w8(32'h37c8f53c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932a2d8),
	.w1(32'hb8ebf3be),
	.w2(32'hb95af336),
	.w3(32'h39754464),
	.w4(32'hb99bc2db),
	.w5(32'hb9df617d),
	.w6(32'h39f3d6d7),
	.w7(32'h3a095b39),
	.w8(32'h3995418e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a356122),
	.w1(32'h38b364e4),
	.w2(32'h3825ed37),
	.w3(32'h3a1ee8c6),
	.w4(32'h399c826b),
	.w5(32'h399410ad),
	.w6(32'h3a133b31),
	.w7(32'h39f065ac),
	.w8(32'hb81b713d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c1eac),
	.w1(32'hb81075f4),
	.w2(32'hb73e6522),
	.w3(32'hb803753c),
	.w4(32'h38d0b9ed),
	.w5(32'hb852ab19),
	.w6(32'h391a36b4),
	.w7(32'h38927892),
	.w8(32'h398abcc1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391ed4ee),
	.w1(32'h36489c55),
	.w2(32'h39a034fe),
	.w3(32'h38d99eec),
	.w4(32'h3894fff0),
	.w5(32'h398a8088),
	.w6(32'h38fb393c),
	.w7(32'h3964d28c),
	.w8(32'hb924e22c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8420923),
	.w1(32'hb9263d46),
	.w2(32'h3a42687e),
	.w3(32'hb822f3b8),
	.w4(32'hb98d9f32),
	.w5(32'h3a13e26b),
	.w6(32'h37fefb61),
	.w7(32'h39493ecb),
	.w8(32'hb94e064e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915bc16),
	.w1(32'h398260c2),
	.w2(32'h39bd93bc),
	.w3(32'hb978eb4b),
	.w4(32'h3946ba49),
	.w5(32'h39afc118),
	.w6(32'h390aa7ac),
	.w7(32'h3970c8d4),
	.w8(32'h3905e11b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68018d),
	.w1(32'h39e0d7e9),
	.w2(32'h398ed578),
	.w3(32'hb9ee0931),
	.w4(32'hb998f806),
	.w5(32'hb9df5b06),
	.w6(32'hba9858aa),
	.w7(32'hba99c222),
	.w8(32'hbabac0d4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb911bb29),
	.w1(32'hb972ee02),
	.w2(32'hb8638d55),
	.w3(32'hb62d22d4),
	.w4(32'hb92480dc),
	.w5(32'hb95e3d19),
	.w6(32'hb8daf7d5),
	.w7(32'hb8aeedc2),
	.w8(32'hb760b92b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee9312),
	.w1(32'h393302ac),
	.w2(32'hba06d862),
	.w3(32'h3a12cd98),
	.w4(32'h396fd4ec),
	.w5(32'hb98f332b),
	.w6(32'h3a5a8128),
	.w7(32'h399c81cc),
	.w8(32'h3971c16e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cdbef),
	.w1(32'hb81e5e5b),
	.w2(32'hb99b54be),
	.w3(32'h3a1a7370),
	.w4(32'hb861e8f2),
	.w5(32'h36ba432b),
	.w6(32'h395dca1d),
	.w7(32'h38b31044),
	.w8(32'hb8201155),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ba094),
	.w1(32'hba305008),
	.w2(32'hb9b3e200),
	.w3(32'hb910f04f),
	.w4(32'hba5b8f5e),
	.w5(32'hb9ff6699),
	.w6(32'hb9b63424),
	.w7(32'hb9e85511),
	.w8(32'hb880109a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9ad8d),
	.w1(32'h39bfe965),
	.w2(32'hb9218f1d),
	.w3(32'h393e734f),
	.w4(32'h38e59c54),
	.w5(32'hba38bbd6),
	.w6(32'h3a1000af),
	.w7(32'h396b6c97),
	.w8(32'hb9d75381),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb848abe7),
	.w1(32'h39406250),
	.w2(32'h3914add8),
	.w3(32'hb889c7f7),
	.w4(32'hb92099e8),
	.w5(32'hb9222bf4),
	.w6(32'h3a307089),
	.w7(32'h39368791),
	.w8(32'h395108e7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f7175),
	.w1(32'h394bf01c),
	.w2(32'hb9921f0d),
	.w3(32'h3a3f5a32),
	.w4(32'h37974366),
	.w5(32'hb95f4892),
	.w6(32'h3a91a92f),
	.w7(32'h3999b869),
	.w8(32'h3a118623),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938f1b8),
	.w1(32'hba3e3624),
	.w2(32'hbaa76f7f),
	.w3(32'hb8ae3b51),
	.w4(32'hba3b8016),
	.w5(32'hba6d67c0),
	.w6(32'hb952f29a),
	.w7(32'hba5e79bd),
	.w8(32'hba2b04f7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3970f643),
	.w1(32'h39fb895d),
	.w2(32'hb914f98f),
	.w3(32'h38b888d4),
	.w4(32'h3a23348a),
	.w5(32'h388b3a81),
	.w6(32'h3a7c1a34),
	.w7(32'hb8ee9e44),
	.w8(32'hb93357d3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8b627),
	.w1(32'h3820a6b8),
	.w2(32'h3a353058),
	.w3(32'h39a87378),
	.w4(32'h3935a970),
	.w5(32'h39e1d22d),
	.w6(32'hb9872aa6),
	.w7(32'h3a7d11cc),
	.w8(32'h39de604c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abece8d),
	.w1(32'h37822dc6),
	.w2(32'hba622dfd),
	.w3(32'h3a92e267),
	.w4(32'h3a126f37),
	.w5(32'hba4d8c37),
	.w6(32'h3ad0fcf1),
	.w7(32'h3a4780fe),
	.w8(32'h39db0234),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b749f5),
	.w1(32'h38d48711),
	.w2(32'hb815e927),
	.w3(32'h37d6d0ad),
	.w4(32'h39185e26),
	.w5(32'hb91cdd4b),
	.w6(32'hb9f2f730),
	.w7(32'hb9b48b35),
	.w8(32'hb99449d7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71018f6),
	.w1(32'h393327bc),
	.w2(32'hb98e8492),
	.w3(32'h38e05fc8),
	.w4(32'hb9c64630),
	.w5(32'hb8e982a4),
	.w6(32'h3a3d24d5),
	.w7(32'hb9a5123b),
	.w8(32'hb975b655),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96cc10),
	.w1(32'h3ab4f5f1),
	.w2(32'h3a43930f),
	.w3(32'hbb092eda),
	.w4(32'hba4d39bf),
	.w5(32'hbb1f745d),
	.w6(32'hbb536144),
	.w7(32'hba726d5a),
	.w8(32'hbaa9cd91),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e73e9),
	.w1(32'h3a9e54f9),
	.w2(32'h39bc8ce0),
	.w3(32'h3a73bd92),
	.w4(32'h3a325520),
	.w5(32'hb900244e),
	.w6(32'h3b17034e),
	.w7(32'h3a5c6ccc),
	.w8(32'hb79fbc8b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa32c94),
	.w1(32'h396f4637),
	.w2(32'hba9498fd),
	.w3(32'h3ad4b4a8),
	.w4(32'h3909aa7f),
	.w5(32'hba315c81),
	.w6(32'hb93a0278),
	.w7(32'hbadb953e),
	.w8(32'hba48138f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce9edf),
	.w1(32'hb8eeb8c0),
	.w2(32'h39e4a115),
	.w3(32'h3856d846),
	.w4(32'hb9d8a92e),
	.w5(32'hb8a33b44),
	.w6(32'h39832aab),
	.w7(32'h37bca8b1),
	.w8(32'hb97d0515),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac68595),
	.w1(32'h3a4552dc),
	.w2(32'hb9a63af4),
	.w3(32'h3a98d9d4),
	.w4(32'h3a2ac420),
	.w5(32'hb95c9bb0),
	.w6(32'h3a32b115),
	.w7(32'h38b71962),
	.w8(32'hb99a5d1d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0ffb9),
	.w1(32'hb93f07f3),
	.w2(32'hb9fe2a93),
	.w3(32'h3a05ccff),
	.w4(32'h398dc4ff),
	.w5(32'hba3f7791),
	.w6(32'h390a99ae),
	.w7(32'h3925b14c),
	.w8(32'hb9689065),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83816a9),
	.w1(32'hba11b832),
	.w2(32'hb9deaa0c),
	.w3(32'hb878788d),
	.w4(32'hb9e5e427),
	.w5(32'hb9ef7cd6),
	.w6(32'hb99dc345),
	.w7(32'hb9d8d336),
	.w8(32'hb9fbffb2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba4f69),
	.w1(32'hb95e74fd),
	.w2(32'hb9a9fc5f),
	.w3(32'hb9ef9716),
	.w4(32'hb9cc3476),
	.w5(32'hba04602c),
	.w6(32'hb92f9c2f),
	.w7(32'hb8e998cc),
	.w8(32'h39306557),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8def59),
	.w1(32'h3901b899),
	.w2(32'hba3c5507),
	.w3(32'h3ada19a8),
	.w4(32'h3a357275),
	.w5(32'hb9636ed8),
	.w6(32'h3b0769b2),
	.w7(32'h3a6e95a2),
	.w8(32'h39395928),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eba1f),
	.w1(32'h3a14be73),
	.w2(32'hba205148),
	.w3(32'h3a4124f1),
	.w4(32'h3a54c56d),
	.w5(32'hb9795733),
	.w6(32'h3a8b04c9),
	.w7(32'h39827502),
	.w8(32'hb9fda142),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c50b2f),
	.w1(32'hba544b1e),
	.w2(32'hba703810),
	.w3(32'hb989694b),
	.w4(32'hba624880),
	.w5(32'hba9b20ee),
	.w6(32'hb948cc04),
	.w7(32'hba01248f),
	.w8(32'hba85b8fa),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d03a47),
	.w1(32'h3acb02de),
	.w2(32'h39f4b90b),
	.w3(32'h39cc64c2),
	.w4(32'h3af33523),
	.w5(32'h39f8df25),
	.w6(32'h3a0309b7),
	.w7(32'hb9294963),
	.w8(32'h396ddb70),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a3a280),
	.w1(32'hba3bd496),
	.w2(32'hba13d4c7),
	.w3(32'hb9d51089),
	.w4(32'hba593417),
	.w5(32'hba412ab5),
	.w6(32'hb9a71958),
	.w7(32'hb9faae7a),
	.w8(32'hba80ad1f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7941f),
	.w1(32'hb9bdf92e),
	.w2(32'hba080ae3),
	.w3(32'h3a475dcc),
	.w4(32'hb6a7ab4a),
	.w5(32'hba3f2fd7),
	.w6(32'h39adca1b),
	.w7(32'h38bff296),
	.w8(32'hba1d0673),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a533e),
	.w1(32'h373ad723),
	.w2(32'hba405455),
	.w3(32'hb9713f1d),
	.w4(32'h39407ea8),
	.w5(32'hb9effd8f),
	.w6(32'h3987f542),
	.w7(32'hb999de1c),
	.w8(32'hb9fb136e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30afde),
	.w1(32'hb9887236),
	.w2(32'hba13d42d),
	.w3(32'hb9db20e6),
	.w4(32'hb8290d47),
	.w5(32'hb9da1000),
	.w6(32'hb898e799),
	.w7(32'hba0d212d),
	.w8(32'hb92a42d0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cdd30d),
	.w1(32'hb9dc1619),
	.w2(32'hb9a13bc2),
	.w3(32'h38b431be),
	.w4(32'hb9d39d1d),
	.w5(32'hb9d0317e),
	.w6(32'hb9afcbba),
	.w7(32'hb9e52f27),
	.w8(32'hb971d2a3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb870b3f3),
	.w1(32'hb9be50e8),
	.w2(32'hb9c3f52d),
	.w3(32'hb98b9dbc),
	.w4(32'hb9e4e899),
	.w5(32'hb9f9562b),
	.w6(32'hb99b7572),
	.w7(32'hba211e88),
	.w8(32'hb97f0415),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98bb4b4),
	.w1(32'hb9f59075),
	.w2(32'hba1e8067),
	.w3(32'hb99c4897),
	.w4(32'h39a83a79),
	.w5(32'h39b885b1),
	.w6(32'hb983e0e0),
	.w7(32'hba241d6e),
	.w8(32'h38c6d4aa),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8baee24),
	.w1(32'hba6f4094),
	.w2(32'hba9b614c),
	.w3(32'h3a2636cc),
	.w4(32'hb9c49daf),
	.w5(32'hbacbea34),
	.w6(32'h39f9a97b),
	.w7(32'hb94289f7),
	.w8(32'hba15b44b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e113cb),
	.w1(32'h397dac13),
	.w2(32'h38f0f61f),
	.w3(32'hba0d1b62),
	.w4(32'h398c9d0d),
	.w5(32'h38323298),
	.w6(32'h39e9a880),
	.w7(32'h395f9146),
	.w8(32'hb838296d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e41bb),
	.w1(32'h39791792),
	.w2(32'hb9a1ff1a),
	.w3(32'h3aa2fd01),
	.w4(32'h39fb3fe9),
	.w5(32'h38d84b6b),
	.w6(32'h39e1fa27),
	.w7(32'h38a43d5b),
	.w8(32'h36ea7a3f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efa7e1),
	.w1(32'hba4253f8),
	.w2(32'hba754cdb),
	.w3(32'h3920eead),
	.w4(32'hba224549),
	.w5(32'hba87bca0),
	.w6(32'hb9e4e073),
	.w7(32'hba6b48fa),
	.w8(32'hba604bff),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94fdc5c),
	.w1(32'h38faa35c),
	.w2(32'hb9da4969),
	.w3(32'hb96a67f8),
	.w4(32'h3a204c08),
	.w5(32'h3a1f984f),
	.w6(32'hb8a0972f),
	.w7(32'h39b38b6f),
	.w8(32'h39561840),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388ec7ce),
	.w1(32'hb9302fd8),
	.w2(32'hb954a54e),
	.w3(32'h3a078366),
	.w4(32'hb92cc28b),
	.w5(32'hb97f6f9f),
	.w6(32'h3903ec99),
	.w7(32'hb91152ef),
	.w8(32'h3851e19b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937419f),
	.w1(32'hb9a7cdae),
	.w2(32'hb8e3d7df),
	.w3(32'hb97b104f),
	.w4(32'hb9963ec1),
	.w5(32'hb971a3e1),
	.w6(32'hb95826da),
	.w7(32'hb93faf6a),
	.w8(32'h38c53be6),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0b298),
	.w1(32'hb94b7e53),
	.w2(32'hb9f0e26c),
	.w3(32'h38d15edf),
	.w4(32'hb991b60c),
	.w5(32'hb9db42d1),
	.w6(32'h37fb27e5),
	.w7(32'hb997995e),
	.w8(32'hb98b3593),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a02f57),
	.w1(32'h38a14dbe),
	.w2(32'h39a5bf37),
	.w3(32'h381e8408),
	.w4(32'hb87cdc00),
	.w5(32'h3910e3c4),
	.w6(32'h37da9c96),
	.w7(32'hb7549e70),
	.w8(32'h393e45a6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98f89f),
	.w1(32'h3a13a8b4),
	.w2(32'hb9cf1806),
	.w3(32'h3a84a7b0),
	.w4(32'h3a2029c3),
	.w5(32'h393c7ef8),
	.w6(32'h3a7da5dd),
	.w7(32'h39fd944d),
	.w8(32'hb8913841),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba6333),
	.w1(32'hb8e97331),
	.w2(32'hb896a784),
	.w3(32'hb6a160fb),
	.w4(32'hb88e1337),
	.w5(32'hb7bf78d7),
	.w6(32'hb9a2afca),
	.w7(32'hb999eddc),
	.w8(32'hb9a0640c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ab7cf1),
	.w1(32'hb956efee),
	.w2(32'hb991c177),
	.w3(32'h3806e225),
	.w4(32'hb998d9fa),
	.w5(32'hb98b7f49),
	.w6(32'hb8f83e14),
	.w7(32'hb9958ef7),
	.w8(32'hb9f4eaaa),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c52afe),
	.w1(32'hb9718742),
	.w2(32'hb9f95b8c),
	.w3(32'hb9b98602),
	.w4(32'hb92a146c),
	.w5(32'hb95466f2),
	.w6(32'hb8bf1b42),
	.w7(32'hb98b84bb),
	.w8(32'hb72a545a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa1a67),
	.w1(32'h39c68be1),
	.w2(32'hb8b0108c),
	.w3(32'h39d047e7),
	.w4(32'h398a3e2d),
	.w5(32'hb88733d5),
	.w6(32'h3a712097),
	.w7(32'h39ec0138),
	.w8(32'h37f8c828),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ff871),
	.w1(32'hb9b0d27a),
	.w2(32'hb9cad5bd),
	.w3(32'h3a0f11b1),
	.w4(32'hb95b6b53),
	.w5(32'hb9abf5ae),
	.w6(32'hb78a529c),
	.w7(32'hb861f732),
	.w8(32'hb9381ffd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01a168),
	.w1(32'hb7c6fa21),
	.w2(32'hb9dc57e7),
	.w3(32'h3a20c6a8),
	.w4(32'h38c6798f),
	.w5(32'hba168a28),
	.w6(32'h3a16a3b7),
	.w7(32'h380de956),
	.w8(32'hb9d7c12b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08f913),
	.w1(32'h3920c88e),
	.w2(32'hba319508),
	.w3(32'h39b267ce),
	.w4(32'h3974dbee),
	.w5(32'hb9de5524),
	.w6(32'h39eac50c),
	.w7(32'h372eb298),
	.w8(32'hb9887324),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8827b5),
	.w1(32'h3a47a38b),
	.w2(32'hb9855160),
	.w3(32'h3988b013),
	.w4(32'h399476ca),
	.w5(32'hb9b441ce),
	.w6(32'hb926a282),
	.w7(32'hb9e7655a),
	.w8(32'hb9a62e7a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a173635),
	.w1(32'h382891a0),
	.w2(32'hb9a52e6b),
	.w3(32'h3966eb13),
	.w4(32'hb96cc718),
	.w5(32'hb9edb3fe),
	.w6(32'hb9b21397),
	.w7(32'hba21d76e),
	.w8(32'hba48a046),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3840e795),
	.w1(32'h3971fed5),
	.w2(32'hb81a725e),
	.w3(32'h38590e6b),
	.w4(32'hb9211642),
	.w5(32'hb8a7056d),
	.w6(32'h3a2cc8e6),
	.w7(32'h3916b0c7),
	.w8(32'h39302518),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8021fd),
	.w1(32'h39ace044),
	.w2(32'hb9de5f66),
	.w3(32'h3a83fe8d),
	.w4(32'h39ef10f6),
	.w5(32'hb98ceca6),
	.w6(32'h3a86d0e3),
	.w7(32'h39ad9b8d),
	.w8(32'hb9a34e85),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d29bf0),
	.w1(32'hb8820b77),
	.w2(32'hb9ad14e3),
	.w3(32'h3966fbe4),
	.w4(32'h385e6940),
	.w5(32'hb8e83104),
	.w6(32'h39907d84),
	.w7(32'h377a1102),
	.w8(32'hb93654a2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b981df),
	.w1(32'hb9cd8198),
	.w2(32'hba9b0fae),
	.w3(32'h3946ecaa),
	.w4(32'hb9b218cb),
	.w5(32'hbad57d4a),
	.w6(32'hb90a3120),
	.w7(32'hba625524),
	.w8(32'hba6b6ecd),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82a7b2c),
	.w1(32'hb7511330),
	.w2(32'hb9cbe8fb),
	.w3(32'hba2e9df9),
	.w4(32'hb8a8e467),
	.w5(32'h3985659a),
	.w6(32'h38c51ffa),
	.w7(32'hb9cda525),
	.w8(32'h389dc296),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993402b),
	.w1(32'hb8ec5b68),
	.w2(32'hb8b1790a),
	.w3(32'h3a0efea3),
	.w4(32'hb882bd2d),
	.w5(32'hb837bfd8),
	.w6(32'hb8b762ed),
	.w7(32'hb88bce38),
	.w8(32'hb8b0d845),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91450b5),
	.w1(32'hb6fcc884),
	.w2(32'h38c306bb),
	.w3(32'hb9362580),
	.w4(32'hb9835fe9),
	.w5(32'hb90d8a9b),
	.w6(32'h38dda606),
	.w7(32'h38dccf7b),
	.w8(32'hb873cfb0),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38be9961),
	.w1(32'hb9bab7cd),
	.w2(32'hb9a8e719),
	.w3(32'hb81b9884),
	.w4(32'hb9af9b41),
	.w5(32'hb982c03e),
	.w6(32'hba01d377),
	.w7(32'hb9d2f66b),
	.w8(32'hb9c36c5d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae8c78),
	.w1(32'h39ced886),
	.w2(32'hb9e0aaa8),
	.w3(32'h38c461cc),
	.w4(32'h391c81e3),
	.w5(32'hb9d15fe3),
	.w6(32'hb8830d79),
	.w7(32'hb9bd7c82),
	.w8(32'hb995a240),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5be697),
	.w1(32'h39d8efa4),
	.w2(32'hb97f01cb),
	.w3(32'h3a9593b5),
	.w4(32'h39937efb),
	.w5(32'hb9f4960b),
	.w6(32'h3a275052),
	.w7(32'hb7d00bc9),
	.w8(32'hba46debf),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37008a5e),
	.w1(32'h38f242f9),
	.w2(32'h39389170),
	.w3(32'hb8092d1c),
	.w4(32'h388a31a5),
	.w5(32'hb8e43fa3),
	.w6(32'h38b877fb),
	.w7(32'h391040c2),
	.w8(32'h378870d6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d33c9),
	.w1(32'hb9ef0513),
	.w2(32'hbab909f5),
	.w3(32'h3a6c492d),
	.w4(32'h39e8b143),
	.w5(32'hb8827555),
	.w6(32'h3a515b46),
	.w7(32'h399a7903),
	.w8(32'hba0f2d1c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bdad01),
	.w1(32'h390d02f1),
	.w2(32'hb861b892),
	.w3(32'h3a64f6cd),
	.w4(32'h39e42b19),
	.w5(32'h39801d5e),
	.w6(32'h3aaa64ab),
	.w7(32'h3a85c3c4),
	.w8(32'h3a6644ec),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1fbc6),
	.w1(32'h39886b44),
	.w2(32'hb9bc2dff),
	.w3(32'h3aae3275),
	.w4(32'h3a05f5d5),
	.w5(32'hb97a7cda),
	.w6(32'h3aab95db),
	.w7(32'h3a549c6c),
	.w8(32'h38b6bbe4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3825db4f),
	.w1(32'hba09265a),
	.w2(32'hba691ab1),
	.w3(32'h39a3f504),
	.w4(32'hb927caab),
	.w5(32'hba1ed0d3),
	.w6(32'h3a52be70),
	.w7(32'h392be315),
	.w8(32'hb9b50a8b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24fd66),
	.w1(32'hb9bed4c1),
	.w2(32'h389cfc98),
	.w3(32'hba7b97b4),
	.w4(32'hba7d5231),
	.w5(32'hb7529c1e),
	.w6(32'hb9420bdb),
	.w7(32'hb9ea19de),
	.w8(32'hb98ee56d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c2090),
	.w1(32'h3a0d23c4),
	.w2(32'hb9653539),
	.w3(32'h393134f6),
	.w4(32'h3a1055bd),
	.w5(32'hb91cbca9),
	.w6(32'h3a6c9bc3),
	.w7(32'h3a780821),
	.w8(32'h3984e364),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7301e),
	.w1(32'h37f99787),
	.w2(32'hba898276),
	.w3(32'h3985277d),
	.w4(32'h38294164),
	.w5(32'hb9e12464),
	.w6(32'h391c914e),
	.w7(32'hb9bc6118),
	.w8(32'hba18f385),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7815869),
	.w1(32'hb8ab473e),
	.w2(32'hb8a64a34),
	.w3(32'hba655b83),
	.w4(32'hba3c316c),
	.w5(32'hba72541a),
	.w6(32'hbaa0e0f8),
	.w7(32'hba93d102),
	.w8(32'hb9a0778f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e47368),
	.w1(32'hb84217d8),
	.w2(32'hb8d73352),
	.w3(32'hb9401c88),
	.w4(32'hb9a946d4),
	.w5(32'hba0a6817),
	.w6(32'h395fe31f),
	.w7(32'h389b3e94),
	.w8(32'h38843b2e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a43dea),
	.w1(32'h388b0260),
	.w2(32'h389511b5),
	.w3(32'h38a75f5e),
	.w4(32'h38b23ac7),
	.w5(32'h3830cb07),
	.w6(32'h367cf13b),
	.w7(32'h386766a2),
	.w8(32'h3856841d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7983e38),
	.w1(32'hb8ae8e20),
	.w2(32'hb89c4d5c),
	.w3(32'hb8c29378),
	.w4(32'hb8696d4e),
	.w5(32'hb80f0065),
	.w6(32'hb8a8b4d9),
	.w7(32'hb7fadb46),
	.w8(32'hb875cb82),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e35d6),
	.w1(32'h39b078da),
	.w2(32'hba093b54),
	.w3(32'h3a99e0e8),
	.w4(32'h3a1bf781),
	.w5(32'hb9acc162),
	.w6(32'h3a76afe7),
	.w7(32'h3a087e6b),
	.w8(32'hb939df53),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998ef6b),
	.w1(32'hb981e418),
	.w2(32'hb92fef2c),
	.w3(32'hb935debb),
	.w4(32'hb8e7c3dc),
	.w5(32'hb9b940b0),
	.w6(32'hb96717c3),
	.w7(32'h38ef38b3),
	.w8(32'h392b1d7c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eac74),
	.w1(32'hb94881aa),
	.w2(32'hba532093),
	.w3(32'h39fa6051),
	.w4(32'hb702e8f4),
	.w5(32'hba078f44),
	.w6(32'h397eba2f),
	.w7(32'hb9227d86),
	.w8(32'hba2b8ab0),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aa0a0a),
	.w1(32'h392e8218),
	.w2(32'h382b4917),
	.w3(32'hb8b04dd6),
	.w4(32'h3991b662),
	.w5(32'hb78c8879),
	.w6(32'h37d635bb),
	.w7(32'h397c7147),
	.w8(32'hb8919522),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a3ff79),
	.w1(32'hb871dafc),
	.w2(32'h3949303c),
	.w3(32'hb8ce8fad),
	.w4(32'h380a4b64),
	.w5(32'h39168cfe),
	.w6(32'h38ee02f5),
	.w7(32'hb7f20409),
	.w8(32'hb95eab3f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f3479),
	.w1(32'hb83de8cc),
	.w2(32'hb756e40e),
	.w3(32'h39922cf1),
	.w4(32'hb8d48786),
	.w5(32'hb8e39ad2),
	.w6(32'hb81b2a70),
	.w7(32'h371285e3),
	.w8(32'hb8ce4716),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92bce38),
	.w1(32'hb7e0e32d),
	.w2(32'h38785d08),
	.w3(32'hb8de95aa),
	.w4(32'h38a9b8ca),
	.w5(32'h3880fb25),
	.w6(32'h38909092),
	.w7(32'h3913b992),
	.w8(32'h393b1603),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2476ce),
	.w1(32'h388460e7),
	.w2(32'hba4215a4),
	.w3(32'h3a72bdf6),
	.w4(32'h383847a6),
	.w5(32'hba237d42),
	.w6(32'h3a9d6e50),
	.w7(32'h3a0be0a0),
	.w8(32'hb9144b23),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a460d43),
	.w1(32'hb992a6f4),
	.w2(32'hba991762),
	.w3(32'h3aaf58d4),
	.w4(32'h39a68087),
	.w5(32'hba0e177c),
	.w6(32'h3ada5ff0),
	.w7(32'h3a277b5d),
	.w8(32'h3a28f460),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cfdef2),
	.w1(32'hba51f56e),
	.w2(32'hba039a17),
	.w3(32'hb9e21d2b),
	.w4(32'hba594302),
	.w5(32'hb9f3c5ed),
	.w6(32'hb9d8e99f),
	.w7(32'hb91b09aa),
	.w8(32'hba0ea812),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40d9fe),
	.w1(32'h39fb7df8),
	.w2(32'hb9a78576),
	.w3(32'h39f5f7b6),
	.w4(32'h394a860e),
	.w5(32'hb93f7f33),
	.w6(32'h3a583c39),
	.w7(32'h39f6e822),
	.w8(32'hb9a18a76),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902ed58),
	.w1(32'hb976b9d2),
	.w2(32'hb94f9fae),
	.w3(32'h38370535),
	.w4(32'hb9b6f7d1),
	.w5(32'hb9c9c980),
	.w6(32'hb804af4b),
	.w7(32'hb93c8222),
	.w8(32'hb8880ceb),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ae79c),
	.w1(32'h3a825445),
	.w2(32'hbabcbf71),
	.w3(32'h3a811ea4),
	.w4(32'h39bdfa41),
	.w5(32'hbb045ffc),
	.w6(32'h3a886737),
	.w7(32'hba5054b2),
	.w8(32'hbaa3b10e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b2a8b),
	.w1(32'h3a0cad9e),
	.w2(32'h379d19a7),
	.w3(32'h3a11df81),
	.w4(32'h3a02fe61),
	.w5(32'h385e27df),
	.w6(32'h3a844e2a),
	.w7(32'h3a3ea68a),
	.w8(32'h39989634),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59a4ec),
	.w1(32'hb91659ea),
	.w2(32'hbaad7732),
	.w3(32'h39f0c3fc),
	.w4(32'hb952616a),
	.w5(32'hba482d0c),
	.w6(32'h3a8eb593),
	.w7(32'h39865aec),
	.w8(32'hb9610024),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3848b140),
	.w1(32'h38d08b98),
	.w2(32'h38c4a20c),
	.w3(32'h39511e19),
	.w4(32'hb700da11),
	.w5(32'hb93a1a4f),
	.w6(32'h39d08295),
	.w7(32'h39968fa0),
	.w8(32'h37c8970c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3af7eb),
	.w1(32'hb873346b),
	.w2(32'hb9bd2708),
	.w3(32'h3a4d9f6e),
	.w4(32'h39a83d13),
	.w5(32'h39226418),
	.w6(32'h3a1b828b),
	.w7(32'h389611be),
	.w8(32'h3940f85e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9332fa2),
	.w1(32'h387350cb),
	.w2(32'h38f96766),
	.w3(32'hb932d893),
	.w4(32'h3898a590),
	.w5(32'h38b46c7a),
	.w6(32'h38acec4d),
	.w7(32'h38912ada),
	.w8(32'h38dc3af4),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c89b02),
	.w1(32'h38900e42),
	.w2(32'h39190f83),
	.w3(32'h39495556),
	.w4(32'hb8cf9ab7),
	.w5(32'hb915cdd8),
	.w6(32'h39dbc49c),
	.w7(32'h39b7313a),
	.w8(32'h391ab1c7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3958abe0),
	.w1(32'h3a09ff6f),
	.w2(32'h38c3f097),
	.w3(32'h38b8375f),
	.w4(32'h3a68e323),
	.w5(32'h39d192f8),
	.w6(32'h3a055375),
	.w7(32'h3987fa77),
	.w8(32'h37e3867b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6635e),
	.w1(32'hb753f4ac),
	.w2(32'hb9b3d5e3),
	.w3(32'h39d6624d),
	.w4(32'hb8ed4f66),
	.w5(32'hba16dd8f),
	.w6(32'h3a0258b7),
	.w7(32'h38411098),
	.w8(32'hb9f57f87),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9172e31),
	.w1(32'h370618ed),
	.w2(32'hb919999e),
	.w3(32'hb8f2cda6),
	.w4(32'hb69b8c65),
	.w5(32'h38c5c308),
	.w6(32'h38e4d185),
	.w7(32'hb91fd8b4),
	.w8(32'hb9a1134e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999772d),
	.w1(32'h393b9364),
	.w2(32'hb8ea6201),
	.w3(32'hb89ae457),
	.w4(32'h3951930c),
	.w5(32'h38173fd2),
	.w6(32'hb5ef673b),
	.w7(32'hb96b5fb4),
	.w8(32'hb959a70a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980923f),
	.w1(32'hb917e097),
	.w2(32'hb83a7995),
	.w3(32'hb9699046),
	.w4(32'hb8f77f42),
	.w5(32'hb87cfc58),
	.w6(32'h38c97c11),
	.w7(32'h3979a4dc),
	.w8(32'h39889e89),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f1fbd),
	.w1(32'h3a006792),
	.w2(32'h371afdc4),
	.w3(32'h39ff04f5),
	.w4(32'hb80d5a09),
	.w5(32'hba1cfbb0),
	.w6(32'hba2c980b),
	.w7(32'hba392ff1),
	.w8(32'hba8208de),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37855d52),
	.w1(32'h39499ee7),
	.w2(32'h39c0f104),
	.w3(32'h380fc310),
	.w4(32'hb8f031d8),
	.w5(32'h39d39073),
	.w6(32'h3a179236),
	.w7(32'h3985f906),
	.w8(32'h3903c627),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce3833),
	.w1(32'hb98954f5),
	.w2(32'hb999f61e),
	.w3(32'h3921f15c),
	.w4(32'hb9a462de),
	.w5(32'hb9c73b8a),
	.w6(32'hb9ce3fee),
	.w7(32'hb9d44069),
	.w8(32'hb95e79ae),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eed25),
	.w1(32'h3ac9e435),
	.w2(32'hba8b7ba0),
	.w3(32'h3b3c1b9e),
	.w4(32'h3afcea41),
	.w5(32'hb97c8a3e),
	.w6(32'h3b20ac7b),
	.w7(32'h3a5726ae),
	.w8(32'h38b5352a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bd834),
	.w1(32'hba36cb17),
	.w2(32'hba769650),
	.w3(32'h3966a724),
	.w4(32'hbaa3277b),
	.w5(32'hba6f2af9),
	.w6(32'hb9b0fcd1),
	.w7(32'hbaca7173),
	.w8(32'hba57bb33),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9621bc4),
	.w1(32'hb8cd2e66),
	.w2(32'hb89ce612),
	.w3(32'hb92470c4),
	.w4(32'hb79be616),
	.w5(32'h38aa8080),
	.w6(32'h38b3f444),
	.w7(32'h391a9d5f),
	.w8(32'h39368487),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7534949),
	.w1(32'h38502836),
	.w2(32'h34dcf94a),
	.w3(32'hb88449b6),
	.w4(32'h393d206e),
	.w5(32'hb6aae17c),
	.w6(32'hb7af79de),
	.w7(32'h395543b7),
	.w8(32'h390daf62),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88548cd),
	.w1(32'hb7e84b53),
	.w2(32'hb98dea7d),
	.w3(32'hba08d1e8),
	.w4(32'hb9a47915),
	.w5(32'hb9e52198),
	.w6(32'hba05fe42),
	.w7(32'hb9b95899),
	.w8(32'hb9c3dc43),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cc5bad),
	.w1(32'hb9190362),
	.w2(32'hb9ac0c9e),
	.w3(32'hb8fd8be6),
	.w4(32'hb87f43fb),
	.w5(32'hb933e05f),
	.w6(32'hb8f4dad0),
	.w7(32'hb9419471),
	.w8(32'hb917242e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac807f),
	.w1(32'hb8c582b5),
	.w2(32'hb8bd58db),
	.w3(32'h38c1fec1),
	.w4(32'hb8db4333),
	.w5(32'hb726939c),
	.w6(32'h39131d6c),
	.w7(32'hb9547126),
	.w8(32'hb919e69a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39849c81),
	.w1(32'h396bd650),
	.w2(32'hb9fb98fe),
	.w3(32'h3969dc8e),
	.w4(32'hb858873a),
	.w5(32'hba0d4fb9),
	.w6(32'h39064281),
	.w7(32'hb9de55ce),
	.w8(32'hb9bc00f0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7b5e0),
	.w1(32'h39ff2ce8),
	.w2(32'hba2c6e20),
	.w3(32'h3aa985c2),
	.w4(32'h395ac8e3),
	.w5(32'hba550b8c),
	.w6(32'h3a9e0471),
	.w7(32'h391afa04),
	.w8(32'hba2ec641),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a1bd32),
	.w1(32'h37dd12e4),
	.w2(32'hb79e5e13),
	.w3(32'hb9611ecf),
	.w4(32'h38088e9b),
	.w5(32'hb8a52c12),
	.w6(32'h38916187),
	.w7(32'hb6793ba2),
	.w8(32'hb8c5e20f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a947da3),
	.w1(32'h3a65bece),
	.w2(32'hb985dd69),
	.w3(32'h3ac7bec9),
	.w4(32'h3a07d53f),
	.w5(32'hb984bbee),
	.w6(32'h3af3244f),
	.w7(32'h3a581075),
	.w8(32'h386d7bdc),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9bc4d),
	.w1(32'hb9c09a89),
	.w2(32'hb99c4311),
	.w3(32'h3916e612),
	.w4(32'hb9b33011),
	.w5(32'hba04d8bd),
	.w6(32'hba17c31e),
	.w7(32'hb9d9b65b),
	.w8(32'hba1ee611),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93336ca),
	.w1(32'hb8e00002),
	.w2(32'hb89cf27d),
	.w3(32'hb96208a9),
	.w4(32'hb8150203),
	.w5(32'hb7a68b49),
	.w6(32'hb83fb10f),
	.w7(32'hb8567cfe),
	.w8(32'h37b3c67f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d0d8e9),
	.w1(32'h3744cbf1),
	.w2(32'h37c79155),
	.w3(32'h388b608e),
	.w4(32'h38332e37),
	.w5(32'h38826682),
	.w6(32'hb88c9b82),
	.w7(32'hb7dc5f77),
	.w8(32'hb856ff88),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ce49bc),
	.w1(32'hb782b54f),
	.w2(32'h3799f61c),
	.w3(32'hb8fef735),
	.w4(32'h370c67da),
	.w5(32'h377aca0c),
	.w6(32'hb901aff9),
	.w7(32'h35d9ff3b),
	.w8(32'hb83ac62d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01b653),
	.w1(32'h38352ce1),
	.w2(32'hb9dde37f),
	.w3(32'h39bc7140),
	.w4(32'h38a19a2f),
	.w5(32'hb9ad4549),
	.w6(32'h399f2929),
	.w7(32'hb86aedac),
	.w8(32'hba1b74ad),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dbb19),
	.w1(32'h390806b2),
	.w2(32'h397ccff9),
	.w3(32'hba9948f2),
	.w4(32'hb9cea4e0),
	.w5(32'h39d0d8e1),
	.w6(32'hb86544f4),
	.w7(32'hb9cc2767),
	.w8(32'h38a17b34),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a219585),
	.w1(32'h39a12258),
	.w2(32'hb9540ad8),
	.w3(32'h3a8cf286),
	.w4(32'h39509f9e),
	.w5(32'hb965d12e),
	.w6(32'h3ab0298e),
	.w7(32'h3a46087d),
	.w8(32'h39f8aaf0),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2338e),
	.w1(32'hb91c3229),
	.w2(32'hb8f7ab3d),
	.w3(32'h38c8a06a),
	.w4(32'hb9a2995b),
	.w5(32'hb9b51970),
	.w6(32'hb98e02d8),
	.w7(32'hb969e88c),
	.w8(32'hb9c0d1c4),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab65c07),
	.w1(32'h3aa1e0f8),
	.w2(32'hb90518b5),
	.w3(32'h3a74fa20),
	.w4(32'h3a7e033b),
	.w5(32'hb9916b3f),
	.w6(32'h3ab3b18a),
	.w7(32'h3a02b76c),
	.w8(32'hba3f5ad6),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bec76c),
	.w1(32'h39a8ce97),
	.w2(32'hb998f932),
	.w3(32'h3a14f620),
	.w4(32'h3986bb0f),
	.w5(32'hb94fd1f0),
	.w6(32'h3a62c5e0),
	.w7(32'h3a0849db),
	.w8(32'h38891781),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ecb87),
	.w1(32'h39e8152f),
	.w2(32'hb91ef92d),
	.w3(32'hb8ba23a8),
	.w4(32'h3a09f48b),
	.w5(32'hba058b0a),
	.w6(32'hb77507ad),
	.w7(32'hb9c68eaa),
	.w8(32'hb9a403b1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388f28b7),
	.w1(32'hb9fdfcbc),
	.w2(32'hb9cd89f3),
	.w3(32'hb74dbe0d),
	.w4(32'hb9eb1044),
	.w5(32'hb9c6e650),
	.w6(32'hba135811),
	.w7(32'hb9e99b85),
	.w8(32'hba1d3c16),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00694e),
	.w1(32'h3681eda2),
	.w2(32'h38e4149f),
	.w3(32'hb9fcba32),
	.w4(32'h381d87d3),
	.w5(32'h37c1426b),
	.w6(32'h3872b952),
	.w7(32'h38f0690a),
	.w8(32'h38a550c6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b520d),
	.w1(32'h37238dbd),
	.w2(32'hb98453e9),
	.w3(32'h39386b27),
	.w4(32'hb8ee3226),
	.w5(32'hb9d20e9c),
	.w6(32'h39b66fa4),
	.w7(32'h393f6094),
	.w8(32'hb94b0f46),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f81ca8),
	.w1(32'h39b3adfe),
	.w2(32'hb9eb24bc),
	.w3(32'h3a5b1955),
	.w4(32'h39ce41d5),
	.w5(32'hba0da390),
	.w6(32'h3ab976cd),
	.w7(32'h3a806313),
	.w8(32'h39a96847),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a788b4c),
	.w1(32'hb897ee6a),
	.w2(32'hb9e08d04),
	.w3(32'h3a5ac70a),
	.w4(32'hb68d1f76),
	.w5(32'hb9f8f0ca),
	.w6(32'h3a8bebde),
	.w7(32'h39fb2b64),
	.w8(32'h388b6ac8),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39017657),
	.w1(32'hb685cb17),
	.w2(32'hb81d25a0),
	.w3(32'h397c3908),
	.w4(32'h39196dd7),
	.w5(32'h381a5f52),
	.w6(32'hb91380b4),
	.w7(32'hb9920452),
	.w8(32'hb8647fdf),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cacd08),
	.w1(32'h387d6cf9),
	.w2(32'h39074c2f),
	.w3(32'hb8b62d63),
	.w4(32'h3748c4e5),
	.w5(32'hb7ad176a),
	.w6(32'h376c49f9),
	.w7(32'h38a05d7c),
	.w8(32'h37ed0f82),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399125df),
	.w1(32'hb58764f5),
	.w2(32'hb941f5fc),
	.w3(32'h390c087e),
	.w4(32'h38fead3d),
	.w5(32'hb7d0af41),
	.w6(32'h379674c7),
	.w7(32'hb931d632),
	.w8(32'hb994a23f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9c404),
	.w1(32'hb83aeed8),
	.w2(32'h38c02470),
	.w3(32'hb9854bc9),
	.w4(32'hb93967e6),
	.w5(32'hb8383b8b),
	.w6(32'h38ad2b65),
	.w7(32'h33244be0),
	.w8(32'hb9910368),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe02c1),
	.w1(32'h3a97f239),
	.w2(32'h39d0f05e),
	.w3(32'h3a733abb),
	.w4(32'h3a92b639),
	.w5(32'h39cc1daa),
	.w6(32'h3a2fb419),
	.w7(32'hb9904c8e),
	.w8(32'hb9c912d8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a995af4),
	.w1(32'h39f0f3e3),
	.w2(32'hb961f152),
	.w3(32'h3a9d6927),
	.w4(32'h39791afb),
	.w5(32'hba12fe3a),
	.w6(32'h3a03ee7e),
	.w7(32'h38e4e858),
	.w8(32'hb9d486d3),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f9a38),
	.w1(32'h397c3b81),
	.w2(32'hb875441c),
	.w3(32'hba119dad),
	.w4(32'h38c29023),
	.w5(32'h379f318e),
	.w6(32'hba180932),
	.w7(32'hb9b1e882),
	.w8(32'hb9d2ce73),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac9a43),
	.w1(32'h38881565),
	.w2(32'hb96e8175),
	.w3(32'h3a1de2da),
	.w4(32'h38ec7df1),
	.w5(32'hb9dc1a5f),
	.w6(32'h3a328bb3),
	.w7(32'h3a27ecdb),
	.w8(32'h39103023),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3741b160),
	.w1(32'hb97f7ab8),
	.w2(32'hb9860460),
	.w3(32'hb7c17ff5),
	.w4(32'hb9015471),
	.w5(32'hb903e271),
	.w6(32'hb987bcdc),
	.w7(32'hb98a3120),
	.w8(32'hb98ce78b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952c271),
	.w1(32'hb9a2559a),
	.w2(32'hb9902140),
	.w3(32'hb9101c65),
	.w4(32'hb97c4e6c),
	.w5(32'hb89577e3),
	.w6(32'hb9636862),
	.w7(32'hb994bb81),
	.w8(32'hb9b0af6d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5d122),
	.w1(32'h3885c960),
	.w2(32'h388fd95e),
	.w3(32'hb8084f74),
	.w4(32'h3907d513),
	.w5(32'hb781b674),
	.w6(32'h385d11bb),
	.w7(32'h38f3212b),
	.w8(32'h391b046e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368319d1),
	.w1(32'h393863d4),
	.w2(32'hb706ab86),
	.w3(32'hb918adcc),
	.w4(32'h3970c993),
	.w5(32'hb79fb542),
	.w6(32'h3947328a),
	.w7(32'h378767d8),
	.w8(32'h395b3ee2),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad4aac),
	.w1(32'hb9b78e68),
	.w2(32'hb99a3d49),
	.w3(32'h3886d7cb),
	.w4(32'hb9a7c039),
	.w5(32'hb9a2af09),
	.w6(32'hba0fe2e9),
	.w7(32'hba11d1d4),
	.w8(32'hba1df3a6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86ab2d9),
	.w1(32'hb8c7dca8),
	.w2(32'hba0324cf),
	.w3(32'h38ef5125),
	.w4(32'h3907760d),
	.w5(32'hb8f73b8d),
	.w6(32'h3a56d19a),
	.w7(32'h3910c240),
	.w8(32'hb7fb1ca3),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c40d04),
	.w1(32'h39f73642),
	.w2(32'hb9b74c75),
	.w3(32'h3a3fc569),
	.w4(32'h3981d1f6),
	.w5(32'h360ff5d3),
	.w6(32'h3a98b55d),
	.w7(32'h398ee56d),
	.w8(32'hb964e275),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387f6c7e),
	.w1(32'hb99519cf),
	.w2(32'hb985a5f1),
	.w3(32'h3980a172),
	.w4(32'hb652894d),
	.w5(32'h39a0c518),
	.w6(32'h39aed1e2),
	.w7(32'hb7cc7863),
	.w8(32'h3712368f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82e91d),
	.w1(32'h3a009f46),
	.w2(32'h39835f56),
	.w3(32'h3abace4f),
	.w4(32'h39eb6b6f),
	.w5(32'hb7e3b9a7),
	.w6(32'h3a4cc32a),
	.w7(32'h39c6fee6),
	.w8(32'hb93493dd),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da1d68),
	.w1(32'hb9af13b0),
	.w2(32'hb94bb2a8),
	.w3(32'h377bf6c9),
	.w4(32'hb99f9dc1),
	.w5(32'hb94c7c32),
	.w6(32'h38b5f038),
	.w7(32'hb8cf7f5e),
	.w8(32'h3881ac49),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb859dbc4),
	.w1(32'h37e70fb7),
	.w2(32'h3895f271),
	.w3(32'hb88761e4),
	.w4(32'hb8535b0d),
	.w5(32'hb8491afc),
	.w6(32'h38d34b17),
	.w7(32'h387c35cc),
	.w8(32'h38f8bb85),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49fd35),
	.w1(32'h3974f374),
	.w2(32'hb918ee30),
	.w3(32'h3a0be500),
	.w4(32'h3914a79a),
	.w5(32'hb925ad93),
	.w6(32'h39ab8ed6),
	.w7(32'h389ba0c8),
	.w8(32'hb9cdda75),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92752e6),
	.w1(32'hba13c5b4),
	.w2(32'hba15aad5),
	.w3(32'hb9141a16),
	.w4(32'hb99c9d10),
	.w5(32'hb9d2e87d),
	.w6(32'hb9b52372),
	.w7(32'hb9ac3f78),
	.w8(32'hb9cfb471),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97cb16b),
	.w1(32'h3925ea92),
	.w2(32'h39930900),
	.w3(32'hb821d423),
	.w4(32'h392c476d),
	.w5(32'hb763399a),
	.w6(32'h39b4bb9a),
	.w7(32'h39a0c5be),
	.w8(32'h39183ca1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3884a25c),
	.w1(32'hb7852292),
	.w2(32'h38582730),
	.w3(32'hb8fc6a0b),
	.w4(32'hb8ba3637),
	.w5(32'hb8a25370),
	.w6(32'h38e991f9),
	.w7(32'h38cbde22),
	.w8(32'h3920b2d5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d7d07c),
	.w1(32'hb937afc5),
	.w2(32'hb994a9ce),
	.w3(32'hb7d85ee3),
	.w4(32'hb918cc13),
	.w5(32'hb967587a),
	.w6(32'hb9481c67),
	.w7(32'hb8f25be1),
	.w8(32'h38a25d88),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f5d76),
	.w1(32'hb90c229f),
	.w2(32'hb937113f),
	.w3(32'hb98100cc),
	.w4(32'hb8871ce0),
	.w5(32'hb87dc4bd),
	.w6(32'hb7fc3823),
	.w7(32'hb89bf766),
	.w8(32'hb9129427),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a320372),
	.w1(32'h3a5ed882),
	.w2(32'hba0a4002),
	.w3(32'h3a874402),
	.w4(32'h3aa0493c),
	.w5(32'hb8c82a15),
	.w6(32'h3acb7b3d),
	.w7(32'h3a55119a),
	.w8(32'h3977ca65),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a581f77),
	.w1(32'h38ccf255),
	.w2(32'hb958dc36),
	.w3(32'h3a24fccd),
	.w4(32'h38971a1c),
	.w5(32'hb8ef668a),
	.w6(32'h39e079d4),
	.w7(32'hb8848467),
	.w8(32'hb93351c0),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a2d52),
	.w1(32'h396327f1),
	.w2(32'hba2e0536),
	.w3(32'h3a8db9a9),
	.w4(32'h39ef6c5f),
	.w5(32'hba0674d2),
	.w6(32'h3a4261da),
	.w7(32'h39ac0162),
	.w8(32'hb9b66821),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923468c),
	.w1(32'hb88a686c),
	.w2(32'hb72038b5),
	.w3(32'hb96251e8),
	.w4(32'hb8fa0081),
	.w5(32'hb8e10870),
	.w6(32'hb8c922a4),
	.w7(32'hb93e5b15),
	.w8(32'hb97cac46),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c4961),
	.w1(32'h38413e17),
	.w2(32'h390d432d),
	.w3(32'hb9848a54),
	.w4(32'hb8a493a5),
	.w5(32'hb88095ed),
	.w6(32'h3922dad2),
	.w7(32'h390ef697),
	.w8(32'h39701ffd),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396539da),
	.w1(32'hb8be3d6b),
	.w2(32'hb89ec057),
	.w3(32'h37128537),
	.w4(32'hb8e1afd4),
	.w5(32'hb9028d7f),
	.w6(32'hb8aa89d7),
	.w7(32'hb73c6085),
	.w8(32'h37635bc1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb39a3682),
	.w1(32'hb85eb25b),
	.w2(32'hb76827ac),
	.w3(32'hb9040e9d),
	.w4(32'hb8b67415),
	.w5(32'hb884113a),
	.w6(32'hb84ce8e7),
	.w7(32'hb8439c03),
	.w8(32'hb811a96a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57dc82),
	.w1(32'hb8abf04c),
	.w2(32'hba53b318),
	.w3(32'h39f5f7d1),
	.w4(32'h39bf289d),
	.w5(32'h3931ed37),
	.w6(32'h39d5ec83),
	.w7(32'hb968c264),
	.w8(32'hb9d6a634),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6e708),
	.w1(32'h38ba9ae2),
	.w2(32'hb8da4b3e),
	.w3(32'hb87b4f19),
	.w4(32'hb86e5994),
	.w5(32'hb8cf56b8),
	.w6(32'hb969a34a),
	.w7(32'hb955dbc3),
	.w8(32'hb9a262fa),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e16d97),
	.w1(32'hb92e92bd),
	.w2(32'h36b03c13),
	.w3(32'h393df6e7),
	.w4(32'hb88d4421),
	.w5(32'hb85be935),
	.w6(32'h39980405),
	.w7(32'h391eb613),
	.w8(32'hb942dd86),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393534a1),
	.w1(32'h39113ade),
	.w2(32'h39146aa7),
	.w3(32'h37c009bd),
	.w4(32'h394b7be7),
	.w5(32'h3912298e),
	.w6(32'hb8f45d33),
	.w7(32'hb89cae9c),
	.w8(32'hb9900a28),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b24837),
	.w1(32'hb8f3bf65),
	.w2(32'hb9176182),
	.w3(32'hb880b1e1),
	.w4(32'hb8b56c10),
	.w5(32'hb8ee4c5f),
	.w6(32'hb94e9d23),
	.w7(32'hb9347303),
	.w8(32'hb63a487a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c8e760),
	.w1(32'hba475277),
	.w2(32'hba952dc4),
	.w3(32'h3997dac9),
	.w4(32'hb8a591c0),
	.w5(32'hb8cea622),
	.w6(32'hb81e4bf6),
	.w7(32'hb8c6d595),
	.w8(32'hb99ca756),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f9951),
	.w1(32'hb998ec88),
	.w2(32'hb80ed3d6),
	.w3(32'hb9df2284),
	.w4(32'hb939c818),
	.w5(32'h38a215cf),
	.w6(32'hb9cc7e00),
	.w7(32'hb99a3412),
	.w8(32'hb95f087d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43c909),
	.w1(32'h3a18c030),
	.w2(32'h39643142),
	.w3(32'h3a674265),
	.w4(32'h3a0107b0),
	.w5(32'h3856cb05),
	.w6(32'h3aa3da91),
	.w7(32'h3a18d161),
	.w8(32'h39245764),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385515dc),
	.w1(32'hb86e1a52),
	.w2(32'hb700dbd9),
	.w3(32'hb86bc8f3),
	.w4(32'hb7df993a),
	.w5(32'h37bce223),
	.w6(32'h38382a42),
	.w7(32'h380e3327),
	.w8(32'h38c0aba9),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ddfa37),
	.w1(32'h36351752),
	.w2(32'hb97350bc),
	.w3(32'hba14fa21),
	.w4(32'hba5fb445),
	.w5(32'hb95e6096),
	.w6(32'hbac4d0fd),
	.w7(32'hbabec3d8),
	.w8(32'hba3ec9a2),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule