module layer_10_featuremap_382(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd81c90),
	.w1(32'h3b4a7f68),
	.w2(32'hbbafd758),
	.w3(32'hbbef7d6c),
	.w4(32'h3b74dd7d),
	.w5(32'hbb9f0bd5),
	.w6(32'hbb1c4d94),
	.w7(32'h3b4d5820),
	.w8(32'hbb6f1cc1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c1cc0),
	.w1(32'hbb990964),
	.w2(32'hbacfce8c),
	.w3(32'hbba85bbb),
	.w4(32'hbbd2ff99),
	.w5(32'h3b751d8d),
	.w6(32'hbafc9611),
	.w7(32'hba510511),
	.w8(32'h3b47a8f1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91d3a2),
	.w1(32'hbbb98104),
	.w2(32'hbc686b3e),
	.w3(32'h3b842963),
	.w4(32'hba4a346f),
	.w5(32'hbc6b6e2b),
	.w6(32'h3b86b202),
	.w7(32'h3c6c6f29),
	.w8(32'hbb911825),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989aa2c),
	.w1(32'h3c09911f),
	.w2(32'h3b91f922),
	.w3(32'hba1d3b63),
	.w4(32'h3c235c68),
	.w5(32'h3c7da161),
	.w6(32'hbc942b9f),
	.w7(32'h3adeada5),
	.w8(32'h3a84e3d5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd96cb4),
	.w1(32'h3aa1ecc0),
	.w2(32'h3bd8a067),
	.w3(32'h3bc80ad2),
	.w4(32'h3b593c20),
	.w5(32'h3bb82fde),
	.w6(32'h3a18003b),
	.w7(32'h3b1e1df5),
	.w8(32'h3a1c1553),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b037003),
	.w1(32'h398a1fd4),
	.w2(32'h3b025b8e),
	.w3(32'hbb4fe3a4),
	.w4(32'hbbd33928),
	.w5(32'hbb614da0),
	.w6(32'hba5fbdc8),
	.w7(32'hbbb4cbdb),
	.w8(32'hbc2a8c49),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a3a17),
	.w1(32'hbbb6e7b9),
	.w2(32'hbc9d5c89),
	.w3(32'h3a387f2e),
	.w4(32'hbbd9f4f4),
	.w5(32'h3ba74f46),
	.w6(32'h3aa3ada9),
	.w7(32'h3b61f874),
	.w8(32'h3a230c80),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26cc8a),
	.w1(32'hba6ed721),
	.w2(32'h3ae336a0),
	.w3(32'hbb3a8abe),
	.w4(32'h3c58757d),
	.w5(32'h3c79ad1c),
	.w6(32'hbc1ae824),
	.w7(32'h3c320122),
	.w8(32'h3a6d5d1f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18d625),
	.w1(32'hbc126803),
	.w2(32'hbc4bc332),
	.w3(32'h3b807bba),
	.w4(32'hbab0a3f1),
	.w5(32'h3ce672d1),
	.w6(32'hbbb2a40c),
	.w7(32'h3ba4b486),
	.w8(32'hbb82cb40),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dcde7),
	.w1(32'hbc00e190),
	.w2(32'hbbe85b6a),
	.w3(32'hbc5cafff),
	.w4(32'hbbb36f04),
	.w5(32'h3b4bd013),
	.w6(32'hbce00a7c),
	.w7(32'hbac3cf55),
	.w8(32'h3a977228),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ad84d),
	.w1(32'hbb96c390),
	.w2(32'h3acba629),
	.w3(32'h3a92d950),
	.w4(32'h3b8a5813),
	.w5(32'h3ae7118d),
	.w6(32'h3bc60400),
	.w7(32'h38132d3c),
	.w8(32'h3b1ab292),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2eefca),
	.w1(32'h3b2f77ff),
	.w2(32'hbc3b869f),
	.w3(32'h3b4fb139),
	.w4(32'hbb97b202),
	.w5(32'hbbb31b34),
	.w6(32'h3bcc03fe),
	.w7(32'hbb1e99d9),
	.w8(32'hbba229f4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb204601),
	.w1(32'h3b88fedc),
	.w2(32'hbbb00b95),
	.w3(32'h3b1b14da),
	.w4(32'hbb1696b4),
	.w5(32'h3c166607),
	.w6(32'hbb24eb00),
	.w7(32'h3b8c5e6f),
	.w8(32'hbba33176),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0f455),
	.w1(32'hbb180ebb),
	.w2(32'h3c0405f0),
	.w3(32'h3bb5b6bb),
	.w4(32'hbc354c40),
	.w5(32'hbbff54f9),
	.w6(32'h3bb4872d),
	.w7(32'hbc41a0d8),
	.w8(32'hbb9466b2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cf146),
	.w1(32'h3a6d70e7),
	.w2(32'hbbf73fc4),
	.w3(32'hbc9dee06),
	.w4(32'h3bda7d6b),
	.w5(32'hbc02caf5),
	.w6(32'hbc853985),
	.w7(32'h3b52b164),
	.w8(32'h3b135ee4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc147d37),
	.w1(32'hbc2ad6f4),
	.w2(32'hbc6502ea),
	.w3(32'hbb8f2449),
	.w4(32'hbc1197fb),
	.w5(32'hbb51058b),
	.w6(32'hbbb3bc33),
	.w7(32'h3a178ab0),
	.w8(32'h3a951097),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a986e10),
	.w1(32'h3b19b6da),
	.w2(32'h3b6e39ea),
	.w3(32'h3bd50422),
	.w4(32'hbaca67a5),
	.w5(32'h3b418fb1),
	.w6(32'h3c09e70a),
	.w7(32'hbbaf777e),
	.w8(32'h3b1ff114),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b228e2b),
	.w1(32'h3ae234ba),
	.w2(32'hbb1f16be),
	.w3(32'h3a9f2679),
	.w4(32'h3b82687e),
	.w5(32'hbba6e76c),
	.w6(32'h386c060e),
	.w7(32'h3bc8059b),
	.w8(32'hbc22f935),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa14d1f),
	.w1(32'hbbab1a31),
	.w2(32'hbc53b299),
	.w3(32'hbb4772a7),
	.w4(32'hbc3b5a27),
	.w5(32'h3be763b6),
	.w6(32'hbbe48bfc),
	.w7(32'hba758668),
	.w8(32'h3c3e08c9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fe4ee),
	.w1(32'hba6619dd),
	.w2(32'h3b787650),
	.w3(32'h3c2526fe),
	.w4(32'hbbf89606),
	.w5(32'hba8925b9),
	.w6(32'h3ab96d13),
	.w7(32'hbbb6fa11),
	.w8(32'h3b4e50ac),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb283875),
	.w1(32'h3b61f64c),
	.w2(32'h3a8e5391),
	.w3(32'hbb857137),
	.w4(32'h3b32d5a7),
	.w5(32'h3b54331d),
	.w6(32'hbbbe7269),
	.w7(32'hb9c63441),
	.w8(32'hbb9d9be7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92b4f4),
	.w1(32'h3b6e50e0),
	.w2(32'h3bebca69),
	.w3(32'h3b626002),
	.w4(32'h3a64d807),
	.w5(32'h39a40443),
	.w6(32'hbb1750b4),
	.w7(32'hba31b109),
	.w8(32'h3aceb4cc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c91b9),
	.w1(32'hbbb22941),
	.w2(32'hbc7a03c7),
	.w3(32'hbc42d6d2),
	.w4(32'hbb6c4a77),
	.w5(32'hbc1f5994),
	.w6(32'hbb3cb34f),
	.w7(32'h3b4459cb),
	.w8(32'hbbf808bf),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbe56d),
	.w1(32'hbc418bf8),
	.w2(32'hbc0d3e56),
	.w3(32'hbbd8ec32),
	.w4(32'hbb6e3e8b),
	.w5(32'hbb085525),
	.w6(32'hba3a2358),
	.w7(32'hbb69d478),
	.w8(32'hb98721c4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc157e93),
	.w1(32'hba4c22a6),
	.w2(32'hba2ea564),
	.w3(32'h3a424ed9),
	.w4(32'h3b3490be),
	.w5(32'h3c14ba1b),
	.w6(32'hbbcb5faa),
	.w7(32'h3be10583),
	.w8(32'hb9f2b414),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce1c1c),
	.w1(32'h3be32ee5),
	.w2(32'h3b52404f),
	.w3(32'hbc14259c),
	.w4(32'h3c03f1ec),
	.w5(32'hbb184ee9),
	.w6(32'hbc0e4888),
	.w7(32'h3b983545),
	.w8(32'hbb12a276),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae0dd5),
	.w1(32'hbab26f18),
	.w2(32'hbbb0290e),
	.w3(32'h3b6de877),
	.w4(32'hbb917877),
	.w5(32'h3c8591b4),
	.w6(32'h3b4ce87b),
	.w7(32'h3bc56c0f),
	.w8(32'h3b9c848b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ebead),
	.w1(32'hbba1cd66),
	.w2(32'hba225333),
	.w3(32'h3ae04548),
	.w4(32'hbb9161ad),
	.w5(32'h3aa94b4d),
	.w6(32'hbb6f1bbd),
	.w7(32'hbb32ac71),
	.w8(32'h3a9c49b2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cecd3),
	.w1(32'h394a0c5e),
	.w2(32'h3af2ba29),
	.w3(32'hba8de07a),
	.w4(32'h3b070e03),
	.w5(32'h3b4c3716),
	.w6(32'h3bb25cee),
	.w7(32'h3bd44b71),
	.w8(32'hba741c35),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0171d7),
	.w1(32'h3b70dd3e),
	.w2(32'h3b7864bd),
	.w3(32'hbc77d2b7),
	.w4(32'h3bb564ee),
	.w5(32'h3a989508),
	.w6(32'hbc22bc5e),
	.w7(32'h3aff7dbc),
	.w8(32'hbbe8c163),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae59621),
	.w1(32'h3ac45694),
	.w2(32'h3b27a8c2),
	.w3(32'hbba81616),
	.w4(32'hbaa0340c),
	.w5(32'h3b8e368a),
	.w6(32'hbbe3ac2e),
	.w7(32'hbadaad07),
	.w8(32'hbb641f57),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b0611),
	.w1(32'hbc06c065),
	.w2(32'hbc84a1a2),
	.w3(32'h3b62dc74),
	.w4(32'hbc1d1cd9),
	.w5(32'hbc888289),
	.w6(32'hbaf49c9f),
	.w7(32'hbc03495c),
	.w8(32'hbc8d33f7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb76d1a),
	.w1(32'hbba6f8a6),
	.w2(32'hbbbfaf8b),
	.w3(32'hbbb2a181),
	.w4(32'hbc15a6c3),
	.w5(32'hbbc559c0),
	.w6(32'hbb52fe45),
	.w7(32'h3b6a7a7f),
	.w8(32'hbb16be15),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b0829),
	.w1(32'hbb5c7b67),
	.w2(32'hbb2dcfe0),
	.w3(32'hbbf60cab),
	.w4(32'hbb407df9),
	.w5(32'h3a3bed59),
	.w6(32'hba85035b),
	.w7(32'h3bac5eaf),
	.w8(32'h3b07840d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa74f57),
	.w1(32'h3bc45ed6),
	.w2(32'hbc0fe6eb),
	.w3(32'hba99e1d9),
	.w4(32'hbc8e3d2e),
	.w5(32'hbc9e4893),
	.w6(32'h3baebdfe),
	.w7(32'hbc523cc2),
	.w8(32'hbc18c2f9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdacee0),
	.w1(32'h39df1780),
	.w2(32'hbb56aa6e),
	.w3(32'hbbd9f30d),
	.w4(32'hb8b4f534),
	.w5(32'h3ba376f3),
	.w6(32'h3c63bd45),
	.w7(32'h3be2bde9),
	.w8(32'hbadc5ac3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2e71b),
	.w1(32'hbb3adf74),
	.w2(32'hba0daac6),
	.w3(32'hbc3eb786),
	.w4(32'hbb645130),
	.w5(32'h3c0b46c6),
	.w6(32'hbc209445),
	.w7(32'h3b6b5dbf),
	.w8(32'hba4b8b3c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b6ad3),
	.w1(32'hbba50369),
	.w2(32'hbb942f8e),
	.w3(32'h3a5b61c8),
	.w4(32'hb9f5cfeb),
	.w5(32'h3ba75ca9),
	.w6(32'hbc8cc3c1),
	.w7(32'hbac77094),
	.w8(32'h3ba925ac),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37ab8c),
	.w1(32'hbb714341),
	.w2(32'hbb4c53bd),
	.w3(32'h3c09769b),
	.w4(32'hbc11bbe4),
	.w5(32'hbb8529e1),
	.w6(32'hba630763),
	.w7(32'hbc334b70),
	.w8(32'h3ad7263a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b8708),
	.w1(32'hbb67e131),
	.w2(32'h3abc2233),
	.w3(32'h3ade072b),
	.w4(32'h3991110d),
	.w5(32'h3b910c0e),
	.w6(32'hbadb3f7e),
	.w7(32'hb9c0cdaa),
	.w8(32'h3b6801c1),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0bdf6),
	.w1(32'h3b92c2f8),
	.w2(32'h3c2f7c42),
	.w3(32'h3b0b1e99),
	.w4(32'h3ccb744a),
	.w5(32'hbc2622d7),
	.w6(32'h3b87a842),
	.w7(32'hbc10dc45),
	.w8(32'hbcc001e6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d0449),
	.w1(32'hba107f9d),
	.w2(32'hbb364cab),
	.w3(32'hbcb6511f),
	.w4(32'h3b7da9cf),
	.w5(32'h3bfd3588),
	.w6(32'hbc96454a),
	.w7(32'hbb7a8b53),
	.w8(32'hbba74404),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35eae9),
	.w1(32'hbb87c4ff),
	.w2(32'hbb5c62f6),
	.w3(32'h3b2c7442),
	.w4(32'hbb457f4b),
	.w5(32'h3bc18540),
	.w6(32'hbc0f0fe4),
	.w7(32'hbaf7bd46),
	.w8(32'hbbf21d11),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5edc30),
	.w1(32'hb9deaeca),
	.w2(32'hbc5927ea),
	.w3(32'hbc320c84),
	.w4(32'hbb10afd0),
	.w5(32'hbc3090e8),
	.w6(32'hbbbaa4d9),
	.w7(32'h3afcdbe9),
	.w8(32'hb89c5c41),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb942bcb),
	.w1(32'hbc24aa8f),
	.w2(32'hb9947d3e),
	.w3(32'hbb38dc9d),
	.w4(32'hb9f8bdb5),
	.w5(32'h3d129da3),
	.w6(32'h38974de9),
	.w7(32'h3c4f119f),
	.w8(32'h3c6494be),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb819135),
	.w1(32'hbc419f60),
	.w2(32'hbbf88632),
	.w3(32'hbaff2a04),
	.w4(32'h3b15ded2),
	.w5(32'h3ba74a20),
	.w6(32'hbbaa3650),
	.w7(32'h3b88814f),
	.w8(32'hbc0176d7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe37a09),
	.w1(32'h3ab6db6f),
	.w2(32'hbbf02978),
	.w3(32'hbbff66a0),
	.w4(32'hba7164f6),
	.w5(32'hbbbd5fce),
	.w6(32'hbb9cf2aa),
	.w7(32'h3b19bcc0),
	.w8(32'hbb991ae7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4a946),
	.w1(32'hbab57c06),
	.w2(32'hbb45791f),
	.w3(32'hbb3bb0a3),
	.w4(32'h39016f3f),
	.w5(32'h3ba5b7d0),
	.w6(32'h3bb0a79e),
	.w7(32'h3a0745d1),
	.w8(32'h3b4c75be),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba870c25),
	.w1(32'h3c126e23),
	.w2(32'h3c66230b),
	.w3(32'hba85e016),
	.w4(32'h3c8b278b),
	.w5(32'h3c939717),
	.w6(32'h3a91da4e),
	.w7(32'h3ba4a2f4),
	.w8(32'hbbb37ddc),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb57012),
	.w1(32'h3b876742),
	.w2(32'hbc88b18f),
	.w3(32'h3b26dbe4),
	.w4(32'hbbc48289),
	.w5(32'hbce1d1ee),
	.w6(32'hb98345eb),
	.w7(32'hbc4d410f),
	.w8(32'hbce316bd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fcb09),
	.w1(32'h3a3c3dda),
	.w2(32'hbc01c935),
	.w3(32'hbc119e95),
	.w4(32'h3b3065b7),
	.w5(32'hbbb68c5b),
	.w6(32'h3a5f4fe1),
	.w7(32'h3bc227bb),
	.w8(32'hbbba6194),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd1127),
	.w1(32'hbc15414b),
	.w2(32'hbc159167),
	.w3(32'hbaa030b1),
	.w4(32'hbc224bb0),
	.w5(32'hbb959061),
	.w6(32'h3b1ef4fe),
	.w7(32'hbbd585b0),
	.w8(32'h3bd71a9c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5e313),
	.w1(32'h3b33b755),
	.w2(32'h3bdea3dc),
	.w3(32'hbbe1cfa0),
	.w4(32'h3a8d0191),
	.w5(32'hba543df7),
	.w6(32'hbb86bb00),
	.w7(32'h39f5f21e),
	.w8(32'hbbb0ed12),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb857367),
	.w1(32'h3a2a43ec),
	.w2(32'hbc25386d),
	.w3(32'hbc2757d3),
	.w4(32'hbbdc2175),
	.w5(32'hbc6906cd),
	.w6(32'h3a92a1fb),
	.w7(32'h3b96e9eb),
	.w8(32'hbaddc2d7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09b8dd),
	.w1(32'h392bf018),
	.w2(32'hba1ce602),
	.w3(32'hbb1c5d47),
	.w4(32'hba920b12),
	.w5(32'h3b0a106d),
	.w6(32'h3b41ba9f),
	.w7(32'h3a900396),
	.w8(32'h3b6bdb62),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb385a1c),
	.w1(32'h3b1e0a63),
	.w2(32'h3bf874e0),
	.w3(32'hbacccce0),
	.w4(32'hbb504075),
	.w5(32'h3b977559),
	.w6(32'h3ae1a21e),
	.w7(32'h3b409dc3),
	.w8(32'h3b623119),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a97d5f),
	.w1(32'hbae20433),
	.w2(32'hbbd08a30),
	.w3(32'hbbcc5df5),
	.w4(32'h3ab3776d),
	.w5(32'hbbffe996),
	.w6(32'hbb82a1ef),
	.w7(32'hbb8121a2),
	.w8(32'hbaa610ab),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacc8e1),
	.w1(32'h3beb331f),
	.w2(32'h3bac0b9d),
	.w3(32'h3bd182c0),
	.w4(32'h3aaf378e),
	.w5(32'h3acfde11),
	.w6(32'h3bd329e8),
	.w7(32'h3bb6d1e9),
	.w8(32'hbb5b0c8b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f013d),
	.w1(32'hbba937f5),
	.w2(32'hbbfeca24),
	.w3(32'hbb199733),
	.w4(32'hbc14fdb4),
	.w5(32'hbc506f6c),
	.w6(32'hbb52655e),
	.w7(32'hbbfd6869),
	.w8(32'hba9fd176),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf581e5),
	.w1(32'hbaf5f6a2),
	.w2(32'h3bdd80f7),
	.w3(32'hbaf629a0),
	.w4(32'h3a953958),
	.w5(32'hbb34d37f),
	.w6(32'h3a3ed98c),
	.w7(32'hbc066070),
	.w8(32'h382582a4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb121e8),
	.w1(32'h3abeb87f),
	.w2(32'hbadbe4fa),
	.w3(32'hbb1bc964),
	.w4(32'h3bfa2591),
	.w5(32'hbb49b05d),
	.w6(32'hba88a2dc),
	.w7(32'hbbb7a0bc),
	.w8(32'hbc058d8b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2853a9),
	.w1(32'hbb25a589),
	.w2(32'hbbf417b5),
	.w3(32'hbb9eb0b7),
	.w4(32'hbb3b16f7),
	.w5(32'h3912cb22),
	.w6(32'hbb92c29a),
	.w7(32'h3b32ea63),
	.w8(32'hba88fd0a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1255),
	.w1(32'hb957fb32),
	.w2(32'hbb6bcb16),
	.w3(32'hbb5841a6),
	.w4(32'hbb72962e),
	.w5(32'hbab32a61),
	.w6(32'hb992a10c),
	.w7(32'hbbe1c14b),
	.w8(32'hbb7f2d4b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb908295),
	.w1(32'hba9303c0),
	.w2(32'hbb482364),
	.w3(32'hbbe93d1a),
	.w4(32'hbb4ce8b4),
	.w5(32'hbba515b8),
	.w6(32'hbb5d13dd),
	.w7(32'hbb74bc98),
	.w8(32'h3acd7b38),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf322e),
	.w1(32'hbac24031),
	.w2(32'hbac551b3),
	.w3(32'h3af52046),
	.w4(32'h3aaac701),
	.w5(32'h3af6b3f8),
	.w6(32'h3ad42e00),
	.w7(32'h3b3286be),
	.w8(32'h3ba14a29),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5aeabd),
	.w1(32'h3b9297e8),
	.w2(32'h3b5203a3),
	.w3(32'h3bb7d488),
	.w4(32'h3ba3421f),
	.w5(32'h3c58702b),
	.w6(32'h3c319b26),
	.w7(32'h3b9834f9),
	.w8(32'h39da8918),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0956d9),
	.w1(32'hbb68f238),
	.w2(32'hbbb6ac3e),
	.w3(32'h3c0affd5),
	.w4(32'hbb3ec89f),
	.w5(32'h3b70872b),
	.w6(32'hbb0c4bad),
	.w7(32'hba846a0b),
	.w8(32'hbb0d0ef3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65593a),
	.w1(32'hbba202cb),
	.w2(32'hbb9d0b4e),
	.w3(32'h3b691a34),
	.w4(32'hbb4bdbb3),
	.w5(32'h3b03de7d),
	.w6(32'hbb5835fe),
	.w7(32'h3c0e91d4),
	.w8(32'hbc9717ad),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93ef11),
	.w1(32'h3b89a74b),
	.w2(32'hbb8d4d57),
	.w3(32'hbc237ab0),
	.w4(32'hbaf18961),
	.w5(32'h3b085d11),
	.w6(32'hbbd53d22),
	.w7(32'h3abd2920),
	.w8(32'h3b203679),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97817c),
	.w1(32'hbb83754c),
	.w2(32'hbb43cd3e),
	.w3(32'hbc3dfd67),
	.w4(32'h3af18162),
	.w5(32'h3a3da1b7),
	.w6(32'hbc39ef57),
	.w7(32'h3a6ae005),
	.w8(32'h3a6167de),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385b80b4),
	.w1(32'h35c60093),
	.w2(32'h370d7a6f),
	.w3(32'h3803a46e),
	.w4(32'hb817df23),
	.w5(32'hb7d78faf),
	.w6(32'h38429871),
	.w7(32'hb72ec690),
	.w8(32'h371b6585),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eb8938),
	.w1(32'h387c817a),
	.w2(32'h38880423),
	.w3(32'h3699679b),
	.w4(32'h37611aab),
	.w5(32'h37813c76),
	.w6(32'h38048a06),
	.w7(32'h384ffb03),
	.w8(32'h3889044d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3802e0c5),
	.w1(32'h38886a88),
	.w2(32'h3899e375),
	.w3(32'hb509a2e3),
	.w4(32'hb792762c),
	.w5(32'hb8a051c1),
	.w6(32'h3829dbd8),
	.w7(32'h36faa51e),
	.w8(32'hb8ed963b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82c520),
	.w1(32'h3989a771),
	.w2(32'hbabf53ac),
	.w3(32'h3a4ca62f),
	.w4(32'h3869b0ed),
	.w5(32'hba127216),
	.w6(32'h3a2e81ac),
	.w7(32'hba3e9714),
	.w8(32'hbadca972),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8afbd60),
	.w1(32'hb8959961),
	.w2(32'hb869100f),
	.w3(32'h3763f152),
	.w4(32'hb7712901),
	.w5(32'hb8141989),
	.w6(32'h3928fdfa),
	.w7(32'h38deed39),
	.w8(32'h38c008ca),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b262079),
	.w1(32'h3a8065a0),
	.w2(32'hba712d3d),
	.w3(32'h3a2e842d),
	.w4(32'h3a1e7956),
	.w5(32'hbac69111),
	.w6(32'h3a306a3e),
	.w7(32'h39348910),
	.w8(32'hba9f9dc7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc3f60),
	.w1(32'h3a10da3a),
	.w2(32'hbb88effe),
	.w3(32'h3a9a43fe),
	.w4(32'h3ad84ae2),
	.w5(32'hbb1494df),
	.w6(32'h3a969484),
	.w7(32'h3a4ea1f5),
	.w8(32'hbb12167d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26d3a1),
	.w1(32'h3a65768f),
	.w2(32'hba9063b6),
	.w3(32'hbaf272ca),
	.w4(32'h3b239c0d),
	.w5(32'h36b6dd22),
	.w6(32'hbac61f51),
	.w7(32'h3b26449c),
	.w8(32'h3a11ece2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fa0f2),
	.w1(32'hbb20576b),
	.w2(32'hbb83b997),
	.w3(32'hbb28cdec),
	.w4(32'hbad96f63),
	.w5(32'hbb2ee608),
	.w6(32'hba8fb461),
	.w7(32'hbaf961fe),
	.w8(32'hbb926c2e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b9a93),
	.w1(32'h3ac0c034),
	.w2(32'hbb0ed829),
	.w3(32'h3a3486ac),
	.w4(32'hba34429d),
	.w5(32'hbaff5752),
	.w6(32'h39107ef9),
	.w7(32'hb99d53ba),
	.w8(32'hbaa53f0e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56fd62),
	.w1(32'hbaf11ce7),
	.w2(32'hbb02385b),
	.w3(32'hbb36df5d),
	.w4(32'hba4812ca),
	.w5(32'hba8c0b13),
	.w6(32'hbb166b1e),
	.w7(32'hb988567f),
	.w8(32'hba30b8dc),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d4ac5),
	.w1(32'h3b08f603),
	.w2(32'hba9a7cff),
	.w3(32'h3a8eaafa),
	.w4(32'h3a25d799),
	.w5(32'hbaf6ccb9),
	.w6(32'h3b1e4b1d),
	.w7(32'h3aa83598),
	.w8(32'hbaba9269),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f6bbe8),
	.w1(32'h37cbfeac),
	.w2(32'h38b11b27),
	.w3(32'hb8b521f6),
	.w4(32'h37ce5cc2),
	.w5(32'h389896f1),
	.w6(32'hb771c55d),
	.w7(32'h38aa26d9),
	.w8(32'h3909714a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e6e971),
	.w1(32'h36867554),
	.w2(32'hb7934c1c),
	.w3(32'h36c08bc5),
	.w4(32'h37c980c8),
	.w5(32'hb7e91b0b),
	.w6(32'h37c4f419),
	.w7(32'h37a40c13),
	.w8(32'hb5ccfa25),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3736bc34),
	.w1(32'hb832d195),
	.w2(32'h3726e96d),
	.w3(32'h384ff96a),
	.w4(32'hb791f8e9),
	.w5(32'h3799d7ac),
	.w6(32'h37b259b1),
	.w7(32'h3632fdcc),
	.w8(32'hb701a957),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993a480),
	.w1(32'h39839106),
	.w2(32'h3a08792f),
	.w3(32'hb9b4e2cc),
	.w4(32'hb89af09e),
	.w5(32'h3961d420),
	.w6(32'hb9fa7888),
	.w7(32'hb880ba46),
	.w8(32'h39b84c48),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba64546),
	.w1(32'hbb25026e),
	.w2(32'hbaaa9dd7),
	.w3(32'hbb1ffdf0),
	.w4(32'h391b56c7),
	.w5(32'h3a208ccb),
	.w6(32'hbb2d515f),
	.w7(32'hba2eb65b),
	.w8(32'hba1910a9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff0f88),
	.w1(32'h3a7a0af8),
	.w2(32'h3aa0b6dc),
	.w3(32'h3997c416),
	.w4(32'h3a253f78),
	.w5(32'h3a688961),
	.w6(32'h389fb996),
	.w7(32'h3a258b0e),
	.w8(32'h3a75155e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd449b9),
	.w1(32'hbb739727),
	.w2(32'hbab1992b),
	.w3(32'hbb86150e),
	.w4(32'hb857584e),
	.w5(32'hbacc8f37),
	.w6(32'hbac17b5f),
	.w7(32'h3a849ac5),
	.w8(32'hbae6768f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18c5be),
	.w1(32'hb9270516),
	.w2(32'hbb1d2aba),
	.w3(32'h39d76814),
	.w4(32'h3a7f0449),
	.w5(32'hba55cfb9),
	.w6(32'hb9b68281),
	.w7(32'h3a379be4),
	.w8(32'hbac5c292),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c15c1),
	.w1(32'h3b159b56),
	.w2(32'h3b8687e0),
	.w3(32'hbb264859),
	.w4(32'h3a8a550c),
	.w5(32'h3b30cccf),
	.w6(32'hbb3da0ec),
	.w7(32'h3a487192),
	.w8(32'h3b80d9fc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8040f),
	.w1(32'hbb3f863d),
	.w2(32'hbc2fa808),
	.w3(32'hbbbabafd),
	.w4(32'hbb1a9dcc),
	.w5(32'hbc118267),
	.w6(32'hbb231667),
	.w7(32'hbaf5c56f),
	.w8(32'hbbaab2ca),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36b632),
	.w1(32'h3b59636e),
	.w2(32'h3b83caf0),
	.w3(32'h3a7bc2e8),
	.w4(32'h3b325f79),
	.w5(32'h3b57868b),
	.w6(32'hbaf18208),
	.w7(32'h3aaf2147),
	.w8(32'h3afb6c86),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47a486),
	.w1(32'hbc145e82),
	.w2(32'hbbe84e1e),
	.w3(32'hbc0ee19e),
	.w4(32'hbb9b9cf4),
	.w5(32'hba986238),
	.w6(32'hbbb301ec),
	.w7(32'hbb62893e),
	.w8(32'hbbaca373),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b14b5),
	.w1(32'hb9270a1f),
	.w2(32'hbb24902d),
	.w3(32'hba9143b1),
	.w4(32'hb9a9b04f),
	.w5(32'hba994361),
	.w6(32'hba9bba5b),
	.w7(32'h3a9048f5),
	.w8(32'h3a267d71),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8f825),
	.w1(32'hba83f398),
	.w2(32'h3b085b21),
	.w3(32'hbb9bc6d4),
	.w4(32'h39255a25),
	.w5(32'h3b4bfdeb),
	.w6(32'hbb6dc5e9),
	.w7(32'h3ab83910),
	.w8(32'h3b9beee4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada8e0f),
	.w1(32'h39e1c87e),
	.w2(32'hba822f14),
	.w3(32'h3b0f3208),
	.w4(32'h3a9e0b1b),
	.w5(32'hb9aed1a5),
	.w6(32'h3a921790),
	.w7(32'h3834c0ec),
	.w8(32'hba6c3f92),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba90d8),
	.w1(32'hba2b4a85),
	.w2(32'hbba9dfd6),
	.w3(32'hbb7b9629),
	.w4(32'h3afbbb93),
	.w5(32'hbb300aae),
	.w6(32'hba947183),
	.w7(32'h3b14f9b9),
	.w8(32'hbb788932),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbc4d1),
	.w1(32'h3b24d4a9),
	.w2(32'hba050e82),
	.w3(32'h3ad652d7),
	.w4(32'hb9a812ca),
	.w5(32'hbaa871ae),
	.w6(32'h3af5e188),
	.w7(32'hba93a974),
	.w8(32'hbb0a587b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cce68),
	.w1(32'hbb8f31b8),
	.w2(32'hbbeddf75),
	.w3(32'hbb131669),
	.w4(32'hbaf3f2d3),
	.w5(32'hbb8d7ed0),
	.w6(32'h3bafa659),
	.w7(32'h3b88cb68),
	.w8(32'h3a710f22),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcceef74),
	.w1(32'hbba7954d),
	.w2(32'h399ac86e),
	.w3(32'hbc9fc385),
	.w4(32'h3a4d81be),
	.w5(32'h3baa203e),
	.w6(32'hbc44bc55),
	.w7(32'h3ba405ea),
	.w8(32'h3c160596),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e955a),
	.w1(32'hbb42f790),
	.w2(32'hba8d6960),
	.w3(32'hbbb96c72),
	.w4(32'h3b50a8a0),
	.w5(32'hb9648c6a),
	.w6(32'hbb43668b),
	.w7(32'h3b87d787),
	.w8(32'h39a12226),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47238b),
	.w1(32'hbb240d86),
	.w2(32'hbbdd4ab8),
	.w3(32'hbbccd38a),
	.w4(32'hbb0fb216),
	.w5(32'hbc02c2ee),
	.w6(32'hbac92ab3),
	.w7(32'h3a8ecbdd),
	.w8(32'hbbe3d744),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b481ee),
	.w1(32'h3b2f2d08),
	.w2(32'h3941ffa1),
	.w3(32'h398cbfc7),
	.w4(32'h3b4f9628),
	.w5(32'h3a20c1a0),
	.w6(32'h3a905a1a),
	.w7(32'h3b108f44),
	.w8(32'h3a83c8c0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d6489),
	.w1(32'hbb626c13),
	.w2(32'hbb6c7b23),
	.w3(32'hbbaf453e),
	.w4(32'h3a47f7e2),
	.w5(32'hbb1b6926),
	.w6(32'h3a1b0b1d),
	.w7(32'hba9027ca),
	.w8(32'hba901624),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2925bc),
	.w1(32'h3a84a9d3),
	.w2(32'hbb0db3fd),
	.w3(32'hba05af0f),
	.w4(32'h39ab3f97),
	.w5(32'hbb664fd9),
	.w6(32'h3abb94dc),
	.w7(32'h3a2a0f0a),
	.w8(32'hba916dfd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a415f),
	.w1(32'h3989145f),
	.w2(32'h3931b972),
	.w3(32'h3974d6de),
	.w4(32'h366926bc),
	.w5(32'hb66f2854),
	.w6(32'h38b24aa4),
	.w7(32'hb828ec0c),
	.w8(32'hb6cbae87),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad26181),
	.w1(32'hbaa25c16),
	.w2(32'hbb2ec1ba),
	.w3(32'hb9518825),
	.w4(32'hba116834),
	.w5(32'hbad49257),
	.w6(32'hba3dcce8),
	.w7(32'hb83bb562),
	.w8(32'hb94639c5),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb132f91),
	.w1(32'h3b19245b),
	.w2(32'hba13ed5e),
	.w3(32'hbacefca9),
	.w4(32'h3b1a59b7),
	.w5(32'hba97c11f),
	.w6(32'h399e3789),
	.w7(32'h3b1e9241),
	.w8(32'hba568a76),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ea36e),
	.w1(32'h3943ec4a),
	.w2(32'hbaf8a245),
	.w3(32'hb9de5aeb),
	.w4(32'h3b7b196e),
	.w5(32'h3a9ef428),
	.w6(32'h39784d48),
	.w7(32'h3b9a0587),
	.w8(32'h3b1f6b41),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbb7e2),
	.w1(32'hba9fcf2f),
	.w2(32'hb8fa5944),
	.w3(32'hbbd3ab0e),
	.w4(32'h3998da3d),
	.w5(32'h3b172c63),
	.w6(32'hbb805094),
	.w7(32'h3a95ef63),
	.w8(32'h3b910c00),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8bab1),
	.w1(32'hbb6a80fb),
	.w2(32'hba504dbf),
	.w3(32'hbb8e1660),
	.w4(32'hba20fb25),
	.w5(32'h396bae17),
	.w6(32'hbb330c7f),
	.w7(32'hba6749ea),
	.w8(32'hba28ad63),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a1126),
	.w1(32'h3b19a0fb),
	.w2(32'hb9b3088e),
	.w3(32'h3739e4b2),
	.w4(32'h3b056448),
	.w5(32'h3a8aeee1),
	.w6(32'h39ea3da4),
	.w7(32'h3b05f057),
	.w8(32'hba2b89f9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d1284),
	.w1(32'hbb50ee1d),
	.w2(32'hbbd2d304),
	.w3(32'hbb484110),
	.w4(32'hbadc6d26),
	.w5(32'hbb22fb6a),
	.w6(32'hbb851f77),
	.w7(32'hba56a6e0),
	.w8(32'hbae82fb6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb120b43),
	.w1(32'hb9a56629),
	.w2(32'hba34f04d),
	.w3(32'hbab546d6),
	.w4(32'h3a4d2033),
	.w5(32'hba179ae5),
	.w6(32'hb9d2ef6c),
	.w7(32'h3abe7fec),
	.w8(32'hba0f6742),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98443c2),
	.w1(32'hb91fb3e8),
	.w2(32'hb9bff47a),
	.w3(32'hb9eefd2f),
	.w4(32'hb99f404f),
	.w5(32'hb98fa287),
	.w6(32'hba038bd1),
	.w7(32'hb9d7e482),
	.w8(32'hb77ba4d2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a91d8),
	.w1(32'hba6ae082),
	.w2(32'hba4a3add),
	.w3(32'hb9e60573),
	.w4(32'hb9ca8d1f),
	.w5(32'hba0e3dcf),
	.w6(32'hb9a95b1c),
	.w7(32'hba300c97),
	.w8(32'hba281edd),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89b0518),
	.w1(32'hb854a7d6),
	.w2(32'hb7cdb5c3),
	.w3(32'hb736abbb),
	.w4(32'hb83c5157),
	.w5(32'h388b1b62),
	.w6(32'h3810a049),
	.w7(32'h37f6786c),
	.w8(32'h3875b75c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad428cf),
	.w1(32'h3ab2fc2f),
	.w2(32'h3a3decf8),
	.w3(32'h3a8b0240),
	.w4(32'h3a2c1a3d),
	.w5(32'h3a2baf83),
	.w6(32'h3a20ade8),
	.w7(32'h3a1fed39),
	.w8(32'h3945d5c4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba77abb),
	.w1(32'hba5cc331),
	.w2(32'hbb169a32),
	.w3(32'hbb5ffcb6),
	.w4(32'h3b0aff49),
	.w5(32'hb9c01247),
	.w6(32'hbadfcf49),
	.w7(32'h3b3550cb),
	.w8(32'h399ef095),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba253ee8),
	.w1(32'hba3be3aa),
	.w2(32'hbb184b45),
	.w3(32'hba1e33f7),
	.w4(32'hba16e78d),
	.w5(32'hbaa9bd7a),
	.w6(32'hba619f67),
	.w7(32'hba326e67),
	.w8(32'hba80c33e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7543b9),
	.w1(32'h3acb979a),
	.w2(32'hba4606b4),
	.w3(32'hb882524c),
	.w4(32'h3a9d59c3),
	.w5(32'hba2ea3da),
	.w6(32'h392d838f),
	.w7(32'h3a5721e5),
	.w8(32'hbad331cf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca9708),
	.w1(32'hbb773fee),
	.w2(32'hbaa04972),
	.w3(32'hbb843e79),
	.w4(32'hbac39fb4),
	.w5(32'h3aa82806),
	.w6(32'hbb960bfc),
	.w7(32'hbb2a9a63),
	.w8(32'h3a424375),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387bd522),
	.w1(32'hb7152e5b),
	.w2(32'h36ccf2ab),
	.w3(32'h388b0aa3),
	.w4(32'h370f6272),
	.w5(32'h3835b6ca),
	.w6(32'h38afb116),
	.w7(32'h38304919),
	.w8(32'h3809ee85),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394bf680),
	.w1(32'h397609b7),
	.w2(32'h390c5dab),
	.w3(32'h39532bd1),
	.w4(32'h391bf5ba),
	.w5(32'h3864d5e1),
	.w6(32'h39474f55),
	.w7(32'h393c1e5f),
	.w8(32'h3908ab5e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70a640f),
	.w1(32'h386fffcf),
	.w2(32'h38dccc2b),
	.w3(32'hb791c24a),
	.w4(32'h37438cdd),
	.w5(32'h387ed7c6),
	.w6(32'h3866b660),
	.w7(32'h38fdd64a),
	.w8(32'h39090154),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980f7d0),
	.w1(32'h3a3469a1),
	.w2(32'h3a37ce1b),
	.w3(32'h39c3694f),
	.w4(32'h3a919240),
	.w5(32'h39a50617),
	.w6(32'h3a20bcb6),
	.w7(32'h3a7374e5),
	.w8(32'h39ce16ed),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d70543),
	.w1(32'hbb20d875),
	.w2(32'hbbf16b2b),
	.w3(32'h39ec34f8),
	.w4(32'hbba9158f),
	.w5(32'hbbd80434),
	.w6(32'h3b9efa84),
	.w7(32'h39ea5975),
	.w8(32'hbbcddd95),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac35b38),
	.w1(32'hbae79676),
	.w2(32'hbbc2c5e0),
	.w3(32'hbb1d04d1),
	.w4(32'hbad75e90),
	.w5(32'hbb88f8cc),
	.w6(32'hba016336),
	.w7(32'h3ab6cce2),
	.w8(32'hbb3fd141),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5233e6),
	.w1(32'h36781342),
	.w2(32'hba0bb506),
	.w3(32'h39c81ad9),
	.w4(32'h3885aff5),
	.w5(32'hb91c0972),
	.w6(32'h39e7fb83),
	.w7(32'h38ef8bda),
	.w8(32'hb8a55b69),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb041bcf),
	.w1(32'hbab3f02d),
	.w2(32'hbaaf6cbb),
	.w3(32'hba09c5ac),
	.w4(32'hb826418e),
	.w5(32'hb9af01a8),
	.w6(32'hba3e5d12),
	.w7(32'hbab90add),
	.w8(32'hbaff077c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cbb74),
	.w1(32'hb9c32749),
	.w2(32'hb9aeed7c),
	.w3(32'hba3a5e3c),
	.w4(32'h3a09384a),
	.w5(32'h3a279f02),
	.w6(32'hba266b56),
	.w7(32'h3a2214cd),
	.w8(32'h3a154087),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34684f),
	.w1(32'hbab09a05),
	.w2(32'hbb13c719),
	.w3(32'hbb205f5e),
	.w4(32'hb93e37e6),
	.w5(32'hb9efd30f),
	.w6(32'hba91c1e5),
	.w7(32'h39d18816),
	.w8(32'hba433072),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69e8eb),
	.w1(32'hbb5a6c08),
	.w2(32'hbb7bba70),
	.w3(32'hbaab901d),
	.w4(32'hbaa1c4c6),
	.w5(32'hba533035),
	.w6(32'hbab91aae),
	.w7(32'hb9035c6a),
	.w8(32'hbaa32a78),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad37a3b),
	.w1(32'h39eb26d9),
	.w2(32'hbb86dd97),
	.w3(32'hba17c61f),
	.w4(32'hbaa64a67),
	.w5(32'hbb617442),
	.w6(32'hb9c4eb5c),
	.w7(32'hb8bb1bc5),
	.w8(32'hbb65ce4e),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a60d1),
	.w1(32'hba6f9311),
	.w2(32'h39928560),
	.w3(32'hbb4fe35a),
	.w4(32'h3a8e76c1),
	.w5(32'h3a92bc7e),
	.w6(32'hbb1ddbd2),
	.w7(32'h3a8883e9),
	.w8(32'h3a8c9628),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb255316),
	.w1(32'hbaa921c3),
	.w2(32'hbb817d00),
	.w3(32'hbb5aa51a),
	.w4(32'hb9accae2),
	.w5(32'hbac61364),
	.w6(32'hbb074303),
	.w7(32'h3986da4b),
	.w8(32'hba653ac0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c3a75),
	.w1(32'h3a094f8c),
	.w2(32'hbb7b54d7),
	.w3(32'hba359c28),
	.w4(32'h3a205b0f),
	.w5(32'hbb834bc7),
	.w6(32'h399d413a),
	.w7(32'h3acbe5f0),
	.w8(32'hbb969ad5),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ff12b),
	.w1(32'hb94574c2),
	.w2(32'hba2e3927),
	.w3(32'hb9a7ede2),
	.w4(32'h3afb8d93),
	.w5(32'h3a269240),
	.w6(32'hba23e2d1),
	.w7(32'h3aabe63e),
	.w8(32'hba2dfde6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b80ff),
	.w1(32'hba8caffa),
	.w2(32'hbb046cc1),
	.w3(32'hbb8f2c1d),
	.w4(32'hba3d451f),
	.w5(32'hba9b887a),
	.w6(32'hbaec15cd),
	.w7(32'h38ad63c6),
	.w8(32'hbae64d52),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa22961),
	.w1(32'hb9d59813),
	.w2(32'hba8420b3),
	.w3(32'hba8fab04),
	.w4(32'h389ee021),
	.w5(32'hba439ae0),
	.w6(32'hb9f52082),
	.w7(32'h39c61913),
	.w8(32'hb9c9a2d0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e976e),
	.w1(32'hbac32f72),
	.w2(32'h3b54753f),
	.w3(32'hbc154bbc),
	.w4(32'hb94111be),
	.w5(32'h3b268e4b),
	.w6(32'hbbdd03e7),
	.w7(32'h3ab9de78),
	.w8(32'h3b46e439),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b633f),
	.w1(32'hbaae7c01),
	.w2(32'hba8defc1),
	.w3(32'hbaedc48b),
	.w4(32'h3a07cebc),
	.w5(32'h3a2bf381),
	.w6(32'hbaabf041),
	.w7(32'h3a745c13),
	.w8(32'h3a2bea86),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ffdd2f),
	.w1(32'hb78be867),
	.w2(32'hb89ca4f3),
	.w3(32'hb836f6c5),
	.w4(32'hb7a7a93d),
	.w5(32'hb7c77f22),
	.w6(32'h378f202d),
	.w7(32'h38067d82),
	.w8(32'hb81f28d3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75c107f),
	.w1(32'h38423db2),
	.w2(32'h38a1bfe0),
	.w3(32'hb6ab192e),
	.w4(32'h37c19c61),
	.w5(32'h383eb707),
	.w6(32'hb7792e7a),
	.w7(32'hb7a8496c),
	.w8(32'h37fdc322),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39617025),
	.w1(32'h38af7c90),
	.w2(32'h3a5b0357),
	.w3(32'hb96ca07b),
	.w4(32'hb7b8ec7c),
	.w5(32'h3a949231),
	.w6(32'hb9bf3db5),
	.w7(32'hb92c9382),
	.w8(32'h3a1e0cce),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5c2a1),
	.w1(32'hbb45752c),
	.w2(32'hb778988a),
	.w3(32'hbb9c3045),
	.w4(32'h39d2ef15),
	.w5(32'h3807f0fa),
	.w6(32'hbb8234c2),
	.w7(32'hba81f756),
	.w8(32'hba3b7614),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae39f7),
	.w1(32'hbaee1026),
	.w2(32'hbbaaea58),
	.w3(32'hb9c21b06),
	.w4(32'hbaad31e5),
	.w5(32'hbb703d84),
	.w6(32'h3a718116),
	.w7(32'hba774896),
	.w8(32'hbb5de37a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73dec35),
	.w1(32'hb8315ab6),
	.w2(32'hb7d29855),
	.w3(32'h3730483b),
	.w4(32'hb8325c87),
	.w5(32'hb615d481),
	.w6(32'hb839712f),
	.w7(32'hb8316855),
	.w8(32'h36aca8a2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25d7e9),
	.w1(32'hbaed7910),
	.w2(32'hbb984ec4),
	.w3(32'hbb6471b4),
	.w4(32'hba4d54ea),
	.w5(32'hbb4cb58e),
	.w6(32'hbaacdef5),
	.w7(32'h3a122924),
	.w8(32'hbb19d1d3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b498c9),
	.w1(32'hb9bc0ecb),
	.w2(32'h3a43d438),
	.w3(32'h3abbef8d),
	.w4(32'h3a246eab),
	.w5(32'hb9c0de52),
	.w6(32'h3abbecfb),
	.w7(32'h3b310720),
	.w8(32'hbaa3a34b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8324d8),
	.w1(32'h3b583a1d),
	.w2(32'hbb494a73),
	.w3(32'hbac30d00),
	.w4(32'h38bf8fd0),
	.w5(32'hbb93ce08),
	.w6(32'hb836a3c0),
	.w7(32'h39d8d01e),
	.w8(32'hbb805146),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6dd6a),
	.w1(32'hba8e3c3b),
	.w2(32'hba0d9835),
	.w3(32'hbbab8e86),
	.w4(32'h3b0647f9),
	.w5(32'h3aeb0e37),
	.w6(32'hbbb165ab),
	.w7(32'h3a0a5f89),
	.w8(32'h3b02ddc4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ca88a),
	.w1(32'hbb278668),
	.w2(32'hbac984e4),
	.w3(32'hba67b3f1),
	.w4(32'hbaef0aec),
	.w5(32'hba450264),
	.w6(32'hb9e95b7a),
	.w7(32'hbacca266),
	.w8(32'hba214ee3),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb6c2f),
	.w1(32'h3a539274),
	.w2(32'h3a513617),
	.w3(32'h3b364b3d),
	.w4(32'h3ac66b01),
	.w5(32'h3b020143),
	.w6(32'h3b25cf0b),
	.w7(32'h3ae82c03),
	.w8(32'h3ab34f18),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1b5d7),
	.w1(32'hba91e7b5),
	.w2(32'h39e71e3c),
	.w3(32'hbb9f6823),
	.w4(32'h39a43eae),
	.w5(32'h3a8e5fbd),
	.w6(32'hbb674264),
	.w7(32'h3a9c4835),
	.w8(32'h3a74479e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba73733),
	.w1(32'hbb83b2d3),
	.w2(32'hbab39cf0),
	.w3(32'hbb5701fd),
	.w4(32'hbb0a5766),
	.w5(32'hba598f06),
	.w6(32'hbb2ab3fa),
	.w7(32'hbb29a10a),
	.w8(32'hba71212e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cf6017),
	.w1(32'h3adcc448),
	.w2(32'h3b23e84c),
	.w3(32'h38b0e76d),
	.w4(32'h3afcc170),
	.w5(32'h3b357f92),
	.w6(32'hba69ec6d),
	.w7(32'h3a64d5c3),
	.w8(32'h3b2ff3a0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e7045),
	.w1(32'h3a24013f),
	.w2(32'hb99ee1af),
	.w3(32'h39e8fb53),
	.w4(32'h38f07b06),
	.w5(32'hba0ade19),
	.w6(32'h39b2812b),
	.w7(32'hb902832e),
	.w8(32'hb9f746ca),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9949498),
	.w1(32'hb9d12177),
	.w2(32'hb9e8365d),
	.w3(32'hb97617cd),
	.w4(32'hb9b223a4),
	.w5(32'hb9b86851),
	.w6(32'hb98291db),
	.w7(32'hb983dfde),
	.w8(32'hb9a2c37d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb770eea),
	.w1(32'hbae52d68),
	.w2(32'hbb4698c1),
	.w3(32'hbb636303),
	.w4(32'hba5c6ee8),
	.w5(32'hba963ff8),
	.w6(32'hba6a1c38),
	.w7(32'h3a1b34cd),
	.w8(32'h378c7f16),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab3ed6),
	.w1(32'h3a337acb),
	.w2(32'hba7d8e80),
	.w3(32'h3a042f66),
	.w4(32'hb91f4fdb),
	.w5(32'hba757855),
	.w6(32'h3a065007),
	.w7(32'h39efa189),
	.w8(32'h397e2555),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8d616),
	.w1(32'hbab20c53),
	.w2(32'hba22e658),
	.w3(32'hbb90a728),
	.w4(32'hba2be75c),
	.w5(32'h3a9da0d2),
	.w6(32'hbb5ac9d8),
	.w7(32'h3a7fb820),
	.w8(32'h3a24c174),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c9df7),
	.w1(32'hb94492a5),
	.w2(32'hb9878ddc),
	.w3(32'hb9cad4e0),
	.w4(32'hb9723fea),
	.w5(32'hb9aecfac),
	.w6(32'hb9fe35b2),
	.w7(32'hb95b6b4b),
	.w8(32'hb849213b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b932559),
	.w1(32'hba14721d),
	.w2(32'hbac9bfe2),
	.w3(32'h3b87ce3c),
	.w4(32'hbb1f4378),
	.w5(32'hba35a2f2),
	.w6(32'h3b81f38c),
	.w7(32'hbaf04512),
	.w8(32'hba5b686a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923c98d),
	.w1(32'h3899d45f),
	.w2(32'h3732047d),
	.w3(32'hb887dc17),
	.w4(32'hb8cdf051),
	.w5(32'hb91d1f6d),
	.w6(32'h39665988),
	.w7(32'h398b0728),
	.w8(32'hb93620df),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3912b819),
	.w1(32'hb9eba821),
	.w2(32'hba0a9340),
	.w3(32'hb98a1f87),
	.w4(32'hba77d98d),
	.w5(32'hba4c90d3),
	.w6(32'hb8e113ba),
	.w7(32'hba54e306),
	.w8(32'hba6ac4b6),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b0656),
	.w1(32'hbb1b7e8a),
	.w2(32'hbad20ae1),
	.w3(32'hbbd545c5),
	.w4(32'h39f248c8),
	.w5(32'h3a9073e4),
	.w6(32'hbba54994),
	.w7(32'hb98a8411),
	.w8(32'h3ae8e20a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbbe38),
	.w1(32'hba392fdf),
	.w2(32'hbafb5d6b),
	.w3(32'hbbb37b66),
	.w4(32'h3a8a5764),
	.w5(32'hba5860b8),
	.w6(32'hba26d636),
	.w7(32'h3b5f520e),
	.w8(32'hbab5b02c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bffef),
	.w1(32'h3ae58324),
	.w2(32'h3ac4ee8f),
	.w3(32'h3aee6f76),
	.w4(32'h3a3d4db3),
	.w5(32'h3a4132a8),
	.w6(32'h3a85e6d0),
	.w7(32'h3a366ce9),
	.w8(32'h3a7638bb),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf36328),
	.w1(32'hbb555d2f),
	.w2(32'hbae6d14a),
	.w3(32'hbba72f74),
	.w4(32'hba892860),
	.w5(32'hbacb4ce1),
	.w6(32'hba6fc60b),
	.w7(32'h3b08046a),
	.w8(32'hb99a704f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb4067),
	.w1(32'h399237d7),
	.w2(32'hba5c0483),
	.w3(32'hba119184),
	.w4(32'hb9a643ed),
	.w5(32'hb9328c62),
	.w6(32'hb84a65e5),
	.w7(32'h3a2d8937),
	.w8(32'h3a639100),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43bf75),
	.w1(32'hbb11c8fb),
	.w2(32'hbbd7e811),
	.w3(32'hbb5f2ea3),
	.w4(32'hbabdcb99),
	.w5(32'hbb0ca399),
	.w6(32'hbb3a8da1),
	.w7(32'hba8747e6),
	.w8(32'hbb65cf67),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab60ac6),
	.w1(32'hbabdf105),
	.w2(32'hbb40c48f),
	.w3(32'hba8441ca),
	.w4(32'hba1b7a3a),
	.w5(32'hba246a9c),
	.w6(32'hba8d24c2),
	.w7(32'h3766ac0a),
	.w8(32'hb90f6884),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd71fdd),
	.w1(32'hbaab5b30),
	.w2(32'hbb4af788),
	.w3(32'hbbb7c723),
	.w4(32'h3a9ca6d1),
	.w5(32'hba5fe463),
	.w6(32'hba784904),
	.w7(32'h3b9edadb),
	.w8(32'hb9f7b3bc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20e9ac),
	.w1(32'h3989cd2c),
	.w2(32'hb8d0873f),
	.w3(32'hb8a234c0),
	.w4(32'h39df6c2c),
	.w5(32'h39f51d18),
	.w6(32'hb9d1af03),
	.w7(32'h39c5110d),
	.w8(32'h3a8eaab7),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88248e),
	.w1(32'hbadab41c),
	.w2(32'hbb2f6e5e),
	.w3(32'hbb6ae0bb),
	.w4(32'hba482c51),
	.w5(32'hba96fcbf),
	.w6(32'hbb0a03ca),
	.w7(32'hb910d0e7),
	.w8(32'hbae9c30f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3853d04c),
	.w1(32'h386a26d2),
	.w2(32'h38022e08),
	.w3(32'h388c933f),
	.w4(32'h371884fd),
	.w5(32'hb761ca09),
	.w6(32'h38c89d52),
	.w7(32'h37b5c7c0),
	.w8(32'h37d3f913),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef4d12),
	.w1(32'h3a125603),
	.w2(32'h39494a31),
	.w3(32'h3a444bc9),
	.w4(32'h3a3788ee),
	.w5(32'h3a6e7e5f),
	.w6(32'h3a19a65c),
	.w7(32'h39d02bbf),
	.w8(32'h39bf147e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40762b),
	.w1(32'hb95054ef),
	.w2(32'hb76586da),
	.w3(32'hba10007b),
	.w4(32'h3945fcbb),
	.w5(32'h398e4b84),
	.w6(32'hba036027),
	.w7(32'hb7230671),
	.w8(32'h3897e842),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba678c04),
	.w1(32'hbac0699b),
	.w2(32'hbb72e4e2),
	.w3(32'hbafca9b8),
	.w4(32'hbabfd867),
	.w5(32'hba420d00),
	.w6(32'hbadec66b),
	.w7(32'hba0b2b47),
	.w8(32'hb9aff05d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4dd48c7),
	.w1(32'hb753cd20),
	.w2(32'hb7286c92),
	.w3(32'h3616944f),
	.w4(32'h3720aa87),
	.w5(32'hb759ce9f),
	.w6(32'hb69e1e96),
	.w7(32'hb68c3014),
	.w8(32'hb7b45f57),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc74df),
	.w1(32'hb99086a0),
	.w2(32'hb910be4c),
	.w3(32'hb7469365),
	.w4(32'h38579ce8),
	.w5(32'hb7d62e36),
	.w6(32'h38c2cddc),
	.w7(32'h397b50f0),
	.w8(32'hb832e89c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01bb39),
	.w1(32'hba12bb07),
	.w2(32'hba2e72e6),
	.w3(32'hb90d27c9),
	.w4(32'h397bd8eb),
	.w5(32'h38a89a20),
	.w6(32'hba4095f1),
	.w7(32'hb905ad43),
	.w8(32'hba0e9477),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d33a9),
	.w1(32'hbafcac7d),
	.w2(32'hbb82153e),
	.w3(32'h3a16df0d),
	.w4(32'hba24b92a),
	.w5(32'hbb51f600),
	.w6(32'h3ad35e60),
	.w7(32'hbb0fc5f6),
	.w8(32'hbb9fd8c6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79f9a1),
	.w1(32'h3a8c8fa6),
	.w2(32'h38ed1c35),
	.w3(32'hbb818bfc),
	.w4(32'h39550276),
	.w5(32'hbac1170d),
	.w6(32'hba96fb61),
	.w7(32'h3aa77cfb),
	.w8(32'hbab58761),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a955d76),
	.w1(32'hb808071d),
	.w2(32'hba4bccf7),
	.w3(32'h3a8457f2),
	.w4(32'hb90ebcc1),
	.w5(32'hb9e21f79),
	.w6(32'h3a3e0f8b),
	.w7(32'hb841be78),
	.w8(32'hb75bdb42),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb42da5),
	.w1(32'hbb4e73a3),
	.w2(32'hbc57603c),
	.w3(32'hbb287305),
	.w4(32'hba4c37d3),
	.w5(32'hbbf218b7),
	.w6(32'h3a1ac34d),
	.w7(32'h39437d0e),
	.w8(32'hbc53b701),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07737f),
	.w1(32'hbb1d2c35),
	.w2(32'hbb09493d),
	.w3(32'hbbb067bc),
	.w4(32'h3aa2a6f4),
	.w5(32'h3af64d87),
	.w6(32'hbbca13eb),
	.w7(32'h3a3cf55e),
	.w8(32'h3b39ae47),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0732ef),
	.w1(32'h3ab0f060),
	.w2(32'hba584f55),
	.w3(32'h3a873923),
	.w4(32'h39d223c1),
	.w5(32'hbab87beb),
	.w6(32'h3a1eaaaa),
	.w7(32'h382d9c03),
	.w8(32'hba791459),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cf6419),
	.w1(32'h37c3c5f0),
	.w2(32'h3610a172),
	.w3(32'hb80b13ab),
	.w4(32'hb7444312),
	.w5(32'hb820a8fe),
	.w6(32'h378f19c1),
	.w7(32'h35adf19e),
	.w8(32'hb7643ac7),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55be64),
	.w1(32'hb9960c52),
	.w2(32'hb94630f0),
	.w3(32'hb986bd91),
	.w4(32'h39c51fe7),
	.w5(32'hb8db54b2),
	.w6(32'h38cb0f99),
	.w7(32'h397083af),
	.w8(32'h36dbc3e6),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f543fa),
	.w1(32'h387cdefb),
	.w2(32'h384cfa27),
	.w3(32'h382b9108),
	.w4(32'hb802e8fc),
	.w5(32'hb7e67b0b),
	.w6(32'hb67f6db1),
	.w7(32'hb7d62235),
	.w8(32'h376493de),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6e77a),
	.w1(32'hb8fa41e3),
	.w2(32'hbb34c60e),
	.w3(32'hba37450c),
	.w4(32'hbab48445),
	.w5(32'hbb580239),
	.w6(32'h3a93ead4),
	.w7(32'hb807b4d1),
	.w8(32'hbb160703),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28c745),
	.w1(32'hbb15b42c),
	.w2(32'hba9930ff),
	.w3(32'hbab6af35),
	.w4(32'hba0f5f1e),
	.w5(32'h39f04da5),
	.w6(32'h38d09c05),
	.w7(32'hba945e07),
	.w8(32'hbac69ec8),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5db10),
	.w1(32'hbb81182c),
	.w2(32'hbbb0c817),
	.w3(32'hbb2dca21),
	.w4(32'h3a5c22ea),
	.w5(32'hbadb897a),
	.w6(32'hbb026220),
	.w7(32'h3a8060a2),
	.w8(32'hba0a0be4),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba916d26),
	.w1(32'hb9bb471d),
	.w2(32'h3808de23),
	.w3(32'h397f7278),
	.w4(32'h3a171cb5),
	.w5(32'h3a4a6cd9),
	.w6(32'h39c8f7e2),
	.w7(32'h39c9d9e4),
	.w8(32'h360ff47a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88437c7),
	.w1(32'hbb404e6d),
	.w2(32'hbbb31e39),
	.w3(32'hba790fbe),
	.w4(32'hbb47ba3e),
	.w5(32'hbbce643c),
	.w6(32'h39b05469),
	.w7(32'hb9c2f51a),
	.w8(32'hbba12b76),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cb445),
	.w1(32'h3b1de31e),
	.w2(32'h3b7f64f4),
	.w3(32'hba822e4d),
	.w4(32'h3b8085b1),
	.w5(32'h3b9bd811),
	.w6(32'hb98fd71c),
	.w7(32'h3bb78e74),
	.w8(32'h3af32021),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b68d7),
	.w1(32'h3c2db777),
	.w2(32'h3bdf67b4),
	.w3(32'h3b0ef868),
	.w4(32'h3c114fee),
	.w5(32'hbb800a99),
	.w6(32'hbb05950b),
	.w7(32'h3929e8b9),
	.w8(32'hbc010d24),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f72d7),
	.w1(32'hbbd90321),
	.w2(32'hbb94740b),
	.w3(32'hbb820984),
	.w4(32'hbba3ff8d),
	.w5(32'hbad32aba),
	.w6(32'hbc395023),
	.w7(32'hbbd922d5),
	.w8(32'hba6cc389),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafe936),
	.w1(32'hbb0cf143),
	.w2(32'hb9a9d76e),
	.w3(32'hbba85893),
	.w4(32'hbae5972d),
	.w5(32'h3b082eac),
	.w6(32'hbb2dc1af),
	.w7(32'hbbbc42cd),
	.w8(32'hbb59a4b7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc269121),
	.w1(32'h3a394f88),
	.w2(32'h3953cf55),
	.w3(32'hbb45ccee),
	.w4(32'h3b7c83d3),
	.w5(32'h3c695883),
	.w6(32'hbbef9e36),
	.w7(32'h3b4cd259),
	.w8(32'h3c2eb469),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac615a),
	.w1(32'hba0913d7),
	.w2(32'hb9c4c7ca),
	.w3(32'h3b892208),
	.w4(32'h3ba15009),
	.w5(32'hba11dfa0),
	.w6(32'h3ba753b4),
	.w7(32'h3b23c47a),
	.w8(32'hbb99436b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fe565),
	.w1(32'h3bb06a8f),
	.w2(32'h3b183480),
	.w3(32'hbb087f3c),
	.w4(32'h3b07778e),
	.w5(32'hb99f31e8),
	.w6(32'hbbe233eb),
	.w7(32'h3ad6a11c),
	.w8(32'h3acf1643),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98f647),
	.w1(32'hb9891e01),
	.w2(32'hbbba0032),
	.w3(32'h3bd92ff5),
	.w4(32'h3c13185a),
	.w5(32'h3badd5ab),
	.w6(32'h3b9a7a33),
	.w7(32'h3c1fba4d),
	.w8(32'h3c41b485),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47718f),
	.w1(32'h3ae6f05f),
	.w2(32'hbb2f8c2f),
	.w3(32'hbc01d623),
	.w4(32'h3c743de0),
	.w5(32'h3bc04d8c),
	.w6(32'h3ba51183),
	.w7(32'h3c3abc38),
	.w8(32'h3b9ec5b4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc197b80),
	.w1(32'hbb018cab),
	.w2(32'hbbb0ef73),
	.w3(32'hbc83c8a5),
	.w4(32'h3b9d8b91),
	.w5(32'h3ab68f6a),
	.w6(32'hbc344672),
	.w7(32'h3ba34922),
	.w8(32'h3b631976),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf864b),
	.w1(32'h3b8f0624),
	.w2(32'hbb9331a5),
	.w3(32'hbb300c8b),
	.w4(32'hb99bea1a),
	.w5(32'hbc1772de),
	.w6(32'hbb138fd2),
	.w7(32'hba8c3239),
	.w8(32'hbc021d5d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39631aa0),
	.w1(32'hbb89d064),
	.w2(32'hbb2b589b),
	.w3(32'hbc044b3d),
	.w4(32'hbba69709),
	.w5(32'hbb66e783),
	.w6(32'hbbdc5e94),
	.w7(32'hbb91b986),
	.w8(32'hbad269b9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7c297),
	.w1(32'hbb01a29c),
	.w2(32'hbafaf9ef),
	.w3(32'hbb983574),
	.w4(32'hbb6e99b4),
	.w5(32'hbb73c327),
	.w6(32'hbb913b34),
	.w7(32'hbbba113e),
	.w8(32'hbbd387eb),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35899b08),
	.w1(32'hbba0a73d),
	.w2(32'hbbec4c14),
	.w3(32'hbb1bbc10),
	.w4(32'hbb64986d),
	.w5(32'hbb327d0a),
	.w6(32'hbbefa07e),
	.w7(32'hbab706fd),
	.w8(32'hbbc24b49),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3354f3),
	.w1(32'h394e9e1c),
	.w2(32'hbb6751bb),
	.w3(32'hbb2ad106),
	.w4(32'h3b2767bb),
	.w5(32'hbb440c1f),
	.w6(32'hbb459f1c),
	.w7(32'h3b6152dd),
	.w8(32'h3a12c03c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb731cd),
	.w1(32'hb865cd0d),
	.w2(32'hbb4ecba0),
	.w3(32'hbb64d017),
	.w4(32'hba5a2b77),
	.w5(32'h3b1e9332),
	.w6(32'hbaaa4163),
	.w7(32'hb9f17d7e),
	.w8(32'hbc1bf170),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad515e5),
	.w1(32'h3b803c4c),
	.w2(32'hbc5a8adb),
	.w3(32'hbba06a9a),
	.w4(32'h3c465e15),
	.w5(32'hbbba79b1),
	.w6(32'hbbdb57b5),
	.w7(32'h3c535d28),
	.w8(32'h3bac4824),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98dcfc),
	.w1(32'h3bea0a0e),
	.w2(32'hbbc920f4),
	.w3(32'hbbfa777c),
	.w4(32'h3bdccd43),
	.w5(32'hbb8b80ea),
	.w6(32'hba90043d),
	.w7(32'h3be72ac9),
	.w8(32'h3bb18228),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d2ded),
	.w1(32'h3ad37172),
	.w2(32'h3b309a57),
	.w3(32'hbbcb4084),
	.w4(32'hbaa0d26d),
	.w5(32'h3b061fc0),
	.w6(32'h3ae14b5c),
	.w7(32'h3a70bc28),
	.w8(32'h3b95d31e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2760d0),
	.w1(32'h3c24add9),
	.w2(32'hbad9a6f6),
	.w3(32'h3c012d0e),
	.w4(32'h3c5f7191),
	.w5(32'h3b128e6b),
	.w6(32'h3ba3e3d3),
	.w7(32'h3c5e94c5),
	.w8(32'h3bfa4f2f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c5164),
	.w1(32'hbc5d9418),
	.w2(32'hbc2832d4),
	.w3(32'hbbf2a40c),
	.w4(32'hbc8457f3),
	.w5(32'hbc38ceb8),
	.w6(32'h3a69d0df),
	.w7(32'hbc302108),
	.w8(32'hbc58353f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90340d),
	.w1(32'hb9583b73),
	.w2(32'hb9fc4f93),
	.w3(32'h3bb007c1),
	.w4(32'hbafbe163),
	.w5(32'h3b86e17d),
	.w6(32'h3afa3767),
	.w7(32'hbaa6c8c1),
	.w8(32'hbba48156),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf51a2),
	.w1(32'h3bef634a),
	.w2(32'h3c81758e),
	.w3(32'hbad7284c),
	.w4(32'h3b405562),
	.w5(32'h3c07f68e),
	.w6(32'hbc129d4f),
	.w7(32'hbbe79b7e),
	.w8(32'hbbd6690f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1742c9),
	.w1(32'h3bb79a1b),
	.w2(32'h3c2dc6d6),
	.w3(32'h3b2d927c),
	.w4(32'h3ba5b2c3),
	.w5(32'h3bb6daf0),
	.w6(32'hbc7ced74),
	.w7(32'hbb6875c3),
	.w8(32'hbc5269d7),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24f0d7),
	.w1(32'hb9e15ed5),
	.w2(32'hbb0f7387),
	.w3(32'h3bd5b405),
	.w4(32'h3b5a47e2),
	.w5(32'h3a028344),
	.w6(32'hbc005efd),
	.w7(32'h3b2ec112),
	.w8(32'hba0d326c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa5635),
	.w1(32'hbb5deec8),
	.w2(32'hbb0742c7),
	.w3(32'hb9f87db8),
	.w4(32'hbc4410ce),
	.w5(32'hbbaa84b3),
	.w6(32'hb9d7d969),
	.w7(32'hbc6e8648),
	.w8(32'hbacc33f3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc16cb5),
	.w1(32'hba5f7747),
	.w2(32'hbbbb65df),
	.w3(32'h3b99bdc6),
	.w4(32'hbbbac2f6),
	.w5(32'hbc0d55a1),
	.w6(32'h3c19318b),
	.w7(32'hba566abf),
	.w8(32'hbb94928c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ae812),
	.w1(32'hbb14a97f),
	.w2(32'h3a2c3ab5),
	.w3(32'hbac46afa),
	.w4(32'hbb438901),
	.w5(32'hbb5aed3d),
	.w6(32'h39a6493a),
	.w7(32'hbae8fefc),
	.w8(32'hbb8307c0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50e876),
	.w1(32'hbc01d2a6),
	.w2(32'hbc0fadeb),
	.w3(32'hbb073cdb),
	.w4(32'hbc4f7d83),
	.w5(32'hbca1110d),
	.w6(32'h3a43e4db),
	.w7(32'hbc27b259),
	.w8(32'hbc16187f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d14af),
	.w1(32'hbb8a8edf),
	.w2(32'hbb9b696d),
	.w3(32'hbc42aee9),
	.w4(32'hbb811cba),
	.w5(32'h3b924c2c),
	.w6(32'hbc167a75),
	.w7(32'hb9b9ef93),
	.w8(32'hba8744d4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03c9b1),
	.w1(32'h3b03b09d),
	.w2(32'h3adc5d30),
	.w3(32'hbb22b61e),
	.w4(32'h3bc95ac3),
	.w5(32'h3b90253a),
	.w6(32'h3b37d198),
	.w7(32'h3b9fd951),
	.w8(32'h3aca353d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b5ebb),
	.w1(32'h3ac3cabd),
	.w2(32'h3ba42c9f),
	.w3(32'h3b830671),
	.w4(32'hbb0e50d8),
	.w5(32'h3b24de30),
	.w6(32'h3a31fa45),
	.w7(32'hbb384427),
	.w8(32'h3a1b88f5),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1439f),
	.w1(32'h3c964c64),
	.w2(32'h3b3b8ef5),
	.w3(32'h3bdc7eb4),
	.w4(32'h3b58f574),
	.w5(32'hbc13f3b2),
	.w6(32'h3bd914a6),
	.w7(32'h3bab4d97),
	.w8(32'h3b74f6d5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3cbfe),
	.w1(32'h3c46e5ee),
	.w2(32'h3c23d1f0),
	.w3(32'h3bc7b73c),
	.w4(32'h3c8c19ac),
	.w5(32'h3c4cd146),
	.w6(32'h3c97fae9),
	.w7(32'h3c462934),
	.w8(32'h3c614114),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f76cb),
	.w1(32'h3b3f9b7c),
	.w2(32'h3b242e28),
	.w3(32'h3a1894f8),
	.w4(32'hbc236b6e),
	.w5(32'hbc39fb85),
	.w6(32'h3bcfda24),
	.w7(32'hbc152ce8),
	.w8(32'hbc618715),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb868ec),
	.w1(32'hbc3d2505),
	.w2(32'hbbe56d8d),
	.w3(32'hbc153cad),
	.w4(32'hbc316141),
	.w5(32'hbbe5c288),
	.w6(32'hbc85282f),
	.w7(32'hbb8cd185),
	.w8(32'hbb7519be),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395185a4),
	.w1(32'h3be60c6f),
	.w2(32'hba2705e1),
	.w3(32'hbb3cf8e0),
	.w4(32'h3c26f23f),
	.w5(32'h3b4e1bcc),
	.w6(32'hbb541b97),
	.w7(32'h3c14f722),
	.w8(32'hbaa3072e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba566bcf),
	.w1(32'hbb1166ec),
	.w2(32'h3b29d709),
	.w3(32'hbc086fd0),
	.w4(32'hbb8d370c),
	.w5(32'h3a864ea7),
	.w6(32'hbbc4ef6e),
	.w7(32'hbbbff8df),
	.w8(32'hbb916710),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17083d),
	.w1(32'h3b1405e2),
	.w2(32'h3bc18b8e),
	.w3(32'h3bff3fc9),
	.w4(32'hbb843ec4),
	.w5(32'hbbbf7d80),
	.w6(32'hbb3336db),
	.w7(32'hb9b03054),
	.w8(32'hbb7bcf16),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b311cc1),
	.w1(32'h3b87289e),
	.w2(32'h3c94993d),
	.w3(32'hbb1a788f),
	.w4(32'hbb729faa),
	.w5(32'h3bb05db4),
	.w6(32'hbb8b7aae),
	.w7(32'hbb7c1cbf),
	.w8(32'hbb9f6b7a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9fb74d),
	.w1(32'hba78eafe),
	.w2(32'h3c149cf0),
	.w3(32'h3c3b777f),
	.w4(32'h3b59a58f),
	.w5(32'h3b0cbbc4),
	.w6(32'hbc1b9f9c),
	.w7(32'h3a87e45b),
	.w8(32'hbb3a7fad),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b1c2f),
	.w1(32'hbc1993b4),
	.w2(32'hbc26ffe0),
	.w3(32'hbb732553),
	.w4(32'hbc62e78c),
	.w5(32'hbc4a8b6e),
	.w6(32'hbadcff34),
	.w7(32'hbc654799),
	.w8(32'hbc174a46),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a84a2),
	.w1(32'hbb8bd740),
	.w2(32'hbb67a90a),
	.w3(32'hbc22e98c),
	.w4(32'hbbf7df79),
	.w5(32'hbaf54180),
	.w6(32'hbb3e5eca),
	.w7(32'hbb67d5b6),
	.w8(32'h3b59b44a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2e11d),
	.w1(32'hbb3b3cec),
	.w2(32'h3b864b17),
	.w3(32'h3b1e600a),
	.w4(32'h3b4efd2d),
	.w5(32'h3c828431),
	.w6(32'h3bb04daa),
	.w7(32'hbad76e0b),
	.w8(32'h3bb907a8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbfe7e),
	.w1(32'hba23e8c6),
	.w2(32'hba1c51bb),
	.w3(32'h3b264a7d),
	.w4(32'h3a9339b8),
	.w5(32'h3a79d3b2),
	.w6(32'hbba88bf1),
	.w7(32'hbb3c9102),
	.w8(32'hba591ac0),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5cf0e),
	.w1(32'hbbcbe4cd),
	.w2(32'h3ac44283),
	.w3(32'hbc123d2d),
	.w4(32'hbbbffeb2),
	.w5(32'h3b90abfb),
	.w6(32'hbc3383ad),
	.w7(32'hbb513138),
	.w8(32'h3b8e1120),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9af0d),
	.w1(32'hbb25dc87),
	.w2(32'h3c3b6bf9),
	.w3(32'h3b060868),
	.w4(32'hbc261cd7),
	.w5(32'h3b3011e3),
	.w6(32'h3aa1346e),
	.w7(32'hbc0b2997),
	.w8(32'hbad68c52),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52d5dc),
	.w1(32'h3c72d905),
	.w2(32'h3c9c80ff),
	.w3(32'h3c5bcbaa),
	.w4(32'h3b8d1d04),
	.w5(32'hbafa5486),
	.w6(32'hb9a08213),
	.w7(32'hbc0185d2),
	.w8(32'hbcb57bac),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48b181),
	.w1(32'hbc711fd7),
	.w2(32'hbc742aae),
	.w3(32'hbbe530d3),
	.w4(32'hbbd50efa),
	.w5(32'hbb53f388),
	.w6(32'hbcc25e3f),
	.w7(32'h398abc53),
	.w8(32'h3c31665d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b95d0),
	.w1(32'h3c0705c9),
	.w2(32'h3bf25a32),
	.w3(32'h3a1409f9),
	.w4(32'h39b6858d),
	.w5(32'hb81da2e5),
	.w6(32'h3c91eb4d),
	.w7(32'h3be9d7c5),
	.w8(32'h3c0e8d96),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8cf58),
	.w1(32'h3b94ecc7),
	.w2(32'h3b63eb08),
	.w3(32'h3c2b3382),
	.w4(32'h3b4a6644),
	.w5(32'h3b7a9b50),
	.w6(32'h3c082c5e),
	.w7(32'h3b1a0903),
	.w8(32'h3b39b74c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baef804),
	.w1(32'hbb8df01b),
	.w2(32'hba4dede3),
	.w3(32'h3c08d0ef),
	.w4(32'hbb54cd3f),
	.w5(32'h3b7fa323),
	.w6(32'h3b621dd0),
	.w7(32'hba4adcce),
	.w8(32'h3bb99f80),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6370d4),
	.w1(32'hbba1c832),
	.w2(32'hbbc568e9),
	.w3(32'h3b4ef848),
	.w4(32'hbbe10097),
	.w5(32'hbb3255b0),
	.w6(32'h3bee0f0f),
	.w7(32'hbba1a155),
	.w8(32'h38099d35),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ecfe6),
	.w1(32'hba9c5594),
	.w2(32'h3bed7024),
	.w3(32'hbaf86a17),
	.w4(32'hbc19f608),
	.w5(32'h3a8b561d),
	.w6(32'hba9e0443),
	.w7(32'hbc21364d),
	.w8(32'hbaea3958),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac2d6c),
	.w1(32'h3aca2dfb),
	.w2(32'h3c23d790),
	.w3(32'h3b90a042),
	.w4(32'hbbaaba3c),
	.w5(32'hbbdb8881),
	.w6(32'hbb003682),
	.w7(32'hbc085d4c),
	.w8(32'hbc402041),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcec824),
	.w1(32'hbb84270e),
	.w2(32'h39275b56),
	.w3(32'hbc097a2e),
	.w4(32'h3be4f03b),
	.w5(32'h3c8126c9),
	.w6(32'hbcab4852),
	.w7(32'hbad15b6c),
	.w8(32'h3b371a80),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21b562),
	.w1(32'h3b5c0cf7),
	.w2(32'h3b9c276e),
	.w3(32'h3c184cd0),
	.w4(32'h3b706640),
	.w5(32'h3be4502b),
	.w6(32'hbbab98b9),
	.w7(32'h3a97cfd8),
	.w8(32'h3b6e20ba),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb415cb),
	.w1(32'hbb862d0f),
	.w2(32'hbacce8ae),
	.w3(32'h3b286c48),
	.w4(32'hbbc78d99),
	.w5(32'hbadfe345),
	.w6(32'h3addaa93),
	.w7(32'hbb8ff64c),
	.w8(32'hbb3d1067),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule