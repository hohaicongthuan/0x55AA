module layer_10_featuremap_276(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade3c67),
	.w1(32'h3a18b827),
	.w2(32'hb9fe5e1c),
	.w3(32'hbaac4034),
	.w4(32'hbb70e66b),
	.w5(32'h3b7db615),
	.w6(32'h3acdb862),
	.w7(32'hbb36cdd6),
	.w8(32'h3b3c4f46),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26ba31),
	.w1(32'h3b982447),
	.w2(32'h3b1d487c),
	.w3(32'h3b5f640c),
	.w4(32'h3af3870a),
	.w5(32'hba880837),
	.w6(32'h3c02c673),
	.w7(32'h3b4d0473),
	.w8(32'h3939fdc0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76857b),
	.w1(32'hbaaffbd1),
	.w2(32'hbb19236c),
	.w3(32'hba8e6e0d),
	.w4(32'h39aa8c7b),
	.w5(32'h3a638240),
	.w6(32'h3b8e4391),
	.w7(32'h394a4160),
	.w8(32'h3ab586f1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2b355),
	.w1(32'h3b1ae74d),
	.w2(32'h3b345123),
	.w3(32'h3b33477a),
	.w4(32'h3b76731e),
	.w5(32'h39e60888),
	.w6(32'h3a93a8e6),
	.w7(32'h3b3ce2d3),
	.w8(32'hba8c130a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02551f),
	.w1(32'hb9870e5f),
	.w2(32'hb9a8eeaa),
	.w3(32'h3a1f6042),
	.w4(32'h3a4c95a0),
	.w5(32'hba9518d8),
	.w6(32'hb9a0d9dd),
	.w7(32'h3a0415e1),
	.w8(32'hbac6c5c4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8821d),
	.w1(32'hb9359efd),
	.w2(32'hba0b476b),
	.w3(32'hb92e0125),
	.w4(32'hbacc2c38),
	.w5(32'h3a78c699),
	.w6(32'hba3c3609),
	.w7(32'hbae104ec),
	.w8(32'h3a8c9436),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e7938),
	.w1(32'h3aeaa949),
	.w2(32'hbb00db54),
	.w3(32'h3b696230),
	.w4(32'h370fc0c8),
	.w5(32'hbb62f561),
	.w6(32'h3b2a84fe),
	.w7(32'hbabed9a2),
	.w8(32'hbb8f4f3a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc154c28),
	.w1(32'hbc22ded0),
	.w2(32'hbbf9c528),
	.w3(32'hbc149303),
	.w4(32'hbb607f78),
	.w5(32'h3abc5943),
	.w6(32'hbc36c5f4),
	.w7(32'hbacee773),
	.w8(32'h3abd6666),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa34e84),
	.w1(32'h3af69495),
	.w2(32'h3b1a1c7f),
	.w3(32'hba5f4c60),
	.w4(32'hb98a9ab2),
	.w5(32'hbb5af225),
	.w6(32'hba6ad5a0),
	.w7(32'hba6ab524),
	.w8(32'hbb88484e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a1664),
	.w1(32'hbaf7fae7),
	.w2(32'h3b497de3),
	.w3(32'h3b919b1f),
	.w4(32'h3b029acb),
	.w5(32'h3b9233f4),
	.w6(32'hbb7fce97),
	.w7(32'hbb7c623c),
	.w8(32'hbb08ca87),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397de68d),
	.w1(32'h39394ec8),
	.w2(32'hbaba8cda),
	.w3(32'hb98a14d6),
	.w4(32'hba575b04),
	.w5(32'h3a3f1632),
	.w6(32'h3a56ca75),
	.w7(32'hb9efd164),
	.w8(32'hba82d530),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51ff3a),
	.w1(32'hb912b19e),
	.w2(32'hbbb3d3cf),
	.w3(32'h3be10b1c),
	.w4(32'hbb13a8d1),
	.w5(32'hbbb001e6),
	.w6(32'h3af192ce),
	.w7(32'hbba6c6b2),
	.w8(32'hbb90be08),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba465f91),
	.w1(32'hbc03bf53),
	.w2(32'hbadfa3a2),
	.w3(32'h3b409bea),
	.w4(32'hbb5486aa),
	.w5(32'h3b09fd87),
	.w6(32'hbbc13c22),
	.w7(32'hbc2d9c2d),
	.w8(32'hbb26c843),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9dd764),
	.w1(32'hbbb07828),
	.w2(32'hbb8ea2af),
	.w3(32'hbaa43347),
	.w4(32'hbadf5a80),
	.w5(32'h3b022d81),
	.w6(32'hbb2bfde3),
	.w7(32'hbb6f2911),
	.w8(32'h39f4bcc1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966356d),
	.w1(32'h3b1e49fd),
	.w2(32'h3b7fd1f4),
	.w3(32'h3b1fc624),
	.w4(32'h3b8d84ca),
	.w5(32'hbb006cf3),
	.w6(32'hbaf86db6),
	.w7(32'hba2c80b3),
	.w8(32'hbb8d5793),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb04286),
	.w1(32'hbb4c9f8d),
	.w2(32'h3a97a861),
	.w3(32'h3a325e16),
	.w4(32'h3b0765d6),
	.w5(32'h3be8692c),
	.w6(32'hbb057f5a),
	.w7(32'h3a342d8c),
	.w8(32'h3b74b35a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ee756),
	.w1(32'h3b4cdb2c),
	.w2(32'h3b1d90b1),
	.w3(32'h3afce61c),
	.w4(32'h3b27d794),
	.w5(32'hb79f0603),
	.w6(32'h3bb7db81),
	.w7(32'h3b502ec6),
	.w8(32'hba231634),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd25478),
	.w1(32'hbc2c2fe7),
	.w2(32'hbbc8ce64),
	.w3(32'hbbbf5b90),
	.w4(32'hbbd23baf),
	.w5(32'h3b4c50c9),
	.w6(32'hbc030be9),
	.w7(32'hbc023a88),
	.w8(32'h3a40ed83),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94725ea),
	.w1(32'hbb891f7f),
	.w2(32'hba104560),
	.w3(32'hb9b4c90f),
	.w4(32'hbb0e8f2a),
	.w5(32'h3b01fdff),
	.w6(32'hbb6d2a2f),
	.w7(32'hbb63b7d9),
	.w8(32'hb98ee3a6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c5676),
	.w1(32'h3950ba34),
	.w2(32'hba062f59),
	.w3(32'h3b06e5a1),
	.w4(32'h3aab2b54),
	.w5(32'hb8130264),
	.w6(32'hba0c776a),
	.w7(32'hb92b077c),
	.w8(32'hba75947f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ec93af),
	.w1(32'hbb34fd99),
	.w2(32'hbaa9b066),
	.w3(32'hba142343),
	.w4(32'h3ab0c10f),
	.w5(32'hbb0a3b74),
	.w6(32'hbab34028),
	.w7(32'h399ba9f9),
	.w8(32'hbab7d844),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd6470),
	.w1(32'h3a911abc),
	.w2(32'h39aede4a),
	.w3(32'h38d93339),
	.w4(32'h3b3b2f03),
	.w5(32'hb6b05e72),
	.w6(32'hba92aa4d),
	.w7(32'h3af220a3),
	.w8(32'hba917aac),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9208ea),
	.w1(32'hbbbf278c),
	.w2(32'h3a2c5902),
	.w3(32'hbbaafdfa),
	.w4(32'h3a66593c),
	.w5(32'h3c14baf7),
	.w6(32'hbbe11064),
	.w7(32'hbb81d1eb),
	.w8(32'h3bcf620d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac83265),
	.w1(32'h3aa90886),
	.w2(32'h3bac9ce6),
	.w3(32'h3b46feb5),
	.w4(32'h3b51ed4a),
	.w5(32'h3b4acc7c),
	.w6(32'hbafc429c),
	.w7(32'hb8cc06e4),
	.w8(32'hbb190ba1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3820e4),
	.w1(32'hba732889),
	.w2(32'hbafd5a2f),
	.w3(32'h3b5ab15d),
	.w4(32'h3ab6f858),
	.w5(32'hb94562c9),
	.w6(32'h3b8209e9),
	.w7(32'hbb3997d4),
	.w8(32'hbc0f633b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ee464),
	.w1(32'h3a340c92),
	.w2(32'h3afcc01e),
	.w3(32'hba92e68c),
	.w4(32'h39cfc5c2),
	.w5(32'hba3939bf),
	.w6(32'hbb12dc54),
	.w7(32'h3a0ffc64),
	.w8(32'hbabd67b3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b474d),
	.w1(32'h3b2bdae7),
	.w2(32'h3ae2f796),
	.w3(32'hba24c929),
	.w4(32'h3aebd167),
	.w5(32'hbacb1598),
	.w6(32'h397c37e6),
	.w7(32'h3ab69cd3),
	.w8(32'hba8701a4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7981b0),
	.w1(32'hbafb1963),
	.w2(32'hb974725b),
	.w3(32'h3b6c00fc),
	.w4(32'hb9fc3526),
	.w5(32'hbb91020e),
	.w6(32'h3a1bdd6e),
	.w7(32'hbb1d9864),
	.w8(32'hbabf181e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9badd5),
	.w1(32'h3bb0b811),
	.w2(32'h3a3e3436),
	.w3(32'h3afe2fed),
	.w4(32'h3ae56148),
	.w5(32'h3ae0b92c),
	.w6(32'h3b3fe24d),
	.w7(32'h3acade01),
	.w8(32'h3b12072a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04a6ef),
	.w1(32'h3bc72d2a),
	.w2(32'h3b8b0e01),
	.w3(32'h3c0a159a),
	.w4(32'h3ab76256),
	.w5(32'h3afe0317),
	.w6(32'h3c090db3),
	.w7(32'h3a40882f),
	.w8(32'hbc03a160),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af06ef1),
	.w1(32'h3bc7e032),
	.w2(32'h3b8198c1),
	.w3(32'h3a4f518f),
	.w4(32'hba994f98),
	.w5(32'h3a153e1c),
	.w6(32'h3a52a329),
	.w7(32'h3914a299),
	.w8(32'h3af2e504),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f650d),
	.w1(32'hbb44c501),
	.w2(32'hbaee0422),
	.w3(32'hba763760),
	.w4(32'hba448da9),
	.w5(32'hba4cd844),
	.w6(32'hba7d3ea0),
	.w7(32'hbaa28e77),
	.w8(32'hbaf86f09),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb438d1d),
	.w1(32'hbb0658a4),
	.w2(32'hba87d36e),
	.w3(32'hbb2fbdbf),
	.w4(32'hba58a321),
	.w5(32'hb9cdc67c),
	.w6(32'hbb1c6e55),
	.w7(32'hbb509222),
	.w8(32'hbb7d2cfb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e2701),
	.w1(32'hbb449555),
	.w2(32'hbb8650ec),
	.w3(32'hba8e730b),
	.w4(32'hbb6bc9f9),
	.w5(32'hbb2eb414),
	.w6(32'hba85bbf4),
	.w7(32'hbbb4672f),
	.w8(32'hbb4d681c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77c38f),
	.w1(32'hba1cefce),
	.w2(32'h39bcea5f),
	.w3(32'h3a60c91e),
	.w4(32'h3aa68206),
	.w5(32'h3a0ea7a3),
	.w6(32'hba1b2e21),
	.w7(32'h3af3106c),
	.w8(32'h3ad76964),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b0c4d),
	.w1(32'hbab6e1bc),
	.w2(32'hbb30d1f1),
	.w3(32'hbafa49e4),
	.w4(32'hbb2efa6a),
	.w5(32'hba76819a),
	.w6(32'h3acc3311),
	.w7(32'hbb61442a),
	.w8(32'hbaf15380),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef4e44),
	.w1(32'hba999c5e),
	.w2(32'hbba3efb8),
	.w3(32'h3b29dcbf),
	.w4(32'hba5fd28e),
	.w5(32'hba8be771),
	.w6(32'h3bc2b04e),
	.w7(32'hbbfeb2ef),
	.w8(32'hba2bc763),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98ba60),
	.w1(32'h3b0a4a3f),
	.w2(32'hbb90aaa0),
	.w3(32'hb92d6919),
	.w4(32'hbb03165f),
	.w5(32'hbc0cab67),
	.w6(32'hbba74821),
	.w7(32'hbbfb840c),
	.w8(32'hbc36762e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c081e28),
	.w1(32'h3bbe28d9),
	.w2(32'hbb665a7e),
	.w3(32'h3bd262d0),
	.w4(32'h3a2587db),
	.w5(32'hbc289783),
	.w6(32'h3b24372e),
	.w7(32'hbb9d1d12),
	.w8(32'hbc4800b2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7ce6c),
	.w1(32'hbb0fbcd9),
	.w2(32'hbaaad071),
	.w3(32'h3b20df20),
	.w4(32'h3ad4fa71),
	.w5(32'h3a06c922),
	.w6(32'hbabab47d),
	.w7(32'h3a4e48a0),
	.w8(32'hbb065fee),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90bda0),
	.w1(32'h3a0f833e),
	.w2(32'h3a1aef6c),
	.w3(32'hbae869be),
	.w4(32'hbb6055e3),
	.w5(32'hbab2979f),
	.w6(32'hbacb7a1e),
	.w7(32'hbaa2a0cd),
	.w8(32'hba02510d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4dfdc0),
	.w1(32'h3a16cc9c),
	.w2(32'h3a4a1730),
	.w3(32'hba9a9165),
	.w4(32'h3a05181c),
	.w5(32'h3ad9bfab),
	.w6(32'h3a0770f2),
	.w7(32'h3aca54ee),
	.w8(32'h398511ce),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82d4ce),
	.w1(32'h3afca1ec),
	.w2(32'h3b107151),
	.w3(32'h3b042697),
	.w4(32'h39d4d580),
	.w5(32'h3b9b02c0),
	.w6(32'hbad0e602),
	.w7(32'hbab04589),
	.w8(32'hb9cf2dae),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d611fc),
	.w1(32'h3a63f740),
	.w2(32'h3bbd8bb9),
	.w3(32'h3bb53e5b),
	.w4(32'h3b762fc6),
	.w5(32'h3b959cc6),
	.w6(32'hba8dc987),
	.w7(32'hba9b479e),
	.w8(32'hba489007),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd081cd),
	.w1(32'hbb81f35b),
	.w2(32'hbb1ea64c),
	.w3(32'hbaa71acf),
	.w4(32'hb93c3c4e),
	.w5(32'h3a83c5be),
	.w6(32'hbbd9f615),
	.w7(32'hbbc8af69),
	.w8(32'hbbf2c72f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bd6b4),
	.w1(32'h39ec843d),
	.w2(32'h3ba3fd12),
	.w3(32'h3abccf4a),
	.w4(32'h3b0ab482),
	.w5(32'h3bbf2b60),
	.w6(32'hbb8382f9),
	.w7(32'hbb08328b),
	.w8(32'hbb3ff226),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5f23c),
	.w1(32'hbb3733a8),
	.w2(32'hba85b8c1),
	.w3(32'hbb2a6963),
	.w4(32'h3a10137e),
	.w5(32'h3980c7a5),
	.w6(32'hbc0618fb),
	.w7(32'hbb8c55fb),
	.w8(32'hbb8bdc6c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91183d),
	.w1(32'hbacf0d72),
	.w2(32'h3afab34a),
	.w3(32'hb9c01e62),
	.w4(32'h3a15a434),
	.w5(32'h3acc7fa0),
	.w6(32'hbb75da30),
	.w7(32'hba8c7cf6),
	.w8(32'h3ab1d6a1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a98952),
	.w1(32'h3ae42b22),
	.w2(32'h3ac196fb),
	.w3(32'hbb08a568),
	.w4(32'hbb867fc7),
	.w5(32'hbab676f4),
	.w6(32'hba9d1379),
	.w7(32'hbb0f40a7),
	.w8(32'hba77c3bb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a037540),
	.w1(32'h3a2de681),
	.w2(32'h3ad19bfe),
	.w3(32'hb91d7eaf),
	.w4(32'h3aecf379),
	.w5(32'h3b5d517a),
	.w6(32'hb998bd1b),
	.w7(32'h3b0002bc),
	.w8(32'h3a1600a3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc643d),
	.w1(32'h3a9279b4),
	.w2(32'h3a6df3a7),
	.w3(32'hbb13c036),
	.w4(32'hbacf930b),
	.w5(32'h38ec7e52),
	.w6(32'hba8ac232),
	.w7(32'h3955ea6b),
	.w8(32'hba654f6a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e16d8),
	.w1(32'hbb9d43f4),
	.w2(32'hbb3311a1),
	.w3(32'hbaa1846c),
	.w4(32'hbab5fb0d),
	.w5(32'h3b79163e),
	.w6(32'hbb545116),
	.w7(32'hbb77dee0),
	.w8(32'hba56a6a3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb478b),
	.w1(32'hbb0c5f5b),
	.w2(32'hbb4f5f15),
	.w3(32'hbb32bd4b),
	.w4(32'hbb1ec127),
	.w5(32'hb9fbdd8a),
	.w6(32'hba5f7b30),
	.w7(32'hbb5cb985),
	.w8(32'hbb58a9c1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0562c6),
	.w1(32'hbc0acc7d),
	.w2(32'hbb4577b7),
	.w3(32'hba3c8160),
	.w4(32'hbae96731),
	.w5(32'h3bb67b99),
	.w6(32'hbbd753cd),
	.w7(32'hbbabf518),
	.w8(32'hb9f0075f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97544e),
	.w1(32'hbb147dd3),
	.w2(32'hba8ad8de),
	.w3(32'h3ac01ec2),
	.w4(32'h3a574456),
	.w5(32'h3abf331f),
	.w6(32'hbaf228da),
	.w7(32'hba6377f8),
	.w8(32'h3ada3006),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4aba6f),
	.w1(32'h387e9715),
	.w2(32'h3aaf6c3e),
	.w3(32'h389e9a6b),
	.w4(32'h39e1fcf9),
	.w5(32'hbade029a),
	.w6(32'h3abb8ab5),
	.w7(32'h3b456c7b),
	.w8(32'hbb41cb73),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42d321),
	.w1(32'hba76dc16),
	.w2(32'hb9a866c7),
	.w3(32'hbb2037f9),
	.w4(32'hbab4868f),
	.w5(32'h3aa9a704),
	.w6(32'hbb76b577),
	.w7(32'hba81ce87),
	.w8(32'h3aff3b97),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12a018),
	.w1(32'h3a515aea),
	.w2(32'hbaa98e4f),
	.w3(32'h3b5a83ab),
	.w4(32'h3a1b86db),
	.w5(32'hbaf24ce3),
	.w6(32'h3b1e3ba9),
	.w7(32'hb9d5bea5),
	.w8(32'hbafc3993),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa45a6f),
	.w1(32'h3a545e11),
	.w2(32'hb7b8de99),
	.w3(32'hba95baa8),
	.w4(32'h3ae86efb),
	.w5(32'hbb4fa5aa),
	.w6(32'hba686402),
	.w7(32'h3abfabf2),
	.w8(32'hbae185ee),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a912d71),
	.w1(32'h39af2389),
	.w2(32'hba9c5060),
	.w3(32'hbacd55b4),
	.w4(32'hb9fe2b1a),
	.w5(32'hb7f3851d),
	.w6(32'h388eea98),
	.w7(32'h3ab029ef),
	.w8(32'h3ac2b1d8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba021a96),
	.w1(32'hbb0f1754),
	.w2(32'h3a39dd25),
	.w3(32'hba2918fb),
	.w4(32'hbb3f2ffa),
	.w5(32'hb995d3fb),
	.w6(32'hbb3327a2),
	.w7(32'hbbbdd3f6),
	.w8(32'hba99aa53),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75d7bb),
	.w1(32'hbac1669f),
	.w2(32'h3b59b8ac),
	.w3(32'hbb8c041e),
	.w4(32'h3af2c26f),
	.w5(32'h3ac57396),
	.w6(32'h3aa18192),
	.w7(32'h3ba1a4c9),
	.w8(32'h3ab866a9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13041e),
	.w1(32'hbb01b59e),
	.w2(32'hba2115e7),
	.w3(32'h3b2af094),
	.w4(32'h3b17ac00),
	.w5(32'hb897a9ca),
	.w6(32'h3a88ea28),
	.w7(32'h3a909d19),
	.w8(32'hba4b9223),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe493a),
	.w1(32'hba96a27b),
	.w2(32'h39646a1d),
	.w3(32'hbabac724),
	.w4(32'hb865101f),
	.w5(32'hba3483f0),
	.w6(32'hbb0b8815),
	.w7(32'h39f72c0f),
	.w8(32'hbafd0434),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb303522),
	.w1(32'hbaa73958),
	.w2(32'hb9b56158),
	.w3(32'h3aed859c),
	.w4(32'h3ac01f76),
	.w5(32'h3b16ea13),
	.w6(32'hba6d93a9),
	.w7(32'h3b0ecdca),
	.w8(32'hb9344bc8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3c7b3),
	.w1(32'h3abe0e3c),
	.w2(32'h3b087919),
	.w3(32'h3b48cb07),
	.w4(32'hb736a180),
	.w5(32'h3b29a0dd),
	.w6(32'h3aed5ac1),
	.w7(32'h3a26cf10),
	.w8(32'h3ae5641d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cc75f),
	.w1(32'hbb7ffc01),
	.w2(32'h3b9221b9),
	.w3(32'h3ab47121),
	.w4(32'h3af5d15f),
	.w5(32'h3bdca44d),
	.w6(32'hbb3bc4b1),
	.w7(32'h3b3a6fc9),
	.w8(32'h3c689482),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb807e337),
	.w1(32'h39b1ff89),
	.w2(32'h3a84b565),
	.w3(32'hb8caa680),
	.w4(32'h3b831206),
	.w5(32'h3bd114ce),
	.w6(32'hbbb959ba),
	.w7(32'hbb27dbe5),
	.w8(32'hbad8ba3c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8a9b9),
	.w1(32'hbc295dd8),
	.w2(32'hbbf85009),
	.w3(32'hbbf5faf3),
	.w4(32'hbbbe05ec),
	.w5(32'hbaa0a697),
	.w6(32'hbc14cc38),
	.w7(32'hbbdeeeed),
	.w8(32'hbbc46f3a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae371a0),
	.w1(32'hbb3ef724),
	.w2(32'hbad29c19),
	.w3(32'h3abb154c),
	.w4(32'hbab29505),
	.w5(32'hbbc22fd4),
	.w6(32'hbc0aa361),
	.w7(32'hbc1fcb24),
	.w8(32'hbc82633b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a147d37),
	.w1(32'h3a3f937a),
	.w2(32'h3a59918c),
	.w3(32'hba23100c),
	.w4(32'h3a2b5a87),
	.w5(32'h3a94888d),
	.w6(32'h38d762d4),
	.w7(32'h3a8c18bc),
	.w8(32'h3b97bbfa),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9eed2d),
	.w1(32'hba690f23),
	.w2(32'h3ac37681),
	.w3(32'h3b5a739c),
	.w4(32'h3ad8b957),
	.w5(32'h3aa64c69),
	.w6(32'h3b8ba241),
	.w7(32'h3a9e26d8),
	.w8(32'h3b601626),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7a722),
	.w1(32'h3ad2974d),
	.w2(32'h3859edb9),
	.w3(32'h3b9531e8),
	.w4(32'h3b8137ef),
	.w5(32'hba9ecdec),
	.w6(32'h3b8819ed),
	.w7(32'hba892547),
	.w8(32'hbb1322f7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fb43a),
	.w1(32'hbbd06ad8),
	.w2(32'hbb9cd472),
	.w3(32'hb983937c),
	.w4(32'hbba582c3),
	.w5(32'h398acf83),
	.w6(32'hbaef61ed),
	.w7(32'hbbb6a9ea),
	.w8(32'hb985be1e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a506d40),
	.w1(32'hbaef6052),
	.w2(32'hbb8285e8),
	.w3(32'h3b166e57),
	.w4(32'hba87c11f),
	.w5(32'hba9ad0f6),
	.w6(32'h3b359f9b),
	.w7(32'hbb3a29ce),
	.w8(32'hbaa2d9d0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3cbb4),
	.w1(32'hbc199154),
	.w2(32'hbbbdef92),
	.w3(32'hbba17b3a),
	.w4(32'hbc018f1b),
	.w5(32'h3ad416f1),
	.w6(32'hbbdcbd51),
	.w7(32'hbc19d6a8),
	.w8(32'h398f7a66),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb337113),
	.w1(32'hbb685a15),
	.w2(32'hbb61b399),
	.w3(32'hbbb42edf),
	.w4(32'hbbbc167e),
	.w5(32'hb974ac85),
	.w6(32'hbbf34b25),
	.w7(32'hbbfa3599),
	.w8(32'hbb6b2211),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a893709),
	.w1(32'hba4d5f10),
	.w2(32'hbaa60d29),
	.w3(32'h3b8ecb90),
	.w4(32'h3addfb8b),
	.w5(32'hba305c3e),
	.w6(32'hbab853cb),
	.w7(32'hbb4e675c),
	.w8(32'hbb81380b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f9e9b),
	.w1(32'hbb06e3dd),
	.w2(32'hbade3b9f),
	.w3(32'hb9cdf0cb),
	.w4(32'h39427896),
	.w5(32'h3b277a2b),
	.w6(32'hbb43ae21),
	.w7(32'hbb3232c8),
	.w8(32'h39c9da19),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd9d27),
	.w1(32'h3a5bbf3a),
	.w2(32'h3bb18ebd),
	.w3(32'h3b5ba33d),
	.w4(32'h3b13d206),
	.w5(32'hb9b55d2e),
	.w6(32'h3b270619),
	.w7(32'h3a973eca),
	.w8(32'h3afd7fb8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7d2cb),
	.w1(32'hba482341),
	.w2(32'hb85ca7ed),
	.w3(32'hba59dd72),
	.w4(32'h3a5a573e),
	.w5(32'hba84a084),
	.w6(32'hbb95fcb0),
	.w7(32'hbb236c27),
	.w8(32'hbba3c960),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70fb93),
	.w1(32'hbba4441c),
	.w2(32'hbb8fc1f0),
	.w3(32'hbaba5ef5),
	.w4(32'hbb87412e),
	.w5(32'hbad90ea1),
	.w6(32'hbb843895),
	.w7(32'hbbb87ad5),
	.w8(32'hbac82769),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ac959d),
	.w1(32'hba470ce4),
	.w2(32'h3a27ee4e),
	.w3(32'hbae42aa5),
	.w4(32'hbb07a4d1),
	.w5(32'h3b2aa522),
	.w6(32'hb9d6a45d),
	.w7(32'hb94d1573),
	.w8(32'h3b693d94),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c182a),
	.w1(32'h3b837cbf),
	.w2(32'h3b7b248e),
	.w3(32'h3b920e1f),
	.w4(32'h3b62c274),
	.w5(32'hbacaf5a9),
	.w6(32'h3b6c257b),
	.w7(32'h3b6d252d),
	.w8(32'hba84120e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f09fb),
	.w1(32'h3a3fb198),
	.w2(32'h3a3c5174),
	.w3(32'hba477c31),
	.w4(32'hb9ea1dc8),
	.w5(32'h3af3f0e0),
	.w6(32'h3acd3f40),
	.w7(32'h3a3e1630),
	.w8(32'h3abb6315),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02b452),
	.w1(32'h3a9f0db0),
	.w2(32'h3a93fc04),
	.w3(32'h3a8338d8),
	.w4(32'h3aab6564),
	.w5(32'hba9a1fb9),
	.w6(32'h3a9ce2b9),
	.w7(32'h3a5434a2),
	.w8(32'h3a00b1c0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee3abe),
	.w1(32'hbacc6cb3),
	.w2(32'hbb91c179),
	.w3(32'hbaa7cf10),
	.w4(32'h394d2a83),
	.w5(32'hba58aa5b),
	.w6(32'hbaa59e60),
	.w7(32'hbbba3104),
	.w8(32'hbbadc216),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a927165),
	.w1(32'h3b07d641),
	.w2(32'h3a8b7b7e),
	.w3(32'h3aaf21f1),
	.w4(32'h3abda1ce),
	.w5(32'h394041a4),
	.w6(32'h38e50f7c),
	.w7(32'h3a06fea4),
	.w8(32'hba12a4b1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1261cb),
	.w1(32'h3abfafb5),
	.w2(32'h3b732fd3),
	.w3(32'hb9f5d4b1),
	.w4(32'h3b6e7664),
	.w5(32'h3b22f6aa),
	.w6(32'h3a672216),
	.w7(32'h3adc35d4),
	.w8(32'hbb0ded95),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82cdd6),
	.w1(32'hb9580703),
	.w2(32'hbadb8162),
	.w3(32'hbb7cedb1),
	.w4(32'hbb800b5f),
	.w5(32'h3baaef48),
	.w6(32'hbbd041e6),
	.w7(32'hbb79c1a4),
	.w8(32'h3ac08578),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3bf34),
	.w1(32'h3b1b2da1),
	.w2(32'h3b02ad83),
	.w3(32'h3a04316a),
	.w4(32'h3a90a51c),
	.w5(32'hbb790248),
	.w6(32'h39726015),
	.w7(32'h3b52da55),
	.w8(32'hbb847b99),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5fa3b),
	.w1(32'hb9a5c5e4),
	.w2(32'h39453b0a),
	.w3(32'h3b8a75c2),
	.w4(32'hbaa021f7),
	.w5(32'h3b99503a),
	.w6(32'h3ad4b35b),
	.w7(32'hbb21fff7),
	.w8(32'h3b638872),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2cca8),
	.w1(32'hbb624275),
	.w2(32'hbb2bb2e0),
	.w3(32'hbb2ca14e),
	.w4(32'hbb02d798),
	.w5(32'hba837e9c),
	.w6(32'hbb70483f),
	.w7(32'hbbb8da05),
	.w8(32'hbb3b3de9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9faab2),
	.w1(32'hbb594e6e),
	.w2(32'hbb386dce),
	.w3(32'hbb0a0799),
	.w4(32'hba97c5c0),
	.w5(32'hbb28ca5e),
	.w6(32'hbb049736),
	.w7(32'hbb827708),
	.w8(32'hbbaf9d8e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb702674),
	.w1(32'hbb2bd3fb),
	.w2(32'h39313b12),
	.w3(32'hbb532ea2),
	.w4(32'hbb32faff),
	.w5(32'h396b5cb4),
	.w6(32'hbb82a019),
	.w7(32'hbb54cc76),
	.w8(32'hbb6784c9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52f8d2),
	.w1(32'hbb5063ae),
	.w2(32'hba7e74ab),
	.w3(32'h3ab4514e),
	.w4(32'h3a55876e),
	.w5(32'hbb19240b),
	.w6(32'hb9d71a83),
	.w7(32'hba9d9f12),
	.w8(32'hbb6a483c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9690f3),
	.w1(32'h3a15c3a5),
	.w2(32'hba8fa3de),
	.w3(32'h3a26a2a8),
	.w4(32'h3a047ffa),
	.w5(32'h3adcb809),
	.w6(32'h3b05e860),
	.w7(32'h3b0e249c),
	.w8(32'hbaf1a7b6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bf66b),
	.w1(32'hba45eae1),
	.w2(32'h3b96039b),
	.w3(32'hbb7aaa41),
	.w4(32'hbab8b710),
	.w5(32'h3c1f5764),
	.w6(32'hbbbe952e),
	.w7(32'hbad6790b),
	.w8(32'h3aacfdf3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb133f7f),
	.w1(32'hbac22acd),
	.w2(32'h3a6af212),
	.w3(32'h3bd11b17),
	.w4(32'h3b8d586b),
	.w5(32'hbc2a845f),
	.w6(32'h3a66584f),
	.w7(32'h3ae4f49d),
	.w8(32'hbbacf960),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93c703),
	.w1(32'hbbaec5e3),
	.w2(32'hbc5acbda),
	.w3(32'hbc47a845),
	.w4(32'hbc08c8fc),
	.w5(32'hbb4ea30c),
	.w6(32'hbabe329d),
	.w7(32'hbc5ab820),
	.w8(32'h3b7d4ba9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94e32f),
	.w1(32'hbb7dfbe2),
	.w2(32'hbc1f59bc),
	.w3(32'hbc0c8657),
	.w4(32'hbc495d7f),
	.w5(32'hbc284573),
	.w6(32'h3b1dd98e),
	.w7(32'hbb46b550),
	.w8(32'hbc814baf),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29e9f2),
	.w1(32'h3b909a84),
	.w2(32'h3bf9f08e),
	.w3(32'h3b98dd66),
	.w4(32'h3a954797),
	.w5(32'hb969c445),
	.w6(32'h3b1340dc),
	.w7(32'hbb70147c),
	.w8(32'hbbfecada),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38d8b2),
	.w1(32'hbb531c2a),
	.w2(32'hbbb33ea4),
	.w3(32'hb8958461),
	.w4(32'hbb2ae7f5),
	.w5(32'hba98b085),
	.w6(32'h3b5ab1d1),
	.w7(32'hbbcf4fba),
	.w8(32'hba4251be),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb817c4b),
	.w1(32'hbb5ac794),
	.w2(32'hbb6e74cb),
	.w3(32'hbb396eea),
	.w4(32'hba705b12),
	.w5(32'h3b22ac3a),
	.w6(32'hba070b1b),
	.w7(32'hba87bf4a),
	.w8(32'h3c0857bf),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ecee9),
	.w1(32'hbc3d8e96),
	.w2(32'hbcb1fb15),
	.w3(32'hbb9f7b83),
	.w4(32'hbc407f98),
	.w5(32'hbb6e1014),
	.w6(32'h3c6a7c23),
	.w7(32'hbc0b7bdc),
	.w8(32'hbb909f8a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af00df6),
	.w1(32'h3b1d820f),
	.w2(32'hbbb21402),
	.w3(32'h3b877e56),
	.w4(32'h390c420f),
	.w5(32'hbc136871),
	.w6(32'h3ba6400b),
	.w7(32'h3aa263e0),
	.w8(32'hbbfdc06d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b5509),
	.w1(32'hb86c9b3f),
	.w2(32'h38c6fcb6),
	.w3(32'hbc259da7),
	.w4(32'hb9e8035b),
	.w5(32'hbaa39d7c),
	.w6(32'h3ad53747),
	.w7(32'hb9c4849c),
	.w8(32'h3bfc1668),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8fc2b),
	.w1(32'h39cc1e38),
	.w2(32'hbbc15ee9),
	.w3(32'h3b87a499),
	.w4(32'hbbad5523),
	.w5(32'h3c1217c0),
	.w6(32'h3cc2c03a),
	.w7(32'h3bf96e62),
	.w8(32'h3b99c594),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b6627),
	.w1(32'h3c0fa235),
	.w2(32'h3c26ceff),
	.w3(32'h3c079e1d),
	.w4(32'h3c1e4015),
	.w5(32'h3c7246f4),
	.w6(32'hba943e06),
	.w7(32'h3b7a5111),
	.w8(32'h3c6b19b7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b9307),
	.w1(32'h3c928ee5),
	.w2(32'h3c653358),
	.w3(32'h3d04d6a6),
	.w4(32'h3c78939a),
	.w5(32'hbbe7879c),
	.w6(32'h3d0a2457),
	.w7(32'h3cb88b53),
	.w8(32'hbbd4ca19),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c365d),
	.w1(32'hba1a6950),
	.w2(32'hbc3b6b8a),
	.w3(32'hbb3c8f66),
	.w4(32'hba2fac71),
	.w5(32'hbbb3a15e),
	.w6(32'h3b6c118a),
	.w7(32'hbafa5e98),
	.w8(32'hba62e03b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c388cb),
	.w1(32'h3baaafc8),
	.w2(32'h3a6915bb),
	.w3(32'hba98d503),
	.w4(32'h3aacabdf),
	.w5(32'h3b9d57a5),
	.w6(32'h3bf8f9c1),
	.w7(32'h3af06594),
	.w8(32'hbb3df6b4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4407d),
	.w1(32'h3bbee8cd),
	.w2(32'h3bb8eaf9),
	.w3(32'hb974cdd6),
	.w4(32'h3b2bc991),
	.w5(32'h3bc42838),
	.w6(32'hbbbb0f53),
	.w7(32'hbb3d0136),
	.w8(32'h3bc06542),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda8c65),
	.w1(32'h3a96ec2c),
	.w2(32'h3af9d3bc),
	.w3(32'h39eedffc),
	.w4(32'h3aea6583),
	.w5(32'h3b8c2844),
	.w6(32'h3b28a134),
	.w7(32'h39944a09),
	.w8(32'hba2ad96e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba72106),
	.w1(32'h3b2990e8),
	.w2(32'h3b312aa3),
	.w3(32'h399fd066),
	.w4(32'h39edb77a),
	.w5(32'hbaa58869),
	.w6(32'h3aa31e07),
	.w7(32'h3ac1ca69),
	.w8(32'hbbcbef22),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fd2a1),
	.w1(32'h3b8723ff),
	.w2(32'h399ba4f6),
	.w3(32'hba2ba97b),
	.w4(32'h3b2f5aa5),
	.w5(32'h39a07fda),
	.w6(32'hbacff378),
	.w7(32'hbb056279),
	.w8(32'hbbba2007),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84cdd5),
	.w1(32'h3a0de495),
	.w2(32'h3c23cf60),
	.w3(32'hbb92a390),
	.w4(32'h3ae8dc8f),
	.w5(32'hbc0122bc),
	.w6(32'hbc22eff9),
	.w7(32'h3b672c5a),
	.w8(32'h39f4dbe1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14944a),
	.w1(32'hbc17bbbe),
	.w2(32'hbbce5ba9),
	.w3(32'hbc0e8a44),
	.w4(32'hbc0ae28a),
	.w5(32'hbba35ca1),
	.w6(32'h3b10917e),
	.w7(32'h3ad81b8f),
	.w8(32'h3ba67e32),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd7288),
	.w1(32'h3be19411),
	.w2(32'hbbaf63f6),
	.w3(32'h3bf19982),
	.w4(32'hbbb0e998),
	.w5(32'h3c4fef96),
	.w6(32'h3c835aff),
	.w7(32'h3bc2e01b),
	.w8(32'h3c308ddd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c5bae),
	.w1(32'h3bc118f5),
	.w2(32'h3bc940ce),
	.w3(32'h3c9b6eb5),
	.w4(32'h3c8ad09e),
	.w5(32'h3b769d43),
	.w6(32'h3c85f837),
	.w7(32'h3c2a4b29),
	.w8(32'hbb29b148),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f3efa),
	.w1(32'h3b0a8b4f),
	.w2(32'h3a72778b),
	.w3(32'hbb8fda80),
	.w4(32'hb9c42c8b),
	.w5(32'hbba69c4c),
	.w6(32'hbb5ff004),
	.w7(32'hba7311b6),
	.w8(32'hbbc5c5e8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b121284),
	.w1(32'hbc509a84),
	.w2(32'hbbb52d4a),
	.w3(32'hbc2e46b2),
	.w4(32'hbb95d25c),
	.w5(32'hba4ea8e9),
	.w6(32'hbc5744d4),
	.w7(32'h3abf1281),
	.w8(32'hbc4334c2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2cff8),
	.w1(32'hbbefc1fc),
	.w2(32'hbc56eb0a),
	.w3(32'h3c573ffe),
	.w4(32'h3c171186),
	.w5(32'hbc418973),
	.w6(32'hbbeb8935),
	.w7(32'hbba6d741),
	.w8(32'hbcaf0151),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc136cb9),
	.w1(32'hbc35528c),
	.w2(32'hba5df8c1),
	.w3(32'hbc0e32c3),
	.w4(32'hbb599a86),
	.w5(32'hb92694df),
	.w6(32'hbc18b9b6),
	.w7(32'hbb964ec0),
	.w8(32'hbbbd631c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48a7d6),
	.w1(32'hbbd48eaf),
	.w2(32'hbc0fe879),
	.w3(32'h3bf5ff8b),
	.w4(32'h3b8b382f),
	.w5(32'hb9b324c2),
	.w6(32'h3bebd474),
	.w7(32'h3bb5406b),
	.w8(32'h3b347787),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5149bf),
	.w1(32'hb8cee0fc),
	.w2(32'h3b29caa1),
	.w3(32'h3ad5458d),
	.w4(32'hbbeb98e6),
	.w5(32'hba6af459),
	.w6(32'h3c21b386),
	.w7(32'h3bbe2477),
	.w8(32'h3a79599f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2fe19),
	.w1(32'hbbc1ed24),
	.w2(32'hbb824f26),
	.w3(32'h3bb3457e),
	.w4(32'h3b1de482),
	.w5(32'hbb8b5bcb),
	.w6(32'h3c30769c),
	.w7(32'h3c219d41),
	.w8(32'hba8848bb),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39124637),
	.w1(32'h3a87ba2f),
	.w2(32'hbbc30f36),
	.w3(32'hbbb449bb),
	.w4(32'hbc024134),
	.w5(32'h3bfebdc6),
	.w6(32'hbb7232cf),
	.w7(32'hbbd38436),
	.w8(32'h3c45b189),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9976674),
	.w1(32'h3b9bd66f),
	.w2(32'hba21a9f6),
	.w3(32'h3c842817),
	.w4(32'h3c493852),
	.w5(32'hba8ecb16),
	.w6(32'h3ce14d54),
	.w7(32'h3c7a8af1),
	.w8(32'hbbd2b369),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a98e4),
	.w1(32'hbbd6814d),
	.w2(32'hbbb6db3b),
	.w3(32'hbae76e27),
	.w4(32'hbc3819c9),
	.w5(32'hbc782ced),
	.w6(32'h39826479),
	.w7(32'hbb867c1f),
	.w8(32'hbbb84118),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb942034),
	.w1(32'h3bab43b5),
	.w2(32'hbb32b78b),
	.w3(32'hbbfce656),
	.w4(32'hbb548675),
	.w5(32'hbb8175e2),
	.w6(32'h3b3b91e5),
	.w7(32'h3acb66f0),
	.w8(32'hbbd3cfcc),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2484f),
	.w1(32'hbc213792),
	.w2(32'hbbf459d6),
	.w3(32'hbc0d0aa5),
	.w4(32'hbbf475ed),
	.w5(32'hbb9fcafa),
	.w6(32'hbbfc26b2),
	.w7(32'hbc2c7f7d),
	.w8(32'hbc1c5e00),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2a4e0),
	.w1(32'hbbf43e2e),
	.w2(32'h3b8d5ee1),
	.w3(32'hbb958f97),
	.w4(32'hbbd75b5e),
	.w5(32'h3c190abf),
	.w6(32'hbc881937),
	.w7(32'hbb59b431),
	.w8(32'h3bc7470e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba206bc),
	.w1(32'h3baf80ea),
	.w2(32'h3b818992),
	.w3(32'h3c34034d),
	.w4(32'h3b3ee4c6),
	.w5(32'hbbedf099),
	.w6(32'h3c43faf1),
	.w7(32'h3bc8aa33),
	.w8(32'hbc371dff),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc811b8e),
	.w1(32'hbc2f1229),
	.w2(32'hbbf53f71),
	.w3(32'hbb9483fc),
	.w4(32'hbc155083),
	.w5(32'h3c2b206d),
	.w6(32'hbb289f57),
	.w7(32'hbb5f6c04),
	.w8(32'h3c2ae342),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c668e70),
	.w1(32'h3bd70689),
	.w2(32'h3be56ba7),
	.w3(32'h3c024d73),
	.w4(32'h3a05e63f),
	.w5(32'hbb2fbe37),
	.w6(32'h39ea5156),
	.w7(32'h3a916c8b),
	.w8(32'hbc0f1a6e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13446e),
	.w1(32'hbb1ea448),
	.w2(32'h3b10a11c),
	.w3(32'hbb319793),
	.w4(32'hba72bf65),
	.w5(32'h3c215c22),
	.w6(32'hbc26d497),
	.w7(32'h3a77e8ce),
	.w8(32'h3b18063b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67e4a8),
	.w1(32'h3b2febe0),
	.w2(32'h3bd150ec),
	.w3(32'h3c589df2),
	.w4(32'h3b910a41),
	.w5(32'hbb2c8828),
	.w6(32'h3c12638b),
	.w7(32'h3bdc8c69),
	.w8(32'hbbe631aa),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59a7c6),
	.w1(32'hb9f64bc3),
	.w2(32'hbae7c547),
	.w3(32'hbb5bdaea),
	.w4(32'hba00b397),
	.w5(32'h3bf532a7),
	.w6(32'hbb4ffb68),
	.w7(32'hbb7ef2c3),
	.w8(32'h3bb4332e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2643f1),
	.w1(32'h3bc21d5b),
	.w2(32'h3b1bf38b),
	.w3(32'h3c1bcfb4),
	.w4(32'h3c02f38c),
	.w5(32'h3b24e5e4),
	.w6(32'h3bc57fc0),
	.w7(32'h3b88cccd),
	.w8(32'hbb6b85e2),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c4673),
	.w1(32'hbb548510),
	.w2(32'h3b6ff424),
	.w3(32'h3b5f76df),
	.w4(32'h3c5ded2a),
	.w5(32'hbc1df1af),
	.w6(32'hbbdc39cb),
	.w7(32'hba630ec7),
	.w8(32'hbc631fe2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0495),
	.w1(32'hbb922049),
	.w2(32'hba91f465),
	.w3(32'h3b17d6ad),
	.w4(32'h39c15fad),
	.w5(32'hbc4791b4),
	.w6(32'hba188345),
	.w7(32'hbb8c5ada),
	.w8(32'hbc5ad4e3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e49c2),
	.w1(32'hbc362d5a),
	.w2(32'hbc5f7d4b),
	.w3(32'hbc1bfb07),
	.w4(32'hbbf85e5f),
	.w5(32'h3b26219f),
	.w6(32'hbbf0545b),
	.w7(32'hbc15043b),
	.w8(32'h3b481bbc),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9be4a1),
	.w1(32'hbbcd26a1),
	.w2(32'hbbb17aad),
	.w3(32'h3b8f4f55),
	.w4(32'hb92812cb),
	.w5(32'hbb07a1b0),
	.w6(32'h3b4ea3a6),
	.w7(32'h3bab8a50),
	.w8(32'h3b9a57c3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc478907),
	.w1(32'hbaf7e766),
	.w2(32'hbc214c60),
	.w3(32'h3c006087),
	.w4(32'hbba8306e),
	.w5(32'hb90433b8),
	.w6(32'h3c92b3bf),
	.w7(32'h3b6805be),
	.w8(32'h3a688882),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a432354),
	.w1(32'h3a8c8534),
	.w2(32'hba80b03c),
	.w3(32'h39b85689),
	.w4(32'hbb0bd553),
	.w5(32'hbbbfb47a),
	.w6(32'h3b0f8ad0),
	.w7(32'h3a927adb),
	.w8(32'h3bdbbb8e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ea98b),
	.w1(32'hbc064b0f),
	.w2(32'hbc1c8e51),
	.w3(32'hbc06df8f),
	.w4(32'hbae90b26),
	.w5(32'hba1badc2),
	.w6(32'h3a76510f),
	.w7(32'h3abe857b),
	.w8(32'hbbbcbe54),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf559d5),
	.w1(32'hbbda0c5e),
	.w2(32'h38c3c0c4),
	.w3(32'h3ba63306),
	.w4(32'hbae091f3),
	.w5(32'h3a3b03ac),
	.w6(32'h3b38352b),
	.w7(32'hbb36f064),
	.w8(32'hbba3bf4b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05c442),
	.w1(32'hbc7745ee),
	.w2(32'hbb1cffb5),
	.w3(32'hbbe34c50),
	.w4(32'h3a62f65c),
	.w5(32'h3be7c30c),
	.w6(32'hbc26e7e0),
	.w7(32'h3c2c1018),
	.w8(32'h3bbaefd4),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c3445),
	.w1(32'h3ba291d7),
	.w2(32'h3c648525),
	.w3(32'h3c1c9692),
	.w4(32'h3bc9bd75),
	.w5(32'hbb0e92ee),
	.w6(32'h3aa00261),
	.w7(32'h3bacd498),
	.w8(32'hbb8f632e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecc06c),
	.w1(32'h36141418),
	.w2(32'h3b0244b6),
	.w3(32'hbb41e91b),
	.w4(32'h3b854b98),
	.w5(32'hbbb62bdf),
	.w6(32'hb9d12faf),
	.w7(32'h3b3ef6db),
	.w8(32'hbc26aa06),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7e588),
	.w1(32'hbc6a0e1d),
	.w2(32'hbbfa05ba),
	.w3(32'h3a52c596),
	.w4(32'hbc006184),
	.w5(32'hba09f8ad),
	.w6(32'h3a5696d6),
	.w7(32'hbbc33a9f),
	.w8(32'hbb19a282),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbd132),
	.w1(32'hbafd18c3),
	.w2(32'h3b091d82),
	.w3(32'h3c24dbc7),
	.w4(32'h3b700982),
	.w5(32'hbbf0b0fa),
	.w6(32'h3b2e4819),
	.w7(32'hbb8a6402),
	.w8(32'hba48dfaf),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf71806),
	.w1(32'h3b4133b2),
	.w2(32'hbc088f09),
	.w3(32'hbaafd6ca),
	.w4(32'hbb9cdb80),
	.w5(32'hbba30625),
	.w6(32'h3cb94a55),
	.w7(32'h3c155fcb),
	.w8(32'h3898a192),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae91bce),
	.w1(32'hbc010ef2),
	.w2(32'hbc21f53d),
	.w3(32'hbc26e9cf),
	.w4(32'hbc45c4c9),
	.w5(32'h3bc98a2f),
	.w6(32'hbb654386),
	.w7(32'hbbde4f99),
	.w8(32'h3c0a34fb),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b308bad),
	.w1(32'h3c46ebd4),
	.w2(32'h3c5da38c),
	.w3(32'h3c92844b),
	.w4(32'h3c5efb68),
	.w5(32'hbbac41ba),
	.w6(32'h3cab7ce6),
	.w7(32'h3ca2eeab),
	.w8(32'hbbc19aef),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb997e90),
	.w1(32'hbbbc1778),
	.w2(32'hbbd9cef1),
	.w3(32'hba885166),
	.w4(32'hbc13a71e),
	.w5(32'hbb67727a),
	.w6(32'h3b00d49d),
	.w7(32'hb98eae18),
	.w8(32'hbc05ac46),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4852ac),
	.w1(32'hbbbc9a93),
	.w2(32'hbb3eea02),
	.w3(32'hbb76c2fb),
	.w4(32'hba0cc983),
	.w5(32'h3c0a1825),
	.w6(32'h3a8acd98),
	.w7(32'h3b090684),
	.w8(32'hba4863ae),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c338d9f),
	.w1(32'h3c378c27),
	.w2(32'h3ca96130),
	.w3(32'h3c3853a7),
	.w4(32'h3bd4d0c9),
	.w5(32'h3c637f6f),
	.w6(32'h3b28686b),
	.w7(32'h3b9802e2),
	.w8(32'h3c056c6f),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00641c),
	.w1(32'h3b05d31f),
	.w2(32'h3c16b4ea),
	.w3(32'h3c592cdd),
	.w4(32'h3cbdc6ae),
	.w5(32'hbba37690),
	.w6(32'h3c053118),
	.w7(32'h3c513c48),
	.w8(32'hb9534eb1),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d781a),
	.w1(32'hbb15949a),
	.w2(32'hbc0054b2),
	.w3(32'hbb495e2e),
	.w4(32'hbad2fc28),
	.w5(32'hbb8e0fee),
	.w6(32'h3b56f807),
	.w7(32'hbb95b0f4),
	.w8(32'hbbdd2edb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd5d6e),
	.w1(32'hbb5ab2db),
	.w2(32'hbb0d6eec),
	.w3(32'h3a8006b3),
	.w4(32'hbbde8be8),
	.w5(32'hbb6ccebe),
	.w6(32'hb9b2d552),
	.w7(32'hbb53ac4c),
	.w8(32'hb9da564f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de2ad4),
	.w1(32'h3a27802f),
	.w2(32'h39f36e6c),
	.w3(32'hbb3344cd),
	.w4(32'h3a2cfeff),
	.w5(32'hba2475e8),
	.w6(32'hbaaa6171),
	.w7(32'hbb076dda),
	.w8(32'hbb61ff96),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b3820),
	.w1(32'hba5bbb94),
	.w2(32'hbb83e6b6),
	.w3(32'hbba78769),
	.w4(32'h3b12c742),
	.w5(32'h3b00b4a3),
	.w6(32'hbb406c87),
	.w7(32'h3b11ee87),
	.w8(32'h3be87682),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f6ff2),
	.w1(32'h3b74d5f9),
	.w2(32'hbad54f61),
	.w3(32'h3b88b36a),
	.w4(32'hba536b4f),
	.w5(32'hbb932e7a),
	.w6(32'h3bd5e895),
	.w7(32'hba0a19bf),
	.w8(32'hbb86e4c9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb68a25),
	.w1(32'h3c34338e),
	.w2(32'h3bbba86a),
	.w3(32'h3b41cf76),
	.w4(32'hbb88259b),
	.w5(32'h3b3bc0de),
	.w6(32'h3c639559),
	.w7(32'h3b8fdcba),
	.w8(32'hbc0d098f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc57958),
	.w1(32'hbb89c8ae),
	.w2(32'hb9668696),
	.w3(32'h3bbdc7ef),
	.w4(32'hb90baf1c),
	.w5(32'hbb1e45d2),
	.w6(32'hbbc6fff9),
	.w7(32'hbbf2065f),
	.w8(32'h3ac58354),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8469c),
	.w1(32'hb9bc2ea5),
	.w2(32'hbb1154af),
	.w3(32'h3a6e96c2),
	.w4(32'hbbc3ecb2),
	.w5(32'h3acb17c1),
	.w6(32'h3b9fa20c),
	.w7(32'hbb83eb40),
	.w8(32'hb92af3e4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cbab8),
	.w1(32'h3bbe88fe),
	.w2(32'h3b5598c2),
	.w3(32'hbad90527),
	.w4(32'h3b07b35f),
	.w5(32'h3b112c92),
	.w6(32'hbc0bd8c8),
	.w7(32'hbc226e42),
	.w8(32'h3a0120df),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e65f5),
	.w1(32'hbbc6688b),
	.w2(32'hbc70ef6e),
	.w3(32'h3ad695e2),
	.w4(32'hbbeaf811),
	.w5(32'h3c53939e),
	.w6(32'h3c7c4a09),
	.w7(32'h3b690ee6),
	.w8(32'h3c314146),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f51b7),
	.w1(32'h3bc81489),
	.w2(32'h3ba2a1d2),
	.w3(32'h3bc6fe78),
	.w4(32'h3c0f8e63),
	.w5(32'h3b4a79ec),
	.w6(32'h3c0ca014),
	.w7(32'h3c2b468a),
	.w8(32'h3b4ae9e4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399aa06e),
	.w1(32'hbaa2ad12),
	.w2(32'hbb906bfe),
	.w3(32'h3ac5bc9f),
	.w4(32'hbbcaea1a),
	.w5(32'hbadf8c76),
	.w6(32'h3b4d8cef),
	.w7(32'h3ac117a4),
	.w8(32'h3b338b61),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37a28d),
	.w1(32'hbc892682),
	.w2(32'hbba83685),
	.w3(32'hba4df80d),
	.w4(32'hba19290d),
	.w5(32'h3bac2b7d),
	.w6(32'hba2ba196),
	.w7(32'hba22a5e0),
	.w8(32'h3c06851b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48625c),
	.w1(32'hba0cba02),
	.w2(32'h3a8ee6ea),
	.w3(32'h3c2f6ff1),
	.w4(32'h3bc61c3f),
	.w5(32'hbc19178f),
	.w6(32'h3ce6f2cb),
	.w7(32'h3c9a57b8),
	.w8(32'hbc4a9c06),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc400b37),
	.w1(32'hbc08eda4),
	.w2(32'hbbcce349),
	.w3(32'hbbb81146),
	.w4(32'hbbdcd5de),
	.w5(32'h3bc8f122),
	.w6(32'hbbf97e63),
	.w7(32'hbc3beb96),
	.w8(32'hbbf1f022),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f32e9),
	.w1(32'hba6d6e27),
	.w2(32'h3c0d7c76),
	.w3(32'h3b198bc6),
	.w4(32'h3c044aa8),
	.w5(32'hbbd82045),
	.w6(32'hbc20fe76),
	.w7(32'h3b28003d),
	.w8(32'hbbed02af),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f50bc),
	.w1(32'hbc6f1eb1),
	.w2(32'hbc408e55),
	.w3(32'hbbec19b1),
	.w4(32'hbb16e682),
	.w5(32'hba244dd0),
	.w6(32'hbc2907c9),
	.w7(32'hbc03a473),
	.w8(32'h39238d1d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40fa49),
	.w1(32'h3b2a16b0),
	.w2(32'h3b2a79b9),
	.w3(32'h3b9c9974),
	.w4(32'hba6919ae),
	.w5(32'h3bd520f4),
	.w6(32'h3c104c4a),
	.w7(32'h3bb3812e),
	.w8(32'hbae8fd1d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8d741),
	.w1(32'h3ba71a5d),
	.w2(32'h3b8de7cf),
	.w3(32'h3b6cc409),
	.w4(32'hba1de85d),
	.w5(32'hb9ec4d08),
	.w6(32'hbb84617b),
	.w7(32'h3a7a04f7),
	.w8(32'h3b93acf0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65e07d),
	.w1(32'hbb97faae),
	.w2(32'hbb82113e),
	.w3(32'hbbb56e1d),
	.w4(32'hbbd38631),
	.w5(32'hbbbab7e9),
	.w6(32'h3aecbeb7),
	.w7(32'h3ad95b05),
	.w8(32'h38252364),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba158883),
	.w1(32'h3b4b5a17),
	.w2(32'hbb7dfc84),
	.w3(32'hbbd50980),
	.w4(32'h3b3ef9be),
	.w5(32'h36a0496c),
	.w6(32'h3ade0359),
	.w7(32'hbb1d0921),
	.w8(32'h3bd9693b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba59c5b),
	.w1(32'hbadb82f7),
	.w2(32'hb9b48a3e),
	.w3(32'hbb6f5327),
	.w4(32'hbb8c6fd9),
	.w5(32'hb9b303fd),
	.w6(32'h3c164e8d),
	.w7(32'h390ae93a),
	.w8(32'hb98914cb),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc18367),
	.w1(32'h3aefcffc),
	.w2(32'h3b335000),
	.w3(32'h3a6d1a6f),
	.w4(32'hbb8f9052),
	.w5(32'hbb1db689),
	.w6(32'h3bbceada),
	.w7(32'hba23ba2a),
	.w8(32'hbba9431b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb183bc7),
	.w1(32'h3aa81188),
	.w2(32'h3b34ae8a),
	.w3(32'hbab21b92),
	.w4(32'hbbfc2657),
	.w5(32'h3be82a93),
	.w6(32'h3a7571d0),
	.w7(32'hba43b925),
	.w8(32'h3ba46491),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b370480),
	.w1(32'h3a8911a9),
	.w2(32'h3bfe8b28),
	.w3(32'h3b2a21d9),
	.w4(32'h3b95d71a),
	.w5(32'h3b8cdc28),
	.w6(32'hbba88435),
	.w7(32'hbac344c0),
	.w8(32'h3bb23e3f),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e33dd),
	.w1(32'h3b41b800),
	.w2(32'hbad1bb6b),
	.w3(32'h3b15f7b3),
	.w4(32'h3b0cb27e),
	.w5(32'hbc1c1fc9),
	.w6(32'h3c19321a),
	.w7(32'hbaa78914),
	.w8(32'hbc0ebc22),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d0620),
	.w1(32'hbad3e0f1),
	.w2(32'hbad98061),
	.w3(32'hba652c85),
	.w4(32'hbad63d87),
	.w5(32'h3bbbd943),
	.w6(32'h3b85a34d),
	.w7(32'h3bbfeee5),
	.w8(32'h3c146933),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba712892),
	.w1(32'hbc56f8a0),
	.w2(32'hbc2db276),
	.w3(32'hbba12a00),
	.w4(32'hbcae3863),
	.w5(32'h3b3a0edf),
	.w6(32'hbca3fe93),
	.w7(32'hbd0aea0c),
	.w8(32'hbc5f7955),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74e9e4),
	.w1(32'hbb2d5e12),
	.w2(32'h3bca3a0f),
	.w3(32'h3bb4ee52),
	.w4(32'h3be080e0),
	.w5(32'h3a17df88),
	.w6(32'hbbc9ec8b),
	.w7(32'h3bf2e744),
	.w8(32'h3b04887c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8d54b),
	.w1(32'hbb070cbd),
	.w2(32'hbba87831),
	.w3(32'h3bdb9784),
	.w4(32'h3bbb53c4),
	.w5(32'hba9bb4f8),
	.w6(32'h3c6d3c72),
	.w7(32'h3ba98b0e),
	.w8(32'hbab307b3),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc2879),
	.w1(32'hba743712),
	.w2(32'h3aa350ac),
	.w3(32'hb8a063d7),
	.w4(32'hbb08cc08),
	.w5(32'hbb01c9e5),
	.w6(32'hba7c2088),
	.w7(32'hb9345db8),
	.w8(32'hbbaed636),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04bef9),
	.w1(32'hb872aaa4),
	.w2(32'hb986b8ac),
	.w3(32'hba9f98b5),
	.w4(32'hbb126a61),
	.w5(32'h3b751439),
	.w6(32'hb9eb8c38),
	.w7(32'hb940b19c),
	.w8(32'hbb86e91a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3987c),
	.w1(32'h39fa4e18),
	.w2(32'h3b84c41b),
	.w3(32'h3b8cd1a2),
	.w4(32'hbb1c332d),
	.w5(32'hbbcbac87),
	.w6(32'h3bc4585e),
	.w7(32'h3b62ed3e),
	.w8(32'hbb766d3d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb677adb),
	.w1(32'hbacd114f),
	.w2(32'hbbb8c97f),
	.w3(32'hbb950768),
	.w4(32'hbb99bfb7),
	.w5(32'hb90efbd1),
	.w6(32'hbab15eb7),
	.w7(32'hbbe177fe),
	.w8(32'h3c0ffe52),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c015a),
	.w1(32'h3aa2f549),
	.w2(32'hbc19b86f),
	.w3(32'hbb7d6c2d),
	.w4(32'hbbb72227),
	.w5(32'h3afab0f7),
	.w6(32'h3bf18abd),
	.w7(32'hbbd0e5ce),
	.w8(32'hba9e5d04),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba890ea4),
	.w1(32'hbc246162),
	.w2(32'hbb9a3c46),
	.w3(32'hbaef196a),
	.w4(32'hbbfcf65b),
	.w5(32'h3bb24bd2),
	.w6(32'hbc466b99),
	.w7(32'hbc15d8f2),
	.w8(32'h39b07b65),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7335ef),
	.w1(32'hb9d6af46),
	.w2(32'hbb9b7b8d),
	.w3(32'hba16a354),
	.w4(32'hbbfa7c96),
	.w5(32'h3a20ce4f),
	.w6(32'h3c04aa85),
	.w7(32'hba96ff84),
	.w8(32'h38deca0a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a8eff),
	.w1(32'hbb6ab13b),
	.w2(32'hbaed5e99),
	.w3(32'hbb18ea7c),
	.w4(32'hb835e9a0),
	.w5(32'hbba768f6),
	.w6(32'hbc04c16e),
	.w7(32'hbb3a9e9b),
	.w8(32'hbb8254db),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb868130),
	.w1(32'hbbc3f0b7),
	.w2(32'hbbe7e49c),
	.w3(32'hbb378199),
	.w4(32'hbb5ee0f7),
	.w5(32'h3b7f4c0a),
	.w6(32'h3b34c9c4),
	.w7(32'hbab79666),
	.w8(32'h3b2434d4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e022e),
	.w1(32'hbb2a9b96),
	.w2(32'h3b227047),
	.w3(32'h3a217041),
	.w4(32'h39b8a499),
	.w5(32'h3c2b3822),
	.w6(32'hbaa0ce19),
	.w7(32'h3b6ada1b),
	.w8(32'h3b1668b7),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa8b97),
	.w1(32'hbb2fe358),
	.w2(32'hbbd02be8),
	.w3(32'h3be0c87e),
	.w4(32'h3c12cd0e),
	.w5(32'hb9a69e87),
	.w6(32'h3b676528),
	.w7(32'hbbad6b78),
	.w8(32'hbb33d978),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a871a3b),
	.w1(32'hbb85e67f),
	.w2(32'hba4aaec7),
	.w3(32'h3bb81daa),
	.w4(32'h3ab1fc92),
	.w5(32'h3b9a04bf),
	.w6(32'hba135a12),
	.w7(32'h3ba44140),
	.w8(32'h3bc82a6e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba945d),
	.w1(32'h3ba9f7fa),
	.w2(32'hbc5e3ecc),
	.w3(32'h3c5c4abc),
	.w4(32'h3a804d79),
	.w5(32'h3bdefca6),
	.w6(32'h3c934ec0),
	.w7(32'hbb81f434),
	.w8(32'hbaa47fd2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0304b4),
	.w1(32'h3a3b9686),
	.w2(32'h3b42d7f3),
	.w3(32'h3b9c6c91),
	.w4(32'h3c398d96),
	.w5(32'hbc169868),
	.w6(32'hbb901c90),
	.w7(32'hb92edc34),
	.w8(32'hbc4405e3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb79edf),
	.w1(32'h3a6e8551),
	.w2(32'h396af198),
	.w3(32'hbbaa1a87),
	.w4(32'h39ef4a6c),
	.w5(32'hb9c7d51d),
	.w6(32'hbbc47849),
	.w7(32'hbba94e0b),
	.w8(32'hbb51c447),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dcde85),
	.w1(32'hbafba786),
	.w2(32'hbb24934e),
	.w3(32'hbb770c4d),
	.w4(32'hbae77542),
	.w5(32'hbb5fbcc5),
	.w6(32'hba7cd02d),
	.w7(32'hbb2c412e),
	.w8(32'hbbc1d1ac),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56f512),
	.w1(32'h3b32f590),
	.w2(32'h3a307d20),
	.w3(32'hbb046106),
	.w4(32'h3bc658c2),
	.w5(32'hbbd9341f),
	.w6(32'hbb9b3018),
	.w7(32'hb978354f),
	.w8(32'hbb95503e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9f718),
	.w1(32'hbb0848b3),
	.w2(32'hb88fddc4),
	.w3(32'h3a6f42de),
	.w4(32'hbb9c686f),
	.w5(32'hbb67e200),
	.w6(32'h3b928226),
	.w7(32'hb9e3fe63),
	.w8(32'hbc03c583),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb64d97),
	.w1(32'hbc3831ee),
	.w2(32'hbb261355),
	.w3(32'hbb8f5702),
	.w4(32'hbc2bee0d),
	.w5(32'h3be798e2),
	.w6(32'hbc92aa02),
	.w7(32'hbc8e2424),
	.w8(32'h3b2a73c8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369ab277),
	.w1(32'hbae6d1fa),
	.w2(32'hbb2adbfb),
	.w3(32'h3bb31fb3),
	.w4(32'h3b8ccb37),
	.w5(32'h3b90942a),
	.w6(32'h3bcb2313),
	.w7(32'h3bc4ae02),
	.w8(32'hbb0995f7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28a3ef),
	.w1(32'hbad02f7c),
	.w2(32'hbb7cf951),
	.w3(32'h39cad698),
	.w4(32'h3ba7d0a7),
	.w5(32'hbc04c687),
	.w6(32'h3aa3907a),
	.w7(32'hbb2e777b),
	.w8(32'hbbaf874e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb482c1b),
	.w1(32'hbbe62c44),
	.w2(32'hbc3d0002),
	.w3(32'hbc167de8),
	.w4(32'hbc3bd9e4),
	.w5(32'h3b41088f),
	.w6(32'hbbde13da),
	.w7(32'hbc363a2f),
	.w8(32'hba963e3a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3a236),
	.w1(32'hbba01c6e),
	.w2(32'hba4e1c8a),
	.w3(32'hbbbd2420),
	.w4(32'h3b310cb2),
	.w5(32'h3a19afa8),
	.w6(32'hbbcf5c8f),
	.w7(32'hbbb50682),
	.w8(32'hbbc04350),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1feb58),
	.w1(32'hbbce5b60),
	.w2(32'hba8c72d7),
	.w3(32'h3c03e2a8),
	.w4(32'h3c33bcd5),
	.w5(32'h3ad86ead),
	.w6(32'h3c54d35d),
	.w7(32'h3c7730fc),
	.w8(32'hb9d77b8a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdb2a4),
	.w1(32'h3b0c7e9a),
	.w2(32'hba1904fd),
	.w3(32'h3be86801),
	.w4(32'hbbdc0e71),
	.w5(32'hbbc48441),
	.w6(32'h3c960106),
	.w7(32'hbaa7a26c),
	.w8(32'h3bc0e765),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90e9f0),
	.w1(32'hbb0358f7),
	.w2(32'h38c1bdd1),
	.w3(32'hbbb847db),
	.w4(32'hbc18ac9c),
	.w5(32'hba22c312),
	.w6(32'h3aebfb8e),
	.w7(32'h3b075fd9),
	.w8(32'h3b894a1d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3969eb),
	.w1(32'h3a85618b),
	.w2(32'h3a1a2f46),
	.w3(32'h3981ce6e),
	.w4(32'hbb534430),
	.w5(32'hbbcd5569),
	.w6(32'h3bfb84b9),
	.w7(32'h3be20eff),
	.w8(32'hbbc715a5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2fa1a),
	.w1(32'h3a57fd68),
	.w2(32'hbbd8e9e3),
	.w3(32'hbb2b62e1),
	.w4(32'hbb8829ab),
	.w5(32'hbc81fea7),
	.w6(32'h3c548eb4),
	.w7(32'h3a075eb6),
	.w8(32'hbc90d0db),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe85230),
	.w1(32'hbc0e9564),
	.w2(32'h39f37411),
	.w3(32'hbb189f3a),
	.w4(32'hbbdfdc99),
	.w5(32'hbb5f71cd),
	.w6(32'h3a8107b3),
	.w7(32'hbad6d33a),
	.w8(32'hbbc7a6bd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba03742),
	.w1(32'hbc064929),
	.w2(32'hbbde74df),
	.w3(32'hbbedc39e),
	.w4(32'hbbfb6cde),
	.w5(32'hba5a2b9a),
	.w6(32'hbc36ec48),
	.w7(32'hbbc5881c),
	.w8(32'h3b3ef4b7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37f4ce),
	.w1(32'hb9b61033),
	.w2(32'h3abb15e5),
	.w3(32'hba629e1b),
	.w4(32'hb9233c73),
	.w5(32'hbb99c275),
	.w6(32'hba9f3223),
	.w7(32'hbaf3c264),
	.w8(32'h3ba4844c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd78741),
	.w1(32'h3c4f3059),
	.w2(32'hbc43fcf4),
	.w3(32'h3c4352c1),
	.w4(32'hbc5fd0d2),
	.w5(32'h3ac0ce8e),
	.w6(32'h3ca75fd1),
	.w7(32'hbbc728e8),
	.w8(32'h3a3b5f4d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5a2b9),
	.w1(32'h3c26d5f9),
	.w2(32'h3c1c7aaf),
	.w3(32'h3ba287f5),
	.w4(32'h3bb5faad),
	.w5(32'h3a5c8ddd),
	.w6(32'h3c43c37b),
	.w7(32'h3c488879),
	.w8(32'h3b2fb0cd),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f1f12),
	.w1(32'h3ab3fee9),
	.w2(32'hbab44a9b),
	.w3(32'h3ad83a52),
	.w4(32'hbb204644),
	.w5(32'h3bd15901),
	.w6(32'h3bfdc93c),
	.w7(32'h3b8e63c9),
	.w8(32'hbb04f0c6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f1d4e),
	.w1(32'h3a218b41),
	.w2(32'h3ac8247e),
	.w3(32'h3b2c1e4f),
	.w4(32'h3b78e3b7),
	.w5(32'hbb2a311b),
	.w6(32'hbbaf1f8b),
	.w7(32'hb85d4dd8),
	.w8(32'h3bba94bc),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83ae0e),
	.w1(32'h3ae25a5b),
	.w2(32'hb98daa33),
	.w3(32'h3bd45f6f),
	.w4(32'hbbe426b0),
	.w5(32'hbb2bf643),
	.w6(32'h3bd10bc8),
	.w7(32'hb895a89a),
	.w8(32'hbb14c966),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad92c9e),
	.w1(32'hbba416cc),
	.w2(32'hbb728da0),
	.w3(32'hbbddb6f3),
	.w4(32'hbb73f0ef),
	.w5(32'hbbd2e011),
	.w6(32'hbbb66800),
	.w7(32'hbb7e8bf4),
	.w8(32'hbbc95b97),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc845dca),
	.w1(32'hbc900ed6),
	.w2(32'hbbfa7547),
	.w3(32'hbc4bb1d5),
	.w4(32'hbbd62166),
	.w5(32'hba851a94),
	.w6(32'hbc00a2a4),
	.w7(32'hbbf152ea),
	.w8(32'hbc05b3c0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4050b8),
	.w1(32'h38447d0d),
	.w2(32'hbab2eea8),
	.w3(32'h39b8c377),
	.w4(32'hba800b23),
	.w5(32'h3ac93aec),
	.w6(32'hbbcacd98),
	.w7(32'hbb77a3d4),
	.w8(32'h3b165a07),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b0fcd1),
	.w1(32'h3a88471c),
	.w2(32'h3ab001b1),
	.w3(32'hba6351d2),
	.w4(32'h398a9f7b),
	.w5(32'h3b39df36),
	.w6(32'h3b82b64d),
	.w7(32'hbc0411df),
	.w8(32'h3b049ac5),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ce8e3),
	.w1(32'hbc06c38a),
	.w2(32'hbb9317e8),
	.w3(32'hbb25ecee),
	.w4(32'hbb920a29),
	.w5(32'h3a501980),
	.w6(32'hbb4c1561),
	.w7(32'hbba995af),
	.w8(32'h3c116815),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90db31),
	.w1(32'h3b324ba8),
	.w2(32'h3b5e86bf),
	.w3(32'h3c70ab9f),
	.w4(32'h3c154b1c),
	.w5(32'hba969ffd),
	.w6(32'h3b9fde2c),
	.w7(32'h3bdfa6ea),
	.w8(32'hbaed5af8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06cfd3),
	.w1(32'hbaf718d0),
	.w2(32'hba36066a),
	.w3(32'hbace4b40),
	.w4(32'hba9a23ad),
	.w5(32'hb7e351b8),
	.w6(32'h3b3bfc6a),
	.w7(32'hbbbec139),
	.w8(32'hbb8354ec),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22f0d3),
	.w1(32'hbbbdd0aa),
	.w2(32'hb948a142),
	.w3(32'hbb040cc6),
	.w4(32'hbb90462d),
	.w5(32'hb9003cb7),
	.w6(32'hbbbfb0b3),
	.w7(32'hbb8c7c0f),
	.w8(32'hbb41014b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb887264),
	.w1(32'h3ae95c1a),
	.w2(32'hbb7e9145),
	.w3(32'hb92a39e2),
	.w4(32'hbada6f47),
	.w5(32'h3b880794),
	.w6(32'h3c2896f9),
	.w7(32'hbb692ca1),
	.w8(32'hb9a7ab27),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1aa0af),
	.w1(32'hbb9e9770),
	.w2(32'h3b13a8aa),
	.w3(32'hb8339198),
	.w4(32'hb9cd7224),
	.w5(32'hb9bcc6c5),
	.w6(32'hbaa4bedb),
	.w7(32'h3aed9f55),
	.w8(32'h394b0f18),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb166f86),
	.w1(32'hbb6cb547),
	.w2(32'h3b154f9a),
	.w3(32'hbbe2affa),
	.w4(32'hbbbff4a2),
	.w5(32'h3bf246d7),
	.w6(32'hbb0b04ee),
	.w7(32'hbab67470),
	.w8(32'h3b8c6530),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b462be3),
	.w1(32'hbb8a4356),
	.w2(32'h3ae7f7d9),
	.w3(32'hb992f960),
	.w4(32'hba978960),
	.w5(32'hbbf4f9e7),
	.w6(32'hbc26d6ee),
	.w7(32'hbbea3092),
	.w8(32'hbc6fcff1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc023adc),
	.w1(32'hbc611c07),
	.w2(32'hbc101f1b),
	.w3(32'hbc78d1d8),
	.w4(32'hbc0afb74),
	.w5(32'hbb641754),
	.w6(32'hbc94619b),
	.w7(32'hbc54b6c4),
	.w8(32'hbb014c61),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c8937),
	.w1(32'hbc17174d),
	.w2(32'h3c01fdc0),
	.w3(32'h3bf89644),
	.w4(32'h3be405eb),
	.w5(32'h3b68bb90),
	.w6(32'h3b798e54),
	.w7(32'h3b35b910),
	.w8(32'hbba90e52),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe01caa),
	.w1(32'hbaccdbb1),
	.w2(32'hbace35b6),
	.w3(32'hbc029ab5),
	.w4(32'hbb956942),
	.w5(32'h3b5c6336),
	.w6(32'hbc1c7dfc),
	.w7(32'hbbc7eeff),
	.w8(32'hbb02fdd1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bfc43),
	.w1(32'h3b1ad984),
	.w2(32'h3c41d85d),
	.w3(32'h3a9b6c21),
	.w4(32'hbb9325c5),
	.w5(32'hbbb50d8a),
	.w6(32'hbc141ae3),
	.w7(32'hbb13fb6b),
	.w8(32'h3afcfd29),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07fea6),
	.w1(32'hbb8cae79),
	.w2(32'h3b876c90),
	.w3(32'hbc49ba3f),
	.w4(32'hbb55862d),
	.w5(32'hbaee1c5e),
	.w6(32'hbc80f33d),
	.w7(32'hb95c19ca),
	.w8(32'h3b68e582),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62005c),
	.w1(32'hbbbe15b8),
	.w2(32'h3b263b3d),
	.w3(32'h3b0de098),
	.w4(32'h3a15f02e),
	.w5(32'h3b7e8227),
	.w6(32'h3c61b995),
	.w7(32'hbb024da4),
	.w8(32'h3afd0c3f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398227f3),
	.w1(32'hbab49f63),
	.w2(32'h3ae61415),
	.w3(32'h39ba3b8d),
	.w4(32'hba633b17),
	.w5(32'hbbf8f638),
	.w6(32'h3a55247c),
	.w7(32'h3a225ea6),
	.w8(32'hbb9af8c6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb292f0e),
	.w1(32'h39c2b9ae),
	.w2(32'hbb7940f7),
	.w3(32'hbbab089f),
	.w4(32'h3b0125f3),
	.w5(32'h3afc173d),
	.w6(32'hbc0f0873),
	.w7(32'hbbdaf33c),
	.w8(32'h392e67d1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7994e),
	.w1(32'hba2ca7e3),
	.w2(32'h3a684ea1),
	.w3(32'hbb857b46),
	.w4(32'h3b410ba9),
	.w5(32'hbb9bea8e),
	.w6(32'hbb80445f),
	.w7(32'hb6f87111),
	.w8(32'hbb6f79b2),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cad93),
	.w1(32'hbc4fd7b4),
	.w2(32'hbc5a9ecf),
	.w3(32'hbc486edd),
	.w4(32'hbb1fb20b),
	.w5(32'hbb367895),
	.w6(32'hbc9568d6),
	.w7(32'hbc2e010e),
	.w8(32'hb8b3d477),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d8c34),
	.w1(32'h3b545c7e),
	.w2(32'h3ab3ee2f),
	.w3(32'h3bab047c),
	.w4(32'h3b4be335),
	.w5(32'h3b4a3fec),
	.w6(32'h3c636171),
	.w7(32'h3adaf277),
	.w8(32'h378a0609),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82b859),
	.w1(32'hbb5d57bf),
	.w2(32'hbb4ae278),
	.w3(32'hbaecd4f4),
	.w4(32'hba0ba2a0),
	.w5(32'h3adb0fc8),
	.w6(32'h39e736e8),
	.w7(32'hbad0fe2e),
	.w8(32'h3b92eded),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6cbc3),
	.w1(32'h3b1789b4),
	.w2(32'hbb85f771),
	.w3(32'h3b89e2cd),
	.w4(32'hbac287ef),
	.w5(32'h3b3c9356),
	.w6(32'hba280df3),
	.w7(32'hbbee646d),
	.w8(32'h3a782f37),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99a3e4),
	.w1(32'hbb337653),
	.w2(32'hbb67c398),
	.w3(32'hbb967018),
	.w4(32'hbb6c9a5a),
	.w5(32'h3bb2a80d),
	.w6(32'hbc731dd2),
	.w7(32'hbbb7f8e0),
	.w8(32'hbb035886),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c098a4e),
	.w1(32'h3baf8db7),
	.w2(32'h3bbf1ea3),
	.w3(32'h3be25357),
	.w4(32'hbacf91a8),
	.w5(32'h3b554146),
	.w6(32'hbc0e47a7),
	.w7(32'hbbabf261),
	.w8(32'hbac099cc),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad09bf),
	.w1(32'h388ad0cd),
	.w2(32'h3c913e94),
	.w3(32'hbb92e572),
	.w4(32'h3b9a7e6f),
	.w5(32'h3a8c4edf),
	.w6(32'hbc967cbf),
	.w7(32'h3b2fc2c4),
	.w8(32'hbab1bfb7),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ad201),
	.w1(32'hbc0fcddf),
	.w2(32'hbb3e7ed6),
	.w3(32'hbb1e9878),
	.w4(32'hbb8c7661),
	.w5(32'hbb60796d),
	.w6(32'hbc178dbc),
	.w7(32'hbbfcb588),
	.w8(32'h399b2e38),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4671de),
	.w1(32'hbadc67fb),
	.w2(32'h3c1bb8b9),
	.w3(32'hb9928eed),
	.w4(32'h3ba26563),
	.w5(32'h3c4e19f2),
	.w6(32'hbc62ffbc),
	.w7(32'h3bac2095),
	.w8(32'hba2d5399),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule