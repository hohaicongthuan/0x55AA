module layer_10_featuremap_107(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ce850),
	.w1(32'h3892dc66),
	.w2(32'h39938771),
	.w3(32'h3a141e55),
	.w4(32'hb8d3c1fb),
	.w5(32'hb937bef9),
	.w6(32'h3886df75),
	.w7(32'h39f84c1d),
	.w8(32'h3a86d72b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d871e),
	.w1(32'h39ea6f97),
	.w2(32'h3ad9e13b),
	.w3(32'h3b80f7ac),
	.w4(32'hbb35fc0c),
	.w5(32'hba4529c7),
	.w6(32'h3b22d4e7),
	.w7(32'h3ac5c237),
	.w8(32'h3b32a04c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39941427),
	.w1(32'h39a4ae32),
	.w2(32'h3951bf57),
	.w3(32'h398e61b9),
	.w4(32'h39d73ca1),
	.w5(32'h39a52f0e),
	.w6(32'hb8ab11f4),
	.w7(32'hb8944770),
	.w8(32'h3887327e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87a4b2),
	.w1(32'hbaaba334),
	.w2(32'hbaceee41),
	.w3(32'hb878858a),
	.w4(32'h3aaa3c36),
	.w5(32'h3aa1a05d),
	.w6(32'hb885cdb7),
	.w7(32'hb9ad553c),
	.w8(32'h3966884e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b0def),
	.w1(32'hb9dcaecf),
	.w2(32'h3a9e5b29),
	.w3(32'hba56e887),
	.w4(32'hba239473),
	.w5(32'h3a23822f),
	.w6(32'hba47a5c7),
	.w7(32'hb9fac056),
	.w8(32'hba0cff8b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ec036),
	.w1(32'h3acddea7),
	.w2(32'h3a37c28f),
	.w3(32'h39fbe1aa),
	.w4(32'h3ad90528),
	.w5(32'h3a901b7f),
	.w6(32'h3aa36725),
	.w7(32'h3a7e3bf2),
	.w8(32'h3a2cd224),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba522a71),
	.w1(32'h3b9018e6),
	.w2(32'h3c6ce587),
	.w3(32'hbb0790d3),
	.w4(32'h3b921b76),
	.w5(32'h3c07dac3),
	.w6(32'h3b837aa9),
	.w7(32'h3abb6ae2),
	.w8(32'h3c0943cc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1ec8c),
	.w1(32'h3c723f84),
	.w2(32'h3b8f96e8),
	.w3(32'h3c89104c),
	.w4(32'h3c86b45b),
	.w5(32'h3b60d8db),
	.w6(32'h3c236692),
	.w7(32'h3b08c653),
	.w8(32'hb92e7acf),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fcb23b),
	.w1(32'h392bd104),
	.w2(32'h3a738148),
	.w3(32'h39b0943a),
	.w4(32'h3a5e7e62),
	.w5(32'h39bd35a9),
	.w6(32'h36d2d1ca),
	.w7(32'h3a2f5a45),
	.w8(32'h3a064d8d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf66fc),
	.w1(32'hbb6b4a67),
	.w2(32'h3bd2802a),
	.w3(32'hbc0d4c7a),
	.w4(32'hbbab34d9),
	.w5(32'hb8c060ba),
	.w6(32'h3c21fe41),
	.w7(32'h3c4ecde7),
	.w8(32'h3ca1577c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49f144),
	.w1(32'h385cc28c),
	.w2(32'h3a4ef9d8),
	.w3(32'hb9f8d7ef),
	.w4(32'hba4e44c8),
	.w5(32'hb904dbd4),
	.w6(32'hba2a7582),
	.w7(32'hbad5d760),
	.w8(32'hbac1636d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30036c),
	.w1(32'hbba64857),
	.w2(32'h3c86dbf4),
	.w3(32'hbbd2fba4),
	.w4(32'hbbbd941b),
	.w5(32'h3c204a23),
	.w6(32'h3bab4855),
	.w7(32'hbbd478ce),
	.w8(32'h3c70037d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc020d74),
	.w1(32'h37db3ec0),
	.w2(32'h3bee90d7),
	.w3(32'hbbed169e),
	.w4(32'hbb010cd8),
	.w5(32'h3b9352ee),
	.w6(32'h3c280650),
	.w7(32'h3c3c68f0),
	.w8(32'h3c9377f2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb2f5e),
	.w1(32'h3baeb050),
	.w2(32'h3c01f2a6),
	.w3(32'h3a91c4cc),
	.w4(32'h3ac8edf4),
	.w5(32'h3bb1cb6b),
	.w6(32'h3b237f53),
	.w7(32'h3b5ea857),
	.w8(32'h3bc2a29a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2667af),
	.w1(32'hbaec9b16),
	.w2(32'h3a8dae28),
	.w3(32'hbb8791f5),
	.w4(32'hbbfa8dfa),
	.w5(32'hbb95c79c),
	.w6(32'h3b110e48),
	.w7(32'h3b12ff1c),
	.w8(32'h3b8e957e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a7e81),
	.w1(32'h3c294630),
	.w2(32'h3bf5a05e),
	.w3(32'hbaa32fcf),
	.w4(32'hbb2ea8b3),
	.w5(32'hbab80416),
	.w6(32'h3c45eafe),
	.w7(32'h3c4a5b94),
	.w8(32'h3c5d910a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a420ef5),
	.w1(32'hb983d08c),
	.w2(32'hb939cee9),
	.w3(32'h39c59a0e),
	.w4(32'hba39afbb),
	.w5(32'hba821377),
	.w6(32'hb9559daa),
	.w7(32'hb95e8a5e),
	.w8(32'h38f0c387),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba306465),
	.w1(32'hbb9c6d87),
	.w2(32'h3c25a63a),
	.w3(32'h3bd1a397),
	.w4(32'h3bbfe93d),
	.w5(32'h3c2c7da6),
	.w6(32'h3c8052a8),
	.w7(32'h3c0fd950),
	.w8(32'h3c95d55f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf26a0d),
	.w1(32'hbb32e05b),
	.w2(32'h3ad78aff),
	.w3(32'h3a0614c2),
	.w4(32'h3ac8b95d),
	.w5(32'h3b05d4dc),
	.w6(32'h3c075c12),
	.w7(32'h3bf17cff),
	.w8(32'h3c2fdcb6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c55391),
	.w1(32'h392aefba),
	.w2(32'h398aacc5),
	.w3(32'h379229e7),
	.w4(32'hb90e5a94),
	.w5(32'hb887161f),
	.w6(32'h39e2625e),
	.w7(32'h388a2a1d),
	.w8(32'hb868decd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3890dde2),
	.w1(32'h3974335f),
	.w2(32'hb90a1230),
	.w3(32'h395613da),
	.w4(32'h39f60129),
	.w5(32'h3920b558),
	.w6(32'h397c3360),
	.w7(32'hb9060dc3),
	.w8(32'hba574f64),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc17692),
	.w1(32'hbb6b82e9),
	.w2(32'h39facac6),
	.w3(32'hbbb4e15d),
	.w4(32'hbb6e437f),
	.w5(32'hb9b65e3b),
	.w6(32'hbb9da7e4),
	.w7(32'hbb351716),
	.w8(32'h3a6cfee5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fd652),
	.w1(32'h3b4dd6ea),
	.w2(32'h3c418bf5),
	.w3(32'hbb929e33),
	.w4(32'hbb8d54ce),
	.w5(32'h3c6da34d),
	.w6(32'h3d2b63b9),
	.w7(32'h3d04ab98),
	.w8(32'h3d33671b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc006840),
	.w1(32'hbb3eaf9b),
	.w2(32'h3bcbcc08),
	.w3(32'hbc05e5a7),
	.w4(32'hbbad1981),
	.w5(32'h3ab288a3),
	.w6(32'h3c0d4332),
	.w7(32'h3c25c45b),
	.w8(32'h3c912994),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe73bd),
	.w1(32'hbc0abfc4),
	.w2(32'h3a8bdfac),
	.w3(32'h3a8b5b48),
	.w4(32'hbbe96fd4),
	.w5(32'hbb5aeccc),
	.w6(32'h3c2506b1),
	.w7(32'h3c49956c),
	.w8(32'h3c9d8e12),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc5815),
	.w1(32'hb85db556),
	.w2(32'h38e6e131),
	.w3(32'hba624367),
	.w4(32'h395b5ab2),
	.w5(32'hb875713e),
	.w6(32'hbaea56b8),
	.w7(32'hba58e12d),
	.w8(32'hb9a96fbc),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba382f2f),
	.w1(32'h3a0d97f1),
	.w2(32'h394e1bf6),
	.w3(32'hba881182),
	.w4(32'h39b25738),
	.w5(32'hb8fc7763),
	.w6(32'h3997e613),
	.w7(32'h3908dddd),
	.w8(32'hba0347e1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd06ff39),
	.w1(32'h3932dcd6),
	.w2(32'h3c240e71),
	.w3(32'hbcc14c98),
	.w4(32'h3be6df9e),
	.w5(32'h3bd07910),
	.w6(32'hbd124ba5),
	.w7(32'h3bc65964),
	.w8(32'h3b9ec857),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a45db),
	.w1(32'hbb8f5903),
	.w2(32'h3b35812d),
	.w3(32'hbb264300),
	.w4(32'hbb9db89b),
	.w5(32'h3b37fd34),
	.w6(32'hbabc2e69),
	.w7(32'hbb76d3b5),
	.w8(32'h3a8c392d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf10fa0),
	.w1(32'hbbcd5f4c),
	.w2(32'hba8ccd1d),
	.w3(32'hbc8a500f),
	.w4(32'hb9a83a3b),
	.w5(32'h3b554371),
	.w6(32'hbcadc404),
	.w7(32'h3b128160),
	.w8(32'h3c0cff14),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf1409),
	.w1(32'h39e64579),
	.w2(32'h380bdb56),
	.w3(32'hb84c17da),
	.w4(32'h39aed5fd),
	.w5(32'h38846c41),
	.w6(32'h399fbe60),
	.w7(32'h37a910fd),
	.w8(32'hb9d0a80a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a1453a),
	.w1(32'h398da8b9),
	.w2(32'hb832844e),
	.w3(32'hb90f2a39),
	.w4(32'h38db3d50),
	.w5(32'hb91490e7),
	.w6(32'h398380e9),
	.w7(32'hb7996c9d),
	.w8(32'hb9b88dee),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0b3c8),
	.w1(32'hbad6c796),
	.w2(32'h3b2acad4),
	.w3(32'hbb9e5555),
	.w4(32'hbb2f5e37),
	.w5(32'h3a54cefd),
	.w6(32'h3b7298b2),
	.w7(32'h3b8ccfd5),
	.w8(32'h3bfd8213),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b471d),
	.w1(32'h39b90c23),
	.w2(32'h3b1a4f02),
	.w3(32'h3b3d8abe),
	.w4(32'hba6a59cb),
	.w5(32'h3a4c2438),
	.w6(32'h3b8306f6),
	.w7(32'h3b88b68b),
	.w8(32'h3b881ae4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39407ef4),
	.w1(32'hba661762),
	.w2(32'h380a83f3),
	.w3(32'hbacaf7ea),
	.w4(32'hbac6d4eb),
	.w5(32'hba3d3c14),
	.w6(32'hbac8c47e),
	.w7(32'hba93d9ad),
	.w8(32'h3a6c392d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d2243),
	.w1(32'hbad45880),
	.w2(32'h3ae59d0b),
	.w3(32'hbb2c2253),
	.w4(32'h3a84b5a9),
	.w5(32'h3b1aea1d),
	.w6(32'h3bb446e2),
	.w7(32'hb99772fa),
	.w8(32'hba0f819d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb56836),
	.w1(32'h3b80bb93),
	.w2(32'h3cd7286d),
	.w3(32'hbb792ba5),
	.w4(32'hbbeae180),
	.w5(32'hb8b08d7c),
	.w6(32'h3bf210cb),
	.w7(32'hbbeeb3a0),
	.w8(32'h3ca245ed),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd8ef92),
	.w1(32'hbc352472),
	.w2(32'h3c717a02),
	.w3(32'hbc8e0d41),
	.w4(32'hbc651b9f),
	.w5(32'h3c0d4da9),
	.w6(32'hbbe0a7bf),
	.w7(32'h3c49f8ef),
	.w8(32'h3cef949e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd232b15),
	.w1(32'hbc3729f5),
	.w2(32'h3c819b10),
	.w3(32'hbcbbff48),
	.w4(32'hbbdc14bb),
	.w5(32'h3c876979),
	.w6(32'hbc8f93b1),
	.w7(32'h3c0330b1),
	.w8(32'h3cd3b0a4),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac234ae),
	.w1(32'hb9efb4c3),
	.w2(32'hba60a98e),
	.w3(32'h3a86a9be),
	.w4(32'hbad60b1a),
	.w5(32'hbab15280),
	.w6(32'h3b019e30),
	.w7(32'h3b2cfabd),
	.w8(32'h3ae4c0d6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e671ac),
	.w1(32'h38d7f529),
	.w2(32'h37f77e61),
	.w3(32'h39ef3ae5),
	.w4(32'hb9301d0b),
	.w5(32'hb9b3b96c),
	.w6(32'hb91d2082),
	.w7(32'h37cefaa5),
	.w8(32'hb9deec27),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98155f2),
	.w1(32'hb99ecfb5),
	.w2(32'hba4b10c5),
	.w3(32'hba062986),
	.w4(32'hb9ce4ca3),
	.w5(32'hba8f4186),
	.w6(32'hba199dae),
	.w7(32'hba8a4334),
	.w8(32'hba8fcfee),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb635a51),
	.w1(32'hbb90ed9b),
	.w2(32'h3b813888),
	.w3(32'hbb999c5a),
	.w4(32'hbbcd6f50),
	.w5(32'h3b464fa9),
	.w6(32'hbb916b14),
	.w7(32'hbbc4786a),
	.w8(32'h3ac447a9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb763f),
	.w1(32'hba8b2a42),
	.w2(32'h3bc11e83),
	.w3(32'hbbe066c2),
	.w4(32'hbc1a6f18),
	.w5(32'h3b113845),
	.w6(32'h3c65bf34),
	.w7(32'h3c369525),
	.w8(32'h3cb5c26a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03fdb5),
	.w1(32'hbb873d0d),
	.w2(32'h3b78817b),
	.w3(32'hbbbe7ec3),
	.w4(32'hbbc1495e),
	.w5(32'h39d02f24),
	.w6(32'h3b4ea2eb),
	.w7(32'h3c004e8c),
	.w8(32'h3c8e4145),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52ba25),
	.w1(32'hbc14b774),
	.w2(32'hba594eee),
	.w3(32'hbbbe5347),
	.w4(32'hbbb04c46),
	.w5(32'hb9093494),
	.w6(32'h3c8eaed0),
	.w7(32'h3c74005c),
	.w8(32'h3cb793fc),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986e35e),
	.w1(32'hba482ee5),
	.w2(32'h3ba7b971),
	.w3(32'hbb5aadbe),
	.w4(32'hbbbeb4ba),
	.w5(32'h3a093a3b),
	.w6(32'h3bff48af),
	.w7(32'h3c279b1e),
	.w8(32'h3c80c941),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37fdab),
	.w1(32'hb9fcea4e),
	.w2(32'h3c3e9cc3),
	.w3(32'hbb2b8fb2),
	.w4(32'h3c1228f7),
	.w5(32'h3c3431fb),
	.w6(32'h3cbbd97d),
	.w7(32'h3cb20595),
	.w8(32'h3cd72253),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0108b5),
	.w1(32'h3955784f),
	.w2(32'h3a0438ed),
	.w3(32'h38a930a7),
	.w4(32'h399d6c8b),
	.w5(32'h39b0c29f),
	.w6(32'h38b88cc2),
	.w7(32'h39be5d4d),
	.w8(32'h38a49665),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba208b87),
	.w1(32'h39ec7590),
	.w2(32'hb6a419ed),
	.w3(32'h39f205d4),
	.w4(32'h3ad1a562),
	.w5(32'h3a44132e),
	.w6(32'h3ab7fa66),
	.w7(32'h3aa6f5e5),
	.w8(32'h3a36a233),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986ccf6),
	.w1(32'h38dd41f4),
	.w2(32'h3a119279),
	.w3(32'hb94c0126),
	.w4(32'h39b56abd),
	.w5(32'h39bd02a5),
	.w6(32'h390f66a5),
	.w7(32'h3a041223),
	.w8(32'h39d4953f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb893b45),
	.w1(32'h3b2b6812),
	.w2(32'h3b298cd6),
	.w3(32'hbb3c0583),
	.w4(32'h3b53fec4),
	.w5(32'h3b7cf3de),
	.w6(32'h3b74afbd),
	.w7(32'h3bfec02e),
	.w8(32'h3c46a959),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a247981),
	.w1(32'h3aa976d0),
	.w2(32'h39db3e27),
	.w3(32'h3981be14),
	.w4(32'h3adae938),
	.w5(32'h3b35eecb),
	.w6(32'h3b8b16bc),
	.w7(32'h3b25fa85),
	.w8(32'h3b588c14),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfcba8),
	.w1(32'hbb158729),
	.w2(32'h3ba8dba3),
	.w3(32'hbb82136e),
	.w4(32'hbae38a70),
	.w5(32'h3b47bf16),
	.w6(32'h3c590a40),
	.w7(32'h3c33cb21),
	.w8(32'h3c807878),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbd26b),
	.w1(32'hba6c757a),
	.w2(32'h3abd0d5b),
	.w3(32'hb91de78c),
	.w4(32'h3a365b1a),
	.w5(32'h3b3995a9),
	.w6(32'h3a82d6b0),
	.w7(32'h3ac77c96),
	.w8(32'h3b424c82),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c4e1d6),
	.w1(32'hb8a3c109),
	.w2(32'h3989fad5),
	.w3(32'hba14b13a),
	.w4(32'hba264089),
	.w5(32'hba1a6a21),
	.w6(32'hba371d17),
	.w7(32'hb92bc999),
	.w8(32'hb9d3c378),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a89103),
	.w1(32'h38c30e7e),
	.w2(32'hba08d1c5),
	.w3(32'hba011020),
	.w4(32'h3a3af02b),
	.w5(32'h391ab2c8),
	.w6(32'h3971626f),
	.w7(32'hb82dc6dd),
	.w8(32'hb8f0eb04),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacffcaf),
	.w1(32'hb9e892c6),
	.w2(32'h3a8a2d38),
	.w3(32'hb8dbdee2),
	.w4(32'h3a588bc9),
	.w5(32'h3aaa58fa),
	.w6(32'hb9b2a238),
	.w7(32'h3a3adfde),
	.w8(32'h3aaaeb92),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f23e7),
	.w1(32'hbb1bb35d),
	.w2(32'h39f1b3b5),
	.w3(32'hba8fb02d),
	.w4(32'hbafba64b),
	.w5(32'h3a7feeed),
	.w6(32'hba6da9a0),
	.w7(32'hbae0f1c5),
	.w8(32'h3a9a734d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b4ccf),
	.w1(32'h38a7ef75),
	.w2(32'h3a332313),
	.w3(32'hbaafeef6),
	.w4(32'h39d8eb80),
	.w5(32'h3adfc71b),
	.w6(32'hba93d02f),
	.w7(32'h388a41b3),
	.w8(32'h3aa1dea0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba420552),
	.w1(32'hbb4c9304),
	.w2(32'h3b13a389),
	.w3(32'hbb1ec0ad),
	.w4(32'hbb0281e3),
	.w5(32'h3b829ccc),
	.w6(32'h3b9eab30),
	.w7(32'h3a415e8e),
	.w8(32'h3c02c16d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba356b02),
	.w1(32'h3b62d5c4),
	.w2(32'h3bb7dfee),
	.w3(32'hbad22a33),
	.w4(32'h3aac184b),
	.w5(32'h3ba12848),
	.w6(32'hbb9d8b08),
	.w7(32'hbb65ce39),
	.w8(32'h3b2576b9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39804cd1),
	.w1(32'hba80f822),
	.w2(32'hba1543ed),
	.w3(32'h39292410),
	.w4(32'hba98eb9c),
	.w5(32'hba38daa2),
	.w6(32'hba19b7ee),
	.w7(32'hba919b92),
	.w8(32'hbad35217),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb4401),
	.w1(32'hba2c9742),
	.w2(32'hba46ee23),
	.w3(32'hba8ce67f),
	.w4(32'hb9e23d8e),
	.w5(32'hba1f8e51),
	.w6(32'hba1dea70),
	.w7(32'hb9af191b),
	.w8(32'h3894a0e6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37668253),
	.w1(32'h3901b99c),
	.w2(32'hb780ae4a),
	.w3(32'hb7210bec),
	.w4(32'hb90d154d),
	.w5(32'hb908a879),
	.w6(32'h39cda6e8),
	.w7(32'h3932d783),
	.w8(32'hb9d9cd52),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d75bab),
	.w1(32'hb9ed535b),
	.w2(32'hb9949327),
	.w3(32'h3931882d),
	.w4(32'hb915deb9),
	.w5(32'hb8104b89),
	.w6(32'hba6543dc),
	.w7(32'hb9eaabfe),
	.w8(32'hb7bd3bbb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc805ff),
	.w1(32'h3c0cc079),
	.w2(32'h3c0da6db),
	.w3(32'hbba05fcc),
	.w4(32'hbc88fe34),
	.w5(32'hbc8f9c25),
	.w6(32'h3bf5530d),
	.w7(32'h3be066dd),
	.w8(32'h3c193993),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7103c4),
	.w1(32'hbc61e4c2),
	.w2(32'hbbc5e11b),
	.w3(32'hb526aba0),
	.w4(32'h38c875fa),
	.w5(32'h3be8d8df),
	.w6(32'h3ce8c2c2),
	.w7(32'h3c6cf5e9),
	.w8(32'h3caa5b0e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5eed3),
	.w1(32'hbb9ae4e5),
	.w2(32'h3c0e7ae6),
	.w3(32'hbb0feae1),
	.w4(32'hba88dc47),
	.w5(32'h3c61bbbc),
	.w6(32'h3c91a51b),
	.w7(32'h3c35cf5b),
	.w8(32'h3cceb4ff),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc935a6),
	.w1(32'hbc8eeaf1),
	.w2(32'h3bc6db90),
	.w3(32'hbb921ac0),
	.w4(32'hbc24acc0),
	.w5(32'h3b15ebc3),
	.w6(32'h3c3a6613),
	.w7(32'h3cb21bcb),
	.w8(32'h3d057b4f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a132d9),
	.w1(32'h37abbffa),
	.w2(32'hb9d8ae37),
	.w3(32'h39e30083),
	.w4(32'h368bbd74),
	.w5(32'hb9d670b9),
	.w6(32'hb887b5ec),
	.w7(32'h38fa9001),
	.w8(32'h38e1ad8d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b11b9d),
	.w1(32'h3a0da9d8),
	.w2(32'hb959576e),
	.w3(32'h380d5235),
	.w4(32'h3a16a606),
	.w5(32'hb921254b),
	.w6(32'h3903f385),
	.w7(32'hb8bffd18),
	.w8(32'hba0df288),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f128dc),
	.w1(32'h3a33cf17),
	.w2(32'h3973b7e2),
	.w3(32'hb8cb8aae),
	.w4(32'h3a132ccf),
	.w5(32'h3933dad2),
	.w6(32'h39c04ad2),
	.w7(32'h399c1f0d),
	.w8(32'hb9aa6770),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29be85),
	.w1(32'hba80087b),
	.w2(32'h38b71ce2),
	.w3(32'hbb005ca3),
	.w4(32'hbb4e4805),
	.w5(32'hba5012eb),
	.w6(32'h3b25985e),
	.w7(32'h3a5476fb),
	.w8(32'h3a73b827),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92582df),
	.w1(32'h394cc17a),
	.w2(32'hba01afa4),
	.w3(32'hb9611b1c),
	.w4(32'h395ca890),
	.w5(32'hb96b07b1),
	.w6(32'h38f20f83),
	.w7(32'hb8ccdad9),
	.w8(32'hb97a669e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0edc17),
	.w1(32'h3b56ec18),
	.w2(32'h3a84c010),
	.w3(32'hba3a3eb1),
	.w4(32'h3a9ee81d),
	.w5(32'hba881252),
	.w6(32'h3be5b1ec),
	.w7(32'h3baf191b),
	.w8(32'h3bafa0c3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04bab5),
	.w1(32'hb9c83b0d),
	.w2(32'h39a16e5a),
	.w3(32'hbb6cc27e),
	.w4(32'h3b60022e),
	.w5(32'h3b08fae1),
	.w6(32'h3c6e462a),
	.w7(32'h3b965d9b),
	.w8(32'h3bdb732a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f59c9),
	.w1(32'h3ad6d0bd),
	.w2(32'h3ac778d6),
	.w3(32'h3ac587bb),
	.w4(32'h3b3ca923),
	.w5(32'hbacefe61),
	.w6(32'h3bd10420),
	.w7(32'h3c6ba64c),
	.w8(32'h3c4f58b0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03b258),
	.w1(32'hbb344e5c),
	.w2(32'h3b37ad56),
	.w3(32'hbb004f78),
	.w4(32'hbb8dd108),
	.w5(32'h39de13e2),
	.w6(32'h3b8db7f8),
	.w7(32'h3b019cea),
	.w8(32'h3bd1b6cf),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c075711),
	.w1(32'h3bce34b2),
	.w2(32'h3bf8b770),
	.w3(32'hbb91090f),
	.w4(32'hba2193a3),
	.w5(32'hbbb8c6bf),
	.w6(32'h3af2a31d),
	.w7(32'h3b663206),
	.w8(32'h3ba28224),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb803520),
	.w1(32'hba388ea5),
	.w2(32'h3b85152d),
	.w3(32'hbb690477),
	.w4(32'hbaf9c201),
	.w5(32'h39d9c5a9),
	.w6(32'hbb072974),
	.w7(32'h3acb6dd6),
	.w8(32'h3bcecf5e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f447ab),
	.w1(32'h3af3e379),
	.w2(32'h3b863a38),
	.w3(32'hbb213f2e),
	.w4(32'h3b626040),
	.w5(32'h3b927a3f),
	.w6(32'h3bdd41e6),
	.w7(32'h3bd7bc8c),
	.w8(32'h3c254cbb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7ef1d),
	.w1(32'hba0e3546),
	.w2(32'hb9eb5def),
	.w3(32'h39bceeac),
	.w4(32'hba2d8286),
	.w5(32'hba2fa5f3),
	.w6(32'hba03b4e3),
	.w7(32'hb9f65ad6),
	.w8(32'hba0e59e3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920c23f),
	.w1(32'h398826f5),
	.w2(32'hb7be61ce),
	.w3(32'hba0bcd1c),
	.w4(32'h38dda882),
	.w5(32'hb6b8d8e5),
	.w6(32'h38fcb6d7),
	.w7(32'h3997f90e),
	.w8(32'h3a30e563),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964478a),
	.w1(32'hb870e23f),
	.w2(32'hba1ff081),
	.w3(32'hb8762efb),
	.w4(32'hba64360d),
	.w5(32'hba749c96),
	.w6(32'hba5b2ee5),
	.w7(32'hba2729b2),
	.w8(32'hba2a1c58),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc2cb5),
	.w1(32'hba47cf4c),
	.w2(32'hb9fb06a7),
	.w3(32'hba0ab07d),
	.w4(32'h3a2f4363),
	.w5(32'h3a0c5580),
	.w6(32'hba8f9681),
	.w7(32'hb787a96e),
	.w8(32'h3a2a1a43),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb188e95),
	.w1(32'hbb2f63a2),
	.w2(32'h3b2f3c0e),
	.w3(32'h3b05dad4),
	.w4(32'hbb328d44),
	.w5(32'h3ab8f417),
	.w6(32'h3c250db1),
	.w7(32'h3c0eff7d),
	.w8(32'h3c07f364),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b0ced),
	.w1(32'hbb3c8a65),
	.w2(32'h3a223de4),
	.w3(32'hba551f4b),
	.w4(32'hbb3beaeb),
	.w5(32'h3a167c76),
	.w6(32'h38602755),
	.w7(32'hbaa0cc30),
	.w8(32'h3a5b0c6d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba27508),
	.w1(32'hbb7c26c8),
	.w2(32'hbbbd3b57),
	.w3(32'h3b50ab6f),
	.w4(32'hba193941),
	.w5(32'hb9af7c9a),
	.w6(32'h3c0d5086),
	.w7(32'h3ba46e61),
	.w8(32'h3ba15574),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a3054),
	.w1(32'h3a8c6697),
	.w2(32'h3b9248b5),
	.w3(32'h3b8939c0),
	.w4(32'h3bc4c844),
	.w5(32'h3bc0af1c),
	.w6(32'h3ccc4cd5),
	.w7(32'h3c698f0d),
	.w8(32'h3ca0d62d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c4b52),
	.w1(32'hbbad22ce),
	.w2(32'h3bc09858),
	.w3(32'hbc533bdf),
	.w4(32'hbb89671e),
	.w5(32'h3bf5c8cd),
	.w6(32'hbc3d1d70),
	.w7(32'hb8eb1c2d),
	.w8(32'h3c27cc29),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bf4e9),
	.w1(32'h3b87f9c6),
	.w2(32'h3c3e604e),
	.w3(32'hbc2f92c0),
	.w4(32'hbc862bfc),
	.w5(32'hbc41cb98),
	.w6(32'h3c1e4a67),
	.w7(32'h3b94e43b),
	.w8(32'h3c87dbf2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38df90),
	.w1(32'hbbe5edb2),
	.w2(32'h39f4f848),
	.w3(32'hbbc1b85c),
	.w4(32'hba690fdd),
	.w5(32'h3bb16622),
	.w6(32'h3b5b12b5),
	.w7(32'h3bc9ed17),
	.w8(32'h3c2f4aac),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b928a4c),
	.w1(32'h3b749d11),
	.w2(32'h3ba2f0be),
	.w3(32'hbaeacaed),
	.w4(32'hbbebc86f),
	.w5(32'hbb88b608),
	.w6(32'h3c90ff65),
	.w7(32'h3c47353f),
	.w8(32'h3c4b2ac8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b54ac),
	.w1(32'h3af9fed4),
	.w2(32'h3a9fdb7f),
	.w3(32'hbaf776fa),
	.w4(32'hbaf7c54f),
	.w5(32'hbba8cf8d),
	.w6(32'h3b9cfe60),
	.w7(32'h3ba39264),
	.w8(32'h3bcd52f3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd869ee),
	.w1(32'h3b19b2b2),
	.w2(32'h3b8b190c),
	.w3(32'hbbcaaf62),
	.w4(32'hbacf68d6),
	.w5(32'hb9c698d7),
	.w6(32'hbbb56573),
	.w7(32'h3be52e30),
	.w8(32'h3c31fd74),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb024e),
	.w1(32'hb9d7a3cc),
	.w2(32'hb99c9374),
	.w3(32'hb9ea1e42),
	.w4(32'hb9368bc3),
	.w5(32'h3917d523),
	.w6(32'hb9bf5d7b),
	.w7(32'hb86616b0),
	.w8(32'hb9841828),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4fdbb),
	.w1(32'hbbcb76b3),
	.w2(32'h3b95c668),
	.w3(32'hbba6610f),
	.w4(32'hb7fb79de),
	.w5(32'h3ba82eba),
	.w6(32'h3c26663e),
	.w7(32'h3c42e81f),
	.w8(32'h3c9ae0de),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa57b9),
	.w1(32'h3bd44f9a),
	.w2(32'h3c81d73d),
	.w3(32'hbc0198ef),
	.w4(32'h3b6b882e),
	.w5(32'h3b9ed63a),
	.w6(32'h3c35a065),
	.w7(32'h3ca1d2b8),
	.w8(32'h3cd2e05c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b965bea),
	.w1(32'hbc17fb11),
	.w2(32'h3b04ec52),
	.w3(32'h3b813e81),
	.w4(32'h3afd1e19),
	.w5(32'h3c4023f5),
	.w6(32'h3cedd3dc),
	.w7(32'h3b9a098d),
	.w8(32'h3c2c8313),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9604cf),
	.w1(32'hbbd1be17),
	.w2(32'h3c9b3451),
	.w3(32'hbc80eae8),
	.w4(32'hbc08332d),
	.w5(32'h3c0dc292),
	.w6(32'hbb6b63c8),
	.w7(32'h3c1029ed),
	.w8(32'h3c8aee22),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51b840),
	.w1(32'hbbd86301),
	.w2(32'hba17d70b),
	.w3(32'hbb352c78),
	.w4(32'hbaf8087a),
	.w5(32'hba9848cc),
	.w6(32'h3ba72b8e),
	.w7(32'h3c240a22),
	.w8(32'h3c6206d8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c593b44),
	.w1(32'h3bddb6a4),
	.w2(32'h3cb68953),
	.w3(32'hbb886fd1),
	.w4(32'hbb626e31),
	.w5(32'h3a8b2702),
	.w6(32'h3c70e8b5),
	.w7(32'h3b4414e6),
	.w8(32'h3c9cf94b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a059a78),
	.w1(32'h3a3b68ac),
	.w2(32'h3a1e025a),
	.w3(32'h3a12a49e),
	.w4(32'h3a18a3b8),
	.w5(32'h39beb4b5),
	.w6(32'h39d6aa7e),
	.w7(32'h397a30d0),
	.w8(32'h38a48d81),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c519f7f),
	.w1(32'h3bad3077),
	.w2(32'h3c6bd619),
	.w3(32'h3b1cd917),
	.w4(32'h3b5486b5),
	.w5(32'h3cac6cee),
	.w6(32'h3c4f6cf6),
	.w7(32'h3b6292f1),
	.w8(32'h3c18b5db),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4086b),
	.w1(32'hba4ab4e6),
	.w2(32'h3c4a060c),
	.w3(32'hbba7d2a0),
	.w4(32'h3bdae1c4),
	.w5(32'h3c533868),
	.w6(32'h3b71c9a9),
	.w7(32'h3c3a7fa3),
	.w8(32'h3c12d41a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f06776),
	.w1(32'h39b313a2),
	.w2(32'h39fe33fc),
	.w3(32'hba1e0c3e),
	.w4(32'h392859c7),
	.w5(32'h39b0a6bd),
	.w6(32'hba90458c),
	.w7(32'hba219120),
	.w8(32'hb93df207),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20ff59),
	.w1(32'h3a2e9f19),
	.w2(32'hbaf86f48),
	.w3(32'h3af6d283),
	.w4(32'h39055dc4),
	.w5(32'hbace9d12),
	.w6(32'h3b8c65ad),
	.w7(32'h3b3bf0e9),
	.w8(32'h3b15372b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8b64b),
	.w1(32'hbadfdfb1),
	.w2(32'h3b0c2122),
	.w3(32'hbbcd079d),
	.w4(32'hbaa53cd5),
	.w5(32'h3a072df6),
	.w6(32'h3c0b24ec),
	.w7(32'h3c3c17c7),
	.w8(32'h3c59f94b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b2c4e),
	.w1(32'hbaf5a508),
	.w2(32'h3aef3098),
	.w3(32'hbb8566ac),
	.w4(32'hba5d78b7),
	.w5(32'hb8194a75),
	.w6(32'hba6da879),
	.w7(32'h3bbe8b77),
	.w8(32'h3c22b312),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1619df),
	.w1(32'h3b280204),
	.w2(32'h3b997661),
	.w3(32'hbb60d515),
	.w4(32'h3b09e16c),
	.w5(32'h3b822aec),
	.w6(32'hbbaa761a),
	.w7(32'h3c2a7c68),
	.w8(32'h3c5d0b6a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed3fc3),
	.w1(32'hb9d6fcd7),
	.w2(32'h3ae26f30),
	.w3(32'hba5971f8),
	.w4(32'hba39ee48),
	.w5(32'h3b40a81e),
	.w6(32'h3ac04bc3),
	.w7(32'h3bd838e7),
	.w8(32'h3c16f55e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a6840),
	.w1(32'hbc587399),
	.w2(32'hbba057e6),
	.w3(32'h3a3c1eb9),
	.w4(32'h3a33f847),
	.w5(32'h3bb2a7de),
	.w6(32'h3c3c64b0),
	.w7(32'h3b9f8b50),
	.w8(32'h3bd0ce97),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c624fae),
	.w1(32'h3c34de2f),
	.w2(32'h3c12d993),
	.w3(32'h3b03a3a4),
	.w4(32'hbabc491e),
	.w5(32'hbb108692),
	.w6(32'h3be134dd),
	.w7(32'h3b4c17af),
	.w8(32'h3b92ceee),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94132d),
	.w1(32'hbb160e89),
	.w2(32'h3aacd7c8),
	.w3(32'hbaf09eb0),
	.w4(32'hba759901),
	.w5(32'h3a487c8b),
	.w6(32'h3b61f9f9),
	.w7(32'h3bcb6711),
	.w8(32'h3c0652b4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e26fce),
	.w1(32'h3a242859),
	.w2(32'h3a096bb2),
	.w3(32'hba23c9a4),
	.w4(32'h3a397f85),
	.w5(32'h3a1d4cde),
	.w6(32'h3a29e31d),
	.w7(32'h39dd91ea),
	.w8(32'h38e1441b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0db6ae),
	.w1(32'h3acce83f),
	.w2(32'h39ad2c5d),
	.w3(32'h3a7d66c3),
	.w4(32'hb90955f4),
	.w5(32'hb8bdb7fe),
	.w6(32'h3a71145b),
	.w7(32'h39d762bc),
	.w8(32'hb96b562e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d60d5),
	.w1(32'h3a204a2f),
	.w2(32'h39a50dbb),
	.w3(32'h39f88d57),
	.w4(32'h3a8b1c7b),
	.w5(32'h3a194540),
	.w6(32'h3a3fbc5b),
	.w7(32'h396a91b6),
	.w8(32'h3902e5df),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f6851),
	.w1(32'hb99b0fbd),
	.w2(32'hb9f81968),
	.w3(32'h387203cf),
	.w4(32'h3894db7b),
	.w5(32'h37d79f13),
	.w6(32'h391a670e),
	.w7(32'hb9ad41c2),
	.w8(32'hb9834069),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeff2f6),
	.w1(32'hbb8f2fab),
	.w2(32'h3aa64222),
	.w3(32'hbb7d1d2d),
	.w4(32'hbb4a12fd),
	.w5(32'h39d4f8ed),
	.w6(32'h3b420555),
	.w7(32'h3bc2073b),
	.w8(32'h3c269104),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8cf22),
	.w1(32'hb8eca14d),
	.w2(32'h3a6b3b82),
	.w3(32'hba0cd69b),
	.w4(32'hba562c4a),
	.w5(32'h3a2f74cf),
	.w6(32'hba0331d2),
	.w7(32'hba6d8933),
	.w8(32'h3932bb66),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52c5ea),
	.w1(32'h3b7b9155),
	.w2(32'h3bc14b91),
	.w3(32'hba70e3ec),
	.w4(32'h3b3b11cf),
	.w5(32'h3af3dc7a),
	.w6(32'h3bc1f9fe),
	.w7(32'h3bd8896d),
	.w8(32'h3beb8ac7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12844a),
	.w1(32'h3a5d2848),
	.w2(32'h3bec745a),
	.w3(32'hbbe2c46c),
	.w4(32'h3b28a83e),
	.w5(32'h3bd9ac07),
	.w6(32'hbba7eee9),
	.w7(32'h3c2b96d0),
	.w8(32'h3c7c0022),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a81e4e),
	.w1(32'h3a35213b),
	.w2(32'hb97a86cb),
	.w3(32'h391b2fd1),
	.w4(32'hb6d0c476),
	.w5(32'hb9fb70cf),
	.w6(32'hb76e75dd),
	.w7(32'h39506d69),
	.w8(32'h3a5eb349),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c38d0b),
	.w1(32'h3a867d5b),
	.w2(32'h39ca8340),
	.w3(32'hb9385f78),
	.w4(32'h3a97c356),
	.w5(32'h3a2eafe3),
	.w6(32'h3aa28193),
	.w7(32'h3a3fc8b0),
	.w8(32'h3a29bdd5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d18be7),
	.w1(32'h39fba644),
	.w2(32'h3913b8af),
	.w3(32'h3a080b37),
	.w4(32'h39c22aa1),
	.w5(32'h3901052f),
	.w6(32'h39d7dbfc),
	.w7(32'hb9032850),
	.w8(32'hba122f22),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d04de),
	.w1(32'h3a242a99),
	.w2(32'h38a959d5),
	.w3(32'h3abfcf2d),
	.w4(32'h3a838a72),
	.w5(32'h39c1877e),
	.w6(32'h3b63c494),
	.w7(32'h3b6e29b7),
	.w8(32'h3ac9cf87),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a0d3a),
	.w1(32'hbbabe895),
	.w2(32'hbbb74ccc),
	.w3(32'h3ae588c0),
	.w4(32'h3c246744),
	.w5(32'h3b92a680),
	.w6(32'h3c92af40),
	.w7(32'h3beb8b27),
	.w8(32'h3c147cd2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3700d),
	.w1(32'hbbcc6086),
	.w2(32'hb980cc29),
	.w3(32'hbbc74fd1),
	.w4(32'hbb86920a),
	.w5(32'hbaf53ff2),
	.w6(32'h3b798828),
	.w7(32'h3b863681),
	.w8(32'h3be9d9e2),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7ec8c),
	.w1(32'h3a182b1e),
	.w2(32'h3a8ee0f3),
	.w3(32'hbacdd357),
	.w4(32'hbaa842a3),
	.w5(32'h3850cc10),
	.w6(32'h394575d9),
	.w7(32'h39cdd2b7),
	.w8(32'h3aed0180),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58a745),
	.w1(32'hba3efbcd),
	.w2(32'h3a88458d),
	.w3(32'hb97e4a2c),
	.w4(32'hb9e0d67e),
	.w5(32'h3b30849f),
	.w6(32'h3b8e61b1),
	.w7(32'h3998121e),
	.w8(32'h3b1c5f8f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89128c),
	.w1(32'h3aa43129),
	.w2(32'h3a9ff7e1),
	.w3(32'hb9883411),
	.w4(32'h39c100ef),
	.w5(32'h3a80e853),
	.w6(32'h3a846dd9),
	.w7(32'h3b24220f),
	.w8(32'h3b4c7320),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba358f36),
	.w1(32'hbb007d41),
	.w2(32'h3a5e33cd),
	.w3(32'hbb42192a),
	.w4(32'hbb95d6d5),
	.w5(32'hbaafd3e5),
	.w6(32'h3af79d10),
	.w7(32'h3a262ee7),
	.w8(32'h3b0f5bfb),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20c378),
	.w1(32'h3bbf6019),
	.w2(32'h3b5bebc2),
	.w3(32'h3bc0a333),
	.w4(32'hbb0820a3),
	.w5(32'hbb9d0ac5),
	.w6(32'h3b2eaea3),
	.w7(32'h3aad4ff9),
	.w8(32'h3b48e0b3),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95cf57),
	.w1(32'h3b09a0ea),
	.w2(32'h3c62a4f1),
	.w3(32'hbb704f46),
	.w4(32'h3a260e9d),
	.w5(32'h3bbd4769),
	.w6(32'h3c378c6f),
	.w7(32'h3c710445),
	.w8(32'h3c9e863b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb625fb3),
	.w1(32'hbaa31d5c),
	.w2(32'h3b25de78),
	.w3(32'hbb2aa4e6),
	.w4(32'hbb4bc428),
	.w5(32'hba32727c),
	.w6(32'hbaf70594),
	.w7(32'h3b971201),
	.w8(32'h3bd62c34),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2b173),
	.w1(32'h3b597539),
	.w2(32'h3b23302b),
	.w3(32'hbb964e29),
	.w4(32'hbb2348fa),
	.w5(32'hb9fa96cb),
	.w6(32'h3c42385b),
	.w7(32'h3c13429c),
	.w8(32'h3c1b86be),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c4a96),
	.w1(32'h3bb59e48),
	.w2(32'h3bb3a5e5),
	.w3(32'h39e9dfb4),
	.w4(32'h3b28ccb7),
	.w5(32'h3b984102),
	.w6(32'h3c368ab7),
	.w7(32'h3be505f8),
	.w8(32'h3c59bc74),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7bccd),
	.w1(32'hbbf13fe1),
	.w2(32'hbb810e41),
	.w3(32'h3b19fb43),
	.w4(32'hbb10167d),
	.w5(32'hbaa14918),
	.w6(32'h3c12c5f1),
	.w7(32'h3bb6c805),
	.w8(32'h3bc1b100),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3aee0f),
	.w1(32'h3a8e1c0a),
	.w2(32'h3b93e282),
	.w3(32'hbb8cf903),
	.w4(32'hbb2380bc),
	.w5(32'h3915e1db),
	.w6(32'h3b9c2758),
	.w7(32'h3bc79152),
	.w8(32'h3c0d465f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec6683),
	.w1(32'hba69422e),
	.w2(32'h3a1e835c),
	.w3(32'hbab1e02e),
	.w4(32'hb9befa01),
	.w5(32'h3a112995),
	.w6(32'h3aa97f71),
	.w7(32'h3affbb2b),
	.w8(32'h3b5a76e9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd435ae),
	.w1(32'hb9c6030c),
	.w2(32'h3b374c47),
	.w3(32'hbc762a15),
	.w4(32'h3bb1f334),
	.w5(32'h3c4416de),
	.w6(32'hbc829f10),
	.w7(32'h3c76c1f0),
	.w8(32'h3c8f1126),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b422144),
	.w1(32'h3aa8ddb6),
	.w2(32'h39201830),
	.w3(32'h3b6a3f0c),
	.w4(32'h3ab77359),
	.w5(32'h394e90f7),
	.w6(32'h3c0871df),
	.w7(32'h3babcc2c),
	.w8(32'h3ba15795),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33ab4cdc),
	.w1(32'h39339c25),
	.w2(32'h392dfbf7),
	.w3(32'hb8e949a5),
	.w4(32'h38827d7b),
	.w5(32'hb9141784),
	.w6(32'h391c0bad),
	.w7(32'h37f8e59c),
	.w8(32'hb8c3fb28),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940d2d0),
	.w1(32'h38880f47),
	.w2(32'hb7b5ab63),
	.w3(32'hb88adad6),
	.w4(32'h38ea071a),
	.w5(32'hb83d2003),
	.w6(32'hb8590ff3),
	.w7(32'h3717ec61),
	.w8(32'h389800e6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdaed7),
	.w1(32'hbae933a9),
	.w2(32'h3b17a4a4),
	.w3(32'hbafb55e6),
	.w4(32'hbae1175e),
	.w5(32'h3a1b5a5c),
	.w6(32'h3b002afc),
	.w7(32'h3b3f1eb8),
	.w8(32'h3b8160fe),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a1237),
	.w1(32'h3aa683b3),
	.w2(32'h3b08f488),
	.w3(32'h3b7a9e3d),
	.w4(32'hb9b9103b),
	.w5(32'h3a8cd316),
	.w6(32'h3c070d6d),
	.w7(32'h3c4bd67e),
	.w8(32'h3c41b40d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc076990),
	.w1(32'hbbe88827),
	.w2(32'hbb09a7de),
	.w3(32'hba84ee20),
	.w4(32'h39b2c35f),
	.w5(32'hb8d37d5a),
	.w6(32'h3c4bc19a),
	.w7(32'h3c4f4939),
	.w8(32'h3c808100),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382296e1),
	.w1(32'h3884fb22),
	.w2(32'hb83387ad),
	.w3(32'hb6ba70f0),
	.w4(32'h36ae9f7c),
	.w5(32'hb8bc87bd),
	.w6(32'hb817200c),
	.w7(32'hb7e2c779),
	.w8(32'hb8e3f36a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26da94),
	.w1(32'hb9e82147),
	.w2(32'h3b857f84),
	.w3(32'hbbd0e161),
	.w4(32'hbb67c769),
	.w5(32'h36fd2940),
	.w6(32'h3ba41b00),
	.w7(32'h3c1dc840),
	.w8(32'h3c6158c3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cc354),
	.w1(32'hba48df13),
	.w2(32'hba816de3),
	.w3(32'hb9b36211),
	.w4(32'h3a9cb73d),
	.w5(32'hbabc3084),
	.w6(32'h3befb25f),
	.w7(32'h3c153176),
	.w8(32'h3bcd00b2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53f19e),
	.w1(32'h3c1dd51b),
	.w2(32'h3c4c7567),
	.w3(32'h3b1e5c6c),
	.w4(32'hb9a51e05),
	.w5(32'hbb58f537),
	.w6(32'h3c43e31f),
	.w7(32'h3c39f859),
	.w8(32'h3c831ef4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca656d2),
	.w1(32'hb92efd86),
	.w2(32'h3aa67306),
	.w3(32'hbc743637),
	.w4(32'hbb098b69),
	.w5(32'h39888332),
	.w6(32'hbc7b70e9),
	.w7(32'h3c39d51e),
	.w8(32'h3cafe19d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b6741),
	.w1(32'h3a373e44),
	.w2(32'h3a40ee3c),
	.w3(32'h3b803476),
	.w4(32'h3ac55da7),
	.w5(32'h3b134cad),
	.w6(32'h3b2b26e1),
	.w7(32'h3b172b7b),
	.w8(32'h3b1e06c9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba430076),
	.w1(32'hba7f17bb),
	.w2(32'hba29f634),
	.w3(32'hba6d6539),
	.w4(32'hb9fd8b7f),
	.w5(32'hba0ccbf4),
	.w6(32'hba255fd0),
	.w7(32'hba631659),
	.w8(32'hba407e35),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d7cd7),
	.w1(32'hbba62b96),
	.w2(32'h39bfaef3),
	.w3(32'hbc06909b),
	.w4(32'hbb967e8d),
	.w5(32'h39e64a2c),
	.w6(32'hbb97a771),
	.w7(32'h3a3c6d67),
	.w8(32'h3bee7d64),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f0205),
	.w1(32'hbb17b771),
	.w2(32'h3b467036),
	.w3(32'h37e6dee2),
	.w4(32'hbb63fc7f),
	.w5(32'h3a00dbf5),
	.w6(32'h3bdd3a34),
	.w7(32'h3ba3bbfc),
	.w8(32'h3c073e6f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ad202),
	.w1(32'hbb88c906),
	.w2(32'h3b1a1f57),
	.w3(32'hbaefbb7e),
	.w4(32'hbb8ab556),
	.w5(32'h3b11e60b),
	.w6(32'hbb1f8494),
	.w7(32'hb96676fd),
	.w8(32'h3ba6b586),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dea64),
	.w1(32'h3a47b59b),
	.w2(32'h3ad802c1),
	.w3(32'hbb08427d),
	.w4(32'hbaef9aca),
	.w5(32'hba95249a),
	.w6(32'h3b72a1fb),
	.w7(32'h3b40463f),
	.w8(32'h3b7041ec),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f59f9c),
	.w1(32'h392081af),
	.w2(32'h38d12ce8),
	.w3(32'h39c400a4),
	.w4(32'h390ef68f),
	.w5(32'hb92061a7),
	.w6(32'h39c590a9),
	.w7(32'h3a4324a4),
	.w8(32'h3a0da3c0),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc0794),
	.w1(32'hb815c906),
	.w2(32'h3a2e71c3),
	.w3(32'hbb433c25),
	.w4(32'hba18c828),
	.w5(32'h39a06da7),
	.w6(32'h3c269fec),
	.w7(32'h3bcafe92),
	.w8(32'h3c11ae06),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f37d3e),
	.w1(32'h39e191fd),
	.w2(32'h3b7fae0e),
	.w3(32'hba5b6d3e),
	.w4(32'h39f8c534),
	.w5(32'h3998f55e),
	.w6(32'h39b7a8d5),
	.w7(32'h3ae31bba),
	.w8(32'h3b313ed2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39aa60),
	.w1(32'hbb4ca1c5),
	.w2(32'hbac57cef),
	.w3(32'hbb6e615a),
	.w4(32'h3a7aa367),
	.w5(32'h3b115457),
	.w6(32'hbb8d5062),
	.w7(32'h3acf3125),
	.w8(32'h3ba541b9),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06745e),
	.w1(32'hba22ffb6),
	.w2(32'h38a4c6a4),
	.w3(32'hb940a33d),
	.w4(32'hba31809c),
	.w5(32'hb96606dd),
	.w6(32'hb9846770),
	.w7(32'hba130d0a),
	.w8(32'hb9cd2f2f),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05aa53),
	.w1(32'hbbe62b08),
	.w2(32'h3bd5a005),
	.w3(32'hbaa12dde),
	.w4(32'h3a146f99),
	.w5(32'h3c51f991),
	.w6(32'h3ade606f),
	.w7(32'hbb01aa79),
	.w8(32'h3c44ad2e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913e2f2),
	.w1(32'h377f98d3),
	.w2(32'hb70d340b),
	.w3(32'h3826e733),
	.w4(32'hb804feb3),
	.w5(32'hb8272a59),
	.w6(32'hb87a8e5b),
	.w7(32'hb893a5d7),
	.w8(32'hb8eb0274),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39809a4a),
	.w1(32'h385ec310),
	.w2(32'h39c86ddb),
	.w3(32'h388f933e),
	.w4(32'h374b2293),
	.w5(32'h39ad2d9a),
	.w6(32'h384d2ec5),
	.w7(32'hb7da9e43),
	.w8(32'h39a943d6),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba38e96),
	.w1(32'hbae2fae5),
	.w2(32'h3a0e1ae5),
	.w3(32'hbba0e513),
	.w4(32'hbb63854c),
	.w5(32'hbb316202),
	.w6(32'hbb572d15),
	.w7(32'h3b020a1d),
	.w8(32'h3b8db2a8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc066dee),
	.w1(32'hbbca9f53),
	.w2(32'hb92f5b22),
	.w3(32'hbbdf60fe),
	.w4(32'h391295fc),
	.w5(32'h3c0569f3),
	.w6(32'h3caf12f4),
	.w7(32'h3c24044c),
	.w8(32'h3c912eba),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ddd64),
	.w1(32'hbb878ee5),
	.w2(32'h3b098654),
	.w3(32'hbaaab513),
	.w4(32'hbb391bd7),
	.w5(32'h3b7d574b),
	.w6(32'hba2dc5ea),
	.w7(32'hbacca63a),
	.w8(32'h3b472aa0),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6ea15),
	.w1(32'hb9eb0777),
	.w2(32'h3af6f1be),
	.w3(32'hbb27f145),
	.w4(32'hb99bd562),
	.w5(32'h3a381d5a),
	.w6(32'hbaaf422f),
	.w7(32'h3bcd8129),
	.w8(32'h3c09cd80),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d7fb8),
	.w1(32'hbac9eaa1),
	.w2(32'hba6a9755),
	.w3(32'hbb6769c5),
	.w4(32'h396dd44d),
	.w5(32'hb9ae79d2),
	.w6(32'hbb93f7e9),
	.w7(32'h3916e812),
	.w8(32'h3a51ccb6),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1da7ca),
	.w1(32'hbb98a080),
	.w2(32'h3c0b1fef),
	.w3(32'hbbc37ef8),
	.w4(32'hbbb8c6e1),
	.w5(32'h3ba439cd),
	.w6(32'h3c3eefd1),
	.w7(32'h3c2f3b55),
	.w8(32'h3c9f26ec),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d85cc),
	.w1(32'h3ace361e),
	.w2(32'h3c1687ce),
	.w3(32'hbb0e02f3),
	.w4(32'hbb53eb61),
	.w5(32'h3af56bf9),
	.w6(32'h3c130583),
	.w7(32'h3c08573e),
	.w8(32'h3c6d307b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8c71e),
	.w1(32'hb9dede28),
	.w2(32'h3b8d6f20),
	.w3(32'hbaa63e44),
	.w4(32'h39b7696c),
	.w5(32'h3b4173d2),
	.w6(32'h3c1c65cb),
	.w7(32'h3bf427de),
	.w8(32'h3c479019),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96085c6),
	.w1(32'hb9400a58),
	.w2(32'hb8f55ce8),
	.w3(32'hb94d1e9e),
	.w4(32'hb90a5050),
	.w5(32'hb9243fb1),
	.w6(32'hb9a81c09),
	.w7(32'hb96a3304),
	.w8(32'hb97eb8f5),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1c089),
	.w1(32'h3b9a7a9d),
	.w2(32'h390657cd),
	.w3(32'hb8e06aa0),
	.w4(32'h3a0cab9a),
	.w5(32'hbb6f7e7c),
	.w6(32'h3b217804),
	.w7(32'h3b834ebb),
	.w8(32'h3b547de9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3865a054),
	.w1(32'h387712f8),
	.w2(32'hb92a7877),
	.w3(32'h38a9c5d6),
	.w4(32'h37d63e14),
	.w5(32'hb937c3d3),
	.w6(32'hb8d5d213),
	.w7(32'hb90fc847),
	.w8(32'hb9a679d4),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba906c7d),
	.w1(32'hbabf38f5),
	.w2(32'hb9a88261),
	.w3(32'hba5cf789),
	.w4(32'hba988cee),
	.w5(32'hb92e0bbc),
	.w6(32'h3ae29496),
	.w7(32'h3b0ca9c1),
	.w8(32'h3b88e03a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92861c0),
	.w1(32'hba549683),
	.w2(32'hba59df52),
	.w3(32'h3a9a75d2),
	.w4(32'hb991397e),
	.w5(32'h3886fdd9),
	.w6(32'hba6c59f5),
	.w7(32'hb9386b4c),
	.w8(32'h38b91487),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaf2e4),
	.w1(32'h3b9bc02f),
	.w2(32'h3bebf11e),
	.w3(32'h3acead44),
	.w4(32'hb88e5e08),
	.w5(32'h3aa056e0),
	.w6(32'h3c1fb8b3),
	.w7(32'h3c11a4c7),
	.w8(32'h3c2d7965),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68ec755),
	.w1(32'hb670f91b),
	.w2(32'hb8d17e34),
	.w3(32'h378cf08c),
	.w4(32'hb6c2a5b9),
	.w5(32'hb8bcfaf2),
	.w6(32'hb8368ae7),
	.w7(32'hb8621436),
	.w8(32'hb902294b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7476411),
	.w1(32'hb73badb8),
	.w2(32'hb897144e),
	.w3(32'hb8695043),
	.w4(32'hb5f591c0),
	.w5(32'hb7d50467),
	.w6(32'hb90ab39a),
	.w7(32'hb9271fd9),
	.w8(32'hb9135bf0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb986ccc),
	.w1(32'hb8d9ac15),
	.w2(32'h3abd6b5d),
	.w3(32'hb9dc9590),
	.w4(32'h3a647c0f),
	.w5(32'h3a1f9103),
	.w6(32'hba966e93),
	.w7(32'h3b3d5765),
	.w8(32'h3b8a2680),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a5081),
	.w1(32'hbad4b8a4),
	.w2(32'h3bfefd7c),
	.w3(32'hbb3bb6c0),
	.w4(32'hbb027148),
	.w5(32'h3b9c4d10),
	.w6(32'h3b932fa9),
	.w7(32'h3c0d8a94),
	.w8(32'h3c716680),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf437b3),
	.w1(32'h3b8b53bc),
	.w2(32'h3c0b022f),
	.w3(32'hba9d0994),
	.w4(32'h3b6507de),
	.w5(32'h3ae89398),
	.w6(32'h3b1d80e7),
	.w7(32'hbb282867),
	.w8(32'h3b42c9ad),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b2cda),
	.w1(32'hb9c24472),
	.w2(32'hb955f0dc),
	.w3(32'hb82a4ae3),
	.w4(32'hb9ec92d8),
	.w5(32'h396f6c70),
	.w6(32'h3ad20d94),
	.w7(32'h39668899),
	.w8(32'h3ab9a458),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a1da2),
	.w1(32'hbc4ea997),
	.w2(32'hbae0a788),
	.w3(32'hbc87cd36),
	.w4(32'hbc573bb4),
	.w5(32'hbab965ce),
	.w6(32'h3c1400ec),
	.w7(32'hbb98f39a),
	.w8(32'h3c0b1294),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c3875),
	.w1(32'h3b9375af),
	.w2(32'h3b781138),
	.w3(32'hbc6f34b8),
	.w4(32'hbc319a3d),
	.w5(32'hbc26fdf1),
	.w6(32'hbc423ec2),
	.w7(32'hb931befa),
	.w8(32'h3bdd3072),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02636a),
	.w1(32'h3b000055),
	.w2(32'h3b5d7151),
	.w3(32'hbb11e7fe),
	.w4(32'h3a98e576),
	.w5(32'h3b2b29f5),
	.w6(32'h3a0d12be),
	.w7(32'h3acae865),
	.w8(32'h3b46fbd5),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bb2ebc),
	.w1(32'h383165b9),
	.w2(32'h3758cc30),
	.w3(32'h38bdb0f0),
	.w4(32'h395b8ec2),
	.w5(32'h36d8fcc4),
	.w6(32'hb6fce55d),
	.w7(32'h389316dc),
	.w8(32'hb8428c19),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37486a17),
	.w1(32'h389bf679),
	.w2(32'h3884cce7),
	.w3(32'hb838b981),
	.w4(32'hb7d9486c),
	.w5(32'hb763ec0c),
	.w6(32'hb8b6b051),
	.w7(32'hb91b5a7f),
	.w8(32'hb89e70c0),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb661765d),
	.w1(32'h373ead70),
	.w2(32'hb8cff982),
	.w3(32'hb7423e01),
	.w4(32'h3590bb21),
	.w5(32'hb8e383b0),
	.w6(32'hb8ed1ec2),
	.w7(32'hb8d73495),
	.w8(32'hb95b112a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01d8e0),
	.w1(32'hba915a2d),
	.w2(32'h3bc43109),
	.w3(32'hbb3fc207),
	.w4(32'h3a83387b),
	.w5(32'h3b6ce8c7),
	.w6(32'h3b2e056b),
	.w7(32'h3a56bdde),
	.w8(32'h3b82fc52),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a812d44),
	.w1(32'h3ad9eec7),
	.w2(32'h3b70b18b),
	.w3(32'hbaf3d539),
	.w4(32'h39a78d56),
	.w5(32'h3ba0bbd8),
	.w6(32'h3c44c262),
	.w7(32'h3c1882e4),
	.w8(32'h3c38bf92),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e310f),
	.w1(32'hbb75a211),
	.w2(32'hba73548e),
	.w3(32'h3b366c7b),
	.w4(32'hbbf4ce2a),
	.w5(32'hbb96ece5),
	.w6(32'h3b9b7bb2),
	.w7(32'h3b8d5e37),
	.w8(32'h3c003ddc),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fde7b),
	.w1(32'hbae5ad2f),
	.w2(32'hb94b1d1f),
	.w3(32'h395a9915),
	.w4(32'h3a823c3b),
	.w5(32'h3af0e5ea),
	.w6(32'h3a8aa1e8),
	.w7(32'h3a846654),
	.w8(32'h3b25885b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ff7c),
	.w1(32'hbb450452),
	.w2(32'h3be112e5),
	.w3(32'hbbcc0224),
	.w4(32'hbb93162d),
	.w5(32'h3b8e85c2),
	.w6(32'h3c59bbcb),
	.w7(32'h3c42bdd7),
	.w8(32'h3c9e9564),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb897471c),
	.w1(32'h378a365c),
	.w2(32'h3b75141b),
	.w3(32'hba978326),
	.w4(32'h3b471aa9),
	.w5(32'h3b95bb16),
	.w6(32'h3b659e07),
	.w7(32'h3bd4339c),
	.w8(32'h3b91de25),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36247ad5),
	.w1(32'h35709709),
	.w2(32'hb94a1e79),
	.w3(32'hb65dff7d),
	.w4(32'hb76dbbae),
	.w5(32'hb94a8a2b),
	.w6(32'hb926a06d),
	.w7(32'hb9225eb2),
	.w8(32'hb9a9a774),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eb68e),
	.w1(32'h3b8801e1),
	.w2(32'h3ac174b0),
	.w3(32'hba0925bc),
	.w4(32'hba7fd316),
	.w5(32'h3b545b0d),
	.w6(32'h3a3e1836),
	.w7(32'hbb21274e),
	.w8(32'hbb31224c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e735f2),
	.w1(32'h38462e15),
	.w2(32'hb9ed01a9),
	.w3(32'h38145cfa),
	.w4(32'hb814d64b),
	.w5(32'hba019e58),
	.w6(32'hb9c2b489),
	.w7(32'hb9d0f339),
	.w8(32'hba59843c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b391e),
	.w1(32'hbb2c5ffd),
	.w2(32'h3b9b8406),
	.w3(32'hbc1efa94),
	.w4(32'hba853f0f),
	.w5(32'h3bc20f30),
	.w6(32'h3b8fe914),
	.w7(32'h3c0b97fe),
	.w8(32'h3c666fa6),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab52145),
	.w1(32'hbb62362f),
	.w2(32'h3b477a66),
	.w3(32'h3b95c406),
	.w4(32'hbbd58782),
	.w5(32'h3a896c8a),
	.w6(32'h3c1de707),
	.w7(32'h3bd44ef8),
	.w8(32'h3c4c4705),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fa73d),
	.w1(32'hbb79ee86),
	.w2(32'h3b349daa),
	.w3(32'hbb641b27),
	.w4(32'hbb83c733),
	.w5(32'h3a65c113),
	.w6(32'h3b7bef65),
	.w7(32'h3be422ed),
	.w8(32'h3c42b208),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14a483),
	.w1(32'hbacea871),
	.w2(32'h3b1a6cb0),
	.w3(32'hbb0296dc),
	.w4(32'hbabd97b1),
	.w5(32'h3b1e0ec5),
	.w6(32'hbab2d71b),
	.w7(32'hb9dfc7eb),
	.w8(32'h3b2b8857),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8aa4f),
	.w1(32'h3a2eeab5),
	.w2(32'h3ac4de1e),
	.w3(32'hbbcafd93),
	.w4(32'hbb7ddea9),
	.w5(32'hbb479a07),
	.w6(32'hbb2fdc71),
	.w7(32'h3c0944a8),
	.w8(32'h3c4312c0),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba684cc9),
	.w1(32'hbb0942be),
	.w2(32'h3aed73a5),
	.w3(32'hbb1fc768),
	.w4(32'hbb56e4a1),
	.w5(32'hbae610b7),
	.w6(32'h3bb0b664),
	.w7(32'h3b88aaf8),
	.w8(32'h3b950de7),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7bc1b),
	.w1(32'hbb79aeb3),
	.w2(32'hb972719d),
	.w3(32'hba95ceea),
	.w4(32'h3b0034af),
	.w5(32'h3b6e069f),
	.w6(32'h3c902924),
	.w7(32'h3c88b1d7),
	.w8(32'h3c9f2f4e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cd1c49),
	.w1(32'hb84308b4),
	.w2(32'hb92c4ace),
	.w3(32'hb8bddc93),
	.w4(32'hb81329e1),
	.w5(32'hb938ea50),
	.w6(32'hb908e365),
	.w7(32'hb8c27751),
	.w8(32'hb94b0d35),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9361fd5),
	.w1(32'hb8c7387c),
	.w2(32'h3828ab7c),
	.w3(32'hb8b8832d),
	.w4(32'h3934a7b1),
	.w5(32'h3a1ebb0d),
	.w6(32'hb8cce170),
	.w7(32'hb8e48a4d),
	.w8(32'h38e3fa84),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a933d),
	.w1(32'hbc1890e6),
	.w2(32'h3a4a61ca),
	.w3(32'hbb953073),
	.w4(32'hbbb0db89),
	.w5(32'h3b3d7fc7),
	.w6(32'h3cae6063),
	.w7(32'h3c58012c),
	.w8(32'h3c84d4cf),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30cfe5),
	.w1(32'hbb55e78b),
	.w2(32'h3b7fda6a),
	.w3(32'hbbe94f93),
	.w4(32'hb9d693e0),
	.w5(32'h3c09dba6),
	.w6(32'h3c9b06d6),
	.w7(32'h3c7d08d0),
	.w8(32'h3c9b746d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad03ac),
	.w1(32'hbba97370),
	.w2(32'hbab0bb04),
	.w3(32'hbaa7f16c),
	.w4(32'hbbadce9c),
	.w5(32'hbb59b6be),
	.w6(32'h3c12429b),
	.w7(32'h3bec2c94),
	.w8(32'h3c3b7069),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c034e23),
	.w1(32'h3a7dce30),
	.w2(32'h3bbe778e),
	.w3(32'hbc0086cd),
	.w4(32'hbb5de1f0),
	.w5(32'hbc199532),
	.w6(32'hbb4875e6),
	.w7(32'h3b2862e7),
	.w8(32'h3c1a657d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d0716c),
	.w1(32'h3a450ad8),
	.w2(32'h39e5d486),
	.w3(32'h3a03c0b9),
	.w4(32'h39779b6b),
	.w5(32'h39cd5d9c),
	.w6(32'h3b0bf5e9),
	.w7(32'h3a2f481a),
	.w8(32'hb82359ad),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3975f775),
	.w1(32'h3a2f586e),
	.w2(32'hb962bc68),
	.w3(32'h39797b8d),
	.w4(32'hb90f3844),
	.w5(32'hba93b5b5),
	.w6(32'h3afecced),
	.w7(32'h3989ae61),
	.w8(32'hba241a6c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a42fd),
	.w1(32'hbb983122),
	.w2(32'h3c2fde40),
	.w3(32'hbaf89df9),
	.w4(32'hbb4c80b0),
	.w5(32'h3c37eb1e),
	.w6(32'h3c6785db),
	.w7(32'hbbd1e654),
	.w8(32'h3bc99495),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97140b),
	.w1(32'hbbee339e),
	.w2(32'h3ba4ae36),
	.w3(32'hba85b001),
	.w4(32'h3918ab34),
	.w5(32'h3b6ed8a4),
	.w6(32'h3c7a4087),
	.w7(32'h3ba6c825),
	.w8(32'h3c37c8af),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2044e9),
	.w1(32'h3ba0202f),
	.w2(32'h3ba582c8),
	.w3(32'hbb36e3a4),
	.w4(32'hbb077de6),
	.w5(32'h3b4d3820),
	.w6(32'h3c85ed05),
	.w7(32'h3c194f4a),
	.w8(32'h3c4f2ae1),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc533a67),
	.w1(32'hbbbbc6df),
	.w2(32'h3a84f6e3),
	.w3(32'hbb314f14),
	.w4(32'hba989cab),
	.w5(32'h3b46bf1c),
	.w6(32'h3aa36865),
	.w7(32'h3bd0e2a0),
	.w8(32'h3c1fdce8),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e6cf5),
	.w1(32'h3709a430),
	.w2(32'h3bf8ae86),
	.w3(32'hbb10bc19),
	.w4(32'hbb6fd06e),
	.w5(32'h3a8b1cac),
	.w6(32'hb954be10),
	.w7(32'h3bcb94eb),
	.w8(32'h3c704f05),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f15399),
	.w1(32'hb80a87ca),
	.w2(32'hb8b10f17),
	.w3(32'hb7db1218),
	.w4(32'hb81c6496),
	.w5(32'hb8b95b14),
	.w6(32'hb8b2a345),
	.w7(32'hb8b3120c),
	.w8(32'hb90bdce1),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86c384a),
	.w1(32'hb7ff6d8d),
	.w2(32'hb8cc9d47),
	.w3(32'hb87c06cd),
	.w4(32'hb80b55cc),
	.w5(32'hb8cc913c),
	.w6(32'hb91395b1),
	.w7(32'hb91825d5),
	.w8(32'hb9586c1c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56eec5),
	.w1(32'hbb2eccf9),
	.w2(32'hba86e1e0),
	.w3(32'hbab35a68),
	.w4(32'h39afe21a),
	.w5(32'h3aaab661),
	.w6(32'hbab514c6),
	.w7(32'hba337d26),
	.w8(32'hb763733e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7555bcd),
	.w1(32'h379025ba),
	.w2(32'hb8d7ff49),
	.w3(32'hb7e7da65),
	.w4(32'h36e456bc),
	.w5(32'hb9005785),
	.w6(32'hb91b78a5),
	.w7(32'hb8e64ad0),
	.w8(32'hb9818e97),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaac33),
	.w1(32'hb8ef3814),
	.w2(32'h3ba377ef),
	.w3(32'hbb01b533),
	.w4(32'h3a1b3cbf),
	.w5(32'h3b1efabc),
	.w6(32'h3a85ae8b),
	.w7(32'h3b0380cb),
	.w8(32'h3b0c16d9),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff46bc),
	.w1(32'h3ad3cfea),
	.w2(32'h3af6977f),
	.w3(32'hba5315ad),
	.w4(32'h3b1a120d),
	.w5(32'h3bcb1421),
	.w6(32'h3c4fc6e4),
	.w7(32'h3c1d2ddb),
	.w8(32'h3c2d2e19),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a44ad),
	.w1(32'hbadc025b),
	.w2(32'h3a7be9ff),
	.w3(32'hba2f848b),
	.w4(32'hba67426c),
	.w5(32'h3abfcbaa),
	.w6(32'h3bae4a1a),
	.w7(32'h3bec31be),
	.w8(32'h3c043397),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8329b2a),
	.w1(32'hb87a21d3),
	.w2(32'hb905751e),
	.w3(32'hb73b4a58),
	.w4(32'hb8b617c9),
	.w5(32'hb932b9dd),
	.w6(32'hb8d8641e),
	.w7(32'hb91fadcc),
	.w8(32'hb962f6cc),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1027c7),
	.w1(32'h3a461b84),
	.w2(32'h3c34f636),
	.w3(32'h39d27f29),
	.w4(32'h3ac610ee),
	.w5(32'h3b8edd26),
	.w6(32'h3c9ece29),
	.w7(32'h3c0c6a8c),
	.w8(32'h3c81a643),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae45f06),
	.w1(32'h38d71e6c),
	.w2(32'h3ab586b0),
	.w3(32'hba908390),
	.w4(32'h3a82260d),
	.w5(32'h3a509b12),
	.w6(32'h3bb903f4),
	.w7(32'h3b22feca),
	.w8(32'h3b869c85),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896b948),
	.w1(32'h39e404e4),
	.w2(32'h389f3cf9),
	.w3(32'h39be948b),
	.w4(32'h3a6cc1d3),
	.w5(32'h39993dc5),
	.w6(32'hb86576b0),
	.w7(32'h39c89d7e),
	.w8(32'h3985f6af),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a6338),
	.w1(32'hba8d00eb),
	.w2(32'h3b45470b),
	.w3(32'hbb5d1d6f),
	.w4(32'hbada087e),
	.w5(32'h3a682c49),
	.w6(32'h3bc93e32),
	.w7(32'h3b8d0a8f),
	.w8(32'h3bbe8653),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90450ea),
	.w1(32'hb8c75f1d),
	.w2(32'hb92ee67b),
	.w3(32'hb835bb59),
	.w4(32'hb81bfcd0),
	.w5(32'hb959f1d4),
	.w6(32'hb8d38062),
	.w7(32'hb8b4a23f),
	.w8(32'hb961b497),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e26759),
	.w1(32'h37ce94c4),
	.w2(32'hb997d347),
	.w3(32'h3898c0cb),
	.w4(32'h3940e908),
	.w5(32'hb92703d5),
	.w6(32'h3ab697d1),
	.w7(32'h3a878164),
	.w8(32'h3a289b61),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb899882a),
	.w1(32'hb8750754),
	.w2(32'hb9225122),
	.w3(32'hb89f9280),
	.w4(32'hb8a6d135),
	.w5(32'hb90485a2),
	.w6(32'hb8fc8762),
	.w7(32'hb8dcc4ac),
	.w8(32'hb940e4b3),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cb5729),
	.w1(32'hb8b33c33),
	.w2(32'hb8c69bb2),
	.w3(32'hb838ea7c),
	.w4(32'hb887fb5b),
	.w5(32'hb89901aa),
	.w6(32'hb8962373),
	.w7(32'hb8e04ed4),
	.w8(32'hb91f8b22),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89dd91),
	.w1(32'hbb12cfa3),
	.w2(32'h3aab138b),
	.w3(32'h3a7a05b5),
	.w4(32'h3a9b5dbd),
	.w5(32'h3b389ba9),
	.w6(32'h3ae15189),
	.w7(32'h3b5337f9),
	.w8(32'h3bab8fa0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad113b),
	.w1(32'h3bb51a08),
	.w2(32'h3c108158),
	.w3(32'hbb9e1f07),
	.w4(32'hbbce6b24),
	.w5(32'hbba45235),
	.w6(32'h3bcae8e1),
	.w7(32'h3c0c9ff8),
	.w8(32'h3c82a860),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb046622),
	.w1(32'hbaaf8ef9),
	.w2(32'h3b99f824),
	.w3(32'hbbb83137),
	.w4(32'hbb50eeb0),
	.w5(32'h3a65a1fd),
	.w6(32'h3b5b1960),
	.w7(32'h3b219630),
	.w8(32'h3bbe30af),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3e98c),
	.w1(32'h3af83ce0),
	.w2(32'h3bbc3417),
	.w3(32'hbb9ad747),
	.w4(32'hbb342d2d),
	.w5(32'hbb1c8bc3),
	.w6(32'h3bf8e4fe),
	.w7(32'h3c17caa3),
	.w8(32'h3c20ca33),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe8642),
	.w1(32'hb9b08b78),
	.w2(32'h3929ad4e),
	.w3(32'hb9e70fcf),
	.w4(32'hba015c22),
	.w5(32'hb815fed0),
	.w6(32'hb948567b),
	.w7(32'hb9b4992d),
	.w8(32'hb8cf45b4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384e1c23),
	.w1(32'hb8b9d8be),
	.w2(32'hba611c4d),
	.w3(32'hb886c60c),
	.w4(32'h39711fe3),
	.w5(32'hb9ac709d),
	.w6(32'h395d0e58),
	.w7(32'hb9be20d0),
	.w8(32'hb9f183bf),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382de513),
	.w1(32'h38190000),
	.w2(32'hb8494160),
	.w3(32'h383648d3),
	.w4(32'h37eff55d),
	.w5(32'hb882b15e),
	.w6(32'hb6c8103a),
	.w7(32'hb7a69d73),
	.w8(32'hb8c7870a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886c764),
	.w1(32'hb824a661),
	.w2(32'hb8c681da),
	.w3(32'hb8b53e27),
	.w4(32'hb704f595),
	.w5(32'hb84a9e28),
	.w6(32'hb8bf80b9),
	.w7(32'hb85043db),
	.w8(32'hb8ddf906),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd21f79),
	.w1(32'h3ad8a5a0),
	.w2(32'hb7ab0538),
	.w3(32'hba81e4d3),
	.w4(32'hbb83e4ff),
	.w5(32'hbacb8a10),
	.w6(32'h3bf697ef),
	.w7(32'h3ba3ad35),
	.w8(32'h3bf4a983),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e397d2),
	.w1(32'h39646224),
	.w2(32'h38b5f808),
	.w3(32'h38f1980e),
	.w4(32'h397b9c1c),
	.w5(32'h38de6443),
	.w6(32'h38988244),
	.w7(32'h39084815),
	.w8(32'hb7ae145b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae94ba4),
	.w1(32'hbb7f95e7),
	.w2(32'h3ac15fcb),
	.w3(32'hbacc7d9a),
	.w4(32'hbb546204),
	.w5(32'h3adc7125),
	.w6(32'hbacd23da),
	.w7(32'hbb3de0dd),
	.w8(32'h3af60b2a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba895f53),
	.w1(32'h3ac54156),
	.w2(32'h3aba1a37),
	.w3(32'hb99d9f67),
	.w4(32'hba2e321c),
	.w5(32'h3b0ae2d0),
	.w6(32'hbab281c4),
	.w7(32'h3918a21e),
	.w8(32'h3a8138e5),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c1ffea),
	.w1(32'h384b1069),
	.w2(32'hb7885fc8),
	.w3(32'h38608c26),
	.w4(32'h38ac5b88),
	.w5(32'hb7456232),
	.w6(32'hb7c57247),
	.w7(32'h388421cb),
	.w8(32'hb791c384),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3664923a),
	.w1(32'h3a242c9b),
	.w2(32'h39a19deb),
	.w3(32'hba77614a),
	.w4(32'hb9c4cdee),
	.w5(32'hba5ade9d),
	.w6(32'h3ba6506d),
	.w7(32'h3b8c123f),
	.w8(32'h3b48c81a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a145f75),
	.w1(32'h3a4f96f8),
	.w2(32'h3a316f7a),
	.w3(32'h3888b3fb),
	.w4(32'hb908f9dc),
	.w5(32'h39424387),
	.w6(32'h39e682d8),
	.w7(32'h3a050747),
	.w8(32'h39760dc0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6211b6),
	.w1(32'h3c2b3685),
	.w2(32'h3c0df6ab),
	.w3(32'hbb47583b),
	.w4(32'hbc3f48cf),
	.w5(32'hbc14ce70),
	.w6(32'h3bdc7282),
	.w7(32'h3a9e7788),
	.w8(32'h3bf5f8c3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888dcdd),
	.w1(32'hbb1be966),
	.w2(32'hbb823710),
	.w3(32'hb8f0fd20),
	.w4(32'hbacfa0a9),
	.w5(32'hbb3b69b6),
	.w6(32'hbae1ecf6),
	.w7(32'hbb32a91b),
	.w8(32'hbaeeff14),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5af1cd),
	.w1(32'hbc286639),
	.w2(32'hbb0e3995),
	.w3(32'hbaa3d960),
	.w4(32'hbb230392),
	.w5(32'h3b591419),
	.w6(32'h3c836b66),
	.w7(32'h3c28a7c0),
	.w8(32'h3c3a140a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule