module layer_10_featuremap_475(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4d001),
	.w1(32'hba3a3c98),
	.w2(32'hb911ed8b),
	.w3(32'h380ad21f),
	.w4(32'hba69f241),
	.w5(32'hb91aaa5c),
	.w6(32'hb9d4feda),
	.w7(32'hba6ba776),
	.w8(32'hb93a04c6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb3d0b),
	.w1(32'hba272570),
	.w2(32'h3983c7de),
	.w3(32'h3a28c70e),
	.w4(32'hb9b44829),
	.w5(32'h3a099dfa),
	.w6(32'h39e90543),
	.w7(32'hb9deaf71),
	.w8(32'h39ba4e99),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f115b),
	.w1(32'h381e6e07),
	.w2(32'h38f46819),
	.w3(32'hbae8fdda),
	.w4(32'hb974a15d),
	.w5(32'hb984c12f),
	.w6(32'hba826824),
	.w7(32'h396d24d9),
	.w8(32'h386de3de),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396523c7),
	.w1(32'hba4357eb),
	.w2(32'h39a7e3fa),
	.w3(32'h375fc0bc),
	.w4(32'hb9856c75),
	.w5(32'h3a41104e),
	.w6(32'h3a1224ee),
	.w7(32'hbacc7f91),
	.w8(32'hba74cb43),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3948ecea),
	.w1(32'hba803cf9),
	.w2(32'hba12de5a),
	.w3(32'hba7d42af),
	.w4(32'hb9fa1717),
	.w5(32'hb9fbb03c),
	.w6(32'h37a43d7b),
	.w7(32'hba2a098c),
	.w8(32'hb9456364),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c20f4),
	.w1(32'hb97f6c98),
	.w2(32'h3a27c783),
	.w3(32'hb99d10dd),
	.w4(32'h3a2f0738),
	.w5(32'h3a84befb),
	.w6(32'hb7cdb976),
	.w7(32'h39811c11),
	.w8(32'h39da4637),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ef451),
	.w1(32'hba5d3d18),
	.w2(32'hba9a6d73),
	.w3(32'hb9c66082),
	.w4(32'hb99b8b97),
	.w5(32'hb9e40fd8),
	.w6(32'hba496dfc),
	.w7(32'h398f987a),
	.w8(32'hba1a4e6f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f35ece),
	.w1(32'hba41640f),
	.w2(32'hba8b612a),
	.w3(32'h39a1a0b7),
	.w4(32'hb99d4550),
	.w5(32'hba12b28f),
	.w6(32'hbaa069ce),
	.w7(32'h3a19f39b),
	.w8(32'hb99d8a52),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0db041),
	.w1(32'hba42e6eb),
	.w2(32'hb8d47fa2),
	.w3(32'hbab77922),
	.w4(32'h395eb96a),
	.w5(32'h3a9aab1c),
	.w6(32'hba2c729b),
	.w7(32'h3a28c3ae),
	.w8(32'h396a525e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8dc64),
	.w1(32'hba930433),
	.w2(32'hba42ffb2),
	.w3(32'hb997eb7e),
	.w4(32'hba2504a4),
	.w5(32'hb993cd1c),
	.w6(32'hb9c3c264),
	.w7(32'hb7bd1e5d),
	.w8(32'h39a9214d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccf7a3),
	.w1(32'hb975a8a6),
	.w2(32'hb98079d5),
	.w3(32'h39dfe89e),
	.w4(32'hb91d91b1),
	.w5(32'hba3773b8),
	.w6(32'h3aa5fc98),
	.w7(32'hb8406136),
	.w8(32'hba134d40),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7c1e2),
	.w1(32'h3a2cd6fd),
	.w2(32'h3997a065),
	.w3(32'hba498d0d),
	.w4(32'h3a28961a),
	.w5(32'h3906a283),
	.w6(32'hb9ada43b),
	.w7(32'h3a8d0417),
	.w8(32'h3a363e00),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9416f72),
	.w1(32'h3a07db36),
	.w2(32'hb7f71a44),
	.w3(32'hb9be1ecb),
	.w4(32'h39d9f9d1),
	.w5(32'h3a1dd5b2),
	.w6(32'hba20ae8f),
	.w7(32'hba0e840e),
	.w8(32'hb9795bfa),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d6cee),
	.w1(32'h3aa4303a),
	.w2(32'h3a9b3647),
	.w3(32'hba991fff),
	.w4(32'h3aa329ce),
	.w5(32'h383ef73a),
	.w6(32'hb9829858),
	.w7(32'hb873fb70),
	.w8(32'hb978fc3d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bb7bc),
	.w1(32'h3996551a),
	.w2(32'hb891dd1a),
	.w3(32'hba596ed0),
	.w4(32'h3966d31f),
	.w5(32'h3a081584),
	.w6(32'hba525d4b),
	.w7(32'h3a58cc8a),
	.w8(32'h3aa5d1cf),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39754d88),
	.w1(32'h3a804fc6),
	.w2(32'h3a388940),
	.w3(32'hba085e3a),
	.w4(32'h3a8f43f5),
	.w5(32'h3a0fa449),
	.w6(32'h39efd981),
	.w7(32'h3a8ea09e),
	.w8(32'h3aa97ad3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d37f9),
	.w1(32'hba908500),
	.w2(32'hbabc5f2c),
	.w3(32'h3a34824a),
	.w4(32'hb95387da),
	.w5(32'hba427c30),
	.w6(32'h39c79ae9),
	.w7(32'hba2b65a1),
	.w8(32'hb9f3c2d4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ceff09),
	.w1(32'hba61b111),
	.w2(32'h390d2cdb),
	.w3(32'hba4c6135),
	.w4(32'hb9ebfcfb),
	.w5(32'hba014942),
	.w6(32'hbaa2c9e3),
	.w7(32'hb9cb588d),
	.w8(32'hba57f4d3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87f5667),
	.w1(32'hba57a925),
	.w2(32'hba97a0f2),
	.w3(32'hb94ed411),
	.w4(32'hba3057ba),
	.w5(32'hb9e174b7),
	.w6(32'h38575749),
	.w7(32'hb9845ec4),
	.w8(32'hba4c6d71),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9793adf),
	.w1(32'h3879324d),
	.w2(32'h3941845f),
	.w3(32'hbac22f84),
	.w4(32'h38500fb7),
	.w5(32'h3a87a69e),
	.w6(32'hbaae4178),
	.w7(32'hb6e28581),
	.w8(32'hb991ba05),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7faeb14),
	.w1(32'h38991106),
	.w2(32'h3a29d988),
	.w3(32'hb9113a43),
	.w4(32'h3a85121b),
	.w5(32'h3b0281e7),
	.w6(32'h391a9382),
	.w7(32'h3aa2efa3),
	.w8(32'h3ae71753),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd4e31),
	.w1(32'h3a7f256f),
	.w2(32'hb96ff782),
	.w3(32'h3ac24d84),
	.w4(32'h3a5d384d),
	.w5(32'hb9b9b328),
	.w6(32'h3ac3ecc7),
	.w7(32'h3a34b903),
	.w8(32'hb9c5d364),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b160d50),
	.w1(32'hba325b3a),
	.w2(32'hb8a566b8),
	.w3(32'h3ab42cf9),
	.w4(32'hbab152ec),
	.w5(32'hb99f7d3c),
	.w6(32'h3aa35e53),
	.w7(32'hba9b0ed3),
	.w8(32'hba8c3209),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba334068),
	.w1(32'hba4ba39d),
	.w2(32'hb8c9b71c),
	.w3(32'hba700e4d),
	.w4(32'hbae3bb16),
	.w5(32'hba87046e),
	.w6(32'hba9be95b),
	.w7(32'hba90d790),
	.w8(32'hb91e5099),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db0fc8),
	.w1(32'hba879943),
	.w2(32'hb9cbdcd0),
	.w3(32'hbaac27c1),
	.w4(32'hba96425b),
	.w5(32'hbad354ab),
	.w6(32'hba8d03d2),
	.w7(32'hb9d825a7),
	.w8(32'hbaa94fcc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9894d37),
	.w1(32'hbb046034),
	.w2(32'hbaa8d575),
	.w3(32'h39c22be3),
	.w4(32'hbaf71f3f),
	.w5(32'hbac9c656),
	.w6(32'h38f2969c),
	.w7(32'hbb212f3e),
	.w8(32'hbb0b797a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d2925),
	.w1(32'h39cfd5ab),
	.w2(32'h38e163d5),
	.w3(32'hba5beb8c),
	.w4(32'h3a53493f),
	.w5(32'h3a5d526d),
	.w6(32'hbab5f3de),
	.w7(32'hb9468590),
	.w8(32'hba0fd3a6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb899fc31),
	.w1(32'hb99e3a29),
	.w2(32'h39600765),
	.w3(32'hb94144fe),
	.w4(32'hb9bb0a65),
	.w5(32'h3a119145),
	.w6(32'hbabd0caa),
	.w7(32'h3870f3e3),
	.w8(32'hb9eff965),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6513b8),
	.w1(32'hba7bd172),
	.w2(32'hba3adbfd),
	.w3(32'h39ccb18a),
	.w4(32'hba4c2030),
	.w5(32'hba270d52),
	.w6(32'h3aa35748),
	.w7(32'hb8c1a08f),
	.w8(32'hb9f84b46),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0ec23),
	.w1(32'h3a6dbd24),
	.w2(32'h3ab24575),
	.w3(32'hba8059a0),
	.w4(32'h3a6a0f94),
	.w5(32'h3a87c9c5),
	.w6(32'hbaeb66a1),
	.w7(32'h3a8505d2),
	.w8(32'h3ab26d3a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae77894),
	.w1(32'hbafa88cc),
	.w2(32'hbaeb61fb),
	.w3(32'h3af7ef73),
	.w4(32'hbafb20fd),
	.w5(32'hba441205),
	.w6(32'h3ab80ba5),
	.w7(32'hba8583cc),
	.w8(32'hba883d28),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac426b1),
	.w1(32'h3a061f9d),
	.w2(32'h39d544f5),
	.w3(32'h38311f22),
	.w4(32'h3a69ffb1),
	.w5(32'h3aa98148),
	.w6(32'hba8fd19c),
	.w7(32'h3a5cb1f6),
	.w8(32'h3a45d2fe),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3798b88b),
	.w1(32'hb917fb3e),
	.w2(32'hba8cd8ea),
	.w3(32'hb99e0443),
	.w4(32'h399a7d64),
	.w5(32'h39982605),
	.w6(32'h399221c5),
	.w7(32'h3a09a9b4),
	.w8(32'hba118623),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabda209),
	.w1(32'hba3295fe),
	.w2(32'hb988f89f),
	.w3(32'hba10f8c8),
	.w4(32'hba84359b),
	.w5(32'h3933bedd),
	.w6(32'hba053576),
	.w7(32'hba19af57),
	.w8(32'hba804f6f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72f2e1a),
	.w1(32'h39b1a618),
	.w2(32'h3a918e97),
	.w3(32'hb904f8c9),
	.w4(32'hb9318794),
	.w5(32'h3a331888),
	.w6(32'hba45f011),
	.w7(32'hb71203c0),
	.w8(32'h3a38ef94),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e38ce),
	.w1(32'hba7361d4),
	.w2(32'hba1510b9),
	.w3(32'h3a275df8),
	.w4(32'hba644ab8),
	.w5(32'hb8e47423),
	.w6(32'hb9ac8b2a),
	.w7(32'hba9b4718),
	.w8(32'hba3dfcb1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24c06e),
	.w1(32'hb75dc845),
	.w2(32'h3a6dc96b),
	.w3(32'hba239075),
	.w4(32'h39de4993),
	.w5(32'h3a942670),
	.w6(32'hba3e50b2),
	.w7(32'h3a40a6ad),
	.w8(32'h3a2be3d6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99187b),
	.w1(32'h392e1c6e),
	.w2(32'hba321368),
	.w3(32'h3a387af1),
	.w4(32'h3a82db7d),
	.w5(32'h39946d2b),
	.w6(32'h3a51e46e),
	.w7(32'h3a57eeb3),
	.w8(32'h3a19a83f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bbed8),
	.w1(32'h3883524d),
	.w2(32'hba4514a2),
	.w3(32'hbae1313e),
	.w4(32'hb8e40f05),
	.w5(32'hb9633bda),
	.w6(32'hba2d3046),
	.w7(32'h39c3c8ae),
	.w8(32'h39cefc2a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98749de),
	.w1(32'hba8c8317),
	.w2(32'hba1bda39),
	.w3(32'hb9d6ad21),
	.w4(32'hba66f8bc),
	.w5(32'h391a22e0),
	.w6(32'h3aa3da96),
	.w7(32'hb9afbf82),
	.w8(32'hba397492),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d18b7),
	.w1(32'h39878817),
	.w2(32'h398b1938),
	.w3(32'hba812559),
	.w4(32'hb9d70cec),
	.w5(32'hbadb3720),
	.w6(32'hb96ff529),
	.w7(32'hba28ce0c),
	.w8(32'hba95d4d8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09e6e7),
	.w1(32'h39c7582b),
	.w2(32'h3994284b),
	.w3(32'hbb499252),
	.w4(32'hba3fd17c),
	.w5(32'h3a0849e7),
	.w6(32'hbb36fb48),
	.w7(32'hb9151e55),
	.w8(32'h39b58d18),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba056560),
	.w1(32'hba323d20),
	.w2(32'h39c776c7),
	.w3(32'hba8852ff),
	.w4(32'hb94744fb),
	.w5(32'h3a5ef03c),
	.w6(32'hb92d8609),
	.w7(32'hba84a2f0),
	.w8(32'h39710c7c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2889d3),
	.w1(32'h3908f3bd),
	.w2(32'h3888cde3),
	.w3(32'hb9106ac1),
	.w4(32'h397a83a3),
	.w5(32'hb7813712),
	.w6(32'h39447e10),
	.w7(32'h392c3e1d),
	.w8(32'hb90c34b2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f4ff6),
	.w1(32'hbaa585ed),
	.w2(32'hba0159d5),
	.w3(32'h3980403f),
	.w4(32'hba7d46d3),
	.w5(32'h3a076989),
	.w6(32'h3a96a42d),
	.w7(32'hba2dfb62),
	.w8(32'hba4d3212),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c8e90),
	.w1(32'h3965d206),
	.w2(32'h39f8acfb),
	.w3(32'hba128de1),
	.w4(32'h39c1318b),
	.w5(32'h39a49ba9),
	.w6(32'hba16d224),
	.w7(32'h3a3f6d14),
	.w8(32'h3abe6b73),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eebd94),
	.w1(32'hb8f37b51),
	.w2(32'hb9f1ecea),
	.w3(32'h396d1538),
	.w4(32'h38340833),
	.w5(32'hba38612c),
	.w6(32'h39d62c77),
	.w7(32'hb955b979),
	.w8(32'hb9ed628f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba575b74),
	.w1(32'hb9b66f27),
	.w2(32'hba0e77f7),
	.w3(32'h394c6c12),
	.w4(32'hba0ef19c),
	.w5(32'hb9a7538f),
	.w6(32'hba3d71de),
	.w7(32'hb905696e),
	.w8(32'hb962b83f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b7148),
	.w1(32'hbaf984d0),
	.w2(32'hbaaab857),
	.w3(32'hb997bbc3),
	.w4(32'hbaf25fe1),
	.w5(32'hba64bc7f),
	.w6(32'h3978e2cc),
	.w7(32'hbac68050),
	.w8(32'hba8a1b40),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a6b46),
	.w1(32'hba0d5711),
	.w2(32'hba920dc0),
	.w3(32'h3699bd75),
	.w4(32'hba88a73b),
	.w5(32'hba0014c2),
	.w6(32'hba67c1f5),
	.w7(32'hba1a38af),
	.w8(32'hba70a104),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54a766),
	.w1(32'hbaa3c6ab),
	.w2(32'hba40f853),
	.w3(32'h3a932366),
	.w4(32'hba6303a6),
	.w5(32'hb97166d3),
	.w6(32'h382efaf5),
	.w7(32'hba403573),
	.w8(32'hba08a6b9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae242fb),
	.w1(32'h3a9f69f7),
	.w2(32'h39fc8fd6),
	.w3(32'hba69a08a),
	.w4(32'h3ad8cf0c),
	.w5(32'h3a055757),
	.w6(32'hba971d53),
	.w7(32'h3aea425c),
	.w8(32'h39cd437c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f3aab),
	.w1(32'h3a294143),
	.w2(32'hb80a60d7),
	.w3(32'hb9c3c53f),
	.w4(32'h399a48af),
	.w5(32'hb7252b4c),
	.w6(32'hb8e87f6a),
	.w7(32'h39cc915a),
	.w8(32'hb8c0f738),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45fc16),
	.w1(32'h39d0b858),
	.w2(32'h388f004c),
	.w3(32'hb98f2887),
	.w4(32'h3a98dac6),
	.w5(32'h3a388784),
	.w6(32'hba820928),
	.w7(32'h3aef691f),
	.w8(32'h3a7d2cb0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4e23e),
	.w1(32'hba27c96a),
	.w2(32'hb924cb23),
	.w3(32'hb9223876),
	.w4(32'hba513ab5),
	.w5(32'h3a8b973a),
	.w6(32'h376e9d45),
	.w7(32'hb8aa8d69),
	.w8(32'h3a1f0ce7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b128b41),
	.w1(32'hba330196),
	.w2(32'hb7bfb422),
	.w3(32'h3aedaf26),
	.w4(32'hb9bb3623),
	.w5(32'h3a729cc6),
	.w6(32'h3ac0df1b),
	.w7(32'hbab27149),
	.w8(32'h39f50d08),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f78a1),
	.w1(32'hba115a33),
	.w2(32'hba54eb9a),
	.w3(32'hba7e241d),
	.w4(32'hba22c919),
	.w5(32'hbabb4129),
	.w6(32'hba7340eb),
	.w7(32'hba4c3440),
	.w8(32'hbac65290),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982787e),
	.w1(32'hb9c21482),
	.w2(32'hb881f554),
	.w3(32'hb939a93c),
	.w4(32'hba619791),
	.w5(32'hb95be592),
	.w6(32'hba7b062e),
	.w7(32'hbaa29f03),
	.w8(32'hba8bf18f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94cf42e),
	.w1(32'h3a727c00),
	.w2(32'hba87ec5c),
	.w3(32'hb99a08fc),
	.w4(32'h3a616dd6),
	.w5(32'hbae015c2),
	.w6(32'hb9ed54b1),
	.w7(32'h3a5bee31),
	.w8(32'hba566682),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e81f2a),
	.w1(32'hb9e4c71b),
	.w2(32'hba6657e8),
	.w3(32'hb9ede857),
	.w4(32'h3a00b2e5),
	.w5(32'hba20d494),
	.w6(32'hb9f09fd4),
	.w7(32'hb9e8064a),
	.w8(32'hba6c9c40),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2befd3),
	.w1(32'hba9bb4b3),
	.w2(32'hba0f9cce),
	.w3(32'hb9e84824),
	.w4(32'hba9aef0d),
	.w5(32'hb9cd378f),
	.w6(32'hb9dcb802),
	.w7(32'hbb00f8a4),
	.w8(32'hbb0a355c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ab8f6),
	.w1(32'hb9f2db14),
	.w2(32'hb9d24a26),
	.w3(32'h3a3e0600),
	.w4(32'hb9478a9a),
	.w5(32'h3a58da2d),
	.w6(32'hbad6daee),
	.w7(32'hb9a0de6f),
	.w8(32'h39fd8727),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a57e5f),
	.w1(32'hbaf501d2),
	.w2(32'hb64a3702),
	.w3(32'hba87089d),
	.w4(32'hba8dba63),
	.w5(32'h39a4b32d),
	.w6(32'h39b6df55),
	.w7(32'hba65cbe5),
	.w8(32'h39e0d072),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ee651),
	.w1(32'hb9cdafe2),
	.w2(32'hba6b3c2f),
	.w3(32'hba23c9e6),
	.w4(32'hba31ffe2),
	.w5(32'hba8f3824),
	.w6(32'hb7282ee9),
	.w7(32'hb9d5f90b),
	.w8(32'hba02169e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba393b9b),
	.w1(32'h391a862e),
	.w2(32'hb8b276bb),
	.w3(32'hba607b63),
	.w4(32'h39ce2104),
	.w5(32'hb971dc46),
	.w6(32'hb9a33864),
	.w7(32'h39c0cfc4),
	.w8(32'hb8c8a373),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ddd1a),
	.w1(32'hb8544c7f),
	.w2(32'h3aa54cb1),
	.w3(32'h39835f98),
	.w4(32'h39e9497e),
	.w5(32'h3ae8358d),
	.w6(32'h388bd33c),
	.w7(32'h38bbcdc3),
	.w8(32'h3af6fe32),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0c59b),
	.w1(32'hb959a14d),
	.w2(32'h3a88662e),
	.w3(32'h3a9978f1),
	.w4(32'h3a14818c),
	.w5(32'h3ab5ecfc),
	.w6(32'h3a8e1076),
	.w7(32'h39d3036a),
	.w8(32'h3a5cc9e1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c2c03),
	.w1(32'h398a5cd1),
	.w2(32'h3ab08488),
	.w3(32'h3a17c310),
	.w4(32'h3a02d4ee),
	.w5(32'h3b0bc34b),
	.w6(32'h3a49ffc2),
	.w7(32'h3a9acebe),
	.w8(32'h3ae6628c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ceb1ac),
	.w1(32'hb97c7c5f),
	.w2(32'h37f29335),
	.w3(32'h38e1cfd8),
	.w4(32'hb8fccf54),
	.w5(32'h3aa316c6),
	.w6(32'h39b49a67),
	.w7(32'h3a3a17f8),
	.w8(32'h3abe60de),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c09b25),
	.w1(32'h3bef9124),
	.w2(32'hbae865e4),
	.w3(32'hb98381c8),
	.w4(32'h3bbe273b),
	.w5(32'hbaaa254b),
	.w6(32'h3a33a288),
	.w7(32'h3bd01f06),
	.w8(32'h38071671),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba130233),
	.w1(32'h3b31a37c),
	.w2(32'hbb61b7d0),
	.w3(32'hbb8f84b5),
	.w4(32'hb9c5871c),
	.w5(32'hbbbe960f),
	.w6(32'hbc081e21),
	.w7(32'hbb1e4512),
	.w8(32'hbb621f34),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ead83),
	.w1(32'hba8498f3),
	.w2(32'h3acea7d1),
	.w3(32'hba28d896),
	.w4(32'h3a164cee),
	.w5(32'hbba9837f),
	.w6(32'hba5840b9),
	.w7(32'h3a0a7869),
	.w8(32'hb7bf3e30),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2161e9),
	.w1(32'hbb07b75f),
	.w2(32'hba6f9157),
	.w3(32'hbb109312),
	.w4(32'h3b486829),
	.w5(32'hbbac9be0),
	.w6(32'hbb04130d),
	.w7(32'h3bc13d8f),
	.w8(32'hbb7a69f5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab771e3),
	.w1(32'hbb7a035d),
	.w2(32'h3a344554),
	.w3(32'hba5f6145),
	.w4(32'h3b055660),
	.w5(32'hbb50e787),
	.w6(32'h3b075528),
	.w7(32'h393e700b),
	.w8(32'hba39e5eb),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17eb26),
	.w1(32'hbc06820d),
	.w2(32'hbbe0b386),
	.w3(32'hb9eb704e),
	.w4(32'hbb9541b8),
	.w5(32'hbb0ba2e5),
	.w6(32'h3926a201),
	.w7(32'h3a4f7acb),
	.w8(32'hbab5e48b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba79559),
	.w1(32'hba9f5bd2),
	.w2(32'h3a6d1762),
	.w3(32'hbb7fa745),
	.w4(32'hbb006fd3),
	.w5(32'hbb9b4000),
	.w6(32'hbb46deee),
	.w7(32'h3721bd3c),
	.w8(32'h3b423165),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b645ce5),
	.w1(32'h3b581752),
	.w2(32'h3b498068),
	.w3(32'hba2eb402),
	.w4(32'h3b84c31e),
	.w5(32'h3c5c2304),
	.w6(32'h3b125643),
	.w7(32'h3aa5fe9f),
	.w8(32'hba8ee2c9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc072d55),
	.w1(32'hbac445b2),
	.w2(32'hbaa86944),
	.w3(32'hbb6e67c1),
	.w4(32'h39a73f8c),
	.w5(32'hba3c251f),
	.w6(32'hbbe572da),
	.w7(32'hbbb56f5c),
	.w8(32'hbb179fea),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59be81),
	.w1(32'h3b0dd967),
	.w2(32'hbb4aad55),
	.w3(32'h3b3a1556),
	.w4(32'h39aca9c4),
	.w5(32'hbaf3549e),
	.w6(32'hb8e50487),
	.w7(32'h3aa05006),
	.w8(32'hba874ad8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa31f1),
	.w1(32'hbaa7ab2c),
	.w2(32'hbb07d666),
	.w3(32'hbaaba4bb),
	.w4(32'hba9b6e53),
	.w5(32'h39e4486b),
	.w6(32'h386a1daf),
	.w7(32'h3b69de40),
	.w8(32'hbb33aea2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8181b),
	.w1(32'h3c4964be),
	.w2(32'h3bf57ebc),
	.w3(32'hba96d7fc),
	.w4(32'h3c1c505a),
	.w5(32'h3c2884f4),
	.w6(32'hbbac75ff),
	.w7(32'h3b90b46f),
	.w8(32'h3c0b2bcf),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1db54),
	.w1(32'h3a492198),
	.w2(32'hbb4a70d5),
	.w3(32'h3b55441e),
	.w4(32'h3a8595a6),
	.w5(32'hbb7be6d4),
	.w6(32'h3bd006e2),
	.w7(32'h3ae81313),
	.w8(32'h39a7e10b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab40b4e),
	.w1(32'hbaa75c5c),
	.w2(32'hba29e281),
	.w3(32'hbb4ae218),
	.w4(32'hbb5b762b),
	.w5(32'hbad40585),
	.w6(32'hba7a6afe),
	.w7(32'hbbb3150a),
	.w8(32'hbb7addec),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1da68b),
	.w1(32'h3ba24442),
	.w2(32'hba81a3c8),
	.w3(32'h3a91325e),
	.w4(32'h39fbd79a),
	.w5(32'hba833806),
	.w6(32'hbaa6d999),
	.w7(32'hbb07002a),
	.w8(32'hba58595b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39addd58),
	.w1(32'h3bb7545d),
	.w2(32'h3aeaebaf),
	.w3(32'hbb4048fb),
	.w4(32'h3bd29ab2),
	.w5(32'hbb1e6b19),
	.w6(32'hb9828545),
	.w7(32'h3b9bc930),
	.w8(32'h3a1bd104),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc264c),
	.w1(32'hbb178bbb),
	.w2(32'hbaaa6052),
	.w3(32'h3b288542),
	.w4(32'hbb282e95),
	.w5(32'hbb9964ad),
	.w6(32'h3b334109),
	.w7(32'h39a73647),
	.w8(32'h3b348348),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4978aa),
	.w1(32'h3bc76ed5),
	.w2(32'h3b8d3495),
	.w3(32'h3adc55ee),
	.w4(32'h3b8d583a),
	.w5(32'h3c1cb5a4),
	.w6(32'h3bd8eabd),
	.w7(32'h3ad977fd),
	.w8(32'h3bd8680c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b339df9),
	.w1(32'h3b16756b),
	.w2(32'hbaff5940),
	.w3(32'h3b2e550f),
	.w4(32'h3aec10a4),
	.w5(32'hbbae37e1),
	.w6(32'h3bf00d3b),
	.w7(32'h3a62480a),
	.w8(32'h3ba759b8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb754c07),
	.w1(32'hba346b01),
	.w2(32'hbb0362a2),
	.w3(32'h387d6616),
	.w4(32'h3b80d3d8),
	.w5(32'h3b90bf5e),
	.w6(32'h3bacdef8),
	.w7(32'h3b202518),
	.w8(32'hba2361dc),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb963537),
	.w1(32'hbafffdc4),
	.w2(32'hbb247bf0),
	.w3(32'hbab5803a),
	.w4(32'hbb107e8b),
	.w5(32'hbb55b634),
	.w6(32'hbb8f1c3f),
	.w7(32'h3b506aec),
	.w8(32'hbb6303bb),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2874fc),
	.w1(32'h3b8f69eb),
	.w2(32'hb8833d50),
	.w3(32'hbb21b723),
	.w4(32'h3b7650cb),
	.w5(32'h38b1a49f),
	.w6(32'hb83399d9),
	.w7(32'h3b3433f6),
	.w8(32'h3ab2da6b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f7704),
	.w1(32'hbad2b297),
	.w2(32'hb9de31a1),
	.w3(32'h3af8d1f8),
	.w4(32'hbb5db736),
	.w5(32'hbb1c71be),
	.w6(32'hba088958),
	.w7(32'h39e7ea56),
	.w8(32'h3b5af3a4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc404b),
	.w1(32'h3b833ab5),
	.w2(32'hb99dcea2),
	.w3(32'hbb0895dd),
	.w4(32'h3b0746d5),
	.w5(32'h3ae57f34),
	.w6(32'h3b4a2bf5),
	.w7(32'hbbc31af8),
	.w8(32'hbb8913d8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96260e1),
	.w1(32'h3ac1e1ff),
	.w2(32'h3aa42fcc),
	.w3(32'h3a734bc1),
	.w4(32'h3b1dfcf3),
	.w5(32'hbacf6004),
	.w6(32'h39b29855),
	.w7(32'hbb346e41),
	.w8(32'hbb896af3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdcf42),
	.w1(32'hbba2b40b),
	.w2(32'hbba97b34),
	.w3(32'h3b724b09),
	.w4(32'hbb45b40b),
	.w5(32'hbb845ffb),
	.w6(32'h3b677369),
	.w7(32'h3bb347c9),
	.w8(32'hba4a0c25),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f2e49),
	.w1(32'hbbe2f8fe),
	.w2(32'h3b91782a),
	.w3(32'hbb91f528),
	.w4(32'hbbcadcb7),
	.w5(32'hba9e5897),
	.w6(32'hbbbc5e81),
	.w7(32'hbbf6b42c),
	.w8(32'hbb00517d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35c646),
	.w1(32'hbae43227),
	.w2(32'hbaa39086),
	.w3(32'h3b9aab8e),
	.w4(32'h3b461b73),
	.w5(32'hbc0f82b0),
	.w6(32'hbb297576),
	.w7(32'h3be3d86d),
	.w8(32'h3a2d6af4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba822dee),
	.w1(32'h3b26d32c),
	.w2(32'h3b135fdc),
	.w3(32'hba84429b),
	.w4(32'h3af7358d),
	.w5(32'hba00c44e),
	.w6(32'hba3073af),
	.w7(32'h3bbe6d73),
	.w8(32'hbb24e237),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384d80be),
	.w1(32'h3ab91042),
	.w2(32'hbb4b1784),
	.w3(32'h3b46272f),
	.w4(32'h3af45862),
	.w5(32'h3b0b51d6),
	.w6(32'h3b74b77c),
	.w7(32'h3bc131c5),
	.w8(32'h3bdc75d3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba941880),
	.w1(32'h399898b8),
	.w2(32'h3ac87b10),
	.w3(32'hb917a887),
	.w4(32'hbaa30935),
	.w5(32'hbb7138a2),
	.w6(32'h3b82134a),
	.w7(32'h3ac63db5),
	.w8(32'hba6d0d9f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb099cc0),
	.w1(32'h3a8ccc56),
	.w2(32'h3a4c1d1e),
	.w3(32'h3a353676),
	.w4(32'h3b632ee2),
	.w5(32'h3af0d1bb),
	.w6(32'hb9630783),
	.w7(32'hb983a44e),
	.w8(32'hbb46bb9b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ede78),
	.w1(32'hbb1e8966),
	.w2(32'hbb04d24a),
	.w3(32'h3ae35d06),
	.w4(32'h3a0ff2f2),
	.w5(32'hbb217a94),
	.w6(32'hba168efb),
	.w7(32'hbaa43959),
	.w8(32'hbb9b1e68),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba486c92),
	.w1(32'hbbaf8d0c),
	.w2(32'hbad29483),
	.w3(32'hba005ef6),
	.w4(32'hbb956611),
	.w5(32'hbbcecf11),
	.w6(32'h3a538065),
	.w7(32'hbaa155ba),
	.w8(32'hb9ca379c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c3264),
	.w1(32'h3bce67ec),
	.w2(32'h39f0f53e),
	.w3(32'hbaaa70bf),
	.w4(32'hba1be6f1),
	.w5(32'hbae2745f),
	.w6(32'hbb8e2e55),
	.w7(32'hbb313327),
	.w8(32'hbae786ea),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cdcc6e),
	.w1(32'h397024c1),
	.w2(32'h3b1aa3ad),
	.w3(32'h3a07c4f3),
	.w4(32'hb981cbef),
	.w5(32'h3b947cb7),
	.w6(32'h3a06c604),
	.w7(32'hbbefdca8),
	.w8(32'hbbcf0fac),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b399c12),
	.w1(32'hb9729d64),
	.w2(32'hbb37122d),
	.w3(32'h3c0d5b6a),
	.w4(32'h3b9f208d),
	.w5(32'hba3dc1df),
	.w6(32'h3b1debe9),
	.w7(32'h3bb59a90),
	.w8(32'h3ba63bb7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb1659),
	.w1(32'h3b1ca7df),
	.w2(32'hbb11caf9),
	.w3(32'h3aad207f),
	.w4(32'hbb14369e),
	.w5(32'hbb75e439),
	.w6(32'h3b7589b9),
	.w7(32'hb8112902),
	.w8(32'hba2a5388),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae978e3),
	.w1(32'hb9a8ba41),
	.w2(32'hba9beb0f),
	.w3(32'hbb4f5637),
	.w4(32'hbacbccf6),
	.w5(32'hbba01dcf),
	.w6(32'hb8fce572),
	.w7(32'h3a47bd66),
	.w8(32'hb9c09bad),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98ad9a),
	.w1(32'hba3fe0d0),
	.w2(32'hb8a9f9a0),
	.w3(32'h3b7e9bf5),
	.w4(32'hbb819c36),
	.w5(32'h3b6b32bf),
	.w6(32'h3ada5d33),
	.w7(32'hbb3b3490),
	.w8(32'hbb4136e4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0ce67),
	.w1(32'h3b2c7038),
	.w2(32'h3ae5825a),
	.w3(32'hb9fa2460),
	.w4(32'h3aea153d),
	.w5(32'h3c3c081c),
	.w6(32'hb945eb71),
	.w7(32'hbc1c0579),
	.w8(32'hbab1d8c9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08995f),
	.w1(32'hbaaeb234),
	.w2(32'hbaf035ec),
	.w3(32'h3c153534),
	.w4(32'hbb6585de),
	.w5(32'hbbb41d59),
	.w6(32'h3bc287c2),
	.w7(32'h3adcb3ef),
	.w8(32'h3a4fbcf0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13585b),
	.w1(32'hbb402402),
	.w2(32'h375e3acb),
	.w3(32'hbb841185),
	.w4(32'hbb3d3147),
	.w5(32'hbb6a26ce),
	.w6(32'hbb1a6632),
	.w7(32'hb9ed44b4),
	.w8(32'hbba55447),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0312e0),
	.w1(32'hbb29b666),
	.w2(32'h3a4285af),
	.w3(32'h3b1c3455),
	.w4(32'h3a0ff8bc),
	.w5(32'hbb89f9c1),
	.w6(32'h3af733ec),
	.w7(32'h3b209454),
	.w8(32'hbaa7ea31),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35d867),
	.w1(32'hb9d954aa),
	.w2(32'h3c16a7dc),
	.w3(32'hba08f944),
	.w4(32'hbbac33c2),
	.w5(32'h3ad6ad39),
	.w6(32'h3a8fa1d7),
	.w7(32'hbb45cfd7),
	.w8(32'hbb752aa9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0c753),
	.w1(32'h3b43fc00),
	.w2(32'hb9392ed4),
	.w3(32'hb8a989a3),
	.w4(32'h3ba91596),
	.w5(32'hbb441e22),
	.w6(32'hba83211b),
	.w7(32'h3bba1ed7),
	.w8(32'h3bf31b49),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3877a4),
	.w1(32'h3a83c188),
	.w2(32'h3a029a6a),
	.w3(32'hbae28631),
	.w4(32'hbb4778ab),
	.w5(32'hbab0cb38),
	.w6(32'h3b2cc0b2),
	.w7(32'hba68ee85),
	.w8(32'h3a28eed1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58aec7),
	.w1(32'h3bd1476d),
	.w2(32'h3ae638c9),
	.w3(32'h3b1a9930),
	.w4(32'h3babd6e7),
	.w5(32'hbb4d90c0),
	.w6(32'hb83b58de),
	.w7(32'h3bad7d0f),
	.w8(32'h3bbf73b4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7727fe),
	.w1(32'h3a0e1a09),
	.w2(32'h3b43add1),
	.w3(32'hbaad6d7f),
	.w4(32'hba3b925a),
	.w5(32'h3a14eb5d),
	.w6(32'hbabb7219),
	.w7(32'hbb439f3b),
	.w8(32'hba181b76),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd05b3),
	.w1(32'hba6f4ce9),
	.w2(32'hba6ed665),
	.w3(32'h3b8ab020),
	.w4(32'h3ab35b86),
	.w5(32'hbb7e1e1b),
	.w6(32'h3b9f1638),
	.w7(32'hbab5eae2),
	.w8(32'hbab1943f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8f4a0),
	.w1(32'hbb33f87b),
	.w2(32'h3b8c8fb6),
	.w3(32'h3a5447ba),
	.w4(32'hbb5452f0),
	.w5(32'h3aa17250),
	.w6(32'hbb34406f),
	.w7(32'hbb45c5fc),
	.w8(32'h3b0000c8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00dc1d),
	.w1(32'h3c80b3c7),
	.w2(32'h3bbb3877),
	.w3(32'h3b5c5542),
	.w4(32'h3c1308c4),
	.w5(32'h3c25345b),
	.w6(32'hbafb00a2),
	.w7(32'h3b67d59d),
	.w8(32'h3bb32413),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb062af0),
	.w1(32'hbbb02300),
	.w2(32'hba047e84),
	.w3(32'hbbb7b0ed),
	.w4(32'hbb918f3a),
	.w5(32'hbab960e8),
	.w6(32'hbb566e0f),
	.w7(32'hba9ddad3),
	.w8(32'hbaefaa78),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9827d0),
	.w1(32'h3b028abe),
	.w2(32'hbb3fbef3),
	.w3(32'h3973e13d),
	.w4(32'hbb1b9660),
	.w5(32'hbbf53a1a),
	.w6(32'h3a8e788b),
	.w7(32'hbaeb8acf),
	.w8(32'hbb06f9ee),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8b906),
	.w1(32'hbb6acf50),
	.w2(32'hbb58418a),
	.w3(32'hbadfa567),
	.w4(32'hbb45bac1),
	.w5(32'hbbb49a11),
	.w6(32'hbb6834f7),
	.w7(32'h3a322a48),
	.w8(32'hbbb2ca18),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b294372),
	.w1(32'hb9a4cba5),
	.w2(32'hbb3161f3),
	.w3(32'h3a0e12e9),
	.w4(32'h3b260667),
	.w5(32'hb9a02635),
	.w6(32'hbb2df465),
	.w7(32'hbb2b046c),
	.w8(32'hbaf8f17e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3433d8),
	.w1(32'hbb8d5ef6),
	.w2(32'hbac9f1c4),
	.w3(32'h391a84e3),
	.w4(32'hbb0851a8),
	.w5(32'hbb9adeb0),
	.w6(32'hbaea4594),
	.w7(32'hbabfc58a),
	.w8(32'hbb8dd08e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3eae43),
	.w1(32'hbc14a764),
	.w2(32'hbb4c24c3),
	.w3(32'hbaaeddb9),
	.w4(32'hbbb08ac5),
	.w5(32'hbb2fdccf),
	.w6(32'hbb1874e9),
	.w7(32'hb9e61093),
	.w8(32'h3ab07c54),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7256d),
	.w1(32'hbb73520b),
	.w2(32'h3ad48096),
	.w3(32'h3b93fe22),
	.w4(32'hbb3c33b6),
	.w5(32'hb5225add),
	.w6(32'h3b3e1b7d),
	.w7(32'hb9e3ffdc),
	.w8(32'h3ac4c861),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a178290),
	.w1(32'h3a0258e9),
	.w2(32'h3b693776),
	.w3(32'hba8efe14),
	.w4(32'h3a891cf4),
	.w5(32'h3c4ccdbf),
	.w6(32'hbb0f37c3),
	.w7(32'hbb6bef2c),
	.w8(32'h3ab6d0c4),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acda0b7),
	.w1(32'hba5e8de8),
	.w2(32'h390e6688),
	.w3(32'h3bd81389),
	.w4(32'h3aa864a7),
	.w5(32'hbb34a8f7),
	.w6(32'h3b5d03d7),
	.w7(32'h3b27ed76),
	.w8(32'hbb0ca6f6),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb942926c),
	.w1(32'h3b5414e4),
	.w2(32'hb98617e9),
	.w3(32'h3a39d5cb),
	.w4(32'hbace25f5),
	.w5(32'hbb21aacc),
	.w6(32'h3a93460e),
	.w7(32'hbb06a32d),
	.w8(32'hb9fbc7d7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08f120),
	.w1(32'hbb22e7fa),
	.w2(32'h3bebcbe1),
	.w3(32'hb930faf7),
	.w4(32'hbb9bfced),
	.w5(32'hbaeaf171),
	.w6(32'h3a95d4f0),
	.w7(32'hbb15f2fe),
	.w8(32'h3b04178d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ded14),
	.w1(32'h3b0bb0d6),
	.w2(32'hba960a60),
	.w3(32'hbb39c2ee),
	.w4(32'hb90b7677),
	.w5(32'h39d2932b),
	.w6(32'hbb3b82f7),
	.w7(32'h3a105a93),
	.w8(32'hba93074a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b131c),
	.w1(32'hbabaeae9),
	.w2(32'hbab55537),
	.w3(32'h3b1eb117),
	.w4(32'h3a2b0f1a),
	.w5(32'hba3d0d46),
	.w6(32'h3adf98fd),
	.w7(32'h3b70a463),
	.w8(32'hbaf991f6),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38a368),
	.w1(32'hbb76290c),
	.w2(32'h39ead6ae),
	.w3(32'hb982cf87),
	.w4(32'hba9cb98b),
	.w5(32'hbb9bf423),
	.w6(32'hba5064e0),
	.w7(32'hbb4010ad),
	.w8(32'hbb13e48d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b294cb7),
	.w1(32'h39209fb1),
	.w2(32'h39e667e0),
	.w3(32'hbaef6366),
	.w4(32'h37556657),
	.w5(32'hbb5983c9),
	.w6(32'hbb7f1553),
	.w7(32'hbab81811),
	.w8(32'hba3835f6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c99bb),
	.w1(32'hbb2b7d67),
	.w2(32'h3bfbe761),
	.w3(32'hba0df22b),
	.w4(32'hba9d77b9),
	.w5(32'h398b8440),
	.w6(32'h3b9a3351),
	.w7(32'hbb598cc9),
	.w8(32'h3b8df5c4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb093ae),
	.w1(32'hba3bdee8),
	.w2(32'h3a8f81d0),
	.w3(32'h3aa75e60),
	.w4(32'hbb3c32bc),
	.w5(32'h3b4433d3),
	.w6(32'h3bc51274),
	.w7(32'hba86f0e5),
	.w8(32'hba9baf26),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a5bcd),
	.w1(32'hba940cb6),
	.w2(32'h3ad4c347),
	.w3(32'h3b167aa9),
	.w4(32'hbb2e4389),
	.w5(32'hbb048819),
	.w6(32'h3af711c5),
	.w7(32'hbb8a29df),
	.w8(32'hbb103f42),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea84e2),
	.w1(32'h3b74d718),
	.w2(32'hbb4ced66),
	.w3(32'h39b587b8),
	.w4(32'h3bb8a83b),
	.w5(32'h38a4453b),
	.w6(32'hbb025180),
	.w7(32'h3bc14b1e),
	.w8(32'hb7a2a2f0),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae39468),
	.w1(32'hbb6fca3f),
	.w2(32'hbb6c8cd6),
	.w3(32'hbb428d60),
	.w4(32'hbbf09af9),
	.w5(32'hbbcd7a27),
	.w6(32'hbb4fe1ec),
	.w7(32'hbb94c8cd),
	.w8(32'hbb6afdca),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabbb74),
	.w1(32'h3befc6ff),
	.w2(32'h3bbe21f8),
	.w3(32'hbaf2ce8c),
	.w4(32'h3b24d504),
	.w5(32'h3b4ca737),
	.w6(32'h3889d66e),
	.w7(32'h3a17be03),
	.w8(32'h3b3b83e7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7389d2),
	.w1(32'hb9e22469),
	.w2(32'hbb40a85f),
	.w3(32'h3bdf989e),
	.w4(32'h3bb55a2d),
	.w5(32'hbb8affe6),
	.w6(32'h3bc162c2),
	.w7(32'h3a819303),
	.w8(32'hbb6734fa),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e71951),
	.w1(32'h3b6c28c3),
	.w2(32'hbb87f00a),
	.w3(32'hba59e18f),
	.w4(32'h3bf62774),
	.w5(32'hbbaaf633),
	.w6(32'hb959fe60),
	.w7(32'h3b514ef7),
	.w8(32'hbb690f33),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b134c2f),
	.w1(32'h3b259e99),
	.w2(32'h3abfee40),
	.w3(32'hbb094914),
	.w4(32'h39244eb1),
	.w5(32'hbb2f1351),
	.w6(32'hbb786d7e),
	.w7(32'hb9e70a5f),
	.w8(32'hbb2bf964),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2dee7d),
	.w1(32'h3bfed55e),
	.w2(32'h3b487f6b),
	.w3(32'hb9ff6718),
	.w4(32'h3c08e2a5),
	.w5(32'h3baf98dd),
	.w6(32'hbab38fb6),
	.w7(32'h3b6c9cb8),
	.w8(32'h3b54e219),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e08d8),
	.w1(32'h3b1386c1),
	.w2(32'h3a376ff9),
	.w3(32'h3b8bed4b),
	.w4(32'h3b76abc4),
	.w5(32'hbab19b18),
	.w6(32'h3b32207d),
	.w7(32'h3b1f6c19),
	.w8(32'hbb1c499a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a396748),
	.w1(32'h3c74d082),
	.w2(32'hbb96c4eb),
	.w3(32'hbacb30d3),
	.w4(32'h3c392227),
	.w5(32'hbba51df8),
	.w6(32'hbb026265),
	.w7(32'h3b680811),
	.w8(32'h3b8b3b71),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad49729),
	.w1(32'hbaa677ad),
	.w2(32'hbb6c55df),
	.w3(32'hba1d1a8a),
	.w4(32'hb8e2627b),
	.w5(32'hbb9c70f9),
	.w6(32'hbae45973),
	.w7(32'h3a2c8bd0),
	.w8(32'hbae1ca34),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13c579),
	.w1(32'h3b303053),
	.w2(32'hbba7245d),
	.w3(32'hbb06e174),
	.w4(32'h3b33e14c),
	.w5(32'hbb8860e8),
	.w6(32'hbad504d7),
	.w7(32'h3983abd3),
	.w8(32'hbadc6b35),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac331c0),
	.w1(32'hb99f5c66),
	.w2(32'h3b8804a8),
	.w3(32'h3a6f09bb),
	.w4(32'h3ab5d7cd),
	.w5(32'h39b45764),
	.w6(32'h3b2be702),
	.w7(32'hbba676f8),
	.w8(32'hbb34c432),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a98056),
	.w1(32'h3a8dfc3a),
	.w2(32'hbb7a00b3),
	.w3(32'h3aa4511a),
	.w4(32'h3b08fcf6),
	.w5(32'hbad8dac1),
	.w6(32'hba954e7e),
	.w7(32'hba4eac35),
	.w8(32'hbbb2d718),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcc579),
	.w1(32'hbc36407e),
	.w2(32'hbbba0b14),
	.w3(32'hba87c3e9),
	.w4(32'hba9b3676),
	.w5(32'hbbed5d8f),
	.w6(32'hbb278832),
	.w7(32'hbac63976),
	.w8(32'hbbc9069b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab89e12),
	.w1(32'hbb6e947b),
	.w2(32'h399e1c9f),
	.w3(32'hbb36df43),
	.w4(32'hba8ee33f),
	.w5(32'hb993e808),
	.w6(32'hba137844),
	.w7(32'h39f23d61),
	.w8(32'h3b2ecad7),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a480c08),
	.w1(32'hbbefc9fb),
	.w2(32'hbb134266),
	.w3(32'h3aa3ccd7),
	.w4(32'hba8c262c),
	.w5(32'hbb0a4a69),
	.w6(32'h3b87e942),
	.w7(32'h3a91b25d),
	.w8(32'h3b3290c7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a742db2),
	.w1(32'hba35b3f1),
	.w2(32'hbb11d29c),
	.w3(32'h3b53d608),
	.w4(32'hba86a4a0),
	.w5(32'hbbb5e69d),
	.w6(32'h3b5d6001),
	.w7(32'hba8545ea),
	.w8(32'hbb9cada1),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4de81),
	.w1(32'hbb3abd34),
	.w2(32'hbab99303),
	.w3(32'hbb48212b),
	.w4(32'hbb51a633),
	.w5(32'hbb8d1c7d),
	.w6(32'hbb11565a),
	.w7(32'hbbb5ef4f),
	.w8(32'hbb888a03),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5abe25),
	.w1(32'h3a040eb8),
	.w2(32'hbb9eb607),
	.w3(32'hba93b6ad),
	.w4(32'h3aaa2738),
	.w5(32'hbb29fba2),
	.w6(32'hbc12afa8),
	.w7(32'h3b8a6b55),
	.w8(32'hbb0731fa),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9ae54),
	.w1(32'h3a8633d9),
	.w2(32'hbb1df170),
	.w3(32'hbba2bb0e),
	.w4(32'h3b998dba),
	.w5(32'hba1105a3),
	.w6(32'hbb96fd66),
	.w7(32'hbb615b89),
	.w8(32'h3b9b92e4),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a3bfe),
	.w1(32'hbb6ea797),
	.w2(32'h3a8eaf3a),
	.w3(32'h3a741b5f),
	.w4(32'hbb3c75a0),
	.w5(32'hbb0440f2),
	.w6(32'hb9cf41fd),
	.w7(32'hb8d92acd),
	.w8(32'hbaab4987),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb019be3),
	.w1(32'h3b7c48b4),
	.w2(32'h3b0d5546),
	.w3(32'hbb38a895),
	.w4(32'h394b3c3a),
	.w5(32'h3ba3e6fa),
	.w6(32'hba875b0d),
	.w7(32'h3a27d246),
	.w8(32'hbaaa00e7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf02d44),
	.w1(32'hbabfc427),
	.w2(32'hbb03ecd6),
	.w3(32'h3ae4a3e7),
	.w4(32'h3b8d1672),
	.w5(32'hb9d93251),
	.w6(32'h38c21c11),
	.w7(32'h397e558c),
	.w8(32'hbb80b9ff),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac67c52),
	.w1(32'h3b15dcfd),
	.w2(32'h3b0495c8),
	.w3(32'h3b2ae25e),
	.w4(32'h3b6ce474),
	.w5(32'h3b0c95d1),
	.w6(32'hbadf89ae),
	.w7(32'hba1d2b9a),
	.w8(32'hbb610e4e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb1e69),
	.w1(32'h3b30f261),
	.w2(32'h3a191b1c),
	.w3(32'h3ba3abf2),
	.w4(32'h39fdd8bb),
	.w5(32'hbb106fd2),
	.w6(32'h3b183097),
	.w7(32'hb6ccc6f4),
	.w8(32'hbaf56925),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02c67c),
	.w1(32'hbb2fc06e),
	.w2(32'hbb1d2f89),
	.w3(32'hbb37309f),
	.w4(32'hbb8c7d2c),
	.w5(32'hbb61604c),
	.w6(32'hbaad1cfd),
	.w7(32'hbb8ae14e),
	.w8(32'hbb323832),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac1c84),
	.w1(32'h3af6c979),
	.w2(32'h39aa3254),
	.w3(32'hbbb67099),
	.w4(32'h3adc074e),
	.w5(32'h3a380f8a),
	.w6(32'hbbd68ddb),
	.w7(32'h3a775035),
	.w8(32'h3b11971c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05077e),
	.w1(32'hb9bdfce1),
	.w2(32'h3be17926),
	.w3(32'hb905abb0),
	.w4(32'h3815fbba),
	.w5(32'h3c15985a),
	.w6(32'h3b877cd9),
	.w7(32'hbb819417),
	.w8(32'h3bc7bc9e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af72442),
	.w1(32'h3adc5381),
	.w2(32'h3883fa29),
	.w3(32'h3c074b0e),
	.w4(32'h397c1072),
	.w5(32'h3a9c9807),
	.w6(32'h3b95396d),
	.w7(32'h39c2cabd),
	.w8(32'h3b5f03f8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ee2e1),
	.w1(32'h3b33be88),
	.w2(32'hb8821c22),
	.w3(32'hbba540a0),
	.w4(32'h39f03e47),
	.w5(32'h3b83937d),
	.w6(32'h3b36a6dc),
	.w7(32'h3a2aa7a3),
	.w8(32'h3b429dd2),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c3ad4),
	.w1(32'hba9fbb3c),
	.w2(32'hbb37029e),
	.w3(32'hbada7db1),
	.w4(32'h3ab9db98),
	.w5(32'hbb757a79),
	.w6(32'hba1fc75a),
	.w7(32'h3abad1b7),
	.w8(32'hba18bfca),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c95f0),
	.w1(32'hbabbcb7f),
	.w2(32'hbb5d6dc4),
	.w3(32'hbb513e4b),
	.w4(32'hbb1f91ff),
	.w5(32'hbbb30313),
	.w6(32'hbacc4adc),
	.w7(32'h3a6976c3),
	.w8(32'hbbc314d1),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9b093),
	.w1(32'h3b95caa7),
	.w2(32'h3ca83281),
	.w3(32'hbbdf4911),
	.w4(32'h3b19ce33),
	.w5(32'h3cc21588),
	.w6(32'hbbe66866),
	.w7(32'h39ecbd53),
	.w8(32'h3c760998),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98822f),
	.w1(32'h3b95ec51),
	.w2(32'h39c323ec),
	.w3(32'h3c1777b2),
	.w4(32'h3a9bef0d),
	.w5(32'hbb75c19e),
	.w6(32'h3c25fc77),
	.w7(32'h39a4a7ec),
	.w8(32'hbb348c2e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71b586),
	.w1(32'h3b8c507a),
	.w2(32'hb85beb80),
	.w3(32'h3b734049),
	.w4(32'h3becb703),
	.w5(32'hbbd39794),
	.w6(32'h3b387234),
	.w7(32'h3b050c93),
	.w8(32'hbb3f037d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b0d09f),
	.w1(32'h3a7947f4),
	.w2(32'hb9b818b1),
	.w3(32'hb9d9aa5e),
	.w4(32'hb97daa1e),
	.w5(32'hbb216ce7),
	.w6(32'hbad867c3),
	.w7(32'hba91c9ba),
	.w8(32'h3b954425),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e40f9),
	.w1(32'h39c9db8a),
	.w2(32'h3a877408),
	.w3(32'hb9b664ca),
	.w4(32'h3b4892d2),
	.w5(32'hbadfa34a),
	.w6(32'h3b0a5b6f),
	.w7(32'hbaac40a5),
	.w8(32'h3a0cf44e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1e6fb),
	.w1(32'h3bfdb327),
	.w2(32'h39a7ef95),
	.w3(32'hbae3d351),
	.w4(32'h3be34a87),
	.w5(32'hbb36e479),
	.w6(32'hbb9c776c),
	.w7(32'h3b9937c0),
	.w8(32'h3b54fe71),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8573af),
	.w1(32'hbb8045bd),
	.w2(32'h3a252399),
	.w3(32'h3b499811),
	.w4(32'hbb8b3722),
	.w5(32'h39b0c640),
	.w6(32'h3bb5bbe6),
	.w7(32'h3a3d2679),
	.w8(32'h3b84b097),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39423934),
	.w1(32'h3a9dd15d),
	.w2(32'h3b7b4e46),
	.w3(32'hbaa934e4),
	.w4(32'h3ba1c1c3),
	.w5(32'h36db89d7),
	.w6(32'h3aeb8e70),
	.w7(32'h3bccc8a5),
	.w8(32'hb91dd2df),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73e96e),
	.w1(32'hbac7602a),
	.w2(32'hbb306c3e),
	.w3(32'hba467aee),
	.w4(32'hbac6a594),
	.w5(32'hbb8d864d),
	.w6(32'hbb1c634f),
	.w7(32'hb96e502c),
	.w8(32'hba57348e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f7bf4),
	.w1(32'h3b30e17b),
	.w2(32'hbb2383fc),
	.w3(32'h3b768d05),
	.w4(32'h3bc5dbe2),
	.w5(32'hbb3d9c92),
	.w6(32'h39b18c04),
	.w7(32'h3b0ad648),
	.w8(32'hba6d3e6d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfd27e),
	.w1(32'h3b1813f6),
	.w2(32'hbb41e44c),
	.w3(32'hb9f97fee),
	.w4(32'h3ac09ae9),
	.w5(32'hba06a23f),
	.w6(32'h3b4b1791),
	.w7(32'h39460e84),
	.w8(32'hbaa6468e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb533024),
	.w1(32'h3bdb1492),
	.w2(32'h3ac74ce0),
	.w3(32'hbad00efe),
	.w4(32'h3bc0ef4b),
	.w5(32'h3a8fbfd5),
	.w6(32'h3adf257d),
	.w7(32'h3b643565),
	.w8(32'h3b81f95a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a6d22),
	.w1(32'h3b10df39),
	.w2(32'hb9832613),
	.w3(32'hbb3a1f63),
	.w4(32'h3ab1cae8),
	.w5(32'h3b36269d),
	.w6(32'h3bae156e),
	.w7(32'hbadbbc0a),
	.w8(32'hbb160535),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb001faf),
	.w1(32'hbba8e6d4),
	.w2(32'hbb59ae6c),
	.w3(32'hb88d73d8),
	.w4(32'hbb5ee0d8),
	.w5(32'h3a385208),
	.w6(32'h3ad6c3c5),
	.w7(32'hba8f2c25),
	.w8(32'hb9e44291),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d5286),
	.w1(32'hba171283),
	.w2(32'h3b8a9189),
	.w3(32'hbb175723),
	.w4(32'h39262265),
	.w5(32'hbb37610b),
	.w6(32'hbb6fe850),
	.w7(32'h3bc7c2a8),
	.w8(32'hbb445614),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f7999),
	.w1(32'hbba8137f),
	.w2(32'h3a1c4aab),
	.w3(32'h3aac41e0),
	.w4(32'hbbbc155c),
	.w5(32'h3affbe8f),
	.w6(32'h3b3f9df3),
	.w7(32'hbb64fd76),
	.w8(32'h3a8754fe),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390de421),
	.w1(32'hbb1443c5),
	.w2(32'hbb9606cc),
	.w3(32'hbb66cf92),
	.w4(32'h3a859ec1),
	.w5(32'hbc1b81c8),
	.w6(32'hbb17306e),
	.w7(32'h3bb9161c),
	.w8(32'h3c49425a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83241c),
	.w1(32'hbbfd5ae7),
	.w2(32'h38bf6146),
	.w3(32'hbb5c4a41),
	.w4(32'hbb5da3a2),
	.w5(32'hbb954cc5),
	.w6(32'h3ba0efa2),
	.w7(32'hba05624f),
	.w8(32'h3ab008d7),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40c9b8),
	.w1(32'hb9e0f106),
	.w2(32'hba6b0fd6),
	.w3(32'hbb8cbff4),
	.w4(32'hba7ee080),
	.w5(32'hbb0ea922),
	.w6(32'hb99597c1),
	.w7(32'hbab264bc),
	.w8(32'hb9984238),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ecb11),
	.w1(32'h3910706e),
	.w2(32'h3b161b39),
	.w3(32'hb9bff853),
	.w4(32'hbaf4742b),
	.w5(32'hbabfe799),
	.w6(32'hbac06857),
	.w7(32'h3ae2a256),
	.w8(32'hbb1072ce),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d10d8),
	.w1(32'h39d30b2b),
	.w2(32'hbac77e78),
	.w3(32'h3a04d5f6),
	.w4(32'h3adce097),
	.w5(32'h3b916982),
	.w6(32'h3b05dcfc),
	.w7(32'h3ae23135),
	.w8(32'h3a8c5aec),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d3787),
	.w1(32'h3bca8687),
	.w2(32'h3bab8a20),
	.w3(32'h3b011f1e),
	.w4(32'h3b823b1b),
	.w5(32'h3bb2b6fc),
	.w6(32'hb8e680ed),
	.w7(32'h3b3e9c37),
	.w8(32'h3b9327b4),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8de9fa),
	.w1(32'hb9cc0616),
	.w2(32'h3bb6cc18),
	.w3(32'h3b6632d2),
	.w4(32'hbb1c6c09),
	.w5(32'hb8c7bf4c),
	.w6(32'h3bbc0b7d),
	.w7(32'hbb95247e),
	.w8(32'hbb096a14),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bd706),
	.w1(32'h3aab791f),
	.w2(32'h3ac1eb52),
	.w3(32'h3b8d1068),
	.w4(32'h3b9730ac),
	.w5(32'hbb10a2fc),
	.w6(32'h3af97bff),
	.w7(32'h3b483b18),
	.w8(32'h3b5bb967),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fa6104),
	.w1(32'hbb52af58),
	.w2(32'hb9d37db1),
	.w3(32'hba033d27),
	.w4(32'h3b8a6793),
	.w5(32'hbb407aed),
	.w6(32'h39cd5297),
	.w7(32'h3bbe67df),
	.w8(32'h3b170124),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff9c22),
	.w1(32'hbb5cae9f),
	.w2(32'h3b8dcff5),
	.w3(32'h3b4124ed),
	.w4(32'hbb8686cd),
	.w5(32'hbab438bc),
	.w6(32'h3a882be7),
	.w7(32'hbb2bd10a),
	.w8(32'hbb929714),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b45cd),
	.w1(32'h3b08ed55),
	.w2(32'h3b808600),
	.w3(32'h3bf919cf),
	.w4(32'h3adbd16b),
	.w5(32'h3b5716cb),
	.w6(32'h3ab89ab7),
	.w7(32'h39625957),
	.w8(32'h3a7bd1c6),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b178f23),
	.w1(32'hbb114ca9),
	.w2(32'hba93152e),
	.w3(32'h3a20cb96),
	.w4(32'h3ae46ebf),
	.w5(32'h3a9325f7),
	.w6(32'h3a1e8fee),
	.w7(32'h3b980f5f),
	.w8(32'h3be0c8e2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4004ba),
	.w1(32'h3b253315),
	.w2(32'hbb4cbf7e),
	.w3(32'h3abf7276),
	.w4(32'h3c235675),
	.w5(32'h3c515ed1),
	.w6(32'h3be2a107),
	.w7(32'hba028d26),
	.w8(32'h3afbc105),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7134b),
	.w1(32'hba9d018f),
	.w2(32'hbb13be59),
	.w3(32'h3c44f7db),
	.w4(32'h3b1edc1d),
	.w5(32'h3a0bd177),
	.w6(32'h3b4599ad),
	.w7(32'hbb848d30),
	.w8(32'hbbc1bba0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb9ed0),
	.w1(32'h3b340b4e),
	.w2(32'h3b279978),
	.w3(32'hbb94c82c),
	.w4(32'hbb33af54),
	.w5(32'hbb3b9ed2),
	.w6(32'hbb38d6be),
	.w7(32'hbaac73d0),
	.w8(32'hbb014a6d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1d509),
	.w1(32'hbaefb3ff),
	.w2(32'hbb569fe1),
	.w3(32'hbb31194c),
	.w4(32'h3c218508),
	.w5(32'h3b4cfddf),
	.w6(32'hbab84235),
	.w7(32'hbb8cd54e),
	.w8(32'hbb8dc14c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9044e4),
	.w1(32'h3a29cbcc),
	.w2(32'h3af3ced6),
	.w3(32'hbb0f2a2b),
	.w4(32'h3b32d6e4),
	.w5(32'h3b8e9f6b),
	.w6(32'hbb6409e3),
	.w7(32'hbb123bf4),
	.w8(32'hba5348d6),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7883ee),
	.w1(32'h3b081f5e),
	.w2(32'h3ad535cd),
	.w3(32'h3af49dca),
	.w4(32'h3a844340),
	.w5(32'hbb129615),
	.w6(32'hba183633),
	.w7(32'h3b31d70a),
	.w8(32'hba05edbc),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad59e14),
	.w1(32'h3a2b5340),
	.w2(32'h3af1a1d0),
	.w3(32'hbb30875a),
	.w4(32'h39678f76),
	.w5(32'hbaafa710),
	.w6(32'h3aa44acb),
	.w7(32'h3a83963b),
	.w8(32'h3b634698),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4394a),
	.w1(32'hba2d3e5e),
	.w2(32'hbb22bf77),
	.w3(32'hb9ff6399),
	.w4(32'hbabb08cf),
	.w5(32'hbabc048e),
	.w6(32'hbb46970d),
	.w7(32'h37f7bf77),
	.w8(32'h39accbb4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb485740),
	.w1(32'h3a9228e7),
	.w2(32'h3b398e9c),
	.w3(32'h3acfafbc),
	.w4(32'hbadaeedc),
	.w5(32'hbb11085b),
	.w6(32'h3b377474),
	.w7(32'h3b36822e),
	.w8(32'hbaabe9ea),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48d049),
	.w1(32'h3a1a9ff2),
	.w2(32'h3a6d9d05),
	.w3(32'hb9cf3eb9),
	.w4(32'hbab0cce3),
	.w5(32'hba8cd452),
	.w6(32'h3a59fa22),
	.w7(32'h3ac034cf),
	.w8(32'hb90d0998),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b67cb),
	.w1(32'hbaed3385),
	.w2(32'hbb3377be),
	.w3(32'hbad89124),
	.w4(32'hb902cc11),
	.w5(32'hba6b6710),
	.w6(32'hb9d31d1e),
	.w7(32'h3a02d63d),
	.w8(32'hba86da75),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399738e8),
	.w1(32'hba4dd126),
	.w2(32'hb946b377),
	.w3(32'hb998bbd1),
	.w4(32'hba791461),
	.w5(32'h39db4bf4),
	.w6(32'hbaa4199c),
	.w7(32'h3b4fce21),
	.w8(32'h3bbfa135),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5611b),
	.w1(32'hbb91dfe9),
	.w2(32'h3b00b0ab),
	.w3(32'h3b737c2d),
	.w4(32'h3a197afc),
	.w5(32'h3b2c18a1),
	.w6(32'h3baebe67),
	.w7(32'hbae4f32e),
	.w8(32'hbbdbfc14),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2799e1),
	.w1(32'hbb658ba9),
	.w2(32'hbb3ab67b),
	.w3(32'hb9bd4c35),
	.w4(32'h3c1d9a83),
	.w5(32'h3bfb3b82),
	.w6(32'hbbc027e1),
	.w7(32'hbae4beb8),
	.w8(32'hbaffb19d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac86265),
	.w1(32'hba86a4d4),
	.w2(32'hb9c51651),
	.w3(32'h3a062531),
	.w4(32'hb8cb3889),
	.w5(32'hbae42f53),
	.w6(32'hbac97e9a),
	.w7(32'hba9af6a7),
	.w8(32'hb9bf13ee),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa70c4),
	.w1(32'h3b609ed3),
	.w2(32'h3b921ad6),
	.w3(32'hba6a3dee),
	.w4(32'hbb16eba5),
	.w5(32'hb95cca4b),
	.w6(32'h37e4ed8b),
	.w7(32'h3b82a203),
	.w8(32'h3b4768e7),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbf80f),
	.w1(32'h3b67f07b),
	.w2(32'h3b2b70c7),
	.w3(32'h3b887d2d),
	.w4(32'hba9a312e),
	.w5(32'hba526f7f),
	.w6(32'h3ab6db16),
	.w7(32'h38bd610d),
	.w8(32'h3aa9923f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b96de),
	.w1(32'hb9ef4f88),
	.w2(32'h3a5358c6),
	.w3(32'hbaabe9b1),
	.w4(32'h3a2b69ae),
	.w5(32'h39cc2043),
	.w6(32'h392f1760),
	.w7(32'h3b287583),
	.w8(32'hba97100e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55b520),
	.w1(32'hb9b330ea),
	.w2(32'h3a3953fb),
	.w3(32'hbb1a49f4),
	.w4(32'hbb0abf1b),
	.w5(32'hba9a1769),
	.w6(32'h39fc5b07),
	.w7(32'hbb45bd0d),
	.w8(32'hbacb54f7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb459e59),
	.w1(32'hb89af1c2),
	.w2(32'h3a0f29b8),
	.w3(32'hbabadd10),
	.w4(32'hba877a6c),
	.w5(32'h3a716a26),
	.w6(32'hba5ec1d5),
	.w7(32'h3a21a8fb),
	.w8(32'hba2535fe),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b776559),
	.w1(32'h3b122133),
	.w2(32'h3b1c16e8),
	.w3(32'h381bbfea),
	.w4(32'h39d9c60a),
	.w5(32'h3af539d5),
	.w6(32'hbaa7364e),
	.w7(32'h3b1136a0),
	.w8(32'hba7d17aa),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3294a3),
	.w1(32'hba9272a2),
	.w2(32'h37c31a18),
	.w3(32'h3b47bcc5),
	.w4(32'h3be59729),
	.w5(32'h3c3308f2),
	.w6(32'hb8fa7787),
	.w7(32'h3a9a4043),
	.w8(32'h3aefea80),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77cdea),
	.w1(32'hb989a7a1),
	.w2(32'h3ad434f3),
	.w3(32'h3c00d43c),
	.w4(32'hbb434158),
	.w5(32'hbb12fcf0),
	.w6(32'h3b4d5fef),
	.w7(32'hba9a1574),
	.w8(32'hbb5e34c8),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bfaf1),
	.w1(32'h3a394cc9),
	.w2(32'h397f4856),
	.w3(32'hbb70f517),
	.w4(32'h3b0a6d9c),
	.w5(32'hb9cf87b5),
	.w6(32'hbb7d3533),
	.w7(32'h3afa5bd7),
	.w8(32'hbba277fb),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4dd90b),
	.w1(32'hbb1261bb),
	.w2(32'hba3e4a75),
	.w3(32'h3b31ac7e),
	.w4(32'h3b1db3ed),
	.w5(32'hbb4b1029),
	.w6(32'h3aa811a0),
	.w7(32'hbab7f8c5),
	.w8(32'hbb5227a9),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1321b1),
	.w1(32'h39a5402a),
	.w2(32'hbb3b7ad0),
	.w3(32'hbb96dcd8),
	.w4(32'hb9d5a690),
	.w5(32'hbb7177b5),
	.w6(32'hba1ef72b),
	.w7(32'hbb1ae6cc),
	.w8(32'hbb4536bf),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d74b4),
	.w1(32'h3ab8817a),
	.w2(32'hba835b2f),
	.w3(32'hbb5848ee),
	.w4(32'hb980c514),
	.w5(32'hbb0f786c),
	.w6(32'h3a857338),
	.w7(32'hbb453b55),
	.w8(32'hbbbc21db),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f048ba),
	.w1(32'hbac42870),
	.w2(32'hbac9e878),
	.w3(32'h3853fbb0),
	.w4(32'hba5b74d1),
	.w5(32'hbb0b192c),
	.w6(32'hbb40e20d),
	.w7(32'hbb3a33d8),
	.w8(32'h3950d154),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbad09),
	.w1(32'hb95be2f8),
	.w2(32'h3a56c9e2),
	.w3(32'hbb37aabf),
	.w4(32'h3c1c7610),
	.w5(32'h3beef238),
	.w6(32'h39fb4b79),
	.w7(32'hbb8d08ae),
	.w8(32'hbb3c44a5),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7be3fba),
	.w1(32'h3ad01b76),
	.w2(32'h3938b5cd),
	.w3(32'h3b84ed39),
	.w4(32'hbb92a856),
	.w5(32'hbb612b53),
	.w6(32'hbaf188a2),
	.w7(32'h3b084144),
	.w8(32'h38059f35),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919f2a2),
	.w1(32'hbb93d605),
	.w2(32'hbb258b0e),
	.w3(32'hbb0f9ee0),
	.w4(32'h3bfcca9a),
	.w5(32'h39966f73),
	.w6(32'h38620ea2),
	.w7(32'h3abf698d),
	.w8(32'hbb2dae78),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae48343),
	.w1(32'h3b7e9d29),
	.w2(32'h3a5e0687),
	.w3(32'hbad0d2a6),
	.w4(32'h3afe0b7f),
	.w5(32'hbae4401b),
	.w6(32'hb9f74300),
	.w7(32'h3b0dbc9c),
	.w8(32'hb9adb654),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39931071),
	.w1(32'h3a02f109),
	.w2(32'h3b1792f2),
	.w3(32'hbb578a06),
	.w4(32'hb9e5b7a0),
	.w5(32'h3af219a9),
	.w6(32'hb9fb0332),
	.w7(32'h3a35dfd9),
	.w8(32'h3b62ece1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3901ca),
	.w1(32'hbbada637),
	.w2(32'hbb1a50ee),
	.w3(32'h3a9239a3),
	.w4(32'h3bb5cd39),
	.w5(32'h3b97790d),
	.w6(32'h3be13d54),
	.w7(32'h3b69dfb5),
	.w8(32'h3b709db1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4fb27),
	.w1(32'hb8e577d9),
	.w2(32'h39a2c2f1),
	.w3(32'h3b89a967),
	.w4(32'h39e2bb06),
	.w5(32'h3a9d4bf2),
	.w6(32'h3bf9d5de),
	.w7(32'h3b13dc6e),
	.w8(32'h3b127173),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a993006),
	.w1(32'hb95aefa6),
	.w2(32'hb9aff7bd),
	.w3(32'h38800ab1),
	.w4(32'h3a6f2c53),
	.w5(32'hb9b2a24b),
	.w6(32'h3af49856),
	.w7(32'hbb0ed804),
	.w8(32'hba821a2d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab30c48),
	.w1(32'hba26434a),
	.w2(32'h3b1456f5),
	.w3(32'h3b5245c3),
	.w4(32'h3a91067d),
	.w5(32'h3b19354f),
	.w6(32'hba6daa18),
	.w7(32'hb931a1ff),
	.w8(32'hb8c15bfe),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2c733),
	.w1(32'hbb081e5a),
	.w2(32'hbafa88d0),
	.w3(32'hba42ef4c),
	.w4(32'h3bb312cf),
	.w5(32'h3b9e25f9),
	.w6(32'hbb500dbf),
	.w7(32'hb7ea52e5),
	.w8(32'h3b696564),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea36e4),
	.w1(32'hbb9962f7),
	.w2(32'hbb329c1d),
	.w3(32'h3b36e8b2),
	.w4(32'h3bbfec54),
	.w5(32'h3af32788),
	.w6(32'h3b2b5ce6),
	.w7(32'h3bdcfc01),
	.w8(32'hb8ba1d5e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb966dd8c),
	.w1(32'h3b94b162),
	.w2(32'h3a68acd7),
	.w3(32'h3aaf7801),
	.w4(32'h3aaa3fe8),
	.w5(32'h3a6bcf5d),
	.w6(32'h3b8c6a06),
	.w7(32'hbad69fbc),
	.w8(32'hba522e2b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39e509),
	.w1(32'h3ac6c359),
	.w2(32'hb8d24644),
	.w3(32'h3a120d93),
	.w4(32'h3a79f0b5),
	.w5(32'hba9f055a),
	.w6(32'hbb2639f4),
	.w7(32'hba0307bf),
	.w8(32'hbb961568),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77f46f),
	.w1(32'hbad44cbd),
	.w2(32'hbb2f3481),
	.w3(32'hbb344c6b),
	.w4(32'h3a74107f),
	.w5(32'hbad73d7a),
	.w6(32'hbb9a1925),
	.w7(32'hbb4595b7),
	.w8(32'hbbad74b7),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01c59e),
	.w1(32'h3a92d986),
	.w2(32'hb9b65f3f),
	.w3(32'hbb2fb727),
	.w4(32'hbbc1938a),
	.w5(32'hbb9aca5f),
	.w6(32'hb9f4c24b),
	.w7(32'hba7218f6),
	.w8(32'hbb4b90a7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91b495),
	.w1(32'h3b38460a),
	.w2(32'h3a75a24f),
	.w3(32'hbb54bf8d),
	.w4(32'hba58b249),
	.w5(32'h3afeb4f7),
	.w6(32'hbb37d2bc),
	.w7(32'hb9eedd28),
	.w8(32'hbafef69c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9eeda4),
	.w1(32'hba6afa09),
	.w2(32'hb997af06),
	.w3(32'h3b234651),
	.w4(32'h38eb4ee0),
	.w5(32'hb9c5e920),
	.w6(32'h38ada328),
	.w7(32'h3b8766cc),
	.w8(32'h3b82bc20),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8aef2),
	.w1(32'hbad830eb),
	.w2(32'hba649f6e),
	.w3(32'hbb081b5a),
	.w4(32'h3bd63e4b),
	.w5(32'h3c077ccc),
	.w6(32'h3a610b1c),
	.w7(32'hba0076ad),
	.w8(32'hbba73c35),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab19140),
	.w1(32'h3b72e022),
	.w2(32'h3b6bb14c),
	.w3(32'h3b2f5806),
	.w4(32'hba2b548a),
	.w5(32'h3a97bf54),
	.w6(32'hba6443ae),
	.w7(32'hbb67c6e6),
	.w8(32'hbbbcfa1c),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf58500),
	.w1(32'h39573583),
	.w2(32'h3a3a4057),
	.w3(32'h3bd1723c),
	.w4(32'hbada3617),
	.w5(32'hbadda58d),
	.w6(32'hbb29db0a),
	.w7(32'hb88ea2b4),
	.w8(32'h3b15b08d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1085e7),
	.w1(32'h3b109cb3),
	.w2(32'h3b0fad7d),
	.w3(32'hbb7c814f),
	.w4(32'h3b66d82c),
	.w5(32'h3a5e0da0),
	.w6(32'hbb36c8a4),
	.w7(32'h3b6ab121),
	.w8(32'h392a2b38),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baac648),
	.w1(32'h395b3af5),
	.w2(32'h3ad175ff),
	.w3(32'h3ae2ba57),
	.w4(32'hb9ef9516),
	.w5(32'hb98d3e59),
	.w6(32'h3a99e078),
	.w7(32'h3b01cf73),
	.w8(32'hba3c85fb),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89babd),
	.w1(32'h39b0b090),
	.w2(32'h3b00d8f8),
	.w3(32'hbb3bf60f),
	.w4(32'h3a3ed857),
	.w5(32'hba3f0a1a),
	.w6(32'hbabad111),
	.w7(32'hbb227d5d),
	.w8(32'hba1fbeb2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd7a58),
	.w1(32'hbb401fde),
	.w2(32'h39104e24),
	.w3(32'hbbbaa8e5),
	.w4(32'h3ad24927),
	.w5(32'hba3e68ef),
	.w6(32'hba29ca46),
	.w7(32'h3b3c94bb),
	.w8(32'h3abdbeeb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33e94f),
	.w1(32'hbb5bf12a),
	.w2(32'hba953bc0),
	.w3(32'hbb0af067),
	.w4(32'h3c1b5454),
	.w5(32'h3b413853),
	.w6(32'h3b583b43),
	.w7(32'h3b64ea88),
	.w8(32'h391b2e2c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad40a9f),
	.w1(32'hb9e15e6f),
	.w2(32'hbb081332),
	.w3(32'hbb3cfb84),
	.w4(32'h3c1e74e4),
	.w5(32'h3c46c6f7),
	.w6(32'hb997b66d),
	.w7(32'hb9e9bf98),
	.w8(32'hba9c830f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3354d3),
	.w1(32'hbac79a8c),
	.w2(32'hba6a40fc),
	.w3(32'h3bc5eb4b),
	.w4(32'hbb490ca1),
	.w5(32'hb92566b1),
	.w6(32'hbaabea52),
	.w7(32'hbb18927b),
	.w8(32'hbb16738a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4e4f8),
	.w1(32'hba803aa4),
	.w2(32'h3a85f810),
	.w3(32'h3b8fb5dd),
	.w4(32'h3a36ce34),
	.w5(32'h3b137768),
	.w6(32'h3a203e58),
	.w7(32'hbb9aed6d),
	.w8(32'hbbbfa0d1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972ad7b),
	.w1(32'hbad80876),
	.w2(32'h3a407235),
	.w3(32'h3a52b344),
	.w4(32'h3a85b6e9),
	.w5(32'h3b33b430),
	.w6(32'hbb7f1212),
	.w7(32'hbb284b78),
	.w8(32'hbb065bea),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule