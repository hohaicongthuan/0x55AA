module layer_10_featuremap_358(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfad3ac),
	.w1(32'hbc56687a),
	.w2(32'hbc2561b7),
	.w3(32'hbc44b10d),
	.w4(32'hbc1c2794),
	.w5(32'h3b9b9aa4),
	.w6(32'hbbc9fd31),
	.w7(32'hbbd7c991),
	.w8(32'h3add48ad),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab684ea),
	.w1(32'hbbc24844),
	.w2(32'hbbbeb70b),
	.w3(32'h38c1bd7d),
	.w4(32'hbac76560),
	.w5(32'h3c34a46d),
	.w6(32'hbc828a40),
	.w7(32'hbc031a16),
	.w8(32'h3b40e9b4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb386330),
	.w1(32'h3bae510f),
	.w2(32'h3c1d2c1e),
	.w3(32'h3b485dfb),
	.w4(32'hbb465d3b),
	.w5(32'h3b35ca49),
	.w6(32'hbb4ce602),
	.w7(32'h3ba708df),
	.w8(32'h3aa9e7ac),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07e4a1),
	.w1(32'hba984c2c),
	.w2(32'h3b22419f),
	.w3(32'h3b91617b),
	.w4(32'h3ad1e6ea),
	.w5(32'hbbac64b0),
	.w6(32'hbc33ee1f),
	.w7(32'hbae10975),
	.w8(32'h3c466eff),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50c684),
	.w1(32'hbbf0fd24),
	.w2(32'hbc636497),
	.w3(32'hbabda5be),
	.w4(32'hbbfa958a),
	.w5(32'h3b456126),
	.w6(32'h3a9665a6),
	.w7(32'hbb1ff72a),
	.w8(32'hbb1ff86f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25af2d),
	.w1(32'h3b03ecac),
	.w2(32'h39b0926a),
	.w3(32'hbb50712c),
	.w4(32'hbab6a425),
	.w5(32'hbb1bb1d9),
	.w6(32'h3b3cdf7e),
	.w7(32'h3aa773f6),
	.w8(32'hbaa01922),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09b032),
	.w1(32'hbb467cc5),
	.w2(32'hbb604bb0),
	.w3(32'hbb17f555),
	.w4(32'h3aa183ac),
	.w5(32'hbc363fb6),
	.w6(32'hbb044d46),
	.w7(32'h3a4595ca),
	.w8(32'hbbad152e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9526745),
	.w1(32'h3c0a3f4e),
	.w2(32'h3b86994a),
	.w3(32'hbb889c4f),
	.w4(32'h3b766d81),
	.w5(32'hbbedeff2),
	.w6(32'h3bbe742b),
	.w7(32'h3bb5d38e),
	.w8(32'hbbaf9611),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba91bf1),
	.w1(32'h3a0c2ac0),
	.w2(32'hbb8de40d),
	.w3(32'hbbdfe574),
	.w4(32'hbb9c344a),
	.w5(32'h3bec9447),
	.w6(32'h3b4a89b2),
	.w7(32'hbb1fb7f1),
	.w8(32'h3aad63c3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b849fea),
	.w1(32'h3b217e58),
	.w2(32'h3a988083),
	.w3(32'h3b5f0892),
	.w4(32'h3ae4af24),
	.w5(32'hbabaa434),
	.w6(32'h3be9afdd),
	.w7(32'h3b827ff4),
	.w8(32'hbbd69bde),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392229e2),
	.w1(32'h392bb9c2),
	.w2(32'hbb41fbd1),
	.w3(32'hbbf729ec),
	.w4(32'hbad94e0f),
	.w5(32'h3b8e2ec7),
	.w6(32'h3b3a01fb),
	.w7(32'h3a95840c),
	.w8(32'hbac501ab),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc05dcf),
	.w1(32'h3c37f4ec),
	.w2(32'h3c205981),
	.w3(32'h3b667f66),
	.w4(32'hbbbd8297),
	.w5(32'hbc126a71),
	.w6(32'hbb4973e0),
	.w7(32'h3c0d9cec),
	.w8(32'hba5f44f6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fae07),
	.w1(32'h3c332b11),
	.w2(32'h3b9602c7),
	.w3(32'h3b050ce2),
	.w4(32'h3b386c1a),
	.w5(32'hbb98af91),
	.w6(32'h3c914d24),
	.w7(32'h3ad84826),
	.w8(32'hbb5b8f5c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beef000),
	.w1(32'h3a14795e),
	.w2(32'h3b3415e1),
	.w3(32'h3b871d03),
	.w4(32'hb93b413f),
	.w5(32'h3b43eac2),
	.w6(32'hbb3eb062),
	.w7(32'hbb824b29),
	.w8(32'h3c1a8b6f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fe5df),
	.w1(32'h3bdc30fd),
	.w2(32'h3c11ccbe),
	.w3(32'h3c1fda17),
	.w4(32'h3c2dc52d),
	.w5(32'h3b4413b4),
	.w6(32'h3c662717),
	.w7(32'h3c6b6f14),
	.w8(32'hbbc2fb3c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07bcf5),
	.w1(32'hbbc86ee7),
	.w2(32'hbc14e9fa),
	.w3(32'hbbdc7303),
	.w4(32'hbabf8e52),
	.w5(32'hbb6cd9d8),
	.w6(32'hbb96cdec),
	.w7(32'hbb9a8bcb),
	.w8(32'hbc4581ce),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa70b4f),
	.w1(32'h3b9ea668),
	.w2(32'hbb327249),
	.w3(32'hbc0c029c),
	.w4(32'hbaeec563),
	.w5(32'h3b31afa4),
	.w6(32'hbb28e85e),
	.w7(32'h3a93a365),
	.w8(32'h39496eee),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c6937),
	.w1(32'hbb406f8d),
	.w2(32'hbba74f5c),
	.w3(32'hb7ffc7a4),
	.w4(32'hbb8da314),
	.w5(32'h3c5bbfab),
	.w6(32'hbc1e27bb),
	.w7(32'hbbd41ae7),
	.w8(32'h3bdde8b6),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ea91c),
	.w1(32'h3baa6202),
	.w2(32'h3c300489),
	.w3(32'h3c6d287f),
	.w4(32'h3c4bde07),
	.w5(32'hbb5f6357),
	.w6(32'h3c24a8e2),
	.w7(32'h3bfa5aef),
	.w8(32'h3b4e24dc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad50f70),
	.w1(32'h3a81b8ee),
	.w2(32'hbb056a77),
	.w3(32'h3b982213),
	.w4(32'hbb0d6a91),
	.w5(32'h3b8bc01f),
	.w6(32'h3b0865da),
	.w7(32'hbb102361),
	.w8(32'h3a484f14),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6bdbb),
	.w1(32'h3b715fa1),
	.w2(32'hbb9bc9ee),
	.w3(32'hbadd7e9c),
	.w4(32'hbbc88505),
	.w5(32'h3a5291be),
	.w6(32'h3a1faf2b),
	.w7(32'hbb66f13e),
	.w8(32'hb831eedc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f3fa),
	.w1(32'hbba2e69f),
	.w2(32'hba1ea1ae),
	.w3(32'hbb62c515),
	.w4(32'hbba9dcd9),
	.w5(32'h3b34aa86),
	.w6(32'hbc378c47),
	.w7(32'hbb7b205c),
	.w8(32'hb9161008),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b78cb),
	.w1(32'h3797f816),
	.w2(32'h3b821572),
	.w3(32'h3a345888),
	.w4(32'hba2bda33),
	.w5(32'hbbd0cd70),
	.w6(32'hbbc2ad8c),
	.w7(32'h3b09c2b2),
	.w8(32'hb91a73ae),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fdf6a),
	.w1(32'h3ba2cc07),
	.w2(32'hba0ace53),
	.w3(32'h3b86a3bd),
	.w4(32'h3b67381a),
	.w5(32'h3b18c40a),
	.w6(32'h3cb71403),
	.w7(32'hbbc26b53),
	.w8(32'h3b73db23),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9ad86),
	.w1(32'hb9f8b561),
	.w2(32'h3bdc58c7),
	.w3(32'h3a1bc91b),
	.w4(32'h3b047fb5),
	.w5(32'h3b0d9d53),
	.w6(32'h3ad84474),
	.w7(32'h3b07bd92),
	.w8(32'h3baf2d0d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dcb37),
	.w1(32'h3b7db36d),
	.w2(32'h3bee15ae),
	.w3(32'hbb2414fb),
	.w4(32'h3af849ec),
	.w5(32'hbbf36c12),
	.w6(32'h3c154f10),
	.w7(32'h3b0c9da2),
	.w8(32'hbbbf1917),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6dc67),
	.w1(32'h3aba3876),
	.w2(32'h3b7e1023),
	.w3(32'hbbcb1226),
	.w4(32'h39068ce8),
	.w5(32'h3a4ebf7e),
	.w6(32'h3b53c0b2),
	.w7(32'h3b565304),
	.w8(32'hbb389091),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb896834),
	.w1(32'hbbce9a64),
	.w2(32'hbc1ffc44),
	.w3(32'hbba106b8),
	.w4(32'hbc010c58),
	.w5(32'hbb6715cb),
	.w6(32'hbaacffcd),
	.w7(32'hbbb051ee),
	.w8(32'h3b56615d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bace0a3),
	.w1(32'h3bc18efc),
	.w2(32'h3bae073e),
	.w3(32'h3b7a3403),
	.w4(32'h3bc5c31a),
	.w5(32'h3a4b4d97),
	.w6(32'hba04becf),
	.w7(32'h3b4197b7),
	.w8(32'hba2bc5bc),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be797c1),
	.w1(32'hb8efc4ff),
	.w2(32'h3b5ab7d7),
	.w3(32'hba3c265c),
	.w4(32'hbb5e54bb),
	.w5(32'hbc2432c9),
	.w6(32'hbb011097),
	.w7(32'hb9a92102),
	.w8(32'h3ba98935),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf0ac6),
	.w1(32'hbbc3d044),
	.w2(32'hbc11daa6),
	.w3(32'h3ac4c8ca),
	.w4(32'h3ad11bc7),
	.w5(32'h3b743737),
	.w6(32'h3c7bcc37),
	.w7(32'h3a91807c),
	.w8(32'hbbc8462d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0f862),
	.w1(32'h3b47617b),
	.w2(32'hbbb46fb8),
	.w3(32'h3b51f540),
	.w4(32'hbc0593b0),
	.w5(32'hbbcbf6a8),
	.w6(32'hbca330e9),
	.w7(32'hbc8bdbde),
	.w8(32'h3cc50ecb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5497e),
	.w1(32'hbbcf14d4),
	.w2(32'h3a38578a),
	.w3(32'h3c204b48),
	.w4(32'h3b3becb2),
	.w5(32'h3a9a6573),
	.w6(32'h3bca1b06),
	.w7(32'hbbddfcdf),
	.w8(32'hbb8ee3f9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d180c),
	.w1(32'hbbdbc992),
	.w2(32'h3ac627dc),
	.w3(32'hbb1aeda0),
	.w4(32'hbbcdf7d1),
	.w5(32'h3a9ade9d),
	.w6(32'hbc182721),
	.w7(32'hbbae44e4),
	.w8(32'h3baa4530),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0247ad),
	.w1(32'hba3ebc1b),
	.w2(32'h3b1b5e40),
	.w3(32'h3b347655),
	.w4(32'h3af8575f),
	.w5(32'h3a96de39),
	.w6(32'h3c000ee7),
	.w7(32'hbae41bb4),
	.w8(32'hbb9c6c29),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bd1be),
	.w1(32'hbb5df2ba),
	.w2(32'hbb973855),
	.w3(32'hbc2b986f),
	.w4(32'hbc02c781),
	.w5(32'hbaa0cfdd),
	.w6(32'h3c0ad478),
	.w7(32'hbb774421),
	.w8(32'h3b5c93ee),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabd35d),
	.w1(32'h3a98782e),
	.w2(32'h3af363d3),
	.w3(32'h3b4c7792),
	.w4(32'h3b699cb8),
	.w5(32'h3b05b6b7),
	.w6(32'hbbf3bba9),
	.w7(32'hba15cf11),
	.w8(32'hbc15b185),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2f511),
	.w1(32'h3ae8e297),
	.w2(32'hbabb7565),
	.w3(32'hbc1d7b63),
	.w4(32'hbb319933),
	.w5(32'h3aebb629),
	.w6(32'h3a7f1b3a),
	.w7(32'h3b25a0ba),
	.w8(32'h3989be2d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0ac12),
	.w1(32'hbc21ff7e),
	.w2(32'hbb8154ef),
	.w3(32'hbaa56aeb),
	.w4(32'hbb4f8d55),
	.w5(32'h3c309f87),
	.w6(32'hbafe9ede),
	.w7(32'hbb53aeb2),
	.w8(32'hbad55619),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac84b73),
	.w1(32'hbc1e79ff),
	.w2(32'hbbd933c7),
	.w3(32'hbacf8ff1),
	.w4(32'hbb92555e),
	.w5(32'h3bab798e),
	.w6(32'hbb8c5f04),
	.w7(32'hbbccef47),
	.w8(32'hbb158b71),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd78eb),
	.w1(32'hbc0a5f86),
	.w2(32'h3b29d556),
	.w3(32'h3aec002e),
	.w4(32'hba9e40cc),
	.w5(32'hbb53b940),
	.w6(32'hbbb93c12),
	.w7(32'hbb3eb321),
	.w8(32'hbba1bbfc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac80372),
	.w1(32'h3b356ca0),
	.w2(32'hb9718f9f),
	.w3(32'hbbc8e50d),
	.w4(32'hbbd0af0b),
	.w5(32'hbab79a19),
	.w6(32'h3a59c64f),
	.w7(32'h3a33309c),
	.w8(32'hbb85ba21),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0117b2),
	.w1(32'hbae84c09),
	.w2(32'hbb55a49e),
	.w3(32'hba0c9b43),
	.w4(32'h39c6761a),
	.w5(32'h3bb3543d),
	.w6(32'hbbd075e7),
	.w7(32'h3b156c13),
	.w8(32'hbc0363cf),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2e3ac),
	.w1(32'h3c52f3c7),
	.w2(32'hbbdcd78a),
	.w3(32'hbc0b1d5c),
	.w4(32'h3ba3d9c8),
	.w5(32'hba17d3af),
	.w6(32'h3c8908c9),
	.w7(32'h3ba08f59),
	.w8(32'h3bfdb2ce),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cfd13),
	.w1(32'h3c65b738),
	.w2(32'h3cb14883),
	.w3(32'h3c32e656),
	.w4(32'h3c2b4eaf),
	.w5(32'hbbec17e1),
	.w6(32'h3c0c631c),
	.w7(32'h3c88ae8b),
	.w8(32'hbc680734),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b325095),
	.w1(32'h3b939f84),
	.w2(32'h3b7fff8d),
	.w3(32'hbb8b3832),
	.w4(32'h3adde518),
	.w5(32'hba1c5abf),
	.w6(32'h3beba267),
	.w7(32'h3c14b606),
	.w8(32'hbb97e410),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf17b5d),
	.w1(32'h3c8a491c),
	.w2(32'h3c865e91),
	.w3(32'h3c05d095),
	.w4(32'h3be7ab80),
	.w5(32'hbb9ac7a9),
	.w6(32'h3c0ea7b1),
	.w7(32'h3c8722fe),
	.w8(32'hbb3d3aa6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf421b4),
	.w1(32'hbbfb7b6a),
	.w2(32'hbc577e79),
	.w3(32'hbb0c392e),
	.w4(32'hbbc32ea4),
	.w5(32'hbc773f8a),
	.w6(32'hbb6dedb1),
	.w7(32'hbc18d377),
	.w8(32'hbc1f85e9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e7813),
	.w1(32'h3bb6e476),
	.w2(32'hbb00f606),
	.w3(32'hbb5477d7),
	.w4(32'hbb8830ce),
	.w5(32'h39b90fe1),
	.w6(32'h3ca34f30),
	.w7(32'h3bc66816),
	.w8(32'hbaaae22f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dfe0a),
	.w1(32'hbbfe6a59),
	.w2(32'hbb5e860b),
	.w3(32'hbbb039eb),
	.w4(32'hbc1619f9),
	.w5(32'h3af6d6ca),
	.w6(32'hbc7cce7a),
	.w7(32'hbbda2776),
	.w8(32'h3aa15a6c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88434f),
	.w1(32'hba241968),
	.w2(32'hbb88d5fd),
	.w3(32'h3a82f7c5),
	.w4(32'hbba7a062),
	.w5(32'hbbc0efd7),
	.w6(32'h3cc2e6e8),
	.w7(32'hbbf3d2a7),
	.w8(32'hbc6486ed),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14d205),
	.w1(32'hbc602a90),
	.w2(32'hbc09efbc),
	.w3(32'hbbaa8f17),
	.w4(32'hbb8c2dc7),
	.w5(32'h3b5e3932),
	.w6(32'hbc62853f),
	.w7(32'hbc452b3f),
	.w8(32'hbb1e0bcf),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86abb1),
	.w1(32'h3b5eab11),
	.w2(32'h3b88e263),
	.w3(32'h3b08b869),
	.w4(32'h3b145314),
	.w5(32'h3b828a0a),
	.w6(32'h3afff178),
	.w7(32'h3b83e21a),
	.w8(32'hbbb9720a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac14dff),
	.w1(32'hbbc15ef0),
	.w2(32'hbb6f1cc5),
	.w3(32'hbb814f80),
	.w4(32'hbc10a18b),
	.w5(32'hbbd4b159),
	.w6(32'hbc10b055),
	.w7(32'h37d43755),
	.w8(32'hba28812a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8282e),
	.w1(32'h3bb12a5c),
	.w2(32'h3b25f4b5),
	.w3(32'h3b5fe3b3),
	.w4(32'h3ac5761d),
	.w5(32'h3a75566a),
	.w6(32'h3b65d0e5),
	.w7(32'hba78d0eb),
	.w8(32'hba9275c0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f61da9),
	.w1(32'hbb57ba4b),
	.w2(32'h3b11974c),
	.w3(32'h3bbe069c),
	.w4(32'hbabf2bdf),
	.w5(32'hbb02cc7a),
	.w6(32'h3a8d22af),
	.w7(32'h3b135b09),
	.w8(32'hbbc2e8d7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86e615),
	.w1(32'hbb0eb2f9),
	.w2(32'hba9471a6),
	.w3(32'h39db6bf6),
	.w4(32'hbbc1791d),
	.w5(32'hbaa99594),
	.w6(32'h3b2376f2),
	.w7(32'hbab62ba3),
	.w8(32'hbb66885b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a721f),
	.w1(32'hbc0ff44c),
	.w2(32'hbc00019e),
	.w3(32'hbbacf2ec),
	.w4(32'hbb2d6f54),
	.w5(32'hbb9ef591),
	.w6(32'hbbfc4ab4),
	.w7(32'hba9d9efe),
	.w8(32'hbba29ba5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbda32d),
	.w1(32'hbc04e3dd),
	.w2(32'hbb47a0c9),
	.w3(32'hbbfb7b86),
	.w4(32'hbc3b6423),
	.w5(32'h3b46b40c),
	.w6(32'hbc7233e4),
	.w7(32'hbc0d8a5e),
	.w8(32'h3a450bec),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc54d46),
	.w1(32'h3b4077cb),
	.w2(32'hbbc30bcb),
	.w3(32'h3c26555a),
	.w4(32'h3bb2b6b6),
	.w5(32'hba2d9edd),
	.w6(32'h3c347129),
	.w7(32'h3bee2e56),
	.w8(32'hb920a11a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7cf62),
	.w1(32'hbb74f172),
	.w2(32'h3aa58003),
	.w3(32'hbac51978),
	.w4(32'h3afabe9f),
	.w5(32'hba35f503),
	.w6(32'h3a23a709),
	.w7(32'h3ad52e3b),
	.w8(32'hba24c261),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04afa6),
	.w1(32'h3b0cd7ab),
	.w2(32'hbb069d0e),
	.w3(32'hbb822097),
	.w4(32'h3929d058),
	.w5(32'hbc027d1f),
	.w6(32'hbb9e2ea1),
	.w7(32'hba425a90),
	.w8(32'h3bb5c847),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9189b2),
	.w1(32'h3a7a6faf),
	.w2(32'h38db2115),
	.w3(32'hbbc062b2),
	.w4(32'hba719482),
	.w5(32'hbaba70ae),
	.w6(32'h3b8294bf),
	.w7(32'h3b4fc879),
	.w8(32'hba278ef6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1771f6),
	.w1(32'hbb4d80c2),
	.w2(32'h3bebc1f0),
	.w3(32'h3ac91296),
	.w4(32'hbb175a54),
	.w5(32'h3b6175c9),
	.w6(32'h3b961390),
	.w7(32'h3b865805),
	.w8(32'h3bfe3cbf),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b068360),
	.w1(32'h3aff6806),
	.w2(32'h3bb16323),
	.w3(32'h3bbbbfaa),
	.w4(32'h3b533ef6),
	.w5(32'h3ae93c04),
	.w6(32'h3a4e1601),
	.w7(32'h3bd7af07),
	.w8(32'h3ba87003),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb198b56),
	.w1(32'hba0825ed),
	.w2(32'h3b10ce6b),
	.w3(32'h3ab26427),
	.w4(32'h3aabc130),
	.w5(32'hba9fc5fd),
	.w6(32'hba77a430),
	.w7(32'hbb95f079),
	.w8(32'hbaf489af),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e8631),
	.w1(32'h3bb0e9ca),
	.w2(32'hba2b0450),
	.w3(32'hbbd66600),
	.w4(32'h3b9a6b84),
	.w5(32'hbc2a2d09),
	.w6(32'h3c2c9a32),
	.w7(32'h3c6514a9),
	.w8(32'hbbfd0397),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c212753),
	.w1(32'h3c47f25a),
	.w2(32'hb916bacd),
	.w3(32'h3bd51526),
	.w4(32'h3bbbef65),
	.w5(32'hbb954a71),
	.w6(32'h3cf37049),
	.w7(32'h3bd02443),
	.w8(32'h3aea3c75),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a769d63),
	.w1(32'h3b2877f0),
	.w2(32'hbac4bc40),
	.w3(32'h3c0de851),
	.w4(32'hbb9e24e2),
	.w5(32'hba823434),
	.w6(32'h3c2f75e9),
	.w7(32'hbbecc3ac),
	.w8(32'hbc2c92fa),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b886d8b),
	.w1(32'h3c31fa01),
	.w2(32'h3a59181e),
	.w3(32'hbc142641),
	.w4(32'h3ac4aad8),
	.w5(32'hbb375b3f),
	.w6(32'h3c0b4406),
	.w7(32'h3b3b96d5),
	.w8(32'h3c4aaaea),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be05269),
	.w1(32'h3afb4ad0),
	.w2(32'h3c451162),
	.w3(32'h3a958624),
	.w4(32'h3bab37e5),
	.w5(32'hbad5d881),
	.w6(32'h3bf43b43),
	.w7(32'h3ba05925),
	.w8(32'hbc1bdfa4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1f3ca),
	.w1(32'h3c5ccdf0),
	.w2(32'h3a9af022),
	.w3(32'hbb7858c6),
	.w4(32'h3b4ed05a),
	.w5(32'hbabc7530),
	.w6(32'h3c7f25ee),
	.w7(32'h3c853823),
	.w8(32'hbc2aad80),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe5b79),
	.w1(32'h3a9eef02),
	.w2(32'hbc2d1a00),
	.w3(32'hbc3e6bdd),
	.w4(32'h3a540aa5),
	.w5(32'hbbde9e1f),
	.w6(32'h3b74300b),
	.w7(32'h3a360622),
	.w8(32'hbbde76ae),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a0875),
	.w1(32'hbc86a718),
	.w2(32'hbbbf20ad),
	.w3(32'hbc115c96),
	.w4(32'hbc71cdeb),
	.w5(32'hbbaf0f13),
	.w6(32'hbca1e667),
	.w7(32'hbbec863b),
	.w8(32'hbc377df5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9c4f2),
	.w1(32'hbba04333),
	.w2(32'hbac78d8f),
	.w3(32'hbc49bcf6),
	.w4(32'hbb0abbb0),
	.w5(32'hba7611b0),
	.w6(32'h3a9db35f),
	.w7(32'hba473447),
	.w8(32'hba3f6624),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39670047),
	.w1(32'h3bfead76),
	.w2(32'h3a017a33),
	.w3(32'h3c2078f7),
	.w4(32'h3a801612),
	.w5(32'h3b3bcdf8),
	.w6(32'h3c750070),
	.w7(32'h3b887cdb),
	.w8(32'h3ac246c4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd90f3),
	.w1(32'hba9b4548),
	.w2(32'h3b2ddc9b),
	.w3(32'h3b6654f7),
	.w4(32'h3b94983d),
	.w5(32'hbb9b062b),
	.w6(32'hb9d19c7e),
	.w7(32'hba226da6),
	.w8(32'hbc373a6c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e7894),
	.w1(32'hbb321610),
	.w2(32'hb9b29bf0),
	.w3(32'hbb6beffc),
	.w4(32'hba46cee8),
	.w5(32'h3a87e9cb),
	.w6(32'hbc321f5b),
	.w7(32'hbb58bec1),
	.w8(32'h3b981308),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69929e),
	.w1(32'h3c39b3fb),
	.w2(32'h3c16d92f),
	.w3(32'h3c08c7a4),
	.w4(32'h3c849cc7),
	.w5(32'hbb8ae2fa),
	.w6(32'h3c610ea3),
	.w7(32'h3c9f7c11),
	.w8(32'hbbadabe1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6ba9e),
	.w1(32'h3b9ce3f3),
	.w2(32'hbb412335),
	.w3(32'hbc0c0649),
	.w4(32'hbabe1b8e),
	.w5(32'h3baf6215),
	.w6(32'h3c2e3684),
	.w7(32'h3c095e1e),
	.w8(32'h3c93a555),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dee38),
	.w1(32'h3ca853c3),
	.w2(32'h3a666619),
	.w3(32'h3cc9d3ab),
	.w4(32'h3c07348a),
	.w5(32'hbb27e003),
	.w6(32'h3d0fd0f1),
	.w7(32'h3c2cb22e),
	.w8(32'h3b0b55af),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399109ba),
	.w1(32'hbb707a6b),
	.w2(32'hbb534f1b),
	.w3(32'h3a4037aa),
	.w4(32'h3b3bd599),
	.w5(32'hbbbfa450),
	.w6(32'h3b0b6f8b),
	.w7(32'h3be25d38),
	.w8(32'hb9af3abb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c48a6),
	.w1(32'hbb687452),
	.w2(32'h3ac64f68),
	.w3(32'h3a04f0e5),
	.w4(32'h3b372af3),
	.w5(32'hb99f4482),
	.w6(32'h3b74709c),
	.w7(32'hbbc5f5a3),
	.w8(32'hbb945f82),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae709a),
	.w1(32'h3c2019f3),
	.w2(32'hbb4e7fbc),
	.w3(32'h3bf132a8),
	.w4(32'h3b2b3a61),
	.w5(32'hb97058b3),
	.w6(32'h3c98f7d0),
	.w7(32'h3a818385),
	.w8(32'h3c0f2eb3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc62f9),
	.w1(32'hbb58ab66),
	.w2(32'h3ba2ad09),
	.w3(32'h3b443124),
	.w4(32'h3b374a93),
	.w5(32'hbbaaefa1),
	.w6(32'h3a6fec90),
	.w7(32'hbb4e00a9),
	.w8(32'hbc25d9ab),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe7302),
	.w1(32'h3af87f42),
	.w2(32'hbbe0f1a3),
	.w3(32'hbb0ad84d),
	.w4(32'hbb00b3fa),
	.w5(32'hbb5ebedd),
	.w6(32'h3c0d3d59),
	.w7(32'h3a7b5eee),
	.w8(32'hba75e5c1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0755b2),
	.w1(32'h3c1ae525),
	.w2(32'h3bbf29f7),
	.w3(32'hbbc72352),
	.w4(32'hbb12355a),
	.w5(32'h3a7fa463),
	.w6(32'hbc14d62e),
	.w7(32'h3c7023f0),
	.w8(32'h3ba293e0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a29f4),
	.w1(32'h3b1a5841),
	.w2(32'h3ab8b6e0),
	.w3(32'h3b8539ca),
	.w4(32'h3b2e4930),
	.w5(32'hbb845202),
	.w6(32'hb90da024),
	.w7(32'h3a7e0bbc),
	.w8(32'hbbb5bbc2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa52800),
	.w1(32'hbb296a1d),
	.w2(32'hbb73c535),
	.w3(32'hbbdc0299),
	.w4(32'hbb877dac),
	.w5(32'hbb0520c8),
	.w6(32'hbba410ca),
	.w7(32'hbb1360d1),
	.w8(32'hbbd88b7d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba129394),
	.w1(32'h3af3ec03),
	.w2(32'h3aaa6193),
	.w3(32'hbbc05dcc),
	.w4(32'hbc23dd19),
	.w5(32'hbb1c6559),
	.w6(32'h3b72126c),
	.w7(32'hbb83f0a8),
	.w8(32'hbacb548e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f8dfa),
	.w1(32'h3b901b29),
	.w2(32'hbaddae2a),
	.w3(32'hbbc568ef),
	.w4(32'hbb8d53c0),
	.w5(32'h3b15ed1d),
	.w6(32'h3bab1e8f),
	.w7(32'h3918e544),
	.w8(32'h3bad0c83),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ff765),
	.w1(32'hbbb71764),
	.w2(32'hbbbf0563),
	.w3(32'hb999f83b),
	.w4(32'h37f02772),
	.w5(32'h3adc6cae),
	.w6(32'hba81b0fd),
	.w7(32'hbb9319ee),
	.w8(32'hbbc02d88),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf850b0),
	.w1(32'hbbaa3b2e),
	.w2(32'hbbd38a80),
	.w3(32'h3b261493),
	.w4(32'h3bbe5af4),
	.w5(32'h3c05b463),
	.w6(32'hbcc948b9),
	.w7(32'hbaa6d288),
	.w8(32'h38fb76b5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba915282),
	.w1(32'hbb82b56b),
	.w2(32'hbaadf532),
	.w3(32'h3bdac6a2),
	.w4(32'h3aa268ac),
	.w5(32'hbc147824),
	.w6(32'h3b59a4a0),
	.w7(32'hbaeb84c0),
	.w8(32'hbc2aaeb7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb226c05),
	.w1(32'hbbadba54),
	.w2(32'hbbcd479c),
	.w3(32'hbc226b4e),
	.w4(32'hbb2ecc68),
	.w5(32'hbb4a7617),
	.w6(32'h3ad87e6c),
	.w7(32'h3ac8e150),
	.w8(32'hbcaa41bd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcffbf1),
	.w1(32'h3abb99e0),
	.w2(32'h3ab797c9),
	.w3(32'hbbfca246),
	.w4(32'hbb7a106e),
	.w5(32'hbb6844ff),
	.w6(32'hbc0b6c6d),
	.w7(32'hbc2159da),
	.w8(32'hbc059d55),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe39028),
	.w1(32'hbc6cfc0c),
	.w2(32'hbb8672f2),
	.w3(32'h39ca9589),
	.w4(32'h3b033b7a),
	.w5(32'hbc1489ef),
	.w6(32'hbc87f00b),
	.w7(32'hba15963b),
	.w8(32'h3bd138f1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26155b),
	.w1(32'hbb909436),
	.w2(32'h3a995c32),
	.w3(32'h3c54da17),
	.w4(32'h3b32f7f3),
	.w5(32'h3d0a52dc),
	.w6(32'h3cce3e43),
	.w7(32'hbc0acad7),
	.w8(32'h3d3662ab),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d133c6a),
	.w1(32'h3c709066),
	.w2(32'hbb134fc0),
	.w3(32'h3c8f5bf7),
	.w4(32'hbadbd7ee),
	.w5(32'h3c3dcbb8),
	.w6(32'h3d1134c5),
	.w7(32'h3c44a97a),
	.w8(32'h3c91c2c4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3137ae),
	.w1(32'hb98cbfdd),
	.w2(32'h3b9acaf4),
	.w3(32'h3b67ce2f),
	.w4(32'h3c0ec616),
	.w5(32'hbca86134),
	.w6(32'h3c613e32),
	.w7(32'h3bedbb09),
	.w8(32'hbc3a8137),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33b825),
	.w1(32'hba8a6b44),
	.w2(32'hbc5f2b3a),
	.w3(32'hbb9e0a2b),
	.w4(32'hbc93ba19),
	.w5(32'hbbcfab07),
	.w6(32'h3bc39d9a),
	.w7(32'hbb327520),
	.w8(32'hbba5ceb2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b884a36),
	.w1(32'hb917f328),
	.w2(32'h3af73ad9),
	.w3(32'hba89de46),
	.w4(32'h3abf4eff),
	.w5(32'h3b9b7aa5),
	.w6(32'hbb9e90b8),
	.w7(32'hbb10948d),
	.w8(32'h3afea1d6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95e79c),
	.w1(32'h3a58c924),
	.w2(32'hbaca69b0),
	.w3(32'h3bcd4cc6),
	.w4(32'hba5d9e37),
	.w5(32'hbc8137e0),
	.w6(32'h3b494e30),
	.w7(32'hbb3ad607),
	.w8(32'hbc83e6df),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc964641),
	.w1(32'hbbefe06c),
	.w2(32'hbc44630c),
	.w3(32'hbc1a40b2),
	.w4(32'hbc38007a),
	.w5(32'hbbc9a1ac),
	.w6(32'h3b687fd1),
	.w7(32'hbbacbb66),
	.w8(32'hbc0d7200),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cbebd),
	.w1(32'hbc36ce5f),
	.w2(32'hbbeb2f17),
	.w3(32'hbbd5e910),
	.w4(32'hbb8a30b9),
	.w5(32'h3aedf13c),
	.w6(32'hbc3b4069),
	.w7(32'hbc2a98da),
	.w8(32'h3c4f3739),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcebb47),
	.w1(32'h3bea77a1),
	.w2(32'hbb8d81c4),
	.w3(32'h3b3e7007),
	.w4(32'hbb7536c7),
	.w5(32'h3c2e35a8),
	.w6(32'h3c5108a7),
	.w7(32'h3b03e397),
	.w8(32'hbb1305b3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a4bc9),
	.w1(32'hb8e77ee7),
	.w2(32'hbba9cfc4),
	.w3(32'hbb0d5c57),
	.w4(32'hbb9c1f47),
	.w5(32'hbb24e6cb),
	.w6(32'hb9bc3c35),
	.w7(32'h39fb5169),
	.w8(32'hba981290),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94daa9),
	.w1(32'h3b22512b),
	.w2(32'h3bac6441),
	.w3(32'h3abf8f1e),
	.w4(32'h3bbe6db7),
	.w5(32'h3d8de9ce),
	.w6(32'h3ba6e210),
	.w7(32'h3c13e36b),
	.w8(32'h3dae8e08),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d871fb4),
	.w1(32'hba4b55e7),
	.w2(32'h3cef5bc1),
	.w3(32'h3aef893b),
	.w4(32'h3cc915f3),
	.w5(32'hbb2e78da),
	.w6(32'h3d034fc3),
	.w7(32'h3d40020e),
	.w8(32'hbafc8815),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafe837),
	.w1(32'h3bc92311),
	.w2(32'hbb3a3682),
	.w3(32'h3c201a88),
	.w4(32'h398054a5),
	.w5(32'hbc6711e3),
	.w6(32'h3c2ea626),
	.w7(32'hbb3661ac),
	.w8(32'hbc85d6a9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc410010),
	.w1(32'hbc0f04ef),
	.w2(32'hbb247abd),
	.w3(32'hbc77e64d),
	.w4(32'hbc3af8f7),
	.w5(32'hbc226329),
	.w6(32'hbc69f5ad),
	.w7(32'hbc03ce42),
	.w8(32'hbc131b50),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc15615),
	.w1(32'hbaab54dc),
	.w2(32'hbaecde75),
	.w3(32'hbb95a4ea),
	.w4(32'hbbb99632),
	.w5(32'hb9f226fd),
	.w6(32'hbba4b9df),
	.w7(32'hbbb3ab74),
	.w8(32'hbaefc5c8),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27db6d),
	.w1(32'hba0dd152),
	.w2(32'hbb9a28a6),
	.w3(32'h3aaea437),
	.w4(32'hbb70eb5b),
	.w5(32'h3b885d54),
	.w6(32'hbb869288),
	.w7(32'hbc0bfe70),
	.w8(32'hbaa99639),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba04c91),
	.w1(32'hbbda040e),
	.w2(32'hbba88b51),
	.w3(32'hba53e37f),
	.w4(32'h3a9b6ebe),
	.w5(32'hbb829bb7),
	.w6(32'hbb6bee15),
	.w7(32'hbb52bc43),
	.w8(32'h3b2842ec),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00debf),
	.w1(32'hbbd6d6e0),
	.w2(32'hbaea5744),
	.w3(32'h3918b09d),
	.w4(32'h3bc5e6bc),
	.w5(32'hbb582e15),
	.w6(32'hbb346812),
	.w7(32'hb9e54b59),
	.w8(32'hbb89f553),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb401e0c),
	.w1(32'hbb9281f3),
	.w2(32'hbb858531),
	.w3(32'hba8ce367),
	.w4(32'hbb1a863f),
	.w5(32'hbc6b5ee7),
	.w6(32'hbb962278),
	.w7(32'hbbc6756c),
	.w8(32'hbc2a73a2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5441f6),
	.w1(32'hbbbf5db2),
	.w2(32'hbc278fdd),
	.w3(32'hbc154eca),
	.w4(32'hbc4b804f),
	.w5(32'hb8024ac8),
	.w6(32'hbb9d44d5),
	.w7(32'hbc0e02f9),
	.w8(32'h3bfc063d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb55ce5),
	.w1(32'h39e6bcc7),
	.w2(32'h3ba584a6),
	.w3(32'hbc6f1fe1),
	.w4(32'hbc2f3bf2),
	.w5(32'h3d0a06a0),
	.w6(32'hbba96658),
	.w7(32'hb927b154),
	.w8(32'h3d209d64),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd56126),
	.w1(32'h3be8381e),
	.w2(32'h3c154dbb),
	.w3(32'h3c9409e2),
	.w4(32'h3c6bc130),
	.w5(32'h3cdab4a0),
	.w6(32'h3cbd57c5),
	.w7(32'h3c882556),
	.w8(32'h3d0977e8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb159b5),
	.w1(32'h3c5a5461),
	.w2(32'h3c9843b6),
	.w3(32'h3c9c0357),
	.w4(32'h3ca78916),
	.w5(32'hbbcd24c9),
	.w6(32'h3d07cf98),
	.w7(32'h3cf930b7),
	.w8(32'hbbf3ac4b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb03f30),
	.w1(32'hba3dbe63),
	.w2(32'h3afa71ff),
	.w3(32'h3a5e5d71),
	.w4(32'h3b08c9b4),
	.w5(32'hbbb00dec),
	.w6(32'hbacd146e),
	.w7(32'h39d7af0c),
	.w8(32'hbbb542e2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb494ba9),
	.w1(32'hbbbb889d),
	.w2(32'hbb665c6a),
	.w3(32'hbbfec1a9),
	.w4(32'hbb06a505),
	.w5(32'hbb88ffd2),
	.w6(32'hbbfed968),
	.w7(32'hbbb9f63f),
	.w8(32'hbbcf3269),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc05696),
	.w1(32'h3b827e34),
	.w2(32'h3b5030af),
	.w3(32'hbb55b058),
	.w4(32'hbb02edbb),
	.w5(32'h3b5592f5),
	.w6(32'hbbee5158),
	.w7(32'hbb955a56),
	.w8(32'h3837c8a8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9820f9),
	.w1(32'hbab37a37),
	.w2(32'hb91b7ba8),
	.w3(32'h3a97fa4b),
	.w4(32'h3b83fea1),
	.w5(32'h3b5324a3),
	.w6(32'hbab5f6f6),
	.w7(32'h3a91c60c),
	.w8(32'hbaed15db),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b439602),
	.w1(32'h3ba26db3),
	.w2(32'h3b220637),
	.w3(32'h3b8768c4),
	.w4(32'h3b26425c),
	.w5(32'h3a65fa78),
	.w6(32'hb986885f),
	.w7(32'hbaf814b5),
	.w8(32'hba49ac9b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b9357),
	.w1(32'hbadc49ab),
	.w2(32'hb755b17b),
	.w3(32'hbb4312f4),
	.w4(32'h3a8ad4a4),
	.w5(32'hbb794ea3),
	.w6(32'hbbabd5ab),
	.w7(32'hbae141f8),
	.w8(32'hbacb697c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bd253),
	.w1(32'hbb9b9c98),
	.w2(32'hbbde15ab),
	.w3(32'hbb6b8c6b),
	.w4(32'hbb73aae9),
	.w5(32'h3b49a648),
	.w6(32'hbace2d17),
	.w7(32'hbb5386b0),
	.w8(32'h3b4b2597),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b932a03),
	.w1(32'h3b62d0fe),
	.w2(32'h3b901ce2),
	.w3(32'h3bc47be3),
	.w4(32'h3af5e1eb),
	.w5(32'hbc3060ef),
	.w6(32'h3b9e94e9),
	.w7(32'h3a8da02a),
	.w8(32'hbc2ec04b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc633f9),
	.w1(32'h3c5fec4b),
	.w2(32'h3c0eb9d9),
	.w3(32'h3c982959),
	.w4(32'h3c5f061d),
	.w5(32'hbb9de46f),
	.w6(32'h3c7614b9),
	.w7(32'h3c1593d4),
	.w8(32'hbbb80190),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63940a),
	.w1(32'hbb576008),
	.w2(32'hbb5d49ca),
	.w3(32'hbba5237c),
	.w4(32'hbaf861b9),
	.w5(32'hb9aaecec),
	.w6(32'hbbe69c2f),
	.w7(32'hbb9768ad),
	.w8(32'hba892a72),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6988a),
	.w1(32'h3bb1c454),
	.w2(32'h3b08c6ad),
	.w3(32'h3b2bab87),
	.w4(32'hb93ad8ef),
	.w5(32'h3c04ff88),
	.w6(32'h3b19a894),
	.w7(32'hb9857159),
	.w8(32'h3c393c19),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b5324),
	.w1(32'h3b0da35d),
	.w2(32'h3c0c182d),
	.w3(32'h3b1015a9),
	.w4(32'h3be93587),
	.w5(32'h3ba90bad),
	.w6(32'h3c217305),
	.w7(32'h3c5807c0),
	.w8(32'hb8f87873),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61ae0e),
	.w1(32'h3c183ab7),
	.w2(32'h3cc33383),
	.w3(32'h3bd9c1ff),
	.w4(32'h3ccb42c0),
	.w5(32'hbbf53d53),
	.w6(32'h3a94eb35),
	.w7(32'h3c81505a),
	.w8(32'hbb348077),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb135b11),
	.w1(32'hb966b127),
	.w2(32'hba90103f),
	.w3(32'hbb2801ed),
	.w4(32'hbb521211),
	.w5(32'hba382f1e),
	.w6(32'h3b354b65),
	.w7(32'hb82efcec),
	.w8(32'h3b0e8099),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17b999),
	.w1(32'h3b70d279),
	.w2(32'hbb7abbc9),
	.w3(32'h3b9e6645),
	.w4(32'hb950b700),
	.w5(32'hbaba1ce3),
	.w6(32'h3be1325a),
	.w7(32'h3a444cbb),
	.w8(32'h38c5da37),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38f798),
	.w1(32'h3c129ba7),
	.w2(32'hbade1522),
	.w3(32'h3bab978e),
	.w4(32'hbc0acbc6),
	.w5(32'hbb49954a),
	.w6(32'h3bc435c2),
	.w7(32'hbbc2c858),
	.w8(32'h395307ee),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad699ac),
	.w1(32'h3bf74a45),
	.w2(32'h39057ab8),
	.w3(32'h3bd4cf8f),
	.w4(32'hba131f07),
	.w5(32'hbc2f95d0),
	.w6(32'h3c1d7987),
	.w7(32'h395c098b),
	.w8(32'hbb8eb373),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2233bd),
	.w1(32'hbab115db),
	.w2(32'hbb53c3ee),
	.w3(32'hbb7d0173),
	.w4(32'hbb4c1985),
	.w5(32'hba09818c),
	.w6(32'h3b180196),
	.w7(32'hb9fee373),
	.w8(32'hbae1a8a6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49446a),
	.w1(32'hbac470ef),
	.w2(32'hbb06100a),
	.w3(32'h3a5d6cc9),
	.w4(32'hb92e4025),
	.w5(32'h3c058734),
	.w6(32'h3b578d68),
	.w7(32'hb8825f94),
	.w8(32'h39bb335e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51f14f),
	.w1(32'hbb6f3541),
	.w2(32'hbb6b2db2),
	.w3(32'h39a08989),
	.w4(32'hba8b70de),
	.w5(32'hb9fdb7e2),
	.w6(32'hbaf62f8a),
	.w7(32'hba842862),
	.w8(32'hbbe361e0),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf1fd0),
	.w1(32'h3bfa4639),
	.w2(32'h3c154a7c),
	.w3(32'h3bd51274),
	.w4(32'h3c443209),
	.w5(32'h3bcb8be2),
	.w6(32'h3ab07f71),
	.w7(32'h3af33bb5),
	.w8(32'h3bbc5db5),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c441d20),
	.w1(32'h3c2c0930),
	.w2(32'h3bc31558),
	.w3(32'h3bd0b3fa),
	.w4(32'h3bccb3b7),
	.w5(32'h3b53ed73),
	.w6(32'h3ba6eb11),
	.w7(32'h3b9898dd),
	.w8(32'h3b78ef45),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad93b91),
	.w1(32'h3aea50ec),
	.w2(32'h3bc9be27),
	.w3(32'h3b2c871b),
	.w4(32'h3a8c3ec6),
	.w5(32'hbb296127),
	.w6(32'h3b79de10),
	.w7(32'h3ba94df1),
	.w8(32'hbbaa75e8),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affe592),
	.w1(32'hbace871c),
	.w2(32'hba4cacea),
	.w3(32'hbafcd66b),
	.w4(32'hbacd5dd9),
	.w5(32'h3b55e9c4),
	.w6(32'hbbb2b819),
	.w7(32'hbb850d89),
	.w8(32'h3ac2491d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bca7e),
	.w1(32'hbb98dd81),
	.w2(32'hbbb89cf4),
	.w3(32'h3ba1e168),
	.w4(32'h3b2da0c7),
	.w5(32'hbc038b80),
	.w6(32'h3b009c4d),
	.w7(32'hbaa69197),
	.w8(32'hbb9c6dfd),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02f5a6),
	.w1(32'hbbe4750d),
	.w2(32'hbc450ead),
	.w3(32'hbc01084c),
	.w4(32'hbc35efe8),
	.w5(32'h3be3b618),
	.w6(32'hbac5a415),
	.w7(32'hbc256098),
	.w8(32'h3c31d3ff),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51fc15),
	.w1(32'h3c089c15),
	.w2(32'h3c1e9771),
	.w3(32'h3bbec66f),
	.w4(32'h3bd54679),
	.w5(32'hbb87521b),
	.w6(32'h3c7d81e4),
	.w7(32'h3c42a365),
	.w8(32'hbb8a7cb0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf9cf8),
	.w1(32'hbb5926ac),
	.w2(32'hbb9dd738),
	.w3(32'hbbcbad85),
	.w4(32'hbb5e4cb1),
	.w5(32'hbb868d3b),
	.w6(32'hbbdf9e03),
	.w7(32'hbbd2e4f1),
	.w8(32'hbb715f2f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c6d02),
	.w1(32'hba3aa8e1),
	.w2(32'hbb0f9d12),
	.w3(32'hbb7d2425),
	.w4(32'hbb59e74a),
	.w5(32'hbc45d9c0),
	.w6(32'hbb82295c),
	.w7(32'hbb78772e),
	.w8(32'hbbb3dd6b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cb198),
	.w1(32'hbbb81d68),
	.w2(32'hbc4b80b2),
	.w3(32'hbbab0af3),
	.w4(32'hbc469e4c),
	.w5(32'h3bce41c5),
	.w6(32'h3b758d22),
	.w7(32'hbbb30c58),
	.w8(32'hbae170fd),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe4c58),
	.w1(32'hbc3247f3),
	.w2(32'hbc240647),
	.w3(32'hbb661b5e),
	.w4(32'hbad0350f),
	.w5(32'hbbd5894b),
	.w6(32'hbc247d78),
	.w7(32'hbbe926b7),
	.w8(32'hbbc2448d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4517ec),
	.w1(32'hbb633a54),
	.w2(32'hbaa40430),
	.w3(32'hbc077ed1),
	.w4(32'hbbc11263),
	.w5(32'hbbc3a7e5),
	.w6(32'hbbfb3c10),
	.w7(32'hbc0848e5),
	.w8(32'hbc1a58a8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb582b90),
	.w1(32'hbc3332f1),
	.w2(32'hbc45f62e),
	.w3(32'h3a209114),
	.w4(32'h38c53df4),
	.w5(32'hbc07825c),
	.w6(32'hbc12b54f),
	.w7(32'hbc06494e),
	.w8(32'hbbd7b01d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f2677),
	.w1(32'hbbc21219),
	.w2(32'hbb20183f),
	.w3(32'hbbaadf67),
	.w4(32'hbbcfb2ac),
	.w5(32'h3ce745c7),
	.w6(32'hbb336948),
	.w7(32'hbab50b76),
	.w8(32'h3cfdf492),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd77373),
	.w1(32'hbb0d7759),
	.w2(32'h3ccc6b3a),
	.w3(32'h38fe535e),
	.w4(32'h3caadcfd),
	.w5(32'hba9e0409),
	.w6(32'h3b84f4e0),
	.w7(32'h3ceec164),
	.w8(32'h3a756c55),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46e7ae),
	.w1(32'h3c8083e2),
	.w2(32'hbb752d7f),
	.w3(32'h3c9971e6),
	.w4(32'h3a435da8),
	.w5(32'hbc1359f2),
	.w6(32'h3c968592),
	.w7(32'hbb5f6a99),
	.w8(32'hbc0d145c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb549b60),
	.w1(32'hbb7098ca),
	.w2(32'hbbe8c4f5),
	.w3(32'hbb94e671),
	.w4(32'hbc1191f5),
	.w5(32'h39dbc97a),
	.w6(32'hbbb2b8ea),
	.w7(32'hbba3e38a),
	.w8(32'h3b229d46),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accac85),
	.w1(32'h3b8a5495),
	.w2(32'h3bb3e176),
	.w3(32'h3b096535),
	.w4(32'h3ba6748f),
	.w5(32'hbc055e52),
	.w6(32'h3adfd90e),
	.w7(32'h3ba2b130),
	.w8(32'hbbc385e2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e9951),
	.w1(32'h3b5726d5),
	.w2(32'h3b853f26),
	.w3(32'hbbbdeec7),
	.w4(32'hbc1545cf),
	.w5(32'h3b5407a2),
	.w6(32'hbc0a0175),
	.w7(32'hbc09cdac),
	.w8(32'hbbc9f447),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fad96),
	.w1(32'hbc351f87),
	.w2(32'hbc17249c),
	.w3(32'h3b8536bf),
	.w4(32'h3c2dc5d0),
	.w5(32'hbbca4f61),
	.w6(32'hbc32198c),
	.w7(32'hbba211b4),
	.w8(32'hba4593ff),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebf75e),
	.w1(32'h3c12b02a),
	.w2(32'h3c223711),
	.w3(32'h3baa52f2),
	.w4(32'h3b3b57c6),
	.w5(32'h3a394bfe),
	.w6(32'h3be78c71),
	.w7(32'h3bb09548),
	.w8(32'hba6acf35),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb958e36),
	.w1(32'hbb7c7f2f),
	.w2(32'hbc326aaf),
	.w3(32'h39c63afd),
	.w4(32'hbb95cf3d),
	.w5(32'hbb77f40d),
	.w6(32'h3ba62a59),
	.w7(32'hbb27abda),
	.w8(32'hbb801f63),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ef549),
	.w1(32'hbbd8256e),
	.w2(32'hbbf8eac2),
	.w3(32'hbbfa56bb),
	.w4(32'hbbdf13be),
	.w5(32'h3b248281),
	.w6(32'hbc05b8b9),
	.w7(32'hbbf22b74),
	.w8(32'h3b9254cb),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb998970),
	.w1(32'hbc29e17d),
	.w2(32'hbc3c086d),
	.w3(32'hbb6e39e3),
	.w4(32'hbbb65e80),
	.w5(32'hbbead8a7),
	.w6(32'h394b7fa7),
	.w7(32'hbbe55950),
	.w8(32'hbb6b5c0c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff47d1),
	.w1(32'hbb2ac4f1),
	.w2(32'hbb10d154),
	.w3(32'hbbddb7fd),
	.w4(32'hbbfeea6f),
	.w5(32'hbc683897),
	.w6(32'hbbed6b60),
	.w7(32'hbbd17539),
	.w8(32'hbbe583de),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ae542),
	.w1(32'h3bdc79a5),
	.w2(32'hbaa7fd28),
	.w3(32'hbb736df9),
	.w4(32'hbc21c160),
	.w5(32'h3b59b77d),
	.w6(32'h3b7d9f5d),
	.w7(32'hbb9da03b),
	.w8(32'hbb82e65a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac192dc),
	.w1(32'hbb096e05),
	.w2(32'hbb412534),
	.w3(32'h3bb32e93),
	.w4(32'h3baa8690),
	.w5(32'hbb9815ae),
	.w6(32'hbb4c331f),
	.w7(32'hbb4a9cc0),
	.w8(32'h3af167bd),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdf4ae),
	.w1(32'hbb723b05),
	.w2(32'hbcd7160c),
	.w3(32'hba7ba58b),
	.w4(32'hbcbcc3e7),
	.w5(32'hbb513c78),
	.w6(32'h3c64b4e5),
	.w7(32'hbc6b991f),
	.w8(32'hbbfb2ab4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a9dc8),
	.w1(32'hbb81dcb9),
	.w2(32'hbaf99b70),
	.w3(32'hbb4394f6),
	.w4(32'hbb3a9f35),
	.w5(32'hbb358c08),
	.w6(32'hbaff9e17),
	.w7(32'hbb0f4631),
	.w8(32'h3b1b8ab0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc885ac),
	.w1(32'hbb5baba3),
	.w2(32'hbb91e6b9),
	.w3(32'h3afcb634),
	.w4(32'hbb5a241d),
	.w5(32'h398e5ec0),
	.w6(32'h3bee0710),
	.w7(32'h3b3a8c5c),
	.w8(32'h3b360d86),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2056e9),
	.w1(32'h3be411bd),
	.w2(32'h3c083e7b),
	.w3(32'hb9ee0049),
	.w4(32'h39bdcaf4),
	.w5(32'hbbdd834c),
	.w6(32'h3bae3c7f),
	.w7(32'h3b69a200),
	.w8(32'hbc33b3e7),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09e1b4),
	.w1(32'hbc93ee28),
	.w2(32'hbbbfeafa),
	.w3(32'hbc81cbae),
	.w4(32'hbc10ff6d),
	.w5(32'hbbeece23),
	.w6(32'hbc9d4f07),
	.w7(32'hbc1b6a08),
	.w8(32'h3bed58dc),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf02a5),
	.w1(32'hba5b9f4a),
	.w2(32'hbc108d51),
	.w3(32'h3a4fc98f),
	.w4(32'hbc375a46),
	.w5(32'hbc4b73f0),
	.w6(32'h3ca178b0),
	.w7(32'h3bdec4f5),
	.w8(32'hbc46038b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a160e),
	.w1(32'hbbc943c8),
	.w2(32'hbc4fbf8b),
	.w3(32'hbb87fc48),
	.w4(32'hbc25a323),
	.w5(32'h3c91ed92),
	.w6(32'hbae94cb7),
	.w7(32'hbbf5e9cc),
	.w8(32'h3ca15668),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c606009),
	.w1(32'h3bd764d6),
	.w2(32'h3be00ef8),
	.w3(32'h3bef4c80),
	.w4(32'h3bff494a),
	.w5(32'hbc85aca4),
	.w6(32'h3c993711),
	.w7(32'h3c967cac),
	.w8(32'hbc72a30d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d3e36),
	.w1(32'hbb963c29),
	.w2(32'hba00bfee),
	.w3(32'hbbc75b56),
	.w4(32'hbaaf3f9c),
	.w5(32'h3bd02885),
	.w6(32'hbbe0c13a),
	.w7(32'hbae940fa),
	.w8(32'h3bb9be3f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d202e),
	.w1(32'h3c3c38fa),
	.w2(32'h3c259de8),
	.w3(32'h3c2cf695),
	.w4(32'h3befdc60),
	.w5(32'hbba2dd89),
	.w6(32'h3c0d8bfb),
	.w7(32'h3ba451bb),
	.w8(32'hb83e27fb),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5c924),
	.w1(32'h3b7e6421),
	.w2(32'hbb814cf7),
	.w3(32'h3bb27833),
	.w4(32'hbb8df39a),
	.w5(32'h3b4ff366),
	.w6(32'h3c254010),
	.w7(32'h3b108cff),
	.w8(32'h3bba28b9),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c2d7c),
	.w1(32'h3be35697),
	.w2(32'hbb8d28c5),
	.w3(32'h3a971137),
	.w4(32'hbb538c4a),
	.w5(32'hb7e1616d),
	.w6(32'h3bb1d4b3),
	.w7(32'hbbaae916),
	.w8(32'h3b9857b9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5e272),
	.w1(32'hba8bcded),
	.w2(32'h3b92d5d6),
	.w3(32'hbbb69c6c),
	.w4(32'hbb759055),
	.w5(32'hb9dcf97c),
	.w6(32'h39cf5c87),
	.w7(32'hb973501e),
	.w8(32'hbc2a1d47),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc510349),
	.w1(32'hbc1fbcfb),
	.w2(32'hbc741c23),
	.w3(32'hbb031c22),
	.w4(32'hbc11e03a),
	.w5(32'h3bc6868c),
	.w6(32'hbbdfe9c1),
	.w7(32'hbc57e4c9),
	.w8(32'h3b17c5f1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf98022),
	.w1(32'h3af591d2),
	.w2(32'hba810cdb),
	.w3(32'h3b3428c0),
	.w4(32'hbb5be665),
	.w5(32'hbc01c634),
	.w6(32'hbb33e01b),
	.w7(32'hbb31f0c7),
	.w8(32'hbbcb0cb4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3932eb),
	.w1(32'hbbe73402),
	.w2(32'hbbabbb16),
	.w3(32'hbbf1d428),
	.w4(32'hbb38f5ec),
	.w5(32'hbb6d1d65),
	.w6(32'hbbff28dc),
	.w7(32'hbb9de903),
	.w8(32'hbae8d46b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e8541),
	.w1(32'h3c181d49),
	.w2(32'hbb0fe62a),
	.w3(32'h3b992a2f),
	.w4(32'hbb5fa0cf),
	.w5(32'hba7dda83),
	.w6(32'h3ba3e097),
	.w7(32'hbb86c504),
	.w8(32'hbaba51d9),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0579dd),
	.w1(32'hba9abe7d),
	.w2(32'hb9fda20c),
	.w3(32'hbb160423),
	.w4(32'hb9dc05d8),
	.w5(32'hba160cb2),
	.w6(32'hbaa0beab),
	.w7(32'hb728d01a),
	.w8(32'hbb61bf51),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34577c),
	.w1(32'h3baa9500),
	.w2(32'hbc132a20),
	.w3(32'h3b9a41be),
	.w4(32'hbc07b8d2),
	.w5(32'hbb7c914e),
	.w6(32'h3b2184d0),
	.w7(32'hbbdc5e06),
	.w8(32'hb9e212e9),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc046a23),
	.w1(32'h3b2e581b),
	.w2(32'hbb9fc5fc),
	.w3(32'h3be5fe76),
	.w4(32'hbb4d3095),
	.w5(32'hbca806d7),
	.w6(32'h3c0c6233),
	.w7(32'h3a63b985),
	.w8(32'hbc4ef3be),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c3ddd),
	.w1(32'hb9ba2456),
	.w2(32'hbc10a416),
	.w3(32'hbc2c1d4f),
	.w4(32'hbc727ca0),
	.w5(32'h3a42bf32),
	.w6(32'hb9b3d106),
	.w7(32'hbc0d8677),
	.w8(32'hbb24560b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9f311),
	.w1(32'hbb738425),
	.w2(32'hb9c4cc95),
	.w3(32'h3af33aa9),
	.w4(32'h3ac12a47),
	.w5(32'hbbffe97e),
	.w6(32'hbb6c2427),
	.w7(32'hbad887be),
	.w8(32'hbc275bf5),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bedec),
	.w1(32'hbbe4d3df),
	.w2(32'hbbe6ed8a),
	.w3(32'hbb777812),
	.w4(32'hbb593e50),
	.w5(32'h3aab8626),
	.w6(32'hbbd9f937),
	.w7(32'hbb878235),
	.w8(32'hbba8b10e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc4669),
	.w1(32'h3a95ea4d),
	.w2(32'h3b27e55f),
	.w3(32'h3bd27b94),
	.w4(32'h3c3cdb7e),
	.w5(32'h3b37a0c3),
	.w6(32'hbba486c7),
	.w7(32'hb8f2ca87),
	.w8(32'hba8b97e9),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cee64b),
	.w1(32'h3ab9f90b),
	.w2(32'hbb51a563),
	.w3(32'h3b476488),
	.w4(32'hbb0c37f1),
	.w5(32'hbb9d6f3b),
	.w6(32'h3addba86),
	.w7(32'hbb48af48),
	.w8(32'hbb8aa5f2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8ae5f),
	.w1(32'h3b39e66e),
	.w2(32'h3a79f85c),
	.w3(32'h3b8ab081),
	.w4(32'h3b17e167),
	.w5(32'hbbb088a6),
	.w6(32'h3b054bf5),
	.w7(32'h3a50f2f1),
	.w8(32'hbc3a7ad7),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb02c2c),
	.w1(32'hbb9b9a14),
	.w2(32'hbbc5ec7b),
	.w3(32'hbbecfb02),
	.w4(32'hbb6c5008),
	.w5(32'h3b6a8818),
	.w6(32'hbc2b6317),
	.w7(32'hbc233fbb),
	.w8(32'hba92d224),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb006473),
	.w1(32'hbc0f59af),
	.w2(32'hbbdf18e5),
	.w3(32'hbaded580),
	.w4(32'hbb8256de),
	.w5(32'h3cb8b83c),
	.w6(32'hbbf10e17),
	.w7(32'hbbd6564f),
	.w8(32'h3cb350a7),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce24069),
	.w1(32'hbc7396af),
	.w2(32'h3c881d7f),
	.w3(32'hbca26826),
	.w4(32'h3c0e1fd6),
	.w5(32'h3b712569),
	.w6(32'hbc955157),
	.w7(32'h3c198d0b),
	.w8(32'h3bf1fed0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55f0ae),
	.w1(32'h3b8592cf),
	.w2(32'hbb903fb4),
	.w3(32'h3a937825),
	.w4(32'hbb9e871f),
	.w5(32'h3c1fc490),
	.w6(32'h3b5bdecb),
	.w7(32'hbbcb2821),
	.w8(32'h3c99d74b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81335a),
	.w1(32'hbb692ce1),
	.w2(32'h3b736a89),
	.w3(32'hbbf890cf),
	.w4(32'hbb81f6a3),
	.w5(32'hba922d50),
	.w6(32'h3c0a1022),
	.w7(32'h3c00da2c),
	.w8(32'h3ada1b40),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b8b0a),
	.w1(32'h3b95fce7),
	.w2(32'h3c1ecf75),
	.w3(32'hb98dc262),
	.w4(32'h3abc3a84),
	.w5(32'hbaf29ccb),
	.w6(32'h3bb60321),
	.w7(32'h3c1569e4),
	.w8(32'hbbb4cdfa),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa3bd2),
	.w1(32'hbb60786c),
	.w2(32'h3b480c94),
	.w3(32'hba21e8db),
	.w4(32'h3a0ec2d1),
	.w5(32'h3ad9939b),
	.w6(32'hbb737c6e),
	.w7(32'h39fedfee),
	.w8(32'hbb78127c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0198c),
	.w1(32'hbb83e6bc),
	.w2(32'hbbadb5e7),
	.w3(32'h3a41f3aa),
	.w4(32'h3a6eef48),
	.w5(32'hbbc9f386),
	.w6(32'hbb2fcbae),
	.w7(32'hbba108e2),
	.w8(32'hbc30e756),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13a443),
	.w1(32'hbbac9ec0),
	.w2(32'hbbfc8a54),
	.w3(32'hbab59712),
	.w4(32'hbb9cbcaf),
	.w5(32'h3b995268),
	.w6(32'hbb8f1d5b),
	.w7(32'hbb702be9),
	.w8(32'hbb36b7a4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac5d24),
	.w1(32'hbc2979a0),
	.w2(32'hbbfa9094),
	.w3(32'h3b267a28),
	.w4(32'h3b7f0d11),
	.w5(32'hbc103034),
	.w6(32'hbbc5c781),
	.w7(32'hbb94dadf),
	.w8(32'hbc81843c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15b09c),
	.w1(32'hbbaf26b8),
	.w2(32'hbba36a91),
	.w3(32'hbae32760),
	.w4(32'h3a38c6a1),
	.w5(32'hbae1a717),
	.w6(32'hbbb94323),
	.w7(32'hbc1c11db),
	.w8(32'hbbae0ac7),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1efd2b),
	.w1(32'h3b87aa47),
	.w2(32'hba27ff47),
	.w3(32'h3a4b028a),
	.w4(32'hbb7630db),
	.w5(32'h3b27196a),
	.w6(32'hbab63b8d),
	.w7(32'hbba479d3),
	.w8(32'h3c1c49e1),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a6957),
	.w1(32'h3b7faa7b),
	.w2(32'hbab4987f),
	.w3(32'h3ace44a0),
	.w4(32'hbb0bc1bf),
	.w5(32'h3c25dd38),
	.w6(32'h3c627156),
	.w7(32'h3bd9815a),
	.w8(32'h3bf79939),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d11ef),
	.w1(32'h3b7d85d1),
	.w2(32'h3b5ef781),
	.w3(32'h3b1cdeba),
	.w4(32'h3a628d56),
	.w5(32'h3bd0d4ba),
	.w6(32'h3be2b5f9),
	.w7(32'h3b606791),
	.w8(32'h3c2220ad),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ba50b),
	.w1(32'h3beda5dd),
	.w2(32'h3bcf864f),
	.w3(32'h3bc62006),
	.w4(32'h3bb3855f),
	.w5(32'hbcaa7d9d),
	.w6(32'h3c13829e),
	.w7(32'h3bec9d40),
	.w8(32'hbcdad646),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5ef8e),
	.w1(32'hbc6b6e17),
	.w2(32'hbbe5353c),
	.w3(32'hbc885ba5),
	.w4(32'hbc3a38eb),
	.w5(32'hbac77ed8),
	.w6(32'hbca6bfab),
	.w7(32'hbc411b1a),
	.w8(32'hbb14cb25),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90091e),
	.w1(32'hbb5fb207),
	.w2(32'hbbfa2262),
	.w3(32'h3b9fbee5),
	.w4(32'hbadec15d),
	.w5(32'hbb1697ca),
	.w6(32'h3b73e63b),
	.w7(32'hbb75fc6f),
	.w8(32'hbae955d5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b6598),
	.w1(32'h3b866368),
	.w2(32'h3ad15dae),
	.w3(32'h3b92e66f),
	.w4(32'h3a342b7f),
	.w5(32'h3d5b44a4),
	.w6(32'h3b2a58c3),
	.w7(32'hb9f2cedb),
	.w8(32'h3d584475),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d405b71),
	.w1(32'hbc5362a1),
	.w2(32'h3d21b20b),
	.w3(32'h3a356076),
	.w4(32'h3d2ff2d8),
	.w5(32'h3a8f1713),
	.w6(32'h3b9b8a30),
	.w7(32'h3d360982),
	.w8(32'hbb17a455),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad8131),
	.w1(32'hbb688279),
	.w2(32'hba824e3b),
	.w3(32'h3b8a6800),
	.w4(32'h3ba5cade),
	.w5(32'hbc419843),
	.w6(32'hbb17533e),
	.w7(32'hb9c73e0a),
	.w8(32'hbc525dfe),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc068256),
	.w1(32'h3985a59b),
	.w2(32'h3b845a2e),
	.w3(32'hb988bb0c),
	.w4(32'h3b2f6477),
	.w5(32'h3b649457),
	.w6(32'hbb0233e0),
	.w7(32'h3b4974c1),
	.w8(32'hbb1fe28d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab82586),
	.w1(32'h3b0db77f),
	.w2(32'hbbf67d67),
	.w3(32'h3b8e6821),
	.w4(32'hbbe03df3),
	.w5(32'hbb0f3e32),
	.w6(32'h3a55ab56),
	.w7(32'hbb818527),
	.w8(32'hbacc3ab3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32b4f4),
	.w1(32'h3b0748cc),
	.w2(32'hb7c3c40f),
	.w3(32'h3a8d9ece),
	.w4(32'h3a1e9b72),
	.w5(32'h3a41fa80),
	.w6(32'hbad2543b),
	.w7(32'hbb44d7d8),
	.w8(32'h3ba0132a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c0681),
	.w1(32'h3bc70acb),
	.w2(32'h3b909654),
	.w3(32'h3b9f47c8),
	.w4(32'h3b74fede),
	.w5(32'hbbe45e67),
	.w6(32'h3c10ed56),
	.w7(32'h3bcf77cd),
	.w8(32'hbbb27a45),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9071de),
	.w1(32'hbbd1dd60),
	.w2(32'hbb3123f4),
	.w3(32'hbbe8692a),
	.w4(32'hbb913c6d),
	.w5(32'hbbe084a5),
	.w6(32'hbbd6aa26),
	.w7(32'hbb895b29),
	.w8(32'hbbb3c6ba),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52884b),
	.w1(32'hbaf1d50e),
	.w2(32'hbacad3d8),
	.w3(32'hbbee5bd6),
	.w4(32'h3a52452d),
	.w5(32'h3a871f0c),
	.w6(32'hbbd24a61),
	.w7(32'hbb5f87a1),
	.w8(32'h3b2102d4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e295c3),
	.w1(32'hbad748d5),
	.w2(32'hbb046df9),
	.w3(32'h3b738f0e),
	.w4(32'hb9bb7549),
	.w5(32'hbb85eaf2),
	.w6(32'h3b0919c2),
	.w7(32'hba5dea3d),
	.w8(32'hbc0ea150),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a6625),
	.w1(32'hbb3ffa89),
	.w2(32'hbb27d603),
	.w3(32'h3bcf1f7e),
	.w4(32'h3c19b288),
	.w5(32'hbab6aa92),
	.w6(32'hbc1548e9),
	.w7(32'hbb8847ab),
	.w8(32'hbc1b68b1),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc825681),
	.w1(32'hbc870429),
	.w2(32'hbcc0995b),
	.w3(32'h3a878094),
	.w4(32'hbbad59c8),
	.w5(32'hbc7934a8),
	.w6(32'hbbe8f9e7),
	.w7(32'hbc8a9836),
	.w8(32'hbc583a90),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b8842),
	.w1(32'hbb8028f4),
	.w2(32'hbbf1991f),
	.w3(32'hbc092b44),
	.w4(32'hbc53c809),
	.w5(32'h3b34b485),
	.w6(32'hbbd80c88),
	.w7(32'hbc247005),
	.w8(32'h3a15da2e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35c7de),
	.w1(32'h3b14473e),
	.w2(32'hbacb51a3),
	.w3(32'h3b10e297),
	.w4(32'h3a50b3f2),
	.w5(32'hbc462cd4),
	.w6(32'hb90528e9),
	.w7(32'hbba0859d),
	.w8(32'hbc5f79f5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39ac0c),
	.w1(32'hbba3a6e4),
	.w2(32'hbc34fb48),
	.w3(32'hbbadc236),
	.w4(32'hbc0e103c),
	.w5(32'hbc96d723),
	.w6(32'hba19f8ce),
	.w7(32'hbc11e5d3),
	.w8(32'hbc49ac8d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf60845),
	.w1(32'h3be7f472),
	.w2(32'h3bc44dad),
	.w3(32'hbc01f8e3),
	.w4(32'hbbdbfc1a),
	.w5(32'hbbf36968),
	.w6(32'hb9d56e44),
	.w7(32'h3af73456),
	.w8(32'hbc9cad3d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86bc60),
	.w1(32'hbc801a98),
	.w2(32'hbae9e6ab),
	.w3(32'hb935def7),
	.w4(32'h3be0fbdf),
	.w5(32'hbc2af68b),
	.w6(32'hbc817f52),
	.w7(32'h3c33682f),
	.w8(32'hbcbea689),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fd29b),
	.w1(32'hbc046b33),
	.w2(32'hbb8c5811),
	.w3(32'h3c67647d),
	.w4(32'h3be35aac),
	.w5(32'hbb9d8c86),
	.w6(32'h3b19cf6c),
	.w7(32'h3c11f969),
	.w8(32'hbd1aa6b6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce4c304),
	.w1(32'hbd0487cf),
	.w2(32'h3bd06d8a),
	.w3(32'h3c9aff3c),
	.w4(32'h3cf0d239),
	.w5(32'h3bd53f9f),
	.w6(32'hbc3f8ab0),
	.w7(32'h3ccfe237),
	.w8(32'h3bb6b2f5),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9eb59),
	.w1(32'h3b42a2c8),
	.w2(32'h3b82d71b),
	.w3(32'h3b48a76e),
	.w4(32'h3b3ef934),
	.w5(32'h3b06094c),
	.w6(32'h3c295415),
	.w7(32'h3ac2acc3),
	.w8(32'hbb1db4b1),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb495126),
	.w1(32'hbbfc0628),
	.w2(32'hbb113a10),
	.w3(32'h3b850e55),
	.w4(32'h3b5253df),
	.w5(32'hbba5f1de),
	.w6(32'hb93adce7),
	.w7(32'hbb2a9661),
	.w8(32'hbd64be3d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1e37cd),
	.w1(32'hbd0a0b53),
	.w2(32'h3cd8ac60),
	.w3(32'h3d293f31),
	.w4(32'h3d71d9e2),
	.w5(32'hbb7b10f8),
	.w6(32'hbcec8f80),
	.w7(32'h3d85026e),
	.w8(32'hbc263a43),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e86cf),
	.w1(32'h3ad22f38),
	.w2(32'hba2e177c),
	.w3(32'h3bf55947),
	.w4(32'hba906865),
	.w5(32'hba818357),
	.w6(32'hbb829371),
	.w7(32'h3c33daab),
	.w8(32'hbc667752),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2afae6),
	.w1(32'hbc020946),
	.w2(32'h3b66411b),
	.w3(32'h3bd3ebe3),
	.w4(32'h3c413487),
	.w5(32'hbb5f560f),
	.w6(32'hbb12583e),
	.w7(32'h3c92f64d),
	.w8(32'h3bfd7dae),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7ca19),
	.w1(32'hbc0e1782),
	.w2(32'h3c1eabfb),
	.w3(32'hbabc4aa5),
	.w4(32'h3c204412),
	.w5(32'h3aa80931),
	.w6(32'hbbb1f229),
	.w7(32'h3c95e3f4),
	.w8(32'hbba2fcd2),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb771265),
	.w1(32'hbc06332d),
	.w2(32'hbab1babc),
	.w3(32'hb901abda),
	.w4(32'h3be4c09c),
	.w5(32'hbc04dbe1),
	.w6(32'hbb8507dc),
	.w7(32'h3b07ea74),
	.w8(32'hbca98dda),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6125f),
	.w1(32'hbc899c42),
	.w2(32'h3bab8345),
	.w3(32'hba583553),
	.w4(32'h3ca12d2d),
	.w5(32'hbbd69e83),
	.w6(32'hbc608510),
	.w7(32'h3c95394c),
	.w8(32'h39618665),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4adf4),
	.w1(32'hbb5fd117),
	.w2(32'hbc1b7163),
	.w3(32'hbc6af49b),
	.w4(32'hbc5daec7),
	.w5(32'hba8d2124),
	.w6(32'hbc03a755),
	.w7(32'hbc81391e),
	.w8(32'h3bce0bdf),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f2c3f),
	.w1(32'h3a977725),
	.w2(32'hbb260006),
	.w3(32'h3ac8dbdc),
	.w4(32'hbb571407),
	.w5(32'h3a6834b2),
	.w6(32'h3b50baaf),
	.w7(32'h3b18ed49),
	.w8(32'hbb269687),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e26b7),
	.w1(32'hba66637d),
	.w2(32'hbba946b1),
	.w3(32'h3c519c4d),
	.w4(32'h3b229580),
	.w5(32'h3b819a84),
	.w6(32'h3b9bbce7),
	.w7(32'hbaac56d0),
	.w8(32'h3d339c1a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d273f2d),
	.w1(32'h3c1b85d0),
	.w2(32'hbcb2c400),
	.w3(32'hbd1cef15),
	.w4(32'hbd23cda7),
	.w5(32'hbc5adac6),
	.w6(32'hbc0198a0),
	.w7(32'hbd20f311),
	.w8(32'hbc42e848),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e4a52),
	.w1(32'h3ad106b6),
	.w2(32'h3b3a4a4e),
	.w3(32'hbc023c45),
	.w4(32'hbba71f55),
	.w5(32'hbc2f425d),
	.w6(32'hbaea3fb8),
	.w7(32'hb9886dda),
	.w8(32'hbc9d292c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafa174),
	.w1(32'hbcb75c6b),
	.w2(32'hbaa1528f),
	.w3(32'h3bca0f08),
	.w4(32'h3b0c9e55),
	.w5(32'h3b41ff93),
	.w6(32'hbc9b635b),
	.w7(32'h3c63176a),
	.w8(32'hbb978c68),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf50b60),
	.w1(32'hbc03acee),
	.w2(32'hba6e9e15),
	.w3(32'h3b912946),
	.w4(32'h3c2bae5c),
	.w5(32'h3a8bb232),
	.w6(32'hbbb6f898),
	.w7(32'h3a5a4209),
	.w8(32'h3b8c117e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39c1bd),
	.w1(32'h3ba2a4ce),
	.w2(32'hbbb795bb),
	.w3(32'hba8ea7ff),
	.w4(32'hbcb01847),
	.w5(32'h3b1cc53d),
	.w6(32'h3bc36c4e),
	.w7(32'hbc5220bb),
	.w8(32'hbbc69793),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1b151),
	.w1(32'hbc410c5b),
	.w2(32'h3c00659c),
	.w3(32'h3c730d68),
	.w4(32'h3c409970),
	.w5(32'hbc0659d0),
	.w6(32'h3b920499),
	.w7(32'h3c2acbf7),
	.w8(32'hbca7105d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75998b),
	.w1(32'hbbf02700),
	.w2(32'hbbc91e3c),
	.w3(32'h3bd2d6a6),
	.w4(32'h3c26f580),
	.w5(32'hbc268d8c),
	.w6(32'hbbdfdc6a),
	.w7(32'h3bcc44d3),
	.w8(32'hbd5bdd3b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1a7b16),
	.w1(32'hbd239ed3),
	.w2(32'h3c61112a),
	.w3(32'h3cc0a390),
	.w4(32'h3cf1de11),
	.w5(32'h3b9c7607),
	.w6(32'hbcf1155e),
	.w7(32'h3d1e9cd8),
	.w8(32'hbac37dee),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab38b3c),
	.w1(32'hbb8e1d48),
	.w2(32'hbb16d2ad),
	.w3(32'h3b06ecee),
	.w4(32'h3a8cfc6c),
	.w5(32'h3b34bb81),
	.w6(32'hbc4ad12e),
	.w7(32'hbb5c61bc),
	.w8(32'h3c8148ae),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3da1ca),
	.w1(32'h3cba2b00),
	.w2(32'hbb0a3a9a),
	.w3(32'hbc861d6c),
	.w4(32'hbc7706b5),
	.w5(32'h3bb882b6),
	.w6(32'h3c3f233c),
	.w7(32'hbc28a89c),
	.w8(32'h3ce76e7b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c269dff),
	.w1(32'h3c004b48),
	.w2(32'hbc1a596f),
	.w3(32'hbc48cf76),
	.w4(32'hbc832355),
	.w5(32'h3b793f94),
	.w6(32'h3c685cf0),
	.w7(32'hbc99bb5a),
	.w8(32'h3cdc2a72),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f483e),
	.w1(32'h3c722fe5),
	.w2(32'hbb6181be),
	.w3(32'hbc947302),
	.w4(32'hbb2a4097),
	.w5(32'hbb0af40a),
	.w6(32'hbbd3e694),
	.w7(32'hbc4b0222),
	.w8(32'h3c738bcc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c914f02),
	.w1(32'h3c9cc68b),
	.w2(32'hbc2d4284),
	.w3(32'hbc1ad07f),
	.w4(32'hbc630dc3),
	.w5(32'hbb121c58),
	.w6(32'hba25a05a),
	.w7(32'hbc81ba33),
	.w8(32'hbbcb2a7a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a8fe29),
	.w1(32'hbb6c756f),
	.w2(32'hbbf8fa2d),
	.w3(32'h3adae931),
	.w4(32'h3a2e90b8),
	.w5(32'hbadd8534),
	.w6(32'h3c8707fb),
	.w7(32'h3ba58add),
	.w8(32'hb91127ec),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10e600),
	.w1(32'h3b431fa9),
	.w2(32'h3a6540b3),
	.w3(32'h3964e09c),
	.w4(32'h3c056203),
	.w5(32'hbadcf8ed),
	.w6(32'hbb47cbea),
	.w7(32'h3abc1761),
	.w8(32'hbc6c0989),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38be19),
	.w1(32'hbc4db8a4),
	.w2(32'hbb4babb2),
	.w3(32'h3bcc3f06),
	.w4(32'h3c0aa28b),
	.w5(32'hbae9763c),
	.w6(32'hb9d85707),
	.w7(32'h3a87d569),
	.w8(32'h3b4d9383),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule