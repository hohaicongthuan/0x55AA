module layer_10_featuremap_99(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62cc294),
	.w1(32'hb60cb4dc),
	.w2(32'hb53c6808),
	.w3(32'hb667201f),
	.w4(32'h360e9a66),
	.w5(32'hb692ed9e),
	.w6(32'hb670fc94),
	.w7(32'h36061fe3),
	.w8(32'h37763d3d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dabe7b),
	.w1(32'h38bb1eee),
	.w2(32'hb8c71922),
	.w3(32'h389c62a6),
	.w4(32'h38b0695b),
	.w5(32'hb944f189),
	.w6(32'hb7405355),
	.w7(32'h38f2a9e0),
	.w8(32'hb9aca963),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5fc810b),
	.w1(32'hb59dafa3),
	.w2(32'hb5f571db),
	.w3(32'hb4a79f37),
	.w4(32'h3484c042),
	.w5(32'hb548441b),
	.w6(32'hb6058271),
	.w7(32'hb60c8cc9),
	.w8(32'hb58d3716),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c276a1),
	.w1(32'hb83698fc),
	.w2(32'hb88473dd),
	.w3(32'h385fe735),
	.w4(32'h37e0a417),
	.w5(32'hb7a6c919),
	.w6(32'h3861650e),
	.w7(32'h36ae799c),
	.w8(32'hb7964657),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ab6210),
	.w1(32'h37d674ea),
	.w2(32'h37d10007),
	.w3(32'h37a194d3),
	.w4(32'h37b5cfaf),
	.w5(32'h37ec2b01),
	.w6(32'h37920527),
	.w7(32'h374868ff),
	.w8(32'h36f830c7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c72676),
	.w1(32'hb671d2e5),
	.w2(32'h3527be68),
	.w3(32'hb6bad44a),
	.w4(32'hb6a46e56),
	.w5(32'h364eaf02),
	.w6(32'hb727778d),
	.w7(32'hb5e64465),
	.w8(32'hb6b57714),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380c3b1c),
	.w1(32'hb96186a9),
	.w2(32'h37e7c097),
	.w3(32'hb6b5ec3e),
	.w4(32'hb92a379a),
	.w5(32'h38d16885),
	.w6(32'hb8088686),
	.w7(32'hb8f22885),
	.w8(32'h3936073e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd6851),
	.w1(32'hb96f6840),
	.w2(32'hb9ddce95),
	.w3(32'h39e11ebb),
	.w4(32'h38002e30),
	.w5(32'hb9301ebf),
	.w6(32'h3a58e49d),
	.w7(32'hb8c740ab),
	.w8(32'hb9a7e6be),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb844143d),
	.w1(32'h3716e40c),
	.w2(32'hb7d83fbb),
	.w3(32'hb8ad1ad3),
	.w4(32'hb8e9aab3),
	.w5(32'hb889b35c),
	.w6(32'hb80e7574),
	.w7(32'hb8c939a9),
	.w8(32'hb7ffb5aa),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a3291),
	.w1(32'h39299d5f),
	.w2(32'hb9e30fed),
	.w3(32'h39bc36f7),
	.w4(32'h39023dd9),
	.w5(32'hba0f2bf3),
	.w6(32'h3a1185c2),
	.w7(32'h39ce35ad),
	.w8(32'hba313abd),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92b94b1),
	.w1(32'hb8a453aa),
	.w2(32'h38a7c82f),
	.w3(32'hb9719638),
	.w4(32'hb86fb47a),
	.w5(32'hb763569c),
	.w6(32'hb897edf7),
	.w7(32'hb8a97c7b),
	.w8(32'h387b6bde),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949f0d8),
	.w1(32'hba062d28),
	.w2(32'hb8f3b044),
	.w3(32'h39462c92),
	.w4(32'hb9b28d5b),
	.w5(32'h392602cb),
	.w6(32'hb7cf577f),
	.w7(32'hb9d815fa),
	.w8(32'h3942e34e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd0b78),
	.w1(32'h399e5a0d),
	.w2(32'hb999e4f5),
	.w3(32'h3a18dc81),
	.w4(32'h39679d19),
	.w5(32'hba182024),
	.w6(32'h3a33e5a3),
	.w7(32'h39d2ec3b),
	.w8(32'hba15323c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb845cdd9),
	.w1(32'h37caf46d),
	.w2(32'h39e247f7),
	.w3(32'hb8dc8e96),
	.w4(32'h379be059),
	.w5(32'h39adf094),
	.w6(32'hb91fb926),
	.w7(32'hb83a5ed0),
	.w8(32'h39744fe5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981f923),
	.w1(32'h399a471d),
	.w2(32'hb9707fc8),
	.w3(32'h38de5bd4),
	.w4(32'h38b85f3d),
	.w5(32'hb9c55e92),
	.w6(32'h38e1803a),
	.w7(32'h396824d8),
	.w8(32'hb9d3d4e4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d94146),
	.w1(32'h39a48ad6),
	.w2(32'hb9d62b22),
	.w3(32'h39fc71bc),
	.w4(32'h3983c64b),
	.w5(32'hba0aee6d),
	.w6(32'h3a108ccb),
	.w7(32'h39d16c53),
	.w8(32'hb9f60778),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3822a615),
	.w1(32'h38857f14),
	.w2(32'h38d5ff30),
	.w3(32'hb753435c),
	.w4(32'hb80c0689),
	.w5(32'h391088ba),
	.w6(32'hb8a7f9a6),
	.w7(32'hb7cdf422),
	.w8(32'h393adf2e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa62dd2),
	.w1(32'hb8c55680),
	.w2(32'hba50eaed),
	.w3(32'h3a4d0bcf),
	.w4(32'hb9db2082),
	.w5(32'hba07a133),
	.w6(32'h3a8e07eb),
	.w7(32'h392062b1),
	.w8(32'hb9954a5d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a428ade),
	.w1(32'h37fecd6a),
	.w2(32'hb96c69ad),
	.w3(32'h3a296139),
	.w4(32'hb897b113),
	.w5(32'hb92f4ba6),
	.w6(32'h3a1fbb3d),
	.w7(32'h38c4d436),
	.w8(32'hb93e9283),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5987521),
	.w1(32'hb5a3fcdb),
	.w2(32'hb63109fe),
	.w3(32'h366f323e),
	.w4(32'hb67cb90d),
	.w5(32'hb62a82d3),
	.w6(32'h361468f4),
	.w7(32'hb611dde3),
	.w8(32'hb61040b4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35284b68),
	.w1(32'hb6f43b6c),
	.w2(32'h369a0fb4),
	.w3(32'h3699318f),
	.w4(32'hb66b87c4),
	.w5(32'h36efe761),
	.w6(32'hb5968307),
	.w7(32'h36a95b99),
	.w8(32'h36aad267),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb816c158),
	.w1(32'h38619c0c),
	.w2(32'h380e6480),
	.w3(32'hb8c59d36),
	.w4(32'h38544f24),
	.w5(32'h37d585d8),
	.w6(32'hb8b5cca8),
	.w7(32'h38dc931f),
	.w8(32'h37e2ea56),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21e11d),
	.w1(32'hba507244),
	.w2(32'hbb12d3b8),
	.w3(32'h3aba17cb),
	.w4(32'hbaaff004),
	.w5(32'hbb16cdbc),
	.w6(32'h3abfd6fd),
	.w7(32'h39cdaa4a),
	.w8(32'hbabb397a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392ffcae),
	.w1(32'h39c448ea),
	.w2(32'hb9af4a8d),
	.w3(32'h39b0412d),
	.w4(32'h398c6ebd),
	.w5(32'hba17127b),
	.w6(32'h39f7279f),
	.w7(32'h3a026a26),
	.w8(32'hba4cbad8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900f0c2),
	.w1(32'h385eb50f),
	.w2(32'hba8cbf6c),
	.w3(32'h384af121),
	.w4(32'h38b0d6c1),
	.w5(32'hba9ac0fb),
	.w6(32'h39c7b429),
	.w7(32'h39e27a2f),
	.w8(32'hba9f1df6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb846772f),
	.w1(32'h3892175d),
	.w2(32'h38f4481b),
	.w3(32'h387e61a0),
	.w4(32'h38e7eb2c),
	.w5(32'h389cf4a3),
	.w6(32'h388c94e8),
	.w7(32'h38cd96b8),
	.w8(32'h3859fc61),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66b4629),
	.w1(32'hb7417b16),
	.w2(32'h370ab541),
	.w3(32'hb5b2a993),
	.w4(32'hb6e582ae),
	.w5(32'h377d657c),
	.w6(32'hb79eaa66),
	.w7(32'hb5e4a3ec),
	.w8(32'h377adaf7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92310ad),
	.w1(32'h38d07a66),
	.w2(32'hb88285ac),
	.w3(32'hb8b8e6d6),
	.w4(32'h3939c995),
	.w5(32'hb7aaf259),
	.w6(32'hb9384a0d),
	.w7(32'h398394fc),
	.w8(32'hb81c8ea6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3826ecde),
	.w1(32'hb8f65bc5),
	.w2(32'h38204290),
	.w3(32'h3761a6a1),
	.w4(32'hb79d5218),
	.w5(32'h3978655e),
	.w6(32'hb9614c27),
	.w7(32'hb88c8966),
	.w8(32'h3905c52c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7acb9ed),
	.w1(32'h3a268f8d),
	.w2(32'h380b6bf2),
	.w3(32'h39201f51),
	.w4(32'h3a014957),
	.w5(32'hb9b0891d),
	.w6(32'h39ca98a4),
	.w7(32'h3a1847de),
	.w8(32'hb9fbc38c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c79a94),
	.w1(32'hb56967fb),
	.w2(32'h37247d0c),
	.w3(32'hb5702a18),
	.w4(32'hb5455a9b),
	.w5(32'h37496ed7),
	.w6(32'h35c4a72e),
	.w7(32'h37136263),
	.w8(32'h376d3d4c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75ffbfe),
	.w1(32'hb88d1491),
	.w2(32'h38129d25),
	.w3(32'hb84a33fd),
	.w4(32'hb83e7ec1),
	.w5(32'h388005a6),
	.w6(32'hb814553c),
	.w7(32'hb8012a25),
	.w8(32'h38854a05),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39893068),
	.w1(32'h38ffc51c),
	.w2(32'hb90eee02),
	.w3(32'h399afa23),
	.w4(32'h38ec18ba),
	.w5(32'hb9868362),
	.w6(32'h39c7e3d5),
	.w7(32'h393f8f1c),
	.w8(32'hb988f444),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39017cd2),
	.w1(32'h38b9874c),
	.w2(32'hb91a0b97),
	.w3(32'h398b0fb3),
	.w4(32'h390d847f),
	.w5(32'hb9413766),
	.w6(32'h39bb17d3),
	.w7(32'h39b02045),
	.w8(32'hb96099c2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3798bd81),
	.w1(32'hb7faf37b),
	.w2(32'hb76e2981),
	.w3(32'h379d0ff1),
	.w4(32'hb8187074),
	.w5(32'hb73d7edb),
	.w6(32'hb68542a3),
	.w7(32'hb79c4c37),
	.w8(32'h366c8943),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c1a0f1),
	.w1(32'hb90dcfaf),
	.w2(32'hb92cc1ec),
	.w3(32'h3916686c),
	.w4(32'hb902adf5),
	.w5(32'hb907ca5e),
	.w6(32'h398d01d6),
	.w7(32'h380c12f4),
	.w8(32'hb832f2c3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c5a0d),
	.w1(32'hb957a471),
	.w2(32'hb9f94786),
	.w3(32'h3a108b80),
	.w4(32'hb8b31f7e),
	.w5(32'hb9ef3c7d),
	.w6(32'h39706dfa),
	.w7(32'hb96fa53b),
	.w8(32'hb9cc91af),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96974f),
	.w1(32'h39a8ce61),
	.w2(32'hb8c34894),
	.w3(32'hb9e2ea56),
	.w4(32'h39da2bfd),
	.w5(32'hb9506add),
	.w6(32'hba9d00ca),
	.w7(32'h3a02512a),
	.w8(32'hba07e692),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac15f4),
	.w1(32'h392d9050),
	.w2(32'h38a0f88d),
	.w3(32'hba5ec7c2),
	.w4(32'h3756adb7),
	.w5(32'hb9652298),
	.w6(32'hba851fc2),
	.w7(32'h39966ebe),
	.w8(32'hb9a46c93),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90bdeca),
	.w1(32'h3903c8d8),
	.w2(32'h38a018fd),
	.w3(32'hb95499e6),
	.w4(32'h38839e21),
	.w5(32'hb78d7613),
	.w6(32'hb95985fa),
	.w7(32'h38691499),
	.w8(32'hb8b502f6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f81f3f),
	.w1(32'hb8838ce3),
	.w2(32'hb8555403),
	.w3(32'h37a4ef35),
	.w4(32'hb7ee9890),
	.w5(32'h37549bee),
	.w6(32'h37943b43),
	.w7(32'h3810dc3c),
	.w8(32'h38555e65),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928bb6d),
	.w1(32'h3912f658),
	.w2(32'h37624f36),
	.w3(32'h3929c335),
	.w4(32'h38f7ed58),
	.w5(32'hb689191f),
	.w6(32'h38a1a3f7),
	.w7(32'h3829bf63),
	.w8(32'h36f42ab4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce7112),
	.w1(32'hb921f3ec),
	.w2(32'h398dbf9d),
	.w3(32'h380140e7),
	.w4(32'hb8777d10),
	.w5(32'h39a918a7),
	.w6(32'h37d64845),
	.w7(32'hb8f715e5),
	.w8(32'h393e3e69),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57dbdd),
	.w1(32'h3a1f29a6),
	.w2(32'hba0180e8),
	.w3(32'h3a87bf84),
	.w4(32'h39f123c8),
	.w5(32'hba431d88),
	.w6(32'h3a655069),
	.w7(32'h3a15a870),
	.w8(32'hba0abda7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d9c9a),
	.w1(32'h3a1a3d82),
	.w2(32'hb942bea9),
	.w3(32'h39d86da3),
	.w4(32'h39de0f25),
	.w5(32'hba115648),
	.w6(32'h3a101af7),
	.w7(32'h3a184ebb),
	.w8(32'hba3a197d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9fec6),
	.w1(32'h3a157ba2),
	.w2(32'hba105099),
	.w3(32'h3a0fc958),
	.w4(32'h39c77a34),
	.w5(32'hba730485),
	.w6(32'h3a6c9a3f),
	.w7(32'h3a48419b),
	.w8(32'hba875d17),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c8682),
	.w1(32'h3a5826cf),
	.w2(32'hb9bc8d03),
	.w3(32'h3a5b93cb),
	.w4(32'h3a11e190),
	.w5(32'hba6b6629),
	.w6(32'h3a74b180),
	.w7(32'h3a1afbbd),
	.w8(32'hba757386),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affd383),
	.w1(32'h38f45e1a),
	.w2(32'hba43b818),
	.w3(32'h3afb7175),
	.w4(32'hb89003fc),
	.w5(32'hb9d70ae1),
	.w6(32'h3af44393),
	.w7(32'h39d73d4d),
	.w8(32'hb9bafb29),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e067f9),
	.w1(32'h38b00b6d),
	.w2(32'hb6eeb90d),
	.w3(32'hb7f5d470),
	.w4(32'h3879bbaf),
	.w5(32'hb817f1f7),
	.w6(32'h3763dc68),
	.w7(32'h38ceef93),
	.w8(32'h384ee17c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38562702),
	.w1(32'h390f4598),
	.w2(32'hb9592ad2),
	.w3(32'h38f9fdc6),
	.w4(32'h37ae69f5),
	.w5(32'hb93021ef),
	.w6(32'h39717b4e),
	.w7(32'h38519dc3),
	.w8(32'hb8afeafd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39294954),
	.w1(32'h38fa1c67),
	.w2(32'hb71b83fc),
	.w3(32'h384fa455),
	.w4(32'h38e4f12a),
	.w5(32'h388acbe6),
	.w6(32'hb82d6758),
	.w7(32'hb892bb27),
	.w8(32'h37b7ab17),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3856ae25),
	.w1(32'h391108dd),
	.w2(32'hb9ba3932),
	.w3(32'h39110b76),
	.w4(32'h3908b049),
	.w5(32'hb9fe1a56),
	.w6(32'h39af19b3),
	.w7(32'h39d671d6),
	.w8(32'hb9c54661),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cd593a),
	.w1(32'hb80ffefd),
	.w2(32'hb91c1480),
	.w3(32'h390191bf),
	.w4(32'hb805a1b9),
	.w5(32'hb91953e3),
	.w6(32'h396fc352),
	.w7(32'h38f385b4),
	.w8(32'hb88f1f62),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5901b1),
	.w1(32'hb9dadcb5),
	.w2(32'hba037d2b),
	.w3(32'h3a54be27),
	.w4(32'hb9c0a4c9),
	.w5(32'hba1160d1),
	.w6(32'h3a413ea3),
	.w7(32'hb74e676f),
	.w8(32'hb9c23d7c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3765867c),
	.w1(32'hb8add56e),
	.w2(32'hb88f3688),
	.w3(32'hb7ca847e),
	.w4(32'h379c9949),
	.w5(32'hb76b9c46),
	.w6(32'h37f4de77),
	.w7(32'h38d1394c),
	.w8(32'hb89fea35),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b0b5a8),
	.w1(32'hb61b4059),
	.w2(32'h3754677e),
	.w3(32'h369fa4b5),
	.w4(32'h36064610),
	.w5(32'h373f1b52),
	.w6(32'hb73b093e),
	.w7(32'h3738d62a),
	.w8(32'h36f4070e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6534a0d),
	.w1(32'hb6d5d4c5),
	.w2(32'h34d47b7b),
	.w3(32'h33e97300),
	.w4(32'hb6c5a512),
	.w5(32'h36347fb0),
	.w6(32'hb6789b15),
	.w7(32'hb4e4b3ec),
	.w8(32'h3578ef1d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bffd57),
	.w1(32'h37e3ff10),
	.w2(32'h379cac1a),
	.w3(32'h36e81554),
	.w4(32'h376e6bc1),
	.w5(32'h37fb66a0),
	.w6(32'h370efb01),
	.w7(32'hb608000d),
	.w8(32'hb6c3e206),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82f72f1),
	.w1(32'hb68a52e9),
	.w2(32'h38a31c84),
	.w3(32'hb6270dd8),
	.w4(32'h371f21f2),
	.w5(32'h38837671),
	.w6(32'hb6979eef),
	.w7(32'h38217aa7),
	.w8(32'h384971d7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71cc818),
	.w1(32'h38a8de5a),
	.w2(32'h37af854b),
	.w3(32'hb8eae83a),
	.w4(32'h38047bc9),
	.w5(32'hb7a61856),
	.w6(32'hb8c6b75d),
	.w7(32'hb7c43a18),
	.w8(32'hb7ad5f7c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb2673),
	.w1(32'hb79b712f),
	.w2(32'hb90e93e4),
	.w3(32'h39ba3fe4),
	.w4(32'hb830f66d),
	.w5(32'hb8d2ba2d),
	.w6(32'h3992cf49),
	.w7(32'h381de717),
	.w8(32'h3807f1e6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987d7e3),
	.w1(32'hb9594a51),
	.w2(32'hb9ad4829),
	.w3(32'hb8c2a4c7),
	.w4(32'hb92a7fa7),
	.w5(32'hb99a2494),
	.w6(32'h39862741),
	.w7(32'h39468ab9),
	.w8(32'hb9163d33),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37219466),
	.w1(32'hb6950b7d),
	.w2(32'hb70d7c24),
	.w3(32'h380513fb),
	.w4(32'h3622938a),
	.w5(32'hb60f15c5),
	.w6(32'h383e607a),
	.w7(32'h375df152),
	.w8(32'h37e75d14),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a12b3d),
	.w1(32'h356d4b41),
	.w2(32'hb585618d),
	.w3(32'h3506f9f1),
	.w4(32'h361d3b83),
	.w5(32'hb217f5d8),
	.w6(32'h359c5f11),
	.w7(32'hb5ff4ec2),
	.w8(32'h35661a61),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7411914),
	.w1(32'hb75f20ef),
	.w2(32'h3786aa5d),
	.w3(32'h37098793),
	.w4(32'hb7e210ee),
	.w5(32'h36a119a6),
	.w6(32'hb799ee96),
	.w7(32'h36348073),
	.w8(32'hb52076ed),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7574741),
	.w1(32'hb58408d2),
	.w2(32'h36d83654),
	.w3(32'hb74100c3),
	.w4(32'h357975cb),
	.w5(32'h378210ad),
	.w6(32'hb680a736),
	.w7(32'hb6a1ee73),
	.w8(32'h370be1ed),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c41d4),
	.w1(32'hb98d6dd3),
	.w2(32'hb9746b21),
	.w3(32'h39589102),
	.w4(32'hb946974e),
	.w5(32'hb9b82cab),
	.w6(32'hb8bcbcd9),
	.w7(32'hb908be6f),
	.w8(32'hb94bc440),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3967b4b3),
	.w1(32'h38f60652),
	.w2(32'hba2d505b),
	.w3(32'h39ae5776),
	.w4(32'h391b2669),
	.w5(32'hba61c388),
	.w6(32'h3a5d8a4a),
	.w7(32'h3a2b6727),
	.w8(32'hba7e32df),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995a643),
	.w1(32'hb9ffb8a8),
	.w2(32'hba578240),
	.w3(32'hb903cb48),
	.w4(32'hb9e6762d),
	.w5(32'hba55aada),
	.w6(32'h3a02796b),
	.w7(32'h393c823b),
	.w8(32'hba43b6c4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70f73ed),
	.w1(32'h3a2e15a5),
	.w2(32'hb9f7d250),
	.w3(32'h39fc4544),
	.w4(32'h3a1fb4b3),
	.w5(32'hba2799fd),
	.w6(32'h3a508e11),
	.w7(32'h3a9c667c),
	.w8(32'hba6a20e8),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66e7e19),
	.w1(32'h364c97be),
	.w2(32'h3554bbb8),
	.w3(32'h3628273e),
	.w4(32'h36200d25),
	.w5(32'h35cc7f0e),
	.w6(32'h3699ace4),
	.w7(32'h360bcfbe),
	.w8(32'h36c6416f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb655065d),
	.w1(32'hb6d00f18),
	.w2(32'h36e1b594),
	.w3(32'h35005efa),
	.w4(32'hb65f90a1),
	.w5(32'h37291bdf),
	.w6(32'hb6d6790c),
	.w7(32'hb62bc44d),
	.w8(32'h371a6d13),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ae4484),
	.w1(32'h3509a63a),
	.w2(32'h3704c551),
	.w3(32'hb27d2c1f),
	.w4(32'hb65eb705),
	.w5(32'h3643407b),
	.w6(32'hb5e11b23),
	.w7(32'hb6292d33),
	.w8(32'h370e2c5a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c5e796),
	.w1(32'hb88194e6),
	.w2(32'hb7ccb991),
	.w3(32'h38911849),
	.w4(32'hb7fee647),
	.w5(32'h3581fe6e),
	.w6(32'h389c5e14),
	.w7(32'hb61a9a5c),
	.w8(32'hb77fbcfe),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c903e4),
	.w1(32'h3877d9d9),
	.w2(32'h371034d8),
	.w3(32'h38907d9c),
	.w4(32'h37c0027a),
	.w5(32'hb7f4b97a),
	.w6(32'h3884b18d),
	.w7(32'h3716023f),
	.w8(32'hb825ed34),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53bfc8),
	.w1(32'hb951d25b),
	.w2(32'hb9d5da64),
	.w3(32'h3a432440),
	.w4(32'hb85c9635),
	.w5(32'hb986a128),
	.w6(32'h3a0ce47e),
	.w7(32'h376ef322),
	.w8(32'hb9407135),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5eb2d),
	.w1(32'h38686442),
	.w2(32'hba56e56a),
	.w3(32'h3ab6799b),
	.w4(32'hb842a4be),
	.w5(32'hba7544eb),
	.w6(32'h3aa93332),
	.w7(32'hb8999f06),
	.w8(32'hba17fff9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39807d60),
	.w1(32'h3a0c098b),
	.w2(32'hb9d599e0),
	.w3(32'h39d4f544),
	.w4(32'h39afe070),
	.w5(32'hba3bbb1d),
	.w6(32'h39d6aaad),
	.w7(32'h3a0a98dc),
	.w8(32'hba4d06d3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0234b6),
	.w1(32'h38da9895),
	.w2(32'hb965e7db),
	.w3(32'h39e2b671),
	.w4(32'h378abc73),
	.w5(32'hb9807853),
	.w6(32'h3a070b76),
	.w7(32'h392b64bc),
	.w8(32'hb985fbac),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ef96b),
	.w1(32'h3751dc45),
	.w2(32'hb8db6dd0),
	.w3(32'h390953cc),
	.w4(32'hb8c04373),
	.w5(32'hb979d100),
	.w6(32'h385f6558),
	.w7(32'hb80a932b),
	.w8(32'hb933e6c3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89fa210),
	.w1(32'h367ae801),
	.w2(32'hb92fa550),
	.w3(32'h3677a729),
	.w4(32'hb3bd9dd4),
	.w5(32'hb9805e53),
	.w6(32'h37c36a64),
	.w7(32'h38d41a3e),
	.w8(32'hb9915013),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a549d80),
	.w1(32'h399138b1),
	.w2(32'hb9ac5bf2),
	.w3(32'h3a422ce8),
	.w4(32'hb7a28773),
	.w5(32'hb9982a1f),
	.w6(32'h3a37dbd5),
	.w7(32'h39484c95),
	.w8(32'hb95bcce9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61996b4),
	.w1(32'hb5fb0872),
	.w2(32'h35ff5821),
	.w3(32'hb452461b),
	.w4(32'h34a50ff3),
	.w5(32'h361e6b87),
	.w6(32'hb5ab07cd),
	.w7(32'h362ea326),
	.w8(32'h368877b6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6699116),
	.w1(32'hb533ce61),
	.w2(32'h33232bbf),
	.w3(32'hb5da9cc0),
	.w4(32'h368b6819),
	.w5(32'h350d40e9),
	.w6(32'h33e8a678),
	.w7(32'h35046ea5),
	.w8(32'hb55877cf),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb807d1f8),
	.w1(32'hb7791b4f),
	.w2(32'hb7d268d4),
	.w3(32'hb7b377ef),
	.w4(32'hb70b63b6),
	.w5(32'hb760485d),
	.w6(32'hb863dd02),
	.w7(32'h370b8b05),
	.w8(32'hb825c098),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36180bb6),
	.w1(32'h373e67da),
	.w2(32'h37917252),
	.w3(32'hb6dff204),
	.w4(32'h3711712c),
	.w5(32'h37a1c028),
	.w6(32'hb73c598f),
	.w7(32'h34c06810),
	.w8(32'h376e61d2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5032b8),
	.w1(32'h38e8f2a4),
	.w2(32'hb93e64ba),
	.w3(32'hb95b1c50),
	.w4(32'h38bec7ce),
	.w5(32'hb9a1842f),
	.w6(32'hb923649b),
	.w7(32'h3995189b),
	.w8(32'hba0395a5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379b0afd),
	.w1(32'h379bb101),
	.w2(32'h3762f9c6),
	.w3(32'hb6eff53c),
	.w4(32'h3734f667),
	.w5(32'hb7b8c05f),
	.w6(32'hb75d6bd2),
	.w7(32'h3887de7f),
	.w8(32'hb74b877a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39232660),
	.w1(32'h3964f310),
	.w2(32'hb91d94f6),
	.w3(32'h394831fb),
	.w4(32'h3900e0e4),
	.w5(32'hb97b41f0),
	.w6(32'h39ba572f),
	.w7(32'h397c8789),
	.w8(32'hb9a00a3f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bf35c),
	.w1(32'hb9cbfee6),
	.w2(32'hba6c5ab5),
	.w3(32'h3ad6bf9e),
	.w4(32'hb9d955a9),
	.w5(32'hba59b7c9),
	.w6(32'h3afa6e18),
	.w7(32'hb8e9f4fa),
	.w8(32'hba5721b7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cef179),
	.w1(32'hb88e5373),
	.w2(32'hb5bce25d),
	.w3(32'hb980fd72),
	.w4(32'hb8933e58),
	.w5(32'hb8168229),
	.w6(32'hb9afb4c3),
	.w7(32'hb736ee07),
	.w8(32'h37aaa064),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a018464),
	.w1(32'h39227993),
	.w2(32'hb9d1b4ec),
	.w3(32'h3a33739a),
	.w4(32'hb8d13ff0),
	.w5(32'hb9fc30fe),
	.w6(32'h39b63b75),
	.w7(32'h39c65cd3),
	.w8(32'hb8f60989),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad0569),
	.w1(32'hb897c7a3),
	.w2(32'hb8343176),
	.w3(32'hb994a452),
	.w4(32'hb6b5397d),
	.w5(32'hb9112ea3),
	.w6(32'h37e01fa1),
	.w7(32'h391916aa),
	.w8(32'hb9297812),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad72b7),
	.w1(32'h38900dd2),
	.w2(32'hb9a2d59f),
	.w3(32'h39bd9e50),
	.w4(32'h37a91e67),
	.w5(32'hba0d8c25),
	.w6(32'h3a0d4078),
	.w7(32'h39a6c4fc),
	.w8(32'hba02947c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a6d03),
	.w1(32'hb8f9bf5c),
	.w2(32'hb96a482a),
	.w3(32'hb79b7f13),
	.w4(32'hb94fb530),
	.w5(32'hb99bc019),
	.w6(32'hb8f53b89),
	.w7(32'hb90a2bf3),
	.w8(32'hb93e91dc),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95fcb85),
	.w1(32'h39a7f738),
	.w2(32'hb93c97e3),
	.w3(32'hb964f4b8),
	.w4(32'h3937cf07),
	.w5(32'hb9d54e32),
	.w6(32'hb90263c4),
	.w7(32'h39b98d4d),
	.w8(32'hb9ff9026),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb158e),
	.w1(32'h391475fb),
	.w2(32'h37c344ff),
	.w3(32'h38559890),
	.w4(32'h37bba111),
	.w5(32'h388b8101),
	.w6(32'h39325fb2),
	.w7(32'h388491bd),
	.w8(32'h38a66b4c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cf9c1),
	.w1(32'h39ea8193),
	.w2(32'hba127c69),
	.w3(32'h3a2a6f64),
	.w4(32'h391bfe38),
	.w5(32'hba5cd75f),
	.w6(32'h3a5260ae),
	.w7(32'h38be5196),
	.w8(32'hba80bd90),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89f6c6c),
	.w1(32'hb5abee94),
	.w2(32'hb9a2e630),
	.w3(32'hb92460b8),
	.w4(32'hb996db8e),
	.w5(32'hba48fd81),
	.w6(32'hb90c786a),
	.w7(32'hb982cc8d),
	.w8(32'hba2be4a4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2b605),
	.w1(32'hb910daf7),
	.w2(32'hba761c85),
	.w3(32'h3ae0dde0),
	.w4(32'hb93dfe9e),
	.w5(32'hba39fcd5),
	.w6(32'h3ac7395c),
	.w7(32'h3912e918),
	.w8(32'hba1b76b8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2190da),
	.w1(32'h39c024c6),
	.w2(32'h3a6af4e1),
	.w3(32'hbaaf598c),
	.w4(32'h39170b6b),
	.w5(32'h39fbccf6),
	.w6(32'hbaa0ef8e),
	.w7(32'h3a059c9f),
	.w8(32'hb98bae6c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392ee5e1),
	.w1(32'h39c568d1),
	.w2(32'hba346b90),
	.w3(32'h3a18fe7b),
	.w4(32'h390cf296),
	.w5(32'hba50284b),
	.w6(32'h3a3f795e),
	.w7(32'h3a15a0f1),
	.w8(32'hba66ce22),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a4d87),
	.w1(32'hb79cc52a),
	.w2(32'hb9a93fec),
	.w3(32'h39edef39),
	.w4(32'hb88bc41c),
	.w5(32'hb9697cd7),
	.w6(32'h3a17eebb),
	.w7(32'h39a6e1b2),
	.w8(32'hb912d452),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395bc8dc),
	.w1(32'h39d8e01c),
	.w2(32'h39b1507f),
	.w3(32'h38db13ae),
	.w4(32'h3915f2d8),
	.w5(32'h381f04f3),
	.w6(32'h38f7d47e),
	.w7(32'h383554f8),
	.w8(32'hb95ace06),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa50cbb),
	.w1(32'h397eb32e),
	.w2(32'hba26740b),
	.w3(32'h3adee2fb),
	.w4(32'h387f8214),
	.w5(32'hba0f2047),
	.w6(32'h3a9d6fc8),
	.w7(32'hb82e82df),
	.w8(32'hba1e7121),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9901a0f),
	.w1(32'h39ec6e2a),
	.w2(32'hb8aada5e),
	.w3(32'h3780e612),
	.w4(32'h39c069b8),
	.w5(32'hb8b9cada),
	.w6(32'hb7df7080),
	.w7(32'h39da5187),
	.w8(32'hb900d05d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3793f966),
	.w1(32'h37c635e7),
	.w2(32'h37553860),
	.w3(32'hb7188ea6),
	.w4(32'h35e89198),
	.w5(32'h36d0e343),
	.w6(32'hb7ff6b6c),
	.w7(32'hb7928703),
	.w8(32'hb41793d2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386bf10f),
	.w1(32'h38678678),
	.w2(32'hb7c8a6c0),
	.w3(32'h37d429cf),
	.w4(32'h37373301),
	.w5(32'hb8b08863),
	.w6(32'h394ce887),
	.w7(32'h390fd5e5),
	.w8(32'hb7ebe03c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1edcf6),
	.w1(32'h39ff41fe),
	.w2(32'hb9841462),
	.w3(32'h3a3e097d),
	.w4(32'h39c8f529),
	.w5(32'hba00703b),
	.w6(32'h3a09df56),
	.w7(32'h39ca7964),
	.w8(32'hba0bfe74),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cf922e),
	.w1(32'h3a1b5eee),
	.w2(32'hb9b3bec2),
	.w3(32'h39ab9904),
	.w4(32'h39bf43d0),
	.w5(32'hb9d3334e),
	.w6(32'h3a3afe55),
	.w7(32'h3a19cdf3),
	.w8(32'hb9e811c0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e557a8),
	.w1(32'hb917fc30),
	.w2(32'hb989f398),
	.w3(32'hb991b4e6),
	.w4(32'hb9565be7),
	.w5(32'hb997b25d),
	.w6(32'hb996b5fd),
	.w7(32'h38710d32),
	.w8(32'hb9e1effe),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f2cca4),
	.w1(32'h38d79168),
	.w2(32'hb99b5569),
	.w3(32'hb78101b4),
	.w4(32'hb8288746),
	.w5(32'hb9ca7b95),
	.w6(32'h39842cb1),
	.w7(32'h3995917a),
	.w8(32'hb9ceb381),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366c4fe0),
	.w1(32'hb92c53cf),
	.w2(32'hb93a3842),
	.w3(32'h38bd6907),
	.w4(32'hb9175e51),
	.w5(32'hb8a91615),
	.w6(32'h394633a1),
	.w7(32'h39295803),
	.w8(32'hb8a56894),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395887fd),
	.w1(32'h392a897c),
	.w2(32'hb8de2791),
	.w3(32'h391b922e),
	.w4(32'hb8b93aa9),
	.w5(32'hb946f501),
	.w6(32'h3990eb29),
	.w7(32'h38e7a6d3),
	.w8(32'hb85634ab),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d555d4),
	.w1(32'h396e106a),
	.w2(32'hb9192a4f),
	.w3(32'h389196e9),
	.w4(32'h39576a52),
	.w5(32'hb99089e9),
	.w6(32'h392a3e4e),
	.w7(32'h39a51cb7),
	.w8(32'hb9ac4208),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74cd9d0),
	.w1(32'hb6af2c0d),
	.w2(32'h360e4537),
	.w3(32'hb7527d59),
	.w4(32'hb78dc116),
	.w5(32'h365db275),
	.w6(32'hb769ee6f),
	.w7(32'hb70f3ffd),
	.w8(32'hb6452709),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7565ad5),
	.w1(32'hb6c1759a),
	.w2(32'hb632f896),
	.w3(32'hb502f4d3),
	.w4(32'hb6d7c07c),
	.w5(32'hb6337729),
	.w6(32'hb7335ae8),
	.w7(32'hb70382fe),
	.w8(32'hb6e9dfa4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79342c4),
	.w1(32'hb70b2445),
	.w2(32'hb50ebd04),
	.w3(32'hb73847f9),
	.w4(32'h3697a0ea),
	.w5(32'h371e1316),
	.w6(32'hb72247e4),
	.w7(32'h3597e051),
	.w8(32'h36293fc4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d6acef),
	.w1(32'h37182571),
	.w2(32'h37e0c804),
	.w3(32'hb718d996),
	.w4(32'h375e6194),
	.w5(32'h37c217ad),
	.w6(32'hb60e076a),
	.w7(32'h365ab73e),
	.w8(32'h377044c9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a5d553),
	.w1(32'h39802fa4),
	.w2(32'hb981f795),
	.w3(32'h39082ae2),
	.w4(32'h3914aa0f),
	.w5(32'hb9fa32b0),
	.w6(32'h397a0249),
	.w7(32'h398432f1),
	.w8(32'hba06b86b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ae5814),
	.w1(32'h364d25c7),
	.w2(32'h38a21a5a),
	.w3(32'hb80931e7),
	.w4(32'h36bf8ade),
	.w5(32'h385586ab),
	.w6(32'hb63353a6),
	.w7(32'h37ea609d),
	.w8(32'h379e72e7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3a1aa),
	.w1(32'hb80bc61a),
	.w2(32'hb90e6fd1),
	.w3(32'h39851658),
	.w4(32'hb6dc62d2),
	.w5(32'hb81068f6),
	.w6(32'h39cebb81),
	.w7(32'h38aaa23f),
	.w8(32'h3821082a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba161a66),
	.w1(32'h396dbebd),
	.w2(32'hb94b89eb),
	.w3(32'hb9bd7f60),
	.w4(32'h39655aa6),
	.w5(32'hb9950b41),
	.w6(32'hb9777b8b),
	.w7(32'h3a060c5f),
	.w8(32'hb9ff3973),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362cfbf7),
	.w1(32'h36c49c96),
	.w2(32'hb6c7549d),
	.w3(32'h3720ad24),
	.w4(32'h37894f05),
	.w5(32'h3698859a),
	.w6(32'h3692ae68),
	.w7(32'h37009c84),
	.w8(32'hb58f7d13),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3783754a),
	.w1(32'hb634c13f),
	.w2(32'h375c6f5b),
	.w3(32'h3773b4dc),
	.w4(32'hb6a945be),
	.w5(32'h3797d881),
	.w6(32'h364c958f),
	.w7(32'hb70fad3e),
	.w8(32'h3751eefc),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61bb70e),
	.w1(32'hb667b65b),
	.w2(32'h376c406e),
	.w3(32'hb6ae2c6d),
	.w4(32'hb53b23e4),
	.w5(32'h35e7d1a0),
	.w6(32'h3732db8f),
	.w7(32'h3700c59e),
	.w8(32'h3722703e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0d3ac),
	.w1(32'h38963d18),
	.w2(32'h384792f7),
	.w3(32'hb7c18984),
	.w4(32'h388a933c),
	.w5(32'h37b85de9),
	.w6(32'hb73c4053),
	.w7(32'h38a6c171),
	.w8(32'hb82bb376),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39601448),
	.w1(32'hb85b2593),
	.w2(32'hb995095f),
	.w3(32'h394293e3),
	.w4(32'hb96976c8),
	.w5(32'hb9b0b835),
	.w6(32'h39e79681),
	.w7(32'h38904b7b),
	.w8(32'hb9859264),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a019d3d),
	.w1(32'h38adeeae),
	.w2(32'hb9349394),
	.w3(32'h39ebe371),
	.w4(32'h389bc80e),
	.w5(32'hb94ab71b),
	.w6(32'h3a0d4ffc),
	.w7(32'h396b0fa9),
	.w8(32'hb9697ad9),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38725789),
	.w1(32'hb7f48371),
	.w2(32'hb751d136),
	.w3(32'h389a7740),
	.w4(32'hb7541643),
	.w5(32'h36c3684e),
	.w6(32'h37f2dccc),
	.w7(32'hb77319e8),
	.w8(32'h370a3e06),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90478c9),
	.w1(32'hb8816056),
	.w2(32'hb8e54244),
	.w3(32'hb7204cd4),
	.w4(32'hb85739e9),
	.w5(32'hb902419e),
	.w6(32'h394b948a),
	.w7(32'h3822069b),
	.w8(32'hb9363c63),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb882006f),
	.w1(32'h381d55c3),
	.w2(32'hb79f3c72),
	.w3(32'hb7c64f79),
	.w4(32'h368de6f0),
	.w5(32'hb8e3e9c9),
	.w6(32'hb828ee73),
	.w7(32'h382bdb04),
	.w8(32'hb8e7d8a4),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985aaad),
	.w1(32'hb7b1b26b),
	.w2(32'hb94c62dd),
	.w3(32'h39773c3a),
	.w4(32'hb706a6d6),
	.w5(32'hb943acb2),
	.w6(32'h39bee107),
	.w7(32'h382cb474),
	.w8(32'hb93cf326),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42da1e),
	.w1(32'h38afff3f),
	.w2(32'hb944e616),
	.w3(32'h3a2e608b),
	.w4(32'h38dead08),
	.w5(32'hb949c358),
	.w6(32'h3a45f317),
	.w7(32'h3847a017),
	.w8(32'hb98d7239),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a184b1e),
	.w1(32'h37375fb1),
	.w2(32'hba02bedb),
	.w3(32'h3a18c319),
	.w4(32'hb8342cac),
	.w5(32'hba0cb27c),
	.w6(32'h3a39c98a),
	.w7(32'h398f9a6e),
	.w8(32'hb9aba5fc),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37daad6e),
	.w1(32'h39b80ebd),
	.w2(32'hb8b341c6),
	.w3(32'h38575859),
	.w4(32'h3981b1ed),
	.w5(32'hb96cc770),
	.w6(32'h39271c59),
	.w7(32'h3a0001f5),
	.w8(32'hb9a322b5),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89cf432),
	.w1(32'h39015d68),
	.w2(32'hb990f5d8),
	.w3(32'hb800a635),
	.w4(32'hb80eb7aa),
	.w5(32'hb9c258b9),
	.w6(32'h38f907da),
	.w7(32'h3991b2de),
	.w8(32'hb8a05f35),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15227b),
	.w1(32'hba09a724),
	.w2(32'hb9c0ccb1),
	.w3(32'h3a30f76e),
	.w4(32'hb9839631),
	.w5(32'hb9ca93a6),
	.w6(32'h3a110ed3),
	.w7(32'hb88b24aa),
	.w8(32'hb95d9fa9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39039d19),
	.w1(32'h391a6175),
	.w2(32'hb9318e14),
	.w3(32'h396ad6c4),
	.w4(32'h3882ff0b),
	.w5(32'hb96a6bb5),
	.w6(32'h39c2ed89),
	.w7(32'h399d7cfc),
	.w8(32'hb9ad9ac3),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38978bed),
	.w1(32'h38f8122d),
	.w2(32'hb8bd0514),
	.w3(32'h3906ff9b),
	.w4(32'h38de3eef),
	.w5(32'hb947be51),
	.w6(32'h3921cd58),
	.w7(32'h3921e0f7),
	.w8(32'hb9319fbd),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38be4b21),
	.w1(32'h38bf1f63),
	.w2(32'hb85e8f8b),
	.w3(32'h38dfaea5),
	.w4(32'h3860aa88),
	.w5(32'hb8ca88c5),
	.w6(32'h38fc03c0),
	.w7(32'h3886bc3a),
	.w8(32'hb8dfddf9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f0fac),
	.w1(32'h39ae5e0d),
	.w2(32'hb97b09b0),
	.w3(32'hb907ed01),
	.w4(32'h39794422),
	.w5(32'hba073ff2),
	.w6(32'hb8a2c832),
	.w7(32'h3a08b1f6),
	.w8(32'hba2591fc),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bc154f),
	.w1(32'hb80b77f2),
	.w2(32'hb90ab2dc),
	.w3(32'hb843f2d8),
	.w4(32'hb8020240),
	.w5(32'hb8f10ef2),
	.w6(32'h37c6ef4f),
	.w7(32'h37bb9d91),
	.w8(32'hb90c894d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36802396),
	.w1(32'hb43a51ba),
	.w2(32'h3685bc2c),
	.w3(32'h373637f5),
	.w4(32'h36038d9c),
	.w5(32'h36474eb8),
	.w6(32'hb4274925),
	.w7(32'hb49015d3),
	.w8(32'h3697cb30),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb607cd8c),
	.w1(32'h364f7e8b),
	.w2(32'h36749308),
	.w3(32'hb637ccf7),
	.w4(32'hb6db6223),
	.w5(32'hb445e218),
	.w6(32'h371660cd),
	.w7(32'hb4bf2d9d),
	.w8(32'h35181624),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93aa5bf),
	.w1(32'h393fa6a4),
	.w2(32'hb8293592),
	.w3(32'h38282bdc),
	.w4(32'h39153a2c),
	.w5(32'hb7ccb765),
	.w6(32'h370cdc8a),
	.w7(32'h39915847),
	.w8(32'hb858bd06),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84c7e70),
	.w1(32'h391f9f5b),
	.w2(32'hb948196b),
	.w3(32'hb80328c3),
	.w4(32'h387aa03e),
	.w5(32'hb9dce87c),
	.w6(32'hb69ae79e),
	.w7(32'h38ef7336),
	.w8(32'hba146fa3),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5cafb),
	.w1(32'h3919d80e),
	.w2(32'hb9e24a5d),
	.w3(32'h3a055ba0),
	.w4(32'h38c6a73e),
	.w5(32'hba15f97b),
	.w6(32'h3a1bbb05),
	.w7(32'h396c4c45),
	.w8(32'hba2d2b56),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h358c855e),
	.w1(32'hb6c80e6b),
	.w2(32'hb6eaa3c1),
	.w3(32'h360b1388),
	.w4(32'hb7516d87),
	.w5(32'hb699a194),
	.w6(32'h370f81fe),
	.w7(32'hb72ca492),
	.w8(32'hb6ab7ea7),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c301b2),
	.w1(32'h396bc23a),
	.w2(32'hb99a69e3),
	.w3(32'h39d68f70),
	.w4(32'h39202130),
	.w5(32'hb9e4f45e),
	.w6(32'h39f7c0fe),
	.w7(32'h3963eb80),
	.w8(32'hba04728f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c525e),
	.w1(32'h39902ff7),
	.w2(32'hb9ace87f),
	.w3(32'h39aae0c1),
	.w4(32'h398fbdda),
	.w5(32'hb99b2bba),
	.w6(32'h397d13ba),
	.w7(32'h3969f973),
	.w8(32'hba019d3d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fe4ac),
	.w1(32'hb8bd5073),
	.w2(32'hb956a844),
	.w3(32'h3a017e3e),
	.w4(32'hb94f76f3),
	.w5(32'hb93d628b),
	.w6(32'h3a36c849),
	.w7(32'h393595b8),
	.w8(32'hb864ed67),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957c4e5),
	.w1(32'h398a2c72),
	.w2(32'hb9d84104),
	.w3(32'hb8a777ec),
	.w4(32'h38d0787c),
	.w5(32'hba25d73b),
	.w6(32'h3808f330),
	.w7(32'h38ff5aee),
	.w8(32'hba40c506),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0eecd4),
	.w1(32'h370ce435),
	.w2(32'hb9628816),
	.w3(32'hb991daca),
	.w4(32'hb85b7ac0),
	.w5(32'hb92d519f),
	.w6(32'hb993c513),
	.w7(32'h3693d06a),
	.w8(32'hb965808b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38248005),
	.w1(32'h390a7f65),
	.w2(32'h39bbf5bd),
	.w3(32'hb902b349),
	.w4(32'hb91cb347),
	.w5(32'h38405cbe),
	.w6(32'h37c83c3d),
	.w7(32'hb8ba2d0a),
	.w8(32'hb9826a8c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81af633),
	.w1(32'h39acbeab),
	.w2(32'h390c700d),
	.w3(32'h391d5736),
	.w4(32'h39519f12),
	.w5(32'hb75e1817),
	.w6(32'h39c22c2c),
	.w7(32'h39809501),
	.w8(32'hb8f83bcc),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b4344),
	.w1(32'hb9a538c6),
	.w2(32'h32895231),
	.w3(32'hba16784e),
	.w4(32'hb9a1e0f9),
	.w5(32'hb8a20ca4),
	.w6(32'hba124289),
	.w7(32'hb990af1f),
	.w8(32'hb965858b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90481d2),
	.w1(32'hb7c7ea4f),
	.w2(32'h380ca88b),
	.w3(32'hb8b74f25),
	.w4(32'hb65b03dd),
	.w5(32'h3801ba2e),
	.w6(32'hb901be30),
	.w7(32'hb6a4d8f6),
	.w8(32'hb74b0618),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e06745),
	.w1(32'hb82c4062),
	.w2(32'hb9729cc7),
	.w3(32'h399335cf),
	.w4(32'hb946198c),
	.w5(32'hb96703a5),
	.w6(32'h39481da7),
	.w7(32'h376ab527),
	.w8(32'hb8b881da),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a88fe8),
	.w1(32'hb775073d),
	.w2(32'hb77b391a),
	.w3(32'hb7ea065f),
	.w4(32'hb628ba5a),
	.w5(32'hb726c2ce),
	.w6(32'hb79b70e4),
	.w7(32'h3580e01b),
	.w8(32'hb79c4f67),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39550e85),
	.w1(32'hb8533b80),
	.w2(32'hb9980cf1),
	.w3(32'h396fbfb6),
	.w4(32'hb8823637),
	.w5(32'hb9cf01b1),
	.w6(32'h399722ec),
	.w7(32'h388edec2),
	.w8(32'hb9beec6e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3645d5c6),
	.w1(32'h37e45c5b),
	.w2(32'h37ca84db),
	.w3(32'h3737210a),
	.w4(32'h36e60c91),
	.w5(32'h37cd6b5c),
	.w6(32'h36ca0cc9),
	.w7(32'hb6fce2e5),
	.w8(32'h37a67bce),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c6e96),
	.w1(32'h390a54c1),
	.w2(32'hb7b11787),
	.w3(32'hb87d874f),
	.w4(32'h386c1f1e),
	.w5(32'hb9027c04),
	.w6(32'h383b1123),
	.w7(32'h39213444),
	.w8(32'hb96a06fd),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e37fea),
	.w1(32'hb8a26fa2),
	.w2(32'h378f303a),
	.w3(32'hb8c0857e),
	.w4(32'hb68055a1),
	.w5(32'h386cd548),
	.w6(32'hb8c9f57c),
	.w7(32'hb8815468),
	.w8(32'h3897ad16),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395db595),
	.w1(32'hb824dc2d),
	.w2(32'hb7dff10e),
	.w3(32'h395622b8),
	.w4(32'h37670684),
	.w5(32'h388f309b),
	.w6(32'h3952b890),
	.w7(32'hb77b492f),
	.w8(32'h388e9add),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb742cba4),
	.w1(32'hb6060848),
	.w2(32'hb792a4ed),
	.w3(32'hb69a5175),
	.w4(32'hb75efd4f),
	.w5(32'hb7c2701b),
	.w6(32'hb80e486c),
	.w7(32'hb8082fab),
	.w8(32'h37090789),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382f6ae0),
	.w1(32'hb84f2b0f),
	.w2(32'hb7e79458),
	.w3(32'h388b7f5a),
	.w4(32'h35f0984a),
	.w5(32'hb62971e7),
	.w6(32'h38563d5b),
	.w7(32'h37309367),
	.w8(32'hb8510d92),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d58c8),
	.w1(32'h39698242),
	.w2(32'h39ba2620),
	.w3(32'hb9d85675),
	.w4(32'h370ebd2a),
	.w5(32'h384f696a),
	.w6(32'hb9df4f1b),
	.w7(32'h38d76b6e),
	.w8(32'hb93562ce),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb533a),
	.w1(32'h39ab12a7),
	.w2(32'hba4e3ca1),
	.w3(32'h39634117),
	.w4(32'h38c9dcf0),
	.w5(32'hba93af1c),
	.w6(32'h3a3f819b),
	.w7(32'h39cc0a9a),
	.w8(32'hba6ab746),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb706e9cd),
	.w1(32'hb8021ee2),
	.w2(32'hb7bb5c7a),
	.w3(32'h37f8561e),
	.w4(32'h36e4993d),
	.w5(32'h38b7ca80),
	.w6(32'h37428f00),
	.w7(32'h38b31ec9),
	.w8(32'h38bb94fb),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb819b3d1),
	.w1(32'h399c225e),
	.w2(32'hb830f788),
	.w3(32'h3903e077),
	.w4(32'h39951d42),
	.w5(32'hb99da004),
	.w6(32'h3966e1b2),
	.w7(32'h3990180d),
	.w8(32'hb9e7eec8),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f4e375),
	.w1(32'h38b342d8),
	.w2(32'hb7ded12c),
	.w3(32'h38948d7e),
	.w4(32'h38531cdf),
	.w5(32'hb80d1aee),
	.w6(32'h37e7fb20),
	.w7(32'h3869046b),
	.w8(32'hb82c390f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae6692),
	.w1(32'hb87d9bcd),
	.w2(32'hb982c20c),
	.w3(32'h39baf227),
	.w4(32'hb907b1cd),
	.w5(32'hba064681),
	.w6(32'h39db272b),
	.w7(32'h39406fc3),
	.w8(32'hba0a95b3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c917fd),
	.w1(32'hb69ffc5c),
	.w2(32'hb9e54df9),
	.w3(32'h39cb72bc),
	.w4(32'hb8856e5c),
	.w5(32'hba0507d1),
	.w6(32'h39d10183),
	.w7(32'h37661255),
	.w8(32'hba0666ff),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a283710),
	.w1(32'h39aaa3f2),
	.w2(32'hb899fcf8),
	.w3(32'h3a4a7ec2),
	.w4(32'h3900e9bc),
	.w5(32'hb99bc17b),
	.w6(32'h3a80a6d8),
	.w7(32'h39893395),
	.w8(32'hb94502af),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37688c70),
	.w1(32'h3807bbc0),
	.w2(32'h38510cd3),
	.w3(32'h378f1a72),
	.w4(32'h385a3452),
	.w5(32'h38ad7c60),
	.w6(32'h3878f55b),
	.w7(32'hb6e7d82d),
	.w8(32'h3908aa0b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8608413),
	.w1(32'hb897bc7a),
	.w2(32'h3824528a),
	.w3(32'hb875473e),
	.w4(32'hb6e12960),
	.w5(32'hb8d0ec3e),
	.w6(32'h38557720),
	.w7(32'h3882af64),
	.w8(32'hb83308e9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3623883e),
	.w1(32'h35eb2555),
	.w2(32'h35dbf89d),
	.w3(32'h36da4001),
	.w4(32'h365c3be8),
	.w5(32'h36e48919),
	.w6(32'hb481dfb5),
	.w7(32'hb68ff546),
	.w8(32'h36a60770),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391bb0bf),
	.w1(32'h3731eb92),
	.w2(32'hb8f8a0bd),
	.w3(32'h393012c7),
	.w4(32'h36a75a1e),
	.w5(32'hb9093c6a),
	.w6(32'h39794eb3),
	.w7(32'h389fe80f),
	.w8(32'hb8eba912),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37607c46),
	.w1(32'hb8252377),
	.w2(32'h36eb2f8b),
	.w3(32'h33f6a821),
	.w4(32'hb80c6172),
	.w5(32'h37ca5161),
	.w6(32'hb80cf174),
	.w7(32'hb8451b65),
	.w8(32'hb6cd0b48),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392fdb20),
	.w1(32'h38fa5f12),
	.w2(32'hb926a15c),
	.w3(32'h39934a08),
	.w4(32'h38c7b58b),
	.w5(32'hb98122f1),
	.w6(32'h39bd322a),
	.w7(32'h39646638),
	.w8(32'hb980ab5f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d6ceef),
	.w1(32'hb61c4e7d),
	.w2(32'hb6970f40),
	.w3(32'hb6ec7f4b),
	.w4(32'h35d2aa18),
	.w5(32'h3598d1ee),
	.w6(32'h3526c6af),
	.w7(32'hb6cd6237),
	.w8(32'hb51a9874),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dbf642),
	.w1(32'h37241ced),
	.w2(32'h37ff6ebc),
	.w3(32'h37e40675),
	.w4(32'h371bb1fe),
	.w5(32'h37c292b2),
	.w6(32'h37ed8b2f),
	.w7(32'h381efefe),
	.w8(32'h37f276a2),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e4e2b5),
	.w1(32'hb81896e2),
	.w2(32'hb915e040),
	.w3(32'hb85418ff),
	.w4(32'h37a79f40),
	.w5(32'hb9287223),
	.w6(32'h386f2ad4),
	.w7(32'h38ea53b2),
	.w8(32'hb978138d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37492393),
	.w1(32'hb8145698),
	.w2(32'hb9f0f245),
	.w3(32'hb7c75db9),
	.w4(32'hb7ebcc21),
	.w5(32'hb9fd23c3),
	.w6(32'h38ff0bf7),
	.w7(32'h3a00713c),
	.w8(32'hb9ea3735),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb03dc),
	.w1(32'hb83a84b9),
	.w2(32'hb9511710),
	.w3(32'h392dc82e),
	.w4(32'hb8a2effb),
	.w5(32'hb93502ea),
	.w6(32'h38e896bd),
	.w7(32'hb94d660d),
	.w8(32'hb92614a0),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a5c87),
	.w1(32'hb9122267),
	.w2(32'hb91d4523),
	.w3(32'hb86600d1),
	.w4(32'hb921c229),
	.w5(32'hb917eec4),
	.w6(32'h3856afee),
	.w7(32'hb889d9c5),
	.w8(32'hb8d12a8a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab542e1),
	.w1(32'h399206a2),
	.w2(32'hba15bebb),
	.w3(32'h3ad37e9c),
	.w4(32'h38477410),
	.w5(32'hba2ef3c2),
	.w6(32'h3afd3c57),
	.w7(32'h3a7abda7),
	.w8(32'hb958fdad),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f6771),
	.w1(32'h39e983f1),
	.w2(32'hb6c9beef),
	.w3(32'hb9fe5ea6),
	.w4(32'h3892b87b),
	.w5(32'hb9a613d8),
	.w6(32'hba21c747),
	.w7(32'h38d6f987),
	.w8(32'hba02dabd),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb792c9d8),
	.w1(32'hb815af91),
	.w2(32'h37a28fde),
	.w3(32'h38833a84),
	.w4(32'h373b045b),
	.w5(32'h382e5cd7),
	.w6(32'h3786c22a),
	.w7(32'hb85d387d),
	.w8(32'h381054be),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63c3708),
	.w1(32'hb654d4db),
	.w2(32'h37116b40),
	.w3(32'h356efb9b),
	.w4(32'hb65644bb),
	.w5(32'h373dc1af),
	.w6(32'h3754d1b1),
	.w7(32'h376c5f31),
	.w8(32'h372a974b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77a327b),
	.w1(32'h381d3c1b),
	.w2(32'h38cd203d),
	.w3(32'hb7e21b50),
	.w4(32'h37afdf6b),
	.w5(32'h38417dd7),
	.w6(32'h38996c2c),
	.w7(32'h391321c2),
	.w8(32'h38b41efc),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370e1a8d),
	.w1(32'hb6498baa),
	.w2(32'h362a07e7),
	.w3(32'h3557c988),
	.w4(32'hb6132029),
	.w5(32'hb507ef78),
	.w6(32'hb71c339c),
	.w7(32'hb71c65cd),
	.w8(32'hb5a15f18),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb852f60e),
	.w1(32'hb81858e8),
	.w2(32'hb63001da),
	.w3(32'hb82ffeff),
	.w4(32'hb8b06f7f),
	.w5(32'h3718e5f2),
	.w6(32'h37897d04),
	.w7(32'h3751bb7a),
	.w8(32'h388b78a5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3817be01),
	.w1(32'hb7ccc703),
	.w2(32'hb82d71b7),
	.w3(32'hb933255a),
	.w4(32'hb8caaff4),
	.w5(32'hb9808184),
	.w6(32'hb7aa72f2),
	.w7(32'h386156e6),
	.w8(32'hb91c3f70),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e242ec),
	.w1(32'h39c8ae1c),
	.w2(32'hb985d1b7),
	.w3(32'h39c2a2f1),
	.w4(32'h397217e4),
	.w5(32'hba0577b4),
	.w6(32'h39b8ff20),
	.w7(32'h39987801),
	.w8(32'hba0ef523),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c77cd0),
	.w1(32'hb6e8cf65),
	.w2(32'h377f68af),
	.w3(32'hb80e2cab),
	.w4(32'h381c5b44),
	.w5(32'hb82c1303),
	.w6(32'hb6e008bd),
	.w7(32'h389457f1),
	.w8(32'hb873a390),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2f3b3),
	.w1(32'h3985b5e7),
	.w2(32'hb9d0a757),
	.w3(32'h3a03d520),
	.w4(32'h398dd46c),
	.w5(32'hb9f7dac6),
	.w6(32'h3a1b86d8),
	.w7(32'h39e58adf),
	.w8(32'hba100372),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a0a305),
	.w1(32'h39754182),
	.w2(32'hb7b9f263),
	.w3(32'h394f9057),
	.w4(32'h396eedac),
	.w5(32'hb87e22dd),
	.w6(32'h39470ab5),
	.w7(32'h39c905ab),
	.w8(32'hb8fed98f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c21c9b),
	.w1(32'hb610e5aa),
	.w2(32'h363a3681),
	.w3(32'hb642f835),
	.w4(32'h35c4e8c2),
	.w5(32'h36db4c58),
	.w6(32'hb5cec2fc),
	.w7(32'hb615d84d),
	.w8(32'h3701fcc8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390de2c6),
	.w1(32'hb88c44de),
	.w2(32'hb8b7d5bc),
	.w3(32'h38eb9ca5),
	.w4(32'h3526bb5f),
	.w5(32'h37806562),
	.w6(32'h38b15820),
	.w7(32'hb8193e66),
	.w8(32'h381c950b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71c4695),
	.w1(32'hb633aaac),
	.w2(32'h370d5751),
	.w3(32'hb69e6150),
	.w4(32'h350e9d88),
	.w5(32'h3760e739),
	.w6(32'hb3d00122),
	.w7(32'hb64f19bc),
	.w8(32'h378dce61),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3960b85a),
	.w1(32'hb8c67208),
	.w2(32'hb9d62c5c),
	.w3(32'h38e6b5d8),
	.w4(32'hb8eea62b),
	.w5(32'hba053f6d),
	.w6(32'h3a0b4f6f),
	.w7(32'h3974519d),
	.w8(32'hb9f68144),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20a464),
	.w1(32'hb938324a),
	.w2(32'hb9872cac),
	.w3(32'hb9c5a8c1),
	.w4(32'hb9847f97),
	.w5(32'hb9a201cf),
	.w6(32'hb9d716c1),
	.w7(32'hb8f9d8e2),
	.w8(32'hb9b6438b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b681f1),
	.w1(32'h398edbe4),
	.w2(32'hb949538b),
	.w3(32'h3832632a),
	.w4(32'h393fece7),
	.w5(32'hb9bbfcf3),
	.w6(32'h38c11fb8),
	.w7(32'h39ad03a9),
	.w8(32'hb9f9a36c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb890e387),
	.w1(32'hb7492ee2),
	.w2(32'h38954cba),
	.w3(32'hb88db70d),
	.w4(32'hb7e7118a),
	.w5(32'h3889464a),
	.w6(32'hb8c7099e),
	.w7(32'hb7917c50),
	.w8(32'h3841eb0c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dde00f),
	.w1(32'h39be098a),
	.w2(32'hb902934b),
	.w3(32'h36204619),
	.w4(32'h3967cef9),
	.w5(32'hb9f9ede8),
	.w6(32'h3778c952),
	.w7(32'h39c1b6c1),
	.w8(32'hba1dfaef),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398adc48),
	.w1(32'h39047dd0),
	.w2(32'hb93525c8),
	.w3(32'h39bbe070),
	.w4(32'h384fd8f4),
	.w5(32'hb9673ba4),
	.w6(32'h3a07f33d),
	.w7(32'h392442dd),
	.w8(32'hb92c2385),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b1773b),
	.w1(32'h38d5df88),
	.w2(32'hba4353ed),
	.w3(32'h3995ee04),
	.w4(32'hb65729b5),
	.w5(32'hba7e1ffb),
	.w6(32'h39dabfae),
	.w7(32'h398acdfe),
	.w8(32'hba4fa97c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d48130),
	.w1(32'h36089ee0),
	.w2(32'h37ba75c2),
	.w3(32'h37de4d19),
	.w4(32'hb68945cc),
	.w5(32'h3762da55),
	.w6(32'h37343b66),
	.w7(32'h375382b9),
	.w8(32'h3706dceb),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37158f2c),
	.w1(32'h35ab7885),
	.w2(32'h35d1cbde),
	.w3(32'h37105fbe),
	.w4(32'h34cd9f38),
	.w5(32'hb669837d),
	.w6(32'h35ab63a4),
	.w7(32'h3564963c),
	.w8(32'hb6840916),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd1e3f),
	.w1(32'h3a0cb279),
	.w2(32'hb9e4c854),
	.w3(32'h38bc1d67),
	.w4(32'h3933afd4),
	.w5(32'hba33c05a),
	.w6(32'h391cffdd),
	.w7(32'h3a05fb91),
	.w8(32'hba29e8e7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aceeca),
	.w1(32'hb795457d),
	.w2(32'hba510d0a),
	.w3(32'h39a271e0),
	.w4(32'h378d9113),
	.w5(32'hba741689),
	.w6(32'h3a6e7799),
	.w7(32'h3a51d624),
	.w8(32'hba4b2faa),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c11a8),
	.w1(32'h39bdfb59),
	.w2(32'hb9b2bc22),
	.w3(32'h398343c9),
	.w4(32'h398f4b5c),
	.w5(32'hba0afb0b),
	.w6(32'h39d38ec9),
	.w7(32'h39bf4993),
	.w8(32'hba257985),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb653d4a6),
	.w1(32'hb98a28e0),
	.w2(32'hb893e82a),
	.w3(32'h38fcc60d),
	.w4(32'hb9848bfc),
	.w5(32'hb929d5b2),
	.w6(32'hb95d4180),
	.w7(32'hb9834e3b),
	.w8(32'h368021bd),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a032fc),
	.w1(32'h36a132c9),
	.w2(32'h378cbdc6),
	.w3(32'hb7cd934e),
	.w4(32'h36a62537),
	.w5(32'h3815156d),
	.w6(32'hb79bceab),
	.w7(32'h37cf28c2),
	.w8(32'h3843747e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36580bdc),
	.w1(32'hb7f6eadd),
	.w2(32'h373d7461),
	.w3(32'hb4e771f2),
	.w4(32'hb7ad3884),
	.w5(32'h375d0d41),
	.w6(32'h37b518d1),
	.w7(32'hb7657b1c),
	.w8(32'h380d26c2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd9542),
	.w1(32'hb786a480),
	.w2(32'hb9a1ae75),
	.w3(32'h39fbee59),
	.w4(32'hb9239a05),
	.w5(32'hb9809bab),
	.w6(32'h3a027643),
	.w7(32'hb8ac42bf),
	.w8(32'hb8a3739a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a637642),
	.w1(32'hb9e8df26),
	.w2(32'hba141d41),
	.w3(32'h3a3b6aaa),
	.w4(32'hb9eb2c58),
	.w5(32'hb9d4d580),
	.w6(32'h3a3d1fbb),
	.w7(32'h3867728b),
	.w8(32'hb970508c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b0dff),
	.w1(32'h39deac83),
	.w2(32'hb9d26358),
	.w3(32'h3a81028b),
	.w4(32'h39115837),
	.w5(32'hb9f596e8),
	.w6(32'h3a55b11b),
	.w7(32'h39b8799d),
	.w8(32'hb93fac3d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b12fe7),
	.w1(32'hb76ab2f6),
	.w2(32'hb8e6231d),
	.w3(32'hb99697ff),
	.w4(32'hb82bf508),
	.w5(32'hb8fa9747),
	.w6(32'hb9632e67),
	.w7(32'h389876e2),
	.w8(32'hb91f2023),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85e9765),
	.w1(32'h3980becb),
	.w2(32'hb9a181e0),
	.w3(32'h37f36a46),
	.w4(32'h3902fc83),
	.w5(32'hba0270e3),
	.w6(32'h388fe985),
	.w7(32'h398a9070),
	.w8(32'hb9f95534),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7140d51),
	.w1(32'hb45a292c),
	.w2(32'h35af0d56),
	.w3(32'hb6bbebfa),
	.w4(32'hb5a83b54),
	.w5(32'hb44c6298),
	.w6(32'hb6c6c35a),
	.w7(32'hb6fb4e77),
	.w8(32'hb5a98172),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a2ea46),
	.w1(32'hb671a9b5),
	.w2(32'hb49dd82b),
	.w3(32'hb69ee621),
	.w4(32'hb6144d18),
	.w5(32'hb606b58c),
	.w6(32'hb6fe1565),
	.w7(32'hb6836268),
	.w8(32'h36a1ef13),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71f6784),
	.w1(32'hb7718aa9),
	.w2(32'h37806d37),
	.w3(32'hb7ac3f00),
	.w4(32'hb738d86f),
	.w5(32'h3708add2),
	.w6(32'hb74af931),
	.w7(32'h36057a4f),
	.w8(32'h38097a96),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6249cb7),
	.w1(32'h370b48c0),
	.w2(32'h36d61ee4),
	.w3(32'h36679f98),
	.w4(32'h3745273f),
	.w5(32'h372dc5a8),
	.w6(32'h36884660),
	.w7(32'h36f1700c),
	.w8(32'h374e5f40),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a62183),
	.w1(32'h380c6f64),
	.w2(32'h3717980c),
	.w3(32'hb822725c),
	.w4(32'hb65ec2d4),
	.w5(32'hb71059b9),
	.w6(32'hb7e02699),
	.w7(32'h3808466a),
	.w8(32'h36e90f61),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385dd0d2),
	.w1(32'hb892a4a9),
	.w2(32'hb9ac3557),
	.w3(32'h392f6809),
	.w4(32'hb8498ca4),
	.w5(32'hb9b0a081),
	.w6(32'h39d822d4),
	.w7(32'h39a2ee8c),
	.w8(32'hb9a77b14),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8857ebb),
	.w1(32'h3921fe66),
	.w2(32'hb986c835),
	.w3(32'h376e0ddd),
	.w4(32'h39038fb5),
	.w5(32'hb9be6d15),
	.w6(32'h39308d3b),
	.w7(32'h39953d70),
	.w8(32'hb9d11b42),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b1b9ae),
	.w1(32'h369e8e46),
	.w2(32'h36fc0ea3),
	.w3(32'h371e685d),
	.w4(32'h36ac3ca1),
	.w5(32'h37556d40),
	.w6(32'hb6d0fc27),
	.w7(32'hb6302d14),
	.w8(32'h370d3ee3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d96e2),
	.w1(32'h39023e2f),
	.w2(32'hba2c9836),
	.w3(32'h3a8de2a0),
	.w4(32'hb7d001c0),
	.w5(32'hba0ca42d),
	.w6(32'h3a8299ef),
	.w7(32'h3978f747),
	.w8(32'hb9874524),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbe708),
	.w1(32'h37fd9b73),
	.w2(32'hb986602a),
	.w3(32'h39d63f18),
	.w4(32'hb8b0fe6a),
	.w5(32'hb9613019),
	.w6(32'h39da85f8),
	.w7(32'h3839225e),
	.w8(32'hb8e6f3f1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371dd41a),
	.w1(32'h37c02d1e),
	.w2(32'h37d6baba),
	.w3(32'h371f1f98),
	.w4(32'h3798563c),
	.w5(32'h3805f117),
	.w6(32'h37c15a8c),
	.w7(32'h377e5b5a),
	.w8(32'h37b019a0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d32f07),
	.w1(32'hb794ffee),
	.w2(32'hb954d9e3),
	.w3(32'h39aa4e15),
	.w4(32'hb8afbb5d),
	.w5(32'hb93d32a4),
	.w6(32'h39a75c0e),
	.w7(32'h388c4fdc),
	.w8(32'hb8d05fad),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389a5d7f),
	.w1(32'h38924031),
	.w2(32'h379257bc),
	.w3(32'h386f6ef7),
	.w4(32'h386b483b),
	.w5(32'hb50029cb),
	.w6(32'h37c6baf4),
	.w7(32'h377779ce),
	.w8(32'hb6d165f8),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b6121a),
	.w1(32'h38903919),
	.w2(32'h3814a78d),
	.w3(32'hb85647b0),
	.w4(32'h3800a77a),
	.w5(32'hb7000e9a),
	.w6(32'hb8543f9a),
	.w7(32'hb72746d3),
	.w8(32'hb64a6bde),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36db3c6d),
	.w1(32'h374b8625),
	.w2(32'h37849e4c),
	.w3(32'h36a979e5),
	.w4(32'h3741a443),
	.w5(32'h3789b33d),
	.w6(32'hb72725bc),
	.w7(32'hb71fa981),
	.w8(32'h3699e43a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b0278a),
	.w1(32'hb631c945),
	.w2(32'h3695a2b9),
	.w3(32'h36eb095c),
	.w4(32'hb6cdf7cc),
	.w5(32'h3659f181),
	.w6(32'hb6e22414),
	.w7(32'hb79e5d07),
	.w8(32'h36ecf896),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ed8fe),
	.w1(32'h377ed5b6),
	.w2(32'hb87aac53),
	.w3(32'hb84748af),
	.w4(32'h370396ab),
	.w5(32'hb8b102af),
	.w6(32'hb895f44c),
	.w7(32'hb582a5da),
	.w8(32'hb92ec521),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02c3b7),
	.w1(32'h39361359),
	.w2(32'hb98c99ed),
	.w3(32'h3a07ed45),
	.w4(32'h38c8fade),
	.w5(32'hb9f6b188),
	.w6(32'h3a30551c),
	.w7(32'h3990a5db),
	.w8(32'hb9ad7b37),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397566d5),
	.w1(32'h3737016b),
	.w2(32'hb97f7162),
	.w3(32'h399cadb1),
	.w4(32'hb8abf710),
	.w5(32'hb99e2697),
	.w6(32'h39d498c7),
	.w7(32'h389ab6c9),
	.w8(32'hb9579fad),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc043c),
	.w1(32'h37dcb4ae),
	.w2(32'hb9451bd0),
	.w3(32'h39baee56),
	.w4(32'hb89bdae9),
	.w5(32'hb9b01057),
	.w6(32'h39b91a7c),
	.w7(32'h390e7299),
	.w8(32'hb98fcb07),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35381199),
	.w1(32'h379629a6),
	.w2(32'h37d334a6),
	.w3(32'hb6956a90),
	.w4(32'h37bd3f82),
	.w5(32'h37f6725e),
	.w6(32'hb699dc7a),
	.w7(32'h36521486),
	.w8(32'h378eb0ff),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70a1808),
	.w1(32'hb5fab120),
	.w2(32'h36f979cc),
	.w3(32'hb5511f79),
	.w4(32'hafa48160),
	.w5(32'h370d63c5),
	.w6(32'hb6978cc8),
	.w7(32'hb69b3b89),
	.w8(32'h36e5a8a3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3617f3ca),
	.w1(32'hb5867854),
	.w2(32'hb6ca0176),
	.w3(32'hb77ccf3e),
	.w4(32'hb7ee36ff),
	.w5(32'hb6cc2f03),
	.w6(32'h379fa3b0),
	.w7(32'hb7d34869),
	.w8(32'hb65a7b95),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3524eaf8),
	.w1(32'hb51d6743),
	.w2(32'h368020e5),
	.w3(32'hb5a775c8),
	.w4(32'hb5c157c4),
	.w5(32'h36d39998),
	.w6(32'hb6a3f7a6),
	.w7(32'hb65f9f16),
	.w8(32'h36896bba),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b287c),
	.w1(32'hb7927141),
	.w2(32'hb97ba4a9),
	.w3(32'h399b5b5d),
	.w4(32'h373953a2),
	.w5(32'hb9b017d2),
	.w6(32'h39c4de5b),
	.w7(32'h395f3363),
	.w8(32'hb9850ef0),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a7a233),
	.w1(32'h36fd4979),
	.w2(32'h386dd055),
	.w3(32'hb80711bf),
	.w4(32'hb7dacac3),
	.w5(32'h384fcc2d),
	.w6(32'h378d5e5e),
	.w7(32'h38b0347d),
	.w8(32'h37db1d62),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381ba2d6),
	.w1(32'hb79ad525),
	.w2(32'h382290ca),
	.w3(32'h382ba88f),
	.w4(32'h367f9e51),
	.w5(32'h38dbe616),
	.w6(32'h3752aa13),
	.w7(32'hb6104bb8),
	.w8(32'h38b4c4f8),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85e38f7),
	.w1(32'h38715562),
	.w2(32'hb50ccccc),
	.w3(32'hb83f1a53),
	.w4(32'h385a9f23),
	.w5(32'h3791a928),
	.w6(32'h3721efc7),
	.w7(32'h38d18ea8),
	.w8(32'h37f84b5a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cfcc32),
	.w1(32'h377bae9a),
	.w2(32'hb785e3ad),
	.w3(32'h37cbe3b9),
	.w4(32'h3814dcd7),
	.w5(32'hb6c2c852),
	.w6(32'h38a0b8c9),
	.w7(32'h38b5d68e),
	.w8(32'h335efe44),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38682095),
	.w1(32'h38027d1b),
	.w2(32'hb8e80862),
	.w3(32'h38a562f9),
	.w4(32'h36a1883d),
	.w5(32'hb956878a),
	.w6(32'h390c0df0),
	.w7(32'h391da761),
	.w8(32'hb923e8c1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7986ab7),
	.w1(32'h35ff1e7b),
	.w2(32'h37010c8c),
	.w3(32'hb6f0ba31),
	.w4(32'hb4b1a48b),
	.w5(32'h36d5f40e),
	.w6(32'hb6d1af8a),
	.w7(32'h361e1806),
	.w8(32'h3796748d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a117263),
	.w1(32'hb8f8d303),
	.w2(32'hb9974120),
	.w3(32'h3989d18c),
	.w4(32'hb9915939),
	.w5(32'hba01da99),
	.w6(32'h39c11789),
	.w7(32'h3929ab0d),
	.w8(32'hb94c3d70),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83aac45),
	.w1(32'hb7a6c065),
	.w2(32'hb7c3588e),
	.w3(32'hb839db41),
	.w4(32'hb69d09d1),
	.w5(32'hb7b3a629),
	.w6(32'hb7e2a191),
	.w7(32'h3724ce67),
	.w8(32'hb71bac33),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f5590),
	.w1(32'hb9167d11),
	.w2(32'hb950494b),
	.w3(32'hb9a7beed),
	.w4(32'hb8f0d270),
	.w5(32'hb9302ad1),
	.w6(32'hb893a744),
	.w7(32'h39446a0d),
	.w8(32'hb972cb8d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule