module layer_8_featuremap_127(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87bc8e),
	.w1(32'h3bfd2960),
	.w2(32'h3c71aebe),
	.w3(32'hbca17034),
	.w4(32'hbc35b0ef),
	.w5(32'h3bc6e089),
	.w6(32'hbbde4d0f),
	.w7(32'hbbaeec93),
	.w8(32'h3c1d396a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b51a6d),
	.w1(32'h3b31059f),
	.w2(32'h3abdb398),
	.w3(32'hba670204),
	.w4(32'hb902aae2),
	.w5(32'hbac66ad8),
	.w6(32'h3b28192e),
	.w7(32'h3aff52fc),
	.w8(32'hba61e440),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23bcab),
	.w1(32'h3b8ceba9),
	.w2(32'h3b67d985),
	.w3(32'h3b23d1b0),
	.w4(32'h3bb001bb),
	.w5(32'h3b84933c),
	.w6(32'h3bae04a7),
	.w7(32'h3bdd0f15),
	.w8(32'h3b79aa44),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12e11a),
	.w1(32'h3abea258),
	.w2(32'h3b906967),
	.w3(32'h3a42780e),
	.w4(32'h3c44b084),
	.w5(32'h3c7a2d08),
	.w6(32'hbbdcada5),
	.w7(32'h3be005e9),
	.w8(32'h3c524c23),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d143b),
	.w1(32'h3ad3eb70),
	.w2(32'hb9bc9463),
	.w3(32'h3b46951b),
	.w4(32'h3b162c4c),
	.w5(32'hba6a12f4),
	.w6(32'h3b5daa67),
	.w7(32'h3b020e80),
	.w8(32'hbafcace2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50ab95),
	.w1(32'h3ad78240),
	.w2(32'hbc814e72),
	.w3(32'h3c4a157d),
	.w4(32'h3c4b6bcb),
	.w5(32'hb9dc28d4),
	.w6(32'h3bbfdb05),
	.w7(32'h3b91e2c3),
	.w8(32'hbbc572f7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb47561bc),
	.w1(32'h3859c1a8),
	.w2(32'h392578d7),
	.w3(32'hb78c83d4),
	.w4(32'h382ec8c5),
	.w5(32'h38f23528),
	.w6(32'hb817ed01),
	.w7(32'h372c7f49),
	.w8(32'h387a7cbf),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12b51d),
	.w1(32'h3b86eb3d),
	.w2(32'h3bf929ea),
	.w3(32'hbb90fc8c),
	.w4(32'h3a498ebf),
	.w5(32'h3bd4badb),
	.w6(32'hb99e928b),
	.w7(32'h3b9fa52d),
	.w8(32'h3bd7ee55),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce7252),
	.w1(32'h3bdd7b82),
	.w2(32'h3bccc8d2),
	.w3(32'h3ba51f8c),
	.w4(32'h3b9cfff7),
	.w5(32'h3b09a669),
	.w6(32'h3bc2788f),
	.w7(32'h3bc54641),
	.w8(32'h3b67cf7e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fc273),
	.w1(32'h3b353d28),
	.w2(32'h3c45ab80),
	.w3(32'hbc98fd6d),
	.w4(32'hbc00a706),
	.w5(32'h3bdeb708),
	.w6(32'hbc128435),
	.w7(32'h3b923d88),
	.w8(32'h3c4de79d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c141fd4),
	.w1(32'h3c9de4cd),
	.w2(32'h3c879b43),
	.w3(32'hbbaaaf7d),
	.w4(32'h3beadc71),
	.w5(32'h3c466907),
	.w6(32'hbbc0326c),
	.w7(32'hbaec5bf0),
	.w8(32'h3c308ba9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc391ec9),
	.w1(32'h3b246404),
	.w2(32'h3c48482c),
	.w3(32'hbcad0670),
	.w4(32'hbc451bc7),
	.w5(32'h3b32e1bc),
	.w6(32'hbb2f0233),
	.w7(32'hbb089864),
	.w8(32'hb99dee64),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba20941),
	.w1(32'hbb8b4ff0),
	.w2(32'hbb8d99a2),
	.w3(32'h3ae5b686),
	.w4(32'h3a812c3b),
	.w5(32'h3b55ae90),
	.w6(32'h3b791673),
	.w7(32'hbb7f41c2),
	.w8(32'h3b0e7c13),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb2fd0),
	.w1(32'h3b68bf7d),
	.w2(32'hbb83f643),
	.w3(32'h3b1acb1a),
	.w4(32'hbbc38ae1),
	.w5(32'hbbf52f55),
	.w6(32'h3b1c9281),
	.w7(32'hbbea7546),
	.w8(32'hba920582),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaf211),
	.w1(32'h3bba0516),
	.w2(32'h3a2882cb),
	.w3(32'hbc0f7347),
	.w4(32'hb9b594bf),
	.w5(32'hbbd7d4b3),
	.w6(32'hbaea2211),
	.w7(32'hbb29d2b8),
	.w8(32'hbbb8cee0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac17315),
	.w1(32'h3a2ee465),
	.w2(32'h39ae0f35),
	.w3(32'hbc2f6440),
	.w4(32'hbc8100f5),
	.w5(32'h3cb64d25),
	.w6(32'hbb8fbf60),
	.w7(32'h3cb72501),
	.w8(32'h3d300194),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa3fc3),
	.w1(32'h3cc281cc),
	.w2(32'h386f225d),
	.w3(32'hbbb10c7b),
	.w4(32'h3baeb245),
	.w5(32'hbb991235),
	.w6(32'hbc4f7f06),
	.w7(32'h3c9ac99f),
	.w8(32'h3ba832c5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd02dec5),
	.w1(32'hbbce587f),
	.w2(32'h3cebc48d),
	.w3(32'hbb3cb07e),
	.w4(32'h3cb1a0ab),
	.w5(32'hba974e90),
	.w6(32'h3bce8142),
	.w7(32'h3c7ca515),
	.w8(32'h3dc224a6),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf31d14),
	.w1(32'hbc5d6fed),
	.w2(32'h3d1e956b),
	.w3(32'hbda8c544),
	.w4(32'hbd00e3c9),
	.w5(32'hbc10ae83),
	.w6(32'hb933ae44),
	.w7(32'hbce44c80),
	.w8(32'h3d9e1bce),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd301d03),
	.w1(32'hbb18d9b3),
	.w2(32'h3c84fcca),
	.w3(32'h3c1eea0f),
	.w4(32'hbc520d1a),
	.w5(32'h3cfbb1a7),
	.w6(32'h3c71e0e5),
	.w7(32'h3c891857),
	.w8(32'h3c7af54f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb41770),
	.w1(32'h3c7f8419),
	.w2(32'hbb5ba7bc),
	.w3(32'hbc92619f),
	.w4(32'h3c0adebb),
	.w5(32'hbc9db810),
	.w6(32'h3c345ac8),
	.w7(32'hbc91d109),
	.w8(32'hbd3d92b1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9939ce),
	.w1(32'h3af1adff),
	.w2(32'hbcbc53a1),
	.w3(32'h3c6184cf),
	.w4(32'hbc23783a),
	.w5(32'hbae08587),
	.w6(32'h3bc350e0),
	.w7(32'hbcd89865),
	.w8(32'h3d6ef4c7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80f1ce),
	.w1(32'h3b26a99b),
	.w2(32'h3d764ac6),
	.w3(32'hbd2cc057),
	.w4(32'hbc86c7b6),
	.w5(32'h3d00859a),
	.w6(32'hba542bbf),
	.w7(32'hbcbbb8fa),
	.w8(32'h3c15e19a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05a3ff),
	.w1(32'h3b8fafa6),
	.w2(32'h3be53a76),
	.w3(32'h3aee6470),
	.w4(32'h3c21f81e),
	.w5(32'h3c03e247),
	.w6(32'hbc1d2c99),
	.w7(32'h3c622092),
	.w8(32'h3bf729f6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4f1bb),
	.w1(32'hbbe0d7cc),
	.w2(32'hbbb34df2),
	.w3(32'h3c16931d),
	.w4(32'h3c5be79a),
	.w5(32'h3aa250aa),
	.w6(32'h3bd0a4f9),
	.w7(32'h3b17d993),
	.w8(32'hbbdd6fff),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53cdea),
	.w1(32'h3bff9f6c),
	.w2(32'h3ce730f0),
	.w3(32'hbc6ef546),
	.w4(32'hbc26f021),
	.w5(32'hbbc3376e),
	.w6(32'h3a9fada6),
	.w7(32'h3c82ed25),
	.w8(32'hbc0fd73c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc850024),
	.w1(32'hbc55eaa8),
	.w2(32'h3ba6b43e),
	.w3(32'h3bb80ebc),
	.w4(32'h3b0a0bc4),
	.w5(32'h3c4dc8f8),
	.w6(32'hbbe3665f),
	.w7(32'hbabcdf3b),
	.w8(32'hbd1136d7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb53b9f),
	.w1(32'h3dfbf95a),
	.w2(32'h3c6357ac),
	.w3(32'hbd4689e4),
	.w4(32'h3bc30299),
	.w5(32'h3c9fc2a1),
	.w6(32'hbd4e8f79),
	.w7(32'hbdd0280e),
	.w8(32'hbcdedd17),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d21dcee),
	.w1(32'h3bf77fed),
	.w2(32'h3c0c6aea),
	.w3(32'hbca35bcb),
	.w4(32'hbb1086fa),
	.w5(32'h3bd6d7bd),
	.w6(32'hbb5d3c64),
	.w7(32'h3962e16e),
	.w8(32'hbc4dffec),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7743b3),
	.w1(32'hba2fb77e),
	.w2(32'h3c0e8644),
	.w3(32'h3c1707e7),
	.w4(32'hbc154b08),
	.w5(32'hbbf4872a),
	.w6(32'hbcb61def),
	.w7(32'h3b0edb27),
	.w8(32'hbcd49b5d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba604ea),
	.w1(32'h3c0d1437),
	.w2(32'h3ac6069a),
	.w3(32'hbba79eb4),
	.w4(32'hbb979b81),
	.w5(32'hbb5807a3),
	.w6(32'hbbac5f61),
	.w7(32'hba9da461),
	.w8(32'h3a9b8401),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bee6b),
	.w1(32'h3a6969a1),
	.w2(32'hbc20605f),
	.w3(32'hba1c0024),
	.w4(32'hbc8d4b2d),
	.w5(32'h3c1a4e57),
	.w6(32'h3bd46d57),
	.w7(32'hbd179c2c),
	.w8(32'h3b02e26b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c999e4b),
	.w1(32'hbc543c2b),
	.w2(32'h3a6f943f),
	.w3(32'hbc88f07e),
	.w4(32'h3c665049),
	.w5(32'hbc2660c8),
	.w6(32'hbca7b9d1),
	.w7(32'h3c4c2c6f),
	.w8(32'hbd51e056),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a777e),
	.w1(32'hbb117967),
	.w2(32'hbc0a150b),
	.w3(32'h3c8fb831),
	.w4(32'hbc163605),
	.w5(32'hb9963f99),
	.w6(32'h3c155ccb),
	.w7(32'h3b93c50d),
	.w8(32'h3c66c0bb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd936113),
	.w1(32'hbd66caac),
	.w2(32'h3bb2461e),
	.w3(32'h3a511d40),
	.w4(32'hbb00b962),
	.w5(32'hbc593ff6),
	.w6(32'h3cc03894),
	.w7(32'h3b66e002),
	.w8(32'hbc6c417a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52e7e0),
	.w1(32'h3ccbd400),
	.w2(32'h3cf7559d),
	.w3(32'hbc9ce6c9),
	.w4(32'hbc791f1a),
	.w5(32'hbc45f26f),
	.w6(32'hbbf141ef),
	.w7(32'hbb6e0cde),
	.w8(32'hbd515f7c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb9e913),
	.w1(32'h3c036fa7),
	.w2(32'h3c83f1ce),
	.w3(32'hbb8c74b3),
	.w4(32'hbc3a0d22),
	.w5(32'h3b520e8b),
	.w6(32'hbcf49264),
	.w7(32'hbc663991),
	.w8(32'hbcb9ae36),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbba7f2),
	.w1(32'h3bee4c1e),
	.w2(32'hbc1a8350),
	.w3(32'hbc050ebb),
	.w4(32'h3b2db2e9),
	.w5(32'hbb6525b3),
	.w6(32'hbd00427e),
	.w7(32'h3d084e20),
	.w8(32'hbb9aee6d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0580df),
	.w1(32'hba606394),
	.w2(32'hbafe7f67),
	.w3(32'h3c87faad),
	.w4(32'hbb2fd1c2),
	.w5(32'h3ba305e5),
	.w6(32'h3cb628ef),
	.w7(32'hbb41d5a8),
	.w8(32'h3d7a0bf0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc84bdb),
	.w1(32'hbd06bb49),
	.w2(32'h3c7b52fe),
	.w3(32'h3b4aad58),
	.w4(32'h3c0e136c),
	.w5(32'h3c621dc5),
	.w6(32'hbc55fe27),
	.w7(32'h3aed039b),
	.w8(32'hbc02b07c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7025f9),
	.w1(32'h3c8fe9bc),
	.w2(32'h3c3f62b5),
	.w3(32'hbc72eabf),
	.w4(32'hbc7e3a63),
	.w5(32'h3d19b591),
	.w6(32'hbcb17926),
	.w7(32'h3bd7e00d),
	.w8(32'h3d2621e7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e27783),
	.w1(32'h3c2e9120),
	.w2(32'h3c5fc8c7),
	.w3(32'hbc70dba7),
	.w4(32'h3b7e260b),
	.w5(32'h3b9cdc6c),
	.w6(32'hbc23fdd9),
	.w7(32'hbcf64ee1),
	.w8(32'hbcec1b56),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d17fa00),
	.w1(32'h3c917bbe),
	.w2(32'hba3e2461),
	.w3(32'hbc3c17e4),
	.w4(32'h3a977f1c),
	.w5(32'hbc11bc19),
	.w6(32'hbc2e41b4),
	.w7(32'h3c9773d0),
	.w8(32'hbcf0afb8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe05b5a),
	.w1(32'h3ca07797),
	.w2(32'h3c1eb0fc),
	.w3(32'h3a8aae1a),
	.w4(32'hbb1ce863),
	.w5(32'h3bffba07),
	.w6(32'hbb933567),
	.w7(32'hbc2a7b59),
	.w8(32'h3adb3bc6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65d8b3),
	.w1(32'h3c8b1e35),
	.w2(32'h3cdb4e4e),
	.w3(32'hbcb7596d),
	.w4(32'hbc265d42),
	.w5(32'hbb9fb0a1),
	.w6(32'hbbc2a5d0),
	.w7(32'h3897f63f),
	.w8(32'hbc078bc3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcff767),
	.w1(32'hbc3aef9d),
	.w2(32'h3c2481e7),
	.w3(32'hbc8397ad),
	.w4(32'hbc1a75f1),
	.w5(32'hbc0c330f),
	.w6(32'hbc26dad3),
	.w7(32'hbc8a613b),
	.w8(32'hbcb1b701),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53168c),
	.w1(32'hbac27217),
	.w2(32'h3c3412a2),
	.w3(32'h3b280d89),
	.w4(32'h3b16b60c),
	.w5(32'h3ab00442),
	.w6(32'hbbad13d2),
	.w7(32'hbbe0226c),
	.w8(32'hbcb2ef49),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85e902),
	.w1(32'h3bf98442),
	.w2(32'h3caefd4d),
	.w3(32'hbbe1f1fb),
	.w4(32'hbc7d7e93),
	.w5(32'h3ae8f064),
	.w6(32'hbca80566),
	.w7(32'hbb2a2056),
	.w8(32'hbd213824),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca29211),
	.w1(32'h3c0cab0c),
	.w2(32'hbcfb094f),
	.w3(32'h3baf02b0),
	.w4(32'hbba0ed22),
	.w5(32'h3c61d3bf),
	.w6(32'h3ba24d73),
	.w7(32'hbcd27fcb),
	.w8(32'h3d023981),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf42c95),
	.w1(32'hbccb1a83),
	.w2(32'hbd2648c5),
	.w3(32'hbca0458e),
	.w4(32'hbcbacdb8),
	.w5(32'h3ce3171f),
	.w6(32'hbd03deea),
	.w7(32'hbc8e4ab1),
	.w8(32'h3d632277),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8a999e),
	.w1(32'hbd999ae9),
	.w2(32'hbc9d6d13),
	.w3(32'hbc222dd8),
	.w4(32'hbc96c3dd),
	.w5(32'hbc9c9f49),
	.w6(32'hbb83398c),
	.w7(32'h3a4eb45b),
	.w8(32'hbd205c68),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d51ff39),
	.w1(32'h3d2f0149),
	.w2(32'h3cabdd5c),
	.w3(32'hbc9c7941),
	.w4(32'h3c94d645),
	.w5(32'h3c58c409),
	.w6(32'h3c01f2b0),
	.w7(32'hbc02a906),
	.w8(32'hbce95976),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d50867b),
	.w1(32'h3d33444d),
	.w2(32'h3bcb703b),
	.w3(32'hbacee8a9),
	.w4(32'h3cd5d56d),
	.w5(32'hbcad7eab),
	.w6(32'hbcb51995),
	.w7(32'hbc094262),
	.w8(32'hbb174b04),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd18f51e),
	.w1(32'hbca560f7),
	.w2(32'h3c60678b),
	.w3(32'hbcdac936),
	.w4(32'hbca2caa9),
	.w5(32'hba29f30e),
	.w6(32'h3c55372f),
	.w7(32'hbb1f655d),
	.w8(32'h3c405af8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa39b1),
	.w1(32'h3abb70c9),
	.w2(32'hbb25f288),
	.w3(32'hbaabf57d),
	.w4(32'hbc8bdf9d),
	.w5(32'h3ab0adcd),
	.w6(32'h3a63204e),
	.w7(32'hbaa29476),
	.w8(32'hbce5e67a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd33d89f),
	.w1(32'hbcbd0ba2),
	.w2(32'hbc01e948),
	.w3(32'hbd35aeec),
	.w4(32'hbda137da),
	.w5(32'hbc1e8d74),
	.w6(32'hbca0fa13),
	.w7(32'hbc790899),
	.w8(32'h3d267421),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1cef17),
	.w1(32'hbcf571d5),
	.w2(32'h3c1e2680),
	.w3(32'h3c4047bb),
	.w4(32'h3bbf10e1),
	.w5(32'h3a97aaf2),
	.w6(32'hbba5fa40),
	.w7(32'h3b898d31),
	.w8(32'hbc9638f1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd478d),
	.w1(32'h3c9ab41c),
	.w2(32'h3c98ea55),
	.w3(32'hbc3d969c),
	.w4(32'h3b258a6f),
	.w5(32'hbc2f9c44),
	.w6(32'hbb609534),
	.w7(32'h3c55fb45),
	.w8(32'hbcac3f2f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa33311),
	.w1(32'h3c17364f),
	.w2(32'h3be8aa02),
	.w3(32'h3a9708ca),
	.w4(32'hb9ea3f5d),
	.w5(32'h3c180654),
	.w6(32'h3be1af27),
	.w7(32'hbc66bca8),
	.w8(32'h3b2a75bb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7235f4),
	.w1(32'hb92ea4ec),
	.w2(32'h3bae3be4),
	.w3(32'hbb9f7802),
	.w4(32'hbad684b4),
	.w5(32'hbc0629bc),
	.w6(32'hbaba1c44),
	.w7(32'hbc15f04e),
	.w8(32'h3bf1a5ad),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af498eb),
	.w1(32'hba845bfb),
	.w2(32'hbbf5f813),
	.w3(32'hbbdbeac0),
	.w4(32'hbb21dcae),
	.w5(32'hbb75e73f),
	.w6(32'hbc4f3a97),
	.w7(32'h3c8359d1),
	.w8(32'h3b9acc52),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb965c860),
	.w1(32'hb98ba3f5),
	.w2(32'hba89100c),
	.w3(32'h3b6059b1),
	.w4(32'h3c85f060),
	.w5(32'h3c1aa963),
	.w6(32'h3a9ae166),
	.w7(32'h3bc10ea7),
	.w8(32'hbb0e6574),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8599b8),
	.w1(32'h3c45fd38),
	.w2(32'hbc8aeca2),
	.w3(32'hbc1370de),
	.w4(32'hbd2acec9),
	.w5(32'h3a9cd820),
	.w6(32'hbba9210e),
	.w7(32'h3cc42562),
	.w8(32'h3d832499),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3be5e6),
	.w1(32'h3bcf636c),
	.w2(32'hbc84e9bf),
	.w3(32'h3aa316f6),
	.w4(32'hbc4b5df7),
	.w5(32'hbc01a60d),
	.w6(32'h3c314d6b),
	.w7(32'hbbb6a568),
	.w8(32'h3cf1ac92),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd81393),
	.w1(32'hbcc42962),
	.w2(32'h3c048452),
	.w3(32'hbb509acc),
	.w4(32'h3c53bf9e),
	.w5(32'hbbddb34f),
	.w6(32'hb90b4421),
	.w7(32'hbc6a5ce3),
	.w8(32'hbd14e230),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ae31b),
	.w1(32'h3ca819f0),
	.w2(32'h3c79cb0f),
	.w3(32'hbc1d532e),
	.w4(32'h3c4866a2),
	.w5(32'h3c361825),
	.w6(32'hbcacabae),
	.w7(32'h3c6e8129),
	.w8(32'hbcd332d8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0d05e0),
	.w1(32'h3c64ee91),
	.w2(32'h3ba6e16f),
	.w3(32'h3cdea2ff),
	.w4(32'hbc5910f5),
	.w5(32'hbc3cad4d),
	.w6(32'h3cd7e2fe),
	.w7(32'hbaea4b07),
	.w8(32'h3d1c8430),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87225e),
	.w1(32'hbd47b7fb),
	.w2(32'h3c028b83),
	.w3(32'hbc879f0a),
	.w4(32'hbc622d08),
	.w5(32'hbcdb6526),
	.w6(32'h3c89bc78),
	.w7(32'hbce42cf4),
	.w8(32'hbd50a09c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d30acd0),
	.w1(32'h3c16ce93),
	.w2(32'hbc666b42),
	.w3(32'hbc0f8c98),
	.w4(32'hbc17af1c),
	.w5(32'h3c8434d2),
	.w6(32'h3d0ab75e),
	.w7(32'hbca329dd),
	.w8(32'h3d12fe62),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f6fe9),
	.w1(32'h3cd94e2e),
	.w2(32'h3a61eb5f),
	.w3(32'hbbe86e8a),
	.w4(32'h3c90ee79),
	.w5(32'h3c4588b4),
	.w6(32'h3b83b8c7),
	.w7(32'hbc1e8f67),
	.w8(32'hbcd037eb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb46afe),
	.w1(32'h3caf9216),
	.w2(32'h3b0a0dca),
	.w3(32'hbb9f7c9b),
	.w4(32'h3b813c3e),
	.w5(32'hbc31a632),
	.w6(32'h3c63b818),
	.w7(32'hbcc14108),
	.w8(32'hbd6ffab7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90d176),
	.w1(32'h3d14e608),
	.w2(32'hbc7c93d4),
	.w3(32'h3b1e32c9),
	.w4(32'hbc303f9e),
	.w5(32'hbb3283ce),
	.w6(32'h3baba1bc),
	.w7(32'h3c84903b),
	.w8(32'hbc147eee),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0f00ef),
	.w1(32'h3c279164),
	.w2(32'h3bd95698),
	.w3(32'h3bd9b796),
	.w4(32'hbb67325e),
	.w5(32'h3b74c0d1),
	.w6(32'hbc84bd13),
	.w7(32'hbc52e023),
	.w8(32'h3b928d9e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45fb08),
	.w1(32'hbc09b481),
	.w2(32'h3c4806cd),
	.w3(32'hbc82c287),
	.w4(32'hb7b8a4fc),
	.w5(32'hbb43ddc4),
	.w6(32'h3cb23056),
	.w7(32'hbca7ec1b),
	.w8(32'hbd2745a4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e8201),
	.w1(32'h3c3dad98),
	.w2(32'h3bd7fb9a),
	.w3(32'hbc175acf),
	.w4(32'hbbda26d5),
	.w5(32'h3bc47e55),
	.w6(32'h3c9d6dd0),
	.w7(32'hbbfdd25f),
	.w8(32'h3c0baa3c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a2dd8),
	.w1(32'hbcd3f0ea),
	.w2(32'hbcbd775a),
	.w3(32'h3c4049ed),
	.w4(32'h3be900e8),
	.w5(32'hbba70355),
	.w6(32'hbc81c9e5),
	.w7(32'h3c2c7748),
	.w8(32'h3d2d41d3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9371cd),
	.w1(32'h3b793338),
	.w2(32'h3b5053aa),
	.w3(32'h3b723d80),
	.w4(32'h39ae655a),
	.w5(32'hba9a2e0b),
	.w6(32'hbaa14193),
	.w7(32'h3b411cda),
	.w8(32'hbbd1974b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b872ab7),
	.w1(32'h3cdacf93),
	.w2(32'h3c984c17),
	.w3(32'hbb65499e),
	.w4(32'h3b575830),
	.w5(32'h3be42f79),
	.w6(32'hbbf18290),
	.w7(32'hbb850b17),
	.w8(32'h3bc8a75a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1649ff),
	.w1(32'hbb3a056b),
	.w2(32'h3bf7f83f),
	.w3(32'hbce8b998),
	.w4(32'hbc8fd53c),
	.w5(32'h3b241857),
	.w6(32'hbc7c80d3),
	.w7(32'hbc72f889),
	.w8(32'h3b9963b8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe7e88),
	.w1(32'h3b9bf7b1),
	.w2(32'hbc07b70d),
	.w3(32'h3b762973),
	.w4(32'hbb8e55de),
	.w5(32'hbb98455b),
	.w6(32'h3bda53b4),
	.w7(32'h39f234ac),
	.w8(32'hbbb1c599),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cbfd9),
	.w1(32'hbca6bcf9),
	.w2(32'h3b4cb1da),
	.w3(32'hbb990e24),
	.w4(32'h385a67d8),
	.w5(32'h3b95bdfa),
	.w6(32'hbb328b33),
	.w7(32'h3b0bfb4c),
	.w8(32'h3bab3a8c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c117486),
	.w1(32'h3b8c184c),
	.w2(32'h3c03a6ad),
	.w3(32'hbac7663a),
	.w4(32'hbab90d66),
	.w5(32'h3c1eb992),
	.w6(32'hb9f0158b),
	.w7(32'hb9bb4d7a),
	.w8(32'hbc3dbcbf),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdf553),
	.w1(32'h3c95bf40),
	.w2(32'h3bcab691),
	.w3(32'hbc3d49f5),
	.w4(32'hbb7a9088),
	.w5(32'h3b9fc114),
	.w6(32'hbc269d69),
	.w7(32'hbb8bf741),
	.w8(32'hbbf81160),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03a5d7),
	.w1(32'h3c0b54a1),
	.w2(32'h3a050ba1),
	.w3(32'h3a03facc),
	.w4(32'h3c6c2b26),
	.w5(32'h3cb29076),
	.w6(32'h3b98c5e4),
	.w7(32'h3d09362f),
	.w8(32'h3cee6e9d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aa745),
	.w1(32'h3be05988),
	.w2(32'h3ccc7d2f),
	.w3(32'hbcd522dc),
	.w4(32'hbcc1da95),
	.w5(32'h3b030ede),
	.w6(32'h3bbc362a),
	.w7(32'hbc2881d3),
	.w8(32'h3d1f44e0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbd2a57),
	.w1(32'h3b9f1aad),
	.w2(32'h3ca1a164),
	.w3(32'hbcaca92f),
	.w4(32'h3bf3b4aa),
	.w5(32'h3c4b1491),
	.w6(32'hbc5578ec),
	.w7(32'h3b513f4f),
	.w8(32'h3c77b167),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96826c),
	.w1(32'hbc2ada3b),
	.w2(32'hbaa0c9e3),
	.w3(32'hbb6a7793),
	.w4(32'h3b2d12f5),
	.w5(32'h3bbf9b7d),
	.w6(32'hbb4ca10f),
	.w7(32'h3b0912cc),
	.w8(32'h3b03fb84),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ffa98),
	.w1(32'hbc218856),
	.w2(32'hba1b0a4f),
	.w3(32'h3c0d5cfc),
	.w4(32'hbb8e598f),
	.w5(32'hbb97f0bf),
	.w6(32'hbabe7dad),
	.w7(32'hbb654681),
	.w8(32'hbb710869),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f4da2),
	.w1(32'h3b047624),
	.w2(32'hb8393fed),
	.w3(32'hbb7d337f),
	.w4(32'hb892513b),
	.w5(32'hbb58a051),
	.w6(32'hbb1cae00),
	.w7(32'hb96b2d0c),
	.w8(32'h39bcbb14),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74f76b),
	.w1(32'hbabb8e71),
	.w2(32'h3bafac54),
	.w3(32'hbbded1f6),
	.w4(32'hb7ced8fa),
	.w5(32'h3bdbeebf),
	.w6(32'hbb8e0998),
	.w7(32'hbc511067),
	.w8(32'h3cf908da),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d939f),
	.w1(32'hbccbda91),
	.w2(32'hbbabed4b),
	.w3(32'h3adccaf4),
	.w4(32'hbbbd2b09),
	.w5(32'hbb94ac1a),
	.w6(32'h3c8f7323),
	.w7(32'hbc5ac836),
	.w8(32'h3b191a19),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f44e8),
	.w1(32'h3c2e7b0e),
	.w2(32'hbbb97881),
	.w3(32'hbbbea5f0),
	.w4(32'h39bb11b6),
	.w5(32'h3bf1a56f),
	.w6(32'h3c9433bf),
	.w7(32'hbc1b51de),
	.w8(32'h3bd4f38b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c8598),
	.w1(32'h3c7a114c),
	.w2(32'hbb73ddd5),
	.w3(32'h3c95da07),
	.w4(32'h3c740b95),
	.w5(32'h3b81fa30),
	.w6(32'h3ba77f5d),
	.w7(32'h393b5324),
	.w8(32'hbbd16049),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c7185),
	.w1(32'h3b2747e1),
	.w2(32'h3b28927d),
	.w3(32'hbbb8973b),
	.w4(32'hbac644cd),
	.w5(32'h39cce357),
	.w6(32'h3b8f0044),
	.w7(32'hbb9952a2),
	.w8(32'hbc444db0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94b8c2),
	.w1(32'h389d51e5),
	.w2(32'h3a335946),
	.w3(32'hbc2fa0a7),
	.w4(32'hbc0c287e),
	.w5(32'hbc10d219),
	.w6(32'hbbb151f0),
	.w7(32'h3a9b9b2f),
	.w8(32'hbc1b472b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49c254),
	.w1(32'hbc03725d),
	.w2(32'hbc1762aa),
	.w3(32'hbc9a9bda),
	.w4(32'hbcbb5ac1),
	.w5(32'hbcc1a1a5),
	.w6(32'hbc0f3765),
	.w7(32'hbcbb784e),
	.w8(32'hbcaa1327),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd5d965),
	.w1(32'h3d5c900c),
	.w2(32'h3cb3d87d),
	.w3(32'hbb9fdd65),
	.w4(32'h3babc304),
	.w5(32'h3be29634),
	.w6(32'hbc122549),
	.w7(32'h3ab84134),
	.w8(32'hbcb56161),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89e2e2),
	.w1(32'hbab2c5bf),
	.w2(32'h3bef4db7),
	.w3(32'h3bc6088d),
	.w4(32'hbb133189),
	.w5(32'hbb5c9856),
	.w6(32'hbc6b7ddf),
	.w7(32'h3a589670),
	.w8(32'h3c338649),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2356a),
	.w1(32'hbc1b0fdf),
	.w2(32'h3b8356fd),
	.w3(32'hbac55cef),
	.w4(32'h3b9ffea5),
	.w5(32'h3b439ec4),
	.w6(32'hbad535fa),
	.w7(32'h3b09d14e),
	.w8(32'hbaeca28f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf89ed),
	.w1(32'hbbe7af5c),
	.w2(32'h3c597509),
	.w3(32'h3bd4ffc8),
	.w4(32'h3c4b79ff),
	.w5(32'h3c785643),
	.w6(32'h3a021790),
	.w7(32'h3c11aaa6),
	.w8(32'hbc441b31),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd46865),
	.w1(32'hbc5f7116),
	.w2(32'hbbe8307c),
	.w3(32'h3c233dab),
	.w4(32'hba266608),
	.w5(32'h3ad51866),
	.w6(32'h3a962032),
	.w7(32'h39bc756e),
	.w8(32'h3b487963),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07547a),
	.w1(32'hbac8ef20),
	.w2(32'hbba0eaea),
	.w3(32'h3b5df766),
	.w4(32'hbb18fccf),
	.w5(32'hbbaf5d82),
	.w6(32'h3bb5c5f7),
	.w7(32'hbb9485f4),
	.w8(32'h3ac64d06),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b231f03),
	.w1(32'h3c04d9bd),
	.w2(32'hbbbc14a4),
	.w3(32'hbc0736d2),
	.w4(32'hbc0858a8),
	.w5(32'hbc0a7dfc),
	.w6(32'h3b4d919f),
	.w7(32'hbc744d22),
	.w8(32'hbc6d4d26),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc298bf8),
	.w1(32'hbbb668d9),
	.w2(32'hbb4ac140),
	.w3(32'h3b009117),
	.w4(32'h3c494d8b),
	.w5(32'hbba57036),
	.w6(32'h3b881842),
	.w7(32'h3b1d57ea),
	.w8(32'hbbdee261),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2858e),
	.w1(32'hbba3b35b),
	.w2(32'hbc0bc8f0),
	.w3(32'hbb980fe8),
	.w4(32'h3b7b86de),
	.w5(32'h3b74afa6),
	.w6(32'h3b438f09),
	.w7(32'h39c80576),
	.w8(32'hbab06796),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f37e9),
	.w1(32'hbafb8877),
	.w2(32'h3c5f7878),
	.w3(32'hbb0f0e49),
	.w4(32'h3b88c83c),
	.w5(32'h3c87cb62),
	.w6(32'h3a8c5ac7),
	.w7(32'hbc58837a),
	.w8(32'h3c0a7746),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc902a11),
	.w1(32'hbbaf67fc),
	.w2(32'h3c9662ee),
	.w3(32'h3a53af76),
	.w4(32'h394091da),
	.w5(32'hbba53910),
	.w6(32'hbc1d7697),
	.w7(32'h3959610f),
	.w8(32'hb838a778),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc805d07),
	.w1(32'hbc4332db),
	.w2(32'hba25c63b),
	.w3(32'h3c520e16),
	.w4(32'h3b4d019b),
	.w5(32'hbb5523b1),
	.w6(32'h3c156193),
	.w7(32'h3bb5c0d8),
	.w8(32'hbc3b8878),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadde51f),
	.w1(32'h3b8216fe),
	.w2(32'hbba407e0),
	.w3(32'h3bfbe15e),
	.w4(32'h3a9808a2),
	.w5(32'h3b91192e),
	.w6(32'h3b0e2d2a),
	.w7(32'hbc139294),
	.w8(32'hbc0ff2a6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc70f5),
	.w1(32'h3c2d60b7),
	.w2(32'h3b8d01b8),
	.w3(32'h3a6da9f2),
	.w4(32'h3a23bef4),
	.w5(32'h3ab5f038),
	.w6(32'hbb00bf34),
	.w7(32'hbb5ac369),
	.w8(32'hbc126fd9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee5c08),
	.w1(32'hbbe1f6b0),
	.w2(32'h3a326934),
	.w3(32'h3b3c099a),
	.w4(32'hb9863aed),
	.w5(32'hbc0f67e3),
	.w6(32'hbb93fb44),
	.w7(32'hbad1c456),
	.w8(32'hbc81af8b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9683d),
	.w1(32'hbba04353),
	.w2(32'hb8b98dee),
	.w3(32'h3adc5514),
	.w4(32'h3b9f0d5b),
	.w5(32'hbc17429d),
	.w6(32'h3b45b4c3),
	.w7(32'h3b6f4b50),
	.w8(32'hbbfbc26f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1fcdb),
	.w1(32'hbc16fe66),
	.w2(32'hbbc17845),
	.w3(32'h39f5a7a9),
	.w4(32'hbc17e905),
	.w5(32'hba024e05),
	.w6(32'h3b172efe),
	.w7(32'h3a5ac529),
	.w8(32'hba9b5491),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb193aa9),
	.w1(32'hb991328a),
	.w2(32'hbc4482dd),
	.w3(32'hbc09c86a),
	.w4(32'hbc9aee57),
	.w5(32'hbc8e176e),
	.w6(32'hbbc7b3a9),
	.w7(32'hbc90c371),
	.w8(32'hbc61b981),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a40b8),
	.w1(32'h3cbdf035),
	.w2(32'hbb632e41),
	.w3(32'hbc363363),
	.w4(32'hbb41a2d7),
	.w5(32'h3c3da73f),
	.w6(32'hbbbb719c),
	.w7(32'hbbd9110a),
	.w8(32'h3ca29993),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd4cc66),
	.w1(32'hbb958acd),
	.w2(32'h3a633768),
	.w3(32'hbbb9ce4b),
	.w4(32'hba1a4d6e),
	.w5(32'h3c2f02a7),
	.w6(32'h3aee67d0),
	.w7(32'h3b47d89c),
	.w8(32'h3cb4cf7a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbef3b4),
	.w1(32'hbd00d793),
	.w2(32'hbbeef108),
	.w3(32'h396af789),
	.w4(32'hbb857aed),
	.w5(32'hbb4dd01b),
	.w6(32'hbbf216e9),
	.w7(32'hbbf99a71),
	.w8(32'hbbdc41bc),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa1e3b),
	.w1(32'h3d4837de),
	.w2(32'h3bbf22a0),
	.w3(32'hbca45cbb),
	.w4(32'hbbcbc424),
	.w5(32'h3a1a09c0),
	.w6(32'hbc4f8601),
	.w7(32'hba1ecb02),
	.w8(32'hb9dee83a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58ef38),
	.w1(32'h3bbe8e15),
	.w2(32'hbbd2fe7f),
	.w3(32'h3b525705),
	.w4(32'hbbbcadf1),
	.w5(32'hbbe70964),
	.w6(32'h3a728e01),
	.w7(32'hbc7eda0f),
	.w8(32'hba1a1b30),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90ec6f),
	.w1(32'h3964cfd1),
	.w2(32'hbb4628cc),
	.w3(32'hbc5c370e),
	.w4(32'hbbddeab4),
	.w5(32'hbbf5bb48),
	.w6(32'h3b9339dd),
	.w7(32'hbba0f986),
	.w8(32'hbc005d5d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83f51a),
	.w1(32'hbbab7983),
	.w2(32'h3c522ea8),
	.w3(32'hbbf4ec66),
	.w4(32'h39eb61fc),
	.w5(32'hbb7236b6),
	.w6(32'h39c7375e),
	.w7(32'h3c04ffae),
	.w8(32'h3bc6ef54),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c038162),
	.w1(32'h3adb9c33),
	.w2(32'hbc013e1e),
	.w3(32'hbc0a0920),
	.w4(32'hbb9cd0ac),
	.w5(32'h3c457722),
	.w6(32'hbbbb8d06),
	.w7(32'h3bac40d8),
	.w8(32'h3cd0718b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ee5e1),
	.w1(32'hbc59220c),
	.w2(32'h3b1b17a6),
	.w3(32'h3be91683),
	.w4(32'h3991f3f5),
	.w5(32'hbacfd1f1),
	.w6(32'h3c87a095),
	.w7(32'h3b7b1b9f),
	.w8(32'hbbce285a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02c915),
	.w1(32'h3b83ac76),
	.w2(32'hbb9c52d1),
	.w3(32'h3b5ed71c),
	.w4(32'h3b975ff8),
	.w5(32'h3bc1ebb9),
	.w6(32'h3ad812f2),
	.w7(32'hbbf0bdc3),
	.w8(32'h3c6ed314),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0901b1),
	.w1(32'hbbd4f7db),
	.w2(32'h3bc88ca3),
	.w3(32'hbbe9e325),
	.w4(32'hbb958e1d),
	.w5(32'h3c24433b),
	.w6(32'hbb74fcaf),
	.w7(32'hbc8a1410),
	.w8(32'h3c2007c8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3951ea),
	.w1(32'hbd282d5c),
	.w2(32'hbba31d8b),
	.w3(32'h3cabc7e1),
	.w4(32'hbc251922),
	.w5(32'hbbb25645),
	.w6(32'h3c488fb7),
	.w7(32'hbbae144d),
	.w8(32'hbb9eaf02),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdc6bc),
	.w1(32'hbb7322a6),
	.w2(32'hbb11043d),
	.w3(32'hbb91b824),
	.w4(32'hbc439ecd),
	.w5(32'hbb0a7a22),
	.w6(32'hb72dd5da),
	.w7(32'hbb7a5c4e),
	.w8(32'hbc53bf7c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0497d7),
	.w1(32'hbcb77cf5),
	.w2(32'hbb7bdc53),
	.w3(32'hbb77abc0),
	.w4(32'hbc09fb81),
	.w5(32'hbbcd773b),
	.w6(32'hbc49b79d),
	.w7(32'hbca32a6a),
	.w8(32'hbc47126f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule