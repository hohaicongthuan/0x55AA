module layer_10_featuremap_453(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384746c1),
	.w1(32'h3842a85c),
	.w2(32'hb8a97398),
	.w3(32'h3951c8e8),
	.w4(32'hb8352636),
	.w5(32'hb90c894b),
	.w6(32'h397866b2),
	.w7(32'h386f7713),
	.w8(32'hb872c8c9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fad13c),
	.w1(32'h398f3aae),
	.w2(32'hb9cb5cca),
	.w3(32'h3a03b481),
	.w4(32'h3abaa552),
	.w5(32'h3a9acccf),
	.w6(32'h39427293),
	.w7(32'h39863cee),
	.w8(32'h3a6705d0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3975e12e),
	.w1(32'hb98b1ed0),
	.w2(32'hb99d5f46),
	.w3(32'h39351541),
	.w4(32'hb82c9368),
	.w5(32'h3913f993),
	.w6(32'hb6a33ad9),
	.w7(32'hb81620b9),
	.w8(32'hb936c3b1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2493f5),
	.w1(32'h3a34d576),
	.w2(32'h3a528ec2),
	.w3(32'hb97ff3c4),
	.w4(32'h3a055350),
	.w5(32'h39ae9a10),
	.w6(32'h398ec7de),
	.w7(32'h3a20b3c1),
	.w8(32'h3935e8bc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92bdb29),
	.w1(32'h38be8e54),
	.w2(32'h38a5aeea),
	.w3(32'hb6aa532c),
	.w4(32'hb789e2cd),
	.w5(32'hb779a989),
	.w6(32'h3921b913),
	.w7(32'hb65fe7a5),
	.w8(32'hb921a74c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3868bb78),
	.w1(32'hb98ab531),
	.w2(32'hb978deec),
	.w3(32'h392a0667),
	.w4(32'hb7d1a14c),
	.w5(32'hb985648e),
	.w6(32'hb870307a),
	.w7(32'h381d6d86),
	.w8(32'h381a619c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1df7d6),
	.w1(32'h3b5cfd52),
	.w2(32'h3afe82f7),
	.w3(32'h3b8d8ae3),
	.w4(32'h3b935705),
	.w5(32'hba4b7939),
	.w6(32'h3b7a8634),
	.w7(32'h3a4f912e),
	.w8(32'hbb6d240d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c5d6e),
	.w1(32'hbb44bd4e),
	.w2(32'hbb96fe2e),
	.w3(32'hbb7b644f),
	.w4(32'hbbd3dde7),
	.w5(32'hbb98b671),
	.w6(32'hbb012fcf),
	.w7(32'hbb252d9f),
	.w8(32'hba0d0636),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905d3d8),
	.w1(32'h39f016b5),
	.w2(32'h3a1aaec9),
	.w3(32'hb952a5e6),
	.w4(32'h39e31880),
	.w5(32'h3922c890),
	.w6(32'h38b1fc24),
	.w7(32'h3a007632),
	.w8(32'h3929e01e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9636197),
	.w1(32'hb8f6f9d0),
	.w2(32'hb946ac11),
	.w3(32'h3a10db7e),
	.w4(32'hb7ef3f04),
	.w5(32'hba6c0749),
	.w6(32'hb9afc869),
	.w7(32'hba9057a9),
	.w8(32'hbb32ba1b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73cc972),
	.w1(32'h396f96c3),
	.w2(32'h38fe329a),
	.w3(32'h38ad8d30),
	.w4(32'hb8065874),
	.w5(32'hb8f925f8),
	.w6(32'hb88ec2fb),
	.w7(32'h38d88d04),
	.w8(32'h37846027),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20ba62),
	.w1(32'h3b5a53e1),
	.w2(32'h3ad18b58),
	.w3(32'h3b9cbd52),
	.w4(32'h3bcfd64a),
	.w5(32'h399b4167),
	.w6(32'h3b91ce4c),
	.w7(32'h3b666a51),
	.w8(32'hbb55bfe5),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a216d34),
	.w1(32'h39a7bb69),
	.w2(32'h39ccbe41),
	.w3(32'h39fdc188),
	.w4(32'hba2d3a33),
	.w5(32'hbabf5834),
	.w6(32'h3913b64a),
	.w7(32'hbb0ab1a2),
	.w8(32'hbb6eca00),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a191f1e),
	.w1(32'hba7cda9f),
	.w2(32'hbac19b8d),
	.w3(32'h39fa7bc9),
	.w4(32'hba8e2a8f),
	.w5(32'h392c0ed0),
	.w6(32'h38988b51),
	.w7(32'hbaa86480),
	.w8(32'h388f805a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38be2665),
	.w1(32'h39af3fb6),
	.w2(32'hb9d21708),
	.w3(32'h3a0e3570),
	.w4(32'h3a9cf4ab),
	.w5(32'h3a8ba911),
	.w6(32'h39a76deb),
	.w7(32'h3a2e7f12),
	.w8(32'h3a1e1467),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc568d),
	.w1(32'hba9049b6),
	.w2(32'hbae3f3d5),
	.w3(32'h3a376893),
	.w4(32'hba0e8539),
	.w5(32'hb9c0f290),
	.w6(32'hbb2323df),
	.w7(32'hbb06c862),
	.w8(32'hba973548),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b4b665),
	.w1(32'hb9bd0799),
	.w2(32'hb9dae9e2),
	.w3(32'h39231a57),
	.w4(32'h387399fc),
	.w5(32'h392639ca),
	.w6(32'h3910924d),
	.w7(32'hb884c0c6),
	.w8(32'h38c52a1b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cfb05),
	.w1(32'h3aac8ff7),
	.w2(32'h3b03746b),
	.w3(32'h3a934aa9),
	.w4(32'hbb1bea59),
	.w5(32'hbba4c319),
	.w6(32'h3a11968e),
	.w7(32'hbabe141c),
	.w8(32'hbb4b63ba),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d3a2b),
	.w1(32'h38a1955a),
	.w2(32'h3a32e830),
	.w3(32'h3a069272),
	.w4(32'hbaa9c0b2),
	.w5(32'hbb2847e6),
	.w6(32'h39ffd3c4),
	.w7(32'hbaa47af9),
	.w8(32'hbb249348),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c0615),
	.w1(32'h36207bb0),
	.w2(32'h389d87d9),
	.w3(32'hb9b7e1eb),
	.w4(32'h385ac13a),
	.w5(32'h39a3e883),
	.w6(32'hb9e05062),
	.w7(32'hb987e1ec),
	.w8(32'h397e971e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6bd0a),
	.w1(32'h3911aa3f),
	.w2(32'h38fd355b),
	.w3(32'h38b13f89),
	.w4(32'h3820ea37),
	.w5(32'h392630c4),
	.w6(32'hb82502a0),
	.w7(32'h384a506b),
	.w8(32'h38b4a171),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c60d3),
	.w1(32'hb88fe874),
	.w2(32'h39abb547),
	.w3(32'h3a12511a),
	.w4(32'h380f03d0),
	.w5(32'h3a25a920),
	.w6(32'h3a1c673e),
	.w7(32'h387abd77),
	.w8(32'h39b6118a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8c9b0),
	.w1(32'h3aeee6d4),
	.w2(32'hbb30d393),
	.w3(32'h3a4bd973),
	.w4(32'h3b87191d),
	.w5(32'hbb467f45),
	.w6(32'hbb7cee45),
	.w7(32'hba369d6b),
	.w8(32'hbb675675),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381e62a8),
	.w1(32'hb9746315),
	.w2(32'hba070cf4),
	.w3(32'h38edbd2a),
	.w4(32'hbaa345dd),
	.w5(32'hbaef5908),
	.w6(32'h38e30a70),
	.w7(32'hba0eb6a2),
	.w8(32'hbabecae4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04e391),
	.w1(32'h3b106a16),
	.w2(32'h3a7566f2),
	.w3(32'h39270c7a),
	.w4(32'h3b2e2a26),
	.w5(32'h3b692d60),
	.w6(32'h3a8743b7),
	.w7(32'h3b3baf7b),
	.w8(32'h3b6fa609),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd8b36),
	.w1(32'hb8fb7f3f),
	.w2(32'h37d2527a),
	.w3(32'hb91e18e6),
	.w4(32'hba14a5c0),
	.w5(32'hb64f8f1a),
	.w6(32'hb9e97aab),
	.w7(32'hb9dafa91),
	.w8(32'hb9e0475b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906354c),
	.w1(32'hb9784401),
	.w2(32'hb8d1d3e0),
	.w3(32'hb7c9097e),
	.w4(32'hb862fa38),
	.w5(32'h390df921),
	.w6(32'h379abaf4),
	.w7(32'hb83ee3f5),
	.w8(32'h396d8670),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d4e62),
	.w1(32'hbafbca83),
	.w2(32'h3a3cfc0f),
	.w3(32'hba76774c),
	.w4(32'hbb0330bb),
	.w5(32'h3b26761a),
	.w6(32'hb9c4f186),
	.w7(32'hbb1122c7),
	.w8(32'h3baa0e58),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b9b03),
	.w1(32'h38ecca0f),
	.w2(32'hb967cd85),
	.w3(32'h384438ba),
	.w4(32'h3a0ff515),
	.w5(32'h3a21be33),
	.w6(32'h392dfa5a),
	.w7(32'h399a2d74),
	.w8(32'h397b657e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa438a7),
	.w1(32'h3a73bf77),
	.w2(32'h3b192b8d),
	.w3(32'h3a2ee746),
	.w4(32'h3a80c71b),
	.w5(32'h3b3f33fc),
	.w6(32'h3abe7ce6),
	.w7(32'h39cb3561),
	.w8(32'h3b52e3ca),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c09047),
	.w1(32'hb907cb24),
	.w2(32'hb97d42af),
	.w3(32'h38753955),
	.w4(32'h37c87806),
	.w5(32'h384e434c),
	.w6(32'h3919d3b0),
	.w7(32'hb616e5ad),
	.w8(32'h386077b4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e660db),
	.w1(32'h3954d6ec),
	.w2(32'h38a5ad9b),
	.w3(32'h394f3a24),
	.w4(32'h39b947df),
	.w5(32'hb7016652),
	.w6(32'h38bc226d),
	.w7(32'h399a3c84),
	.w8(32'h39547c69),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5854c6),
	.w1(32'hb8cc3a25),
	.w2(32'hb84028fe),
	.w3(32'h39dd0ddb),
	.w4(32'hb98aab97),
	.w5(32'hba73a9df),
	.w6(32'h3a373970),
	.w7(32'hba1db8b5),
	.w8(32'hba9c7a38),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9879120),
	.w1(32'hb94d7ea3),
	.w2(32'hba60a95e),
	.w3(32'h38defe42),
	.w4(32'h39d70843),
	.w5(32'h3a1ab020),
	.w6(32'h38f60c36),
	.w7(32'h3a4e3372),
	.w8(32'h3a64d794),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3744b124),
	.w1(32'hb75e6150),
	.w2(32'h380c5ae3),
	.w3(32'h3a4d834f),
	.w4(32'h3960a28b),
	.w5(32'h3975165e),
	.w6(32'h3a0a2148),
	.w7(32'hb9c66392),
	.w8(32'hba3176b7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5f12d),
	.w1(32'h3b227f0e),
	.w2(32'h3a3d8547),
	.w3(32'hb97d4995),
	.w4(32'h3a8a34d8),
	.w5(32'hbaa3c8df),
	.w6(32'h37628110),
	.w7(32'h3b065ddd),
	.w8(32'hb9cc7d10),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55953e),
	.w1(32'h3aa5d999),
	.w2(32'hbbb77621),
	.w3(32'h3a47bc19),
	.w4(32'h3c051599),
	.w5(32'h39cf9c0b),
	.w6(32'h393a0ef1),
	.w7(32'h3c32a57d),
	.w8(32'hbbb8fa15),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3889935f),
	.w1(32'h3b53b5d9),
	.w2(32'h3afa25be),
	.w3(32'h3a9230cc),
	.w4(32'h3bd13ffb),
	.w5(32'h3bdc2a35),
	.w6(32'h3a1ed897),
	.w7(32'h3b1684f0),
	.w8(32'h3b6e8be4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56bdbe),
	.w1(32'h3b77e56a),
	.w2(32'h3b8d2715),
	.w3(32'h3abcf26e),
	.w4(32'h3b366187),
	.w5(32'h3b8edce6),
	.w6(32'h3b108453),
	.w7(32'h3a25aa38),
	.w8(32'h3b5a3975),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f037e7),
	.w1(32'h3a2c1519),
	.w2(32'h3a4aa0ac),
	.w3(32'h3799a442),
	.w4(32'h3a9f6256),
	.w5(32'h3ab65ed9),
	.w6(32'h39727537),
	.w7(32'h3aa19e8f),
	.w8(32'h3a5ea7f2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899182c),
	.w1(32'h3982ac4e),
	.w2(32'h3816fa3c),
	.w3(32'h393a70d1),
	.w4(32'h394ff900),
	.w5(32'hb839c84d),
	.w6(32'h391642ae),
	.w7(32'hb87ec0c3),
	.w8(32'hb9c655ed),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2463a),
	.w1(32'hb8d80c34),
	.w2(32'h3854c148),
	.w3(32'h3978b68f),
	.w4(32'hb93f4b7c),
	.w5(32'hb90901c2),
	.w6(32'h38b5687d),
	.w7(32'hb91ab422),
	.w8(32'h38c1b736),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969ed70),
	.w1(32'hb8bfc643),
	.w2(32'hb8196a41),
	.w3(32'h39ec49cc),
	.w4(32'h39a91b77),
	.w5(32'hb8ad079a),
	.w6(32'h3824b64b),
	.w7(32'hb95c1348),
	.w8(32'hba34d227),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389d8820),
	.w1(32'h3adf1a74),
	.w2(32'h3aab39c9),
	.w3(32'h396d4bbf),
	.w4(32'hbb34f700),
	.w5(32'hbb277ad3),
	.w6(32'hbb1975bd),
	.w7(32'hbb77ce3d),
	.w8(32'hbb311b6e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51d84c),
	.w1(32'h3966c26f),
	.w2(32'h39119522),
	.w3(32'hba79a51f),
	.w4(32'h38b82c90),
	.w5(32'h3a974d9e),
	.w6(32'hb8c0a791),
	.w7(32'h39d4bb5e),
	.w8(32'h3adbc617),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5816b),
	.w1(32'hba3cce3d),
	.w2(32'hba5f3402),
	.w3(32'hba84b889),
	.w4(32'hba8b4938),
	.w5(32'hbac12d61),
	.w6(32'h396e9db0),
	.w7(32'h3ad401fd),
	.w8(32'h382cf9e6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8913847),
	.w1(32'hba153657),
	.w2(32'hb997be12),
	.w3(32'h39aab3c0),
	.w4(32'hb81ee10b),
	.w5(32'h3abcd81c),
	.w6(32'h398ef970),
	.w7(32'hb961c108),
	.w8(32'h3a05453a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06670e),
	.w1(32'h3b02ef07),
	.w2(32'h3affb26d),
	.w3(32'h3a5f2a96),
	.w4(32'hba71f424),
	.w5(32'hbb95b924),
	.w6(32'h3a8da123),
	.w7(32'hbac66ea8),
	.w8(32'hbba22c73),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940908f),
	.w1(32'h399c38d2),
	.w2(32'h3922b4c3),
	.w3(32'h394289b5),
	.w4(32'h398ca758),
	.w5(32'h39233c1a),
	.w6(32'h39a9360c),
	.w7(32'h39a28c18),
	.w8(32'h36c5ba8c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e34d5c),
	.w1(32'h394f166a),
	.w2(32'hb7d0b4d5),
	.w3(32'hb8b87a41),
	.w4(32'h39ff41a0),
	.w5(32'h3972b00d),
	.w6(32'hb8d0552e),
	.w7(32'h39c8b5fd),
	.w8(32'h390e3b7a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1d674),
	.w1(32'hb96e23b5),
	.w2(32'hb9b369bf),
	.w3(32'h39131f06),
	.w4(32'hb80b9092),
	.w5(32'hb88b4f77),
	.w6(32'h39de9cc7),
	.w7(32'h38b26093),
	.w8(32'hb9681849),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb5d9a),
	.w1(32'hba8096ad),
	.w2(32'hb9c7bd4d),
	.w3(32'hba9c9cfd),
	.w4(32'hba9f1b7b),
	.w5(32'hba83945e),
	.w6(32'hbaaf1daa),
	.w7(32'hbb000ce8),
	.w8(32'hba3c4bb4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bb871a),
	.w1(32'hb96a9376),
	.w2(32'hb9f7b868),
	.w3(32'hb9cdce0d),
	.w4(32'hb9c9e975),
	.w5(32'hba1d9714),
	.w6(32'hba280ce2),
	.w7(32'hb9b42cb9),
	.w8(32'hb9df3463),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bae448),
	.w1(32'hb9bc0550),
	.w2(32'h3aac3ec7),
	.w3(32'hba2194fd),
	.w4(32'hbae070e4),
	.w5(32'hbb560171),
	.w6(32'h3a5b0e17),
	.w7(32'hbaf9e451),
	.w8(32'hbb467d36),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9993a49),
	.w1(32'h39a13594),
	.w2(32'hb97a860e),
	.w3(32'hba72e05f),
	.w4(32'hba22df04),
	.w5(32'hb8625fd0),
	.w6(32'h3914696e),
	.w7(32'hb7b94b71),
	.w8(32'h3a9dfec2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38168a95),
	.w1(32'h39993dc7),
	.w2(32'h39072dd8),
	.w3(32'h378f0cfc),
	.w4(32'h39072b7d),
	.w5(32'h392c2bda),
	.w6(32'hb88bd7e2),
	.w7(32'hb8a5e37f),
	.w8(32'hb8a8c7f6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88dc047),
	.w1(32'hb96b222a),
	.w2(32'hb99b53cc),
	.w3(32'hb8fada5e),
	.w4(32'hb95a7cf5),
	.w5(32'hb9cc0a6e),
	.w6(32'hb91e6797),
	.w7(32'hb939e50e),
	.w8(32'hb99bf2fb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389eb5a7),
	.w1(32'hb80fc89d),
	.w2(32'h398c05bd),
	.w3(32'hb7a0877f),
	.w4(32'hb950533f),
	.w5(32'h38f1c610),
	.w6(32'h389cb328),
	.w7(32'hb91e87ca),
	.w8(32'h397fcd39),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba8e00),
	.w1(32'hb8101e15),
	.w2(32'hb9ae5c0c),
	.w3(32'h3953a88d),
	.w4(32'h3829f85d),
	.w5(32'hb983728c),
	.w6(32'h39906507),
	.w7(32'hb7b4a584),
	.w8(32'hb9951b9a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39175238),
	.w1(32'h391077fc),
	.w2(32'hb932d9ce),
	.w3(32'h39f22916),
	.w4(32'h39ba2302),
	.w5(32'h3933105e),
	.w6(32'h389475a9),
	.w7(32'h38b8e5fa),
	.w8(32'hb97b14b0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b861ce),
	.w1(32'h3912ea3d),
	.w2(32'h398e855f),
	.w3(32'hb93b0d18),
	.w4(32'hba6123c6),
	.w5(32'hbac165cf),
	.w6(32'hba23c8d5),
	.w7(32'hba5e1c53),
	.w8(32'hbad726eb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba099998),
	.w1(32'h38a737d5),
	.w2(32'h3a7626d8),
	.w3(32'hb9155994),
	.w4(32'hbb0ae6da),
	.w5(32'h3825cad9),
	.w6(32'hbae5539f),
	.w7(32'hbb47674f),
	.w8(32'h3ae0ef2c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fa68c6),
	.w1(32'hb8c25fc9),
	.w2(32'hb95affc3),
	.w3(32'h379c8b4f),
	.w4(32'hb946f188),
	.w5(32'hb99f5b8b),
	.w6(32'hb9053a1f),
	.w7(32'hb81d7611),
	.w8(32'hb878c9da),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902b595),
	.w1(32'h38fdbc31),
	.w2(32'h37ced6d7),
	.w3(32'hb83478e9),
	.w4(32'hb6c7839f),
	.w5(32'hb87ad1ce),
	.w6(32'hb88422f6),
	.w7(32'h37cd7be4),
	.w8(32'hb83cb384),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9017be9),
	.w1(32'h39aac406),
	.w2(32'h3981355e),
	.w3(32'hb8d3f452),
	.w4(32'h3938b883),
	.w5(32'hb89c962c),
	.w6(32'h3802738d),
	.w7(32'h3968e938),
	.w8(32'h38f9b50e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d81f1),
	.w1(32'h39628e89),
	.w2(32'h3966a040),
	.w3(32'h391f89ae),
	.w4(32'h389e20c3),
	.w5(32'hb71e92e4),
	.w6(32'h3943d4f1),
	.w7(32'h3945d2ee),
	.w8(32'h398d8ff5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d52e17),
	.w1(32'hb9ece35a),
	.w2(32'h3ac7bafd),
	.w3(32'h3b94eb1c),
	.w4(32'h3a625691),
	.w5(32'h3b823251),
	.w6(32'h3b0a22ab),
	.w7(32'hbb270469),
	.w8(32'hba874cac),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8c40f),
	.w1(32'hb8e97b33),
	.w2(32'hbb12a5ef),
	.w3(32'h39124c68),
	.w4(32'hbb666ada),
	.w5(32'hbb9a4307),
	.w6(32'h39c43578),
	.w7(32'h39fcb088),
	.w8(32'hba68e40e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5be42),
	.w1(32'hba459060),
	.w2(32'hba7e1ac6),
	.w3(32'hba040e3d),
	.w4(32'hbac00178),
	.w5(32'hbb227942),
	.w6(32'hb9c6ba8a),
	.w7(32'hba60fa9d),
	.w8(32'h39db7b71),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d1e1e),
	.w1(32'h3b47c673),
	.w2(32'h3b0ba4f1),
	.w3(32'h3a4a18c9),
	.w4(32'h3b8815bb),
	.w5(32'h3ba341c2),
	.w6(32'h3ac35b5d),
	.w7(32'h3b060a04),
	.w8(32'h3b55d0ec),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb739bd38),
	.w1(32'h36661a2a),
	.w2(32'hb79e7f0b),
	.w3(32'hb6890bcd),
	.w4(32'h3797986b),
	.w5(32'h3752689f),
	.w6(32'h372af106),
	.w7(32'h380b163b),
	.w8(32'hb72852d5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb656b3c0),
	.w1(32'hb76b315a),
	.w2(32'hb716bd53),
	.w3(32'hb6e9d731),
	.w4(32'hb71b3cac),
	.w5(32'h3820bf48),
	.w6(32'h37882579),
	.w7(32'h37d7afba),
	.w8(32'h387870b8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb769ec25),
	.w1(32'hb6f673d4),
	.w2(32'h3771413b),
	.w3(32'hb784c52e),
	.w4(32'hb74f57f5),
	.w5(32'h371ae669),
	.w6(32'hb763b5aa),
	.w7(32'hb7b73bde),
	.w8(32'h36d38e16),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39937af9),
	.w1(32'h3881b0e5),
	.w2(32'h398e23a7),
	.w3(32'hb7ba6546),
	.w4(32'hb9b72fb3),
	.w5(32'hb9e8ac99),
	.w6(32'h393b68be),
	.w7(32'hba3d63d7),
	.w8(32'hba37674f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d9b444),
	.w1(32'hb7a58d1c),
	.w2(32'h36168cec),
	.w3(32'h36bc91ee),
	.w4(32'h3704de2d),
	.w5(32'h3800d727),
	.w6(32'h37895b5e),
	.w7(32'h37f30d8f),
	.w8(32'h382639cd),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a3dfa),
	.w1(32'h398b44da),
	.w2(32'h39792bf8),
	.w3(32'h394b464f),
	.w4(32'h3a85551a),
	.w5(32'h3a1515be),
	.w6(32'h3a4c23ba),
	.w7(32'h3a13f6a3),
	.w8(32'hba694cf3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00a48c),
	.w1(32'h3aa5d3ee),
	.w2(32'h39a8b96f),
	.w3(32'hba7be28d),
	.w4(32'hba07fa9f),
	.w5(32'hbb3c3547),
	.w6(32'hba98d5a4),
	.w7(32'hba36126a),
	.w8(32'hbb701b9d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6265b),
	.w1(32'h3996dcbe),
	.w2(32'hb9bb2900),
	.w3(32'h388a38d1),
	.w4(32'h3a8a50fe),
	.w5(32'h3a95e49d),
	.w6(32'h398e1afd),
	.w7(32'h3a66eafd),
	.w8(32'h3a668416),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3882808c),
	.w1(32'hb9c3b7b4),
	.w2(32'hb961746e),
	.w3(32'hb9b3a9cc),
	.w4(32'hba7ee61b),
	.w5(32'hbaa480b1),
	.w6(32'hb9f1e166),
	.w7(32'hba8c7989),
	.w8(32'hba3e1629),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39920124),
	.w1(32'hb92b00ce),
	.w2(32'h39f7767f),
	.w3(32'h3b4707d9),
	.w4(32'h3b23d8f9),
	.w5(32'h3ae14284),
	.w6(32'h3b6e0de4),
	.w7(32'h3b0cb92a),
	.w8(32'hb9c0a110),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae2303),
	.w1(32'hb970f131),
	.w2(32'hb9c16043),
	.w3(32'hba3cb3a4),
	.w4(32'hb9bdb202),
	.w5(32'h3a88a0f8),
	.w6(32'hba18cb64),
	.w7(32'hba78b65a),
	.w8(32'h3a9c1824),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cba871),
	.w1(32'h3a0d5d11),
	.w2(32'h39df9e8f),
	.w3(32'h399da235),
	.w4(32'hb83c088d),
	.w5(32'hba9d1015),
	.w6(32'h39426972),
	.w7(32'hb9c2aa71),
	.w8(32'hbac34388),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b946fb),
	.w1(32'hb6ce9da5),
	.w2(32'hb3c8a070),
	.w3(32'h3604d829),
	.w4(32'hb73d1ac4),
	.w5(32'hb6ff02bb),
	.w6(32'h36e5cc95),
	.w7(32'h36c29b97),
	.w8(32'h375db917),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb789d4dc),
	.w1(32'hb80066b9),
	.w2(32'hb5e77417),
	.w3(32'hb778e4b0),
	.w4(32'h3703a8e7),
	.w5(32'h37c1c4ea),
	.w6(32'hb7c67f55),
	.w7(32'hb77b8d5b),
	.w8(32'hb5dadfb9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64e12c7),
	.w1(32'hb575f1f2),
	.w2(32'hb508fc87),
	.w3(32'hb5937354),
	.w4(32'hb4ac4afc),
	.w5(32'hb6534032),
	.w6(32'hb50e51ea),
	.w7(32'h367efbad),
	.w8(32'hb6144909),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ade8a3),
	.w1(32'h3992667e),
	.w2(32'h39b091c8),
	.w3(32'h38c1e140),
	.w4(32'hb6aa191a),
	.w5(32'h38e3fbc4),
	.w6(32'hb815a316),
	.w7(32'hb94e5cc0),
	.w8(32'hb98e67e3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9336d),
	.w1(32'h39c49d19),
	.w2(32'hb9636db6),
	.w3(32'h39d96414),
	.w4(32'h3b4030c6),
	.w5(32'h3b46df7a),
	.w6(32'hb9ab39f2),
	.w7(32'h3aec2908),
	.w8(32'h3ad88cd4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393fce25),
	.w1(32'h399b141d),
	.w2(32'h390eea76),
	.w3(32'hb7bc1c4a),
	.w4(32'h39338876),
	.w5(32'hb76b0f69),
	.w6(32'hb8d6bdc2),
	.w7(32'h38e06a88),
	.w8(32'h37f6212a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bcf91),
	.w1(32'hb8815674),
	.w2(32'hb759c632),
	.w3(32'hb979710f),
	.w4(32'hba2e0420),
	.w5(32'hb9f49bb7),
	.w6(32'h3ace122a),
	.w7(32'h3b29469f),
	.w8(32'h3aa5acaa),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d5ff1),
	.w1(32'hb932d389),
	.w2(32'h3a0cca68),
	.w3(32'hba212f6a),
	.w4(32'hbaae338c),
	.w5(32'hbb3babfd),
	.w6(32'h3977385f),
	.w7(32'hbaa35566),
	.w8(32'hbb1f556b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a357760),
	.w1(32'h3a978b91),
	.w2(32'h3ab943c2),
	.w3(32'h3a7a908c),
	.w4(32'h3b100217),
	.w5(32'h3b399ffd),
	.w6(32'h39b2f890),
	.w7(32'h3a54f3b0),
	.w8(32'h3a9f13d6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba644a3f),
	.w1(32'h3a8e2863),
	.w2(32'h3a5a9410),
	.w3(32'h3a12f289),
	.w4(32'h3bb6920d),
	.w5(32'h3b070ff6),
	.w6(32'h3a92c928),
	.w7(32'h3b5c3582),
	.w8(32'hbb243963),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0f71f),
	.w1(32'h3a0c47d0),
	.w2(32'h3aa5cb5d),
	.w3(32'hb9e05bc5),
	.w4(32'h394f9948),
	.w5(32'h3a031ca1),
	.w6(32'hb9dd1719),
	.w7(32'hb9d473f7),
	.w8(32'h39c23681),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d5616),
	.w1(32'hbafa2ea3),
	.w2(32'hbb01d0ab),
	.w3(32'hba564ab2),
	.w4(32'hbb01f2fa),
	.w5(32'hbb2704c5),
	.w6(32'hb9caceaa),
	.w7(32'hbad34a4d),
	.w8(32'hbaa426a1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3c551),
	.w1(32'hbae0f851),
	.w2(32'hbae34bd5),
	.w3(32'h3ad37b5a),
	.w4(32'h3adbf759),
	.w5(32'h3a9f92a5),
	.w6(32'h3abc567e),
	.w7(32'h3a50fe64),
	.w8(32'h3a5f981e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9980b30),
	.w1(32'h39e36792),
	.w2(32'h3ad81fae),
	.w3(32'h3a808ecc),
	.w4(32'h3b28f042),
	.w5(32'h3b5e06bb),
	.w6(32'h3a56e595),
	.w7(32'h3a7f1334),
	.w8(32'h3a897aa5),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899a031),
	.w1(32'h3853310e),
	.w2(32'hb898e343),
	.w3(32'h37a456c8),
	.w4(32'h37a04412),
	.w5(32'hb8e10c6e),
	.w6(32'h37e17012),
	.w7(32'h37697e74),
	.w8(32'hb8bb8a4b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3285ee),
	.w1(32'h3900d380),
	.w2(32'hb7f0f319),
	.w3(32'h3959ffe5),
	.w4(32'hbab273d7),
	.w5(32'hbb5833d9),
	.w6(32'h3905db85),
	.w7(32'hba88d1d4),
	.w8(32'hbb27e84b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b06a5),
	.w1(32'h3a9fd71e),
	.w2(32'h3aa49c7c),
	.w3(32'h3aa5108c),
	.w4(32'h3baa974a),
	.w5(32'h3b8a371d),
	.w6(32'h3b4d7db0),
	.w7(32'h3b428687),
	.w8(32'h3a44c66b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fb8ad),
	.w1(32'h39f5ed1f),
	.w2(32'hbbb28e7a),
	.w3(32'hbb4bbe6c),
	.w4(32'h3b5e3e17),
	.w5(32'hba993cc5),
	.w6(32'hbb73819d),
	.w7(32'h3c09f2cf),
	.w8(32'hbb56a359),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acaa65d),
	.w1(32'h3b2e3880),
	.w2(32'h3af0c67e),
	.w3(32'h3b0c1314),
	.w4(32'h3bcbc7ba),
	.w5(32'h3b98faef),
	.w6(32'hbaa2cb90),
	.w7(32'h3b66a5e9),
	.w8(32'h3b19bf0e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9789e5b),
	.w1(32'h3a97fd6e),
	.w2(32'h3a132ed2),
	.w3(32'hba186598),
	.w4(32'h3a097108),
	.w5(32'h3a25dd2e),
	.w6(32'h3a6a9f91),
	.w7(32'h3b044e0d),
	.w8(32'h3a86144b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f898f),
	.w1(32'h39d48c0f),
	.w2(32'hbac31375),
	.w3(32'h3a8c2071),
	.w4(32'h3bcd037b),
	.w5(32'h3a4d1cf8),
	.w6(32'h3aa306ac),
	.w7(32'h3bce39f8),
	.w8(32'hbab328d8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c60b2),
	.w1(32'hb872cf16),
	.w2(32'hb937853c),
	.w3(32'hb9098bbf),
	.w4(32'hb83ef926),
	.w5(32'hb98a0beb),
	.w6(32'h37826467),
	.w7(32'h37c063e8),
	.w8(32'hb8fb8243),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1df1cd),
	.w1(32'hbab20f23),
	.w2(32'hbb9e6576),
	.w3(32'hbb217189),
	.w4(32'h3b90d662),
	.w5(32'hba6cbd8a),
	.w6(32'hb95353df),
	.w7(32'h3bedfe2c),
	.w8(32'h3a5fed6b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd6bf0),
	.w1(32'h3938cd0c),
	.w2(32'h3a582645),
	.w3(32'h3a52849d),
	.w4(32'h3aaa849f),
	.w5(32'h3af666de),
	.w6(32'h399b3611),
	.w7(32'h3b0d3eff),
	.w8(32'hb958491b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38298938),
	.w1(32'hb6b8012b),
	.w2(32'hb7ddc4bc),
	.w3(32'h38740bb4),
	.w4(32'h381a77a6),
	.w5(32'h38173762),
	.w6(32'h380521cf),
	.w7(32'h3768cec5),
	.w8(32'h383163a9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396c34be),
	.w1(32'hb950ea5a),
	.w2(32'hbaab145d),
	.w3(32'hb8c5c11b),
	.w4(32'h39f0851e),
	.w5(32'hb9854392),
	.w6(32'hba622051),
	.w7(32'hb7effe40),
	.w8(32'h3a144021),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389c8fda),
	.w1(32'h39971961),
	.w2(32'hb7927042),
	.w3(32'h3a0a31b4),
	.w4(32'hba4a02c3),
	.w5(32'hbb12bb78),
	.w6(32'hb8d26211),
	.w7(32'hbabd97f6),
	.w8(32'hbb4e7394),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39892c22),
	.w1(32'h3a362a74),
	.w2(32'h39e8d6b7),
	.w3(32'hba0b3e47),
	.w4(32'h399c92d6),
	.w5(32'h3a22c2f8),
	.w6(32'h3980df02),
	.w7(32'h3a08974c),
	.w8(32'h3a269ca6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f4049),
	.w1(32'h38d20a3e),
	.w2(32'h3a27ff64),
	.w3(32'h39d01c1f),
	.w4(32'h3a425509),
	.w5(32'h3a825f60),
	.w6(32'h3ac7d5fa),
	.w7(32'hb8b6cccb),
	.w8(32'h3a802e56),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1aa33b),
	.w1(32'h39a44ca3),
	.w2(32'hb95785da),
	.w3(32'h39f13afd),
	.w4(32'h3aca9325),
	.w5(32'h3ab915ef),
	.w6(32'h39d25d58),
	.w7(32'h3a42b025),
	.w8(32'h3a10bad5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11e089),
	.w1(32'h3b6a5c43),
	.w2(32'h3b0b2a13),
	.w3(32'hb9f85df6),
	.w4(32'h3ad25d9d),
	.w5(32'hba8711f6),
	.w6(32'h3b152d22),
	.w7(32'h3ba56846),
	.w8(32'h3b0d3ddb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d8917),
	.w1(32'hbaf7b3dd),
	.w2(32'hbb5a6dca),
	.w3(32'h3a68236a),
	.w4(32'hbaaa4339),
	.w5(32'hba97cb99),
	.w6(32'hbab40aba),
	.w7(32'hbb0e6175),
	.w8(32'hba19599b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9ae8a),
	.w1(32'h38be9ba7),
	.w2(32'h3a224f58),
	.w3(32'hba32162e),
	.w4(32'hba0a24bd),
	.w5(32'h383ede4d),
	.w6(32'hb9ab136e),
	.w7(32'hb92755dc),
	.w8(32'h39c0def9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6713588),
	.w1(32'hb7834956),
	.w2(32'h364760ae),
	.w3(32'h360eb986),
	.w4(32'h33e07dfc),
	.w5(32'h37db300d),
	.w6(32'hb6d28e1b),
	.w7(32'hb7cd4f27),
	.w8(32'h36ab77a0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb947864d),
	.w1(32'hb9ccf226),
	.w2(32'hb9e7e323),
	.w3(32'h38581c6e),
	.w4(32'h389e505b),
	.w5(32'h398c90b6),
	.w6(32'hb7c5b087),
	.w7(32'h39bab4a2),
	.w8(32'h39c23b15),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360070f0),
	.w1(32'h3830abe9),
	.w2(32'h37f3df6a),
	.w3(32'h3769c0e0),
	.w4(32'h385e05e9),
	.w5(32'h37c9490b),
	.w6(32'h3666d6f6),
	.w7(32'h373d522f),
	.w8(32'h3651b3be),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h356b52ad),
	.w1(32'hb72770a6),
	.w2(32'hb5d34c67),
	.w3(32'h36918625),
	.w4(32'hb700e784),
	.w5(32'hb7a92226),
	.w6(32'hb640ba04),
	.w7(32'hb73893d7),
	.w8(32'hb7759640),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6dc1a),
	.w1(32'h39525e01),
	.w2(32'h3a13d415),
	.w3(32'hba1249c7),
	.w4(32'hb9f60000),
	.w5(32'h380ba888),
	.w6(32'hb98b8639),
	.w7(32'h390113f1),
	.w8(32'h3a123e1a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38333952),
	.w1(32'h3767e2b4),
	.w2(32'h38b4b48a),
	.w3(32'h38ea54b3),
	.w4(32'h37ea2e36),
	.w5(32'hb4e08d33),
	.w6(32'hb68ade28),
	.w7(32'hb8b2432a),
	.w8(32'hb8f21fd5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a251ccb),
	.w1(32'h3a7b19e7),
	.w2(32'h39f4f1f4),
	.w3(32'h39679c1b),
	.w4(32'h3aa664b6),
	.w5(32'hba1e6d8f),
	.w6(32'h3a2e52d3),
	.w7(32'h3a4af1c3),
	.w8(32'hbacf324f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3d958),
	.w1(32'h3a9f9678),
	.w2(32'h3a675fd5),
	.w3(32'h3a6cfe7b),
	.w4(32'h3b27e24e),
	.w5(32'h3b455c42),
	.w6(32'h3a323051),
	.w7(32'h3a3f1102),
	.w8(32'h3ac2c687),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70c74da),
	.w1(32'hb72b2e36),
	.w2(32'hb6a7c1bd),
	.w3(32'hb4c2ad9a),
	.w4(32'h37b48e69),
	.w5(32'h37f7f483),
	.w6(32'h36853bda),
	.w7(32'h380ef9ac),
	.w8(32'h3831dc5d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381ea5b8),
	.w1(32'h38804340),
	.w2(32'h3851dafc),
	.w3(32'h37fb0c46),
	.w4(32'hb807c301),
	.w5(32'hb7cfc015),
	.w6(32'h388248f8),
	.w7(32'hb88b0f3b),
	.w8(32'h367cffbb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377ff3cc),
	.w1(32'h37b96f76),
	.w2(32'h375b2472),
	.w3(32'h3721b3ac),
	.w4(32'h378a91b7),
	.w5(32'h378591b9),
	.w6(32'h36f81b53),
	.w7(32'h3744a051),
	.w8(32'h36f6d458),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64b7231),
	.w1(32'h38cfc4a9),
	.w2(32'hb90de33f),
	.w3(32'h3956f4cf),
	.w4(32'h392e5fdd),
	.w5(32'hb98ca823),
	.w6(32'h399bdc1b),
	.w7(32'h3999bda0),
	.w8(32'hb82d3664),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b745b2f),
	.w1(32'h3b2765f7),
	.w2(32'h39b2b10f),
	.w3(32'hb7bf0bdb),
	.w4(32'h3a9d40e8),
	.w5(32'hbc0485d7),
	.w6(32'h3af21cf1),
	.w7(32'h3b28bc45),
	.w8(32'hbaefa97c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a688e),
	.w1(32'hb9bf7f3f),
	.w2(32'h3a6dec58),
	.w3(32'h39b20cf5),
	.w4(32'hbafc962b),
	.w5(32'hbb20ff27),
	.w6(32'h374bbbe2),
	.w7(32'hbb030a24),
	.w8(32'hbb2da731),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38199526),
	.w1(32'h38bd1736),
	.w2(32'h37fa5631),
	.w3(32'h39856bf1),
	.w4(32'h3a09f08e),
	.w5(32'h392b7aae),
	.w6(32'hb89c9d6d),
	.w7(32'h38fb5d8e),
	.w8(32'hb9ddc5c8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52aed3),
	.w1(32'hba9e99c2),
	.w2(32'hbac976b4),
	.w3(32'h388682e6),
	.w4(32'hba536ae9),
	.w5(32'hba2a0dc7),
	.w6(32'h3a31b8ea),
	.w7(32'h390a0014),
	.w8(32'hb96867f6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949ad9c),
	.w1(32'hb77c4a76),
	.w2(32'hb8663d0d),
	.w3(32'h38e3c441),
	.w4(32'h39bab790),
	.w5(32'h3a3ec9ff),
	.w6(32'h3967bde5),
	.w7(32'h39e44c73),
	.w8(32'h3a0cfe41),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380949cd),
	.w1(32'hb9c940b9),
	.w2(32'h3598acb4),
	.w3(32'hb9e640c5),
	.w4(32'hba49517e),
	.w5(32'hb9bb3e98),
	.w6(32'hb987eaab),
	.w7(32'hba870f64),
	.w8(32'hba2131f9),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a30172),
	.w1(32'hba3a050a),
	.w2(32'hba8bf34e),
	.w3(32'h390ef05d),
	.w4(32'h3a1f5d84),
	.w5(32'h3ad1e6aa),
	.w6(32'h39af62a6),
	.w7(32'hb9d67821),
	.w8(32'h3ace8d5a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75bb5d),
	.w1(32'h3a7654d4),
	.w2(32'h3ac80b93),
	.w3(32'h3a718428),
	.w4(32'h398426db),
	.w5(32'hbb166fb1),
	.w6(32'h3a434667),
	.w7(32'hbaae539f),
	.w8(32'hbb3437bf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398441e6),
	.w1(32'h39ac4e50),
	.w2(32'h3a35162f),
	.w3(32'h39fe51cf),
	.w4(32'h3a8883e7),
	.w5(32'h3a9b6bfb),
	.w6(32'h38841b27),
	.w7(32'h39ce1700),
	.w8(32'h3986e51f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cc0a5),
	.w1(32'hb8a013dc),
	.w2(32'hb9eb52c8),
	.w3(32'h3ab26adb),
	.w4(32'h3b2566be),
	.w5(32'h38ccf648),
	.w6(32'h39bab982),
	.w7(32'h395fda9c),
	.w8(32'hba8fbe3a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a015ed),
	.w1(32'h3a8c9ea9),
	.w2(32'h3ac03f4a),
	.w3(32'h399ca1a4),
	.w4(32'h3a4e1050),
	.w5(32'hbab56797),
	.w6(32'h3a06f348),
	.w7(32'h3a5c6533),
	.w8(32'hbadb98dc),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72c91c),
	.w1(32'hb55f6272),
	.w2(32'hb6231e14),
	.w3(32'hba95d78c),
	.w4(32'h399e0eac),
	.w5(32'h39795d32),
	.w6(32'hb9ac792b),
	.w7(32'h3aed46b4),
	.w8(32'h3ae12d02),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa92e1),
	.w1(32'h38b48ade),
	.w2(32'h3a71a0ac),
	.w3(32'h3a027b75),
	.w4(32'h3998b6ce),
	.w5(32'hba383edf),
	.w6(32'h375df60b),
	.w7(32'hba501844),
	.w8(32'hbaeeb96d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df819f),
	.w1(32'hb89c348a),
	.w2(32'hb690f78f),
	.w3(32'hb82ed2f3),
	.w4(32'hb8e4bebc),
	.w5(32'hb82bf070),
	.w6(32'hb875a8a8),
	.w7(32'hb8a2ff7e),
	.w8(32'hb9257c72),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b0316),
	.w1(32'h3abd36af),
	.w2(32'h3afec44e),
	.w3(32'h3a5f7985),
	.w4(32'h3ae1f1db),
	.w5(32'h3b033c66),
	.w6(32'h3a2187b9),
	.w7(32'h3a8c68e8),
	.w8(32'h3aeaff15),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8be7c4a),
	.w1(32'h398234cd),
	.w2(32'h39d71cfd),
	.w3(32'hba276bf4),
	.w4(32'h3a15c4a0),
	.w5(32'h3a1c68d3),
	.w6(32'h3944f0a4),
	.w7(32'h39f13f45),
	.w8(32'h39f561c8),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38572593),
	.w1(32'h37282870),
	.w2(32'hb7132b2f),
	.w3(32'h38d51fac),
	.w4(32'h38ca08ea),
	.w5(32'hb79925eb),
	.w6(32'h38cc0ec1),
	.w7(32'h37e7e90e),
	.w8(32'h374f8bd2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84ef589),
	.w1(32'hb6dcdd0a),
	.w2(32'h383830e4),
	.w3(32'h38782186),
	.w4(32'h3798a416),
	.w5(32'hb7ed113b),
	.w6(32'h37481950),
	.w7(32'hb81e70ca),
	.w8(32'h38994fa7),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941f8ee),
	.w1(32'hb9b7f926),
	.w2(32'hb9a044fa),
	.w3(32'hb8b30dad),
	.w4(32'h39c5010e),
	.w5(32'h3a0e2b75),
	.w6(32'hb81c8491),
	.w7(32'h3a13de55),
	.w8(32'h37b9178d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d44ca),
	.w1(32'h3a212c33),
	.w2(32'hb9837e4f),
	.w3(32'hb9af3819),
	.w4(32'h3b041e39),
	.w5(32'h3b07f2be),
	.w6(32'hba5a5ec5),
	.w7(32'h3abd8b69),
	.w8(32'h39ca7166),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fe9a3),
	.w1(32'h3a2999d6),
	.w2(32'h395ba08c),
	.w3(32'h3a191fa2),
	.w4(32'hb9a84aac),
	.w5(32'hba595d40),
	.w6(32'h3993c7bb),
	.w7(32'hba36f3db),
	.w8(32'hbae04941),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6936679),
	.w1(32'hb78a51a6),
	.w2(32'hb7f68f38),
	.w3(32'hb71acb35),
	.w4(32'hb660e1fc),
	.w5(32'hb781fb7f),
	.w6(32'h378dabb3),
	.w7(32'hb74d4a97),
	.w8(32'hb75c01c5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38754d46),
	.w1(32'hba097dad),
	.w2(32'hb9873d7f),
	.w3(32'hb9ce6ec7),
	.w4(32'hba8d8a6a),
	.w5(32'hba24e3ab),
	.w6(32'hb9d7cd7c),
	.w7(32'hbad30af5),
	.w8(32'hbaf898e5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f9ef3),
	.w1(32'hb993d508),
	.w2(32'hb8b26dbc),
	.w3(32'hb953ccc0),
	.w4(32'hb9c70214),
	.w5(32'hba0341e4),
	.w6(32'h38cfe8cf),
	.w7(32'hb9f8b038),
	.w8(32'hba426c98),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b62845),
	.w1(32'h3a9b4c06),
	.w2(32'hb885a3ee),
	.w3(32'h3a850523),
	.w4(32'h3b796415),
	.w5(32'hb87bd8f6),
	.w6(32'h3a3a966b),
	.w7(32'h3aab5c67),
	.w8(32'hbb38553a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6657ae),
	.w1(32'h3999c7f0),
	.w2(32'h3a8920e3),
	.w3(32'hba3a4f30),
	.w4(32'h3a981e57),
	.w5(32'h3bc02237),
	.w6(32'h3b333740),
	.w7(32'hbab46066),
	.w8(32'h3b7a8c86),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb825a107),
	.w1(32'h3907520c),
	.w2(32'hb909e6e7),
	.w3(32'h39529cc7),
	.w4(32'h3a823d77),
	.w5(32'h3a8b1904),
	.w6(32'h38bd07e6),
	.w7(32'h3a1e3a25),
	.w8(32'h3a9afc73),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925e610),
	.w1(32'hb940a072),
	.w2(32'hb94880c8),
	.w3(32'hb9888e54),
	.w4(32'hb9178a60),
	.w5(32'hb8fb38f8),
	.w6(32'hb7f1272e),
	.w7(32'h386c77ec),
	.w8(32'h388f61f4),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946d6e2),
	.w1(32'h39d9af40),
	.w2(32'h3a50b69d),
	.w3(32'hb9eeaeb3),
	.w4(32'h390df78a),
	.w5(32'h3a2f4eb7),
	.w6(32'h39b74d2d),
	.w7(32'h3a70d1ff),
	.w8(32'h3a75c847),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f7995),
	.w1(32'h39d5c9fa),
	.w2(32'h38fbf7cf),
	.w3(32'hb955288d),
	.w4(32'h3aed7a00),
	.w5(32'h3b240474),
	.w6(32'hba028c2e),
	.w7(32'h3a1ec5d2),
	.w8(32'h3aeccdd7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1d239),
	.w1(32'h3a53b17f),
	.w2(32'h3a57c8db),
	.w3(32'h397af38c),
	.w4(32'h3aa52815),
	.w5(32'h3acf1900),
	.w6(32'h392e5cfc),
	.w7(32'h3a02a22f),
	.w8(32'h3a38e53a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d0ebd),
	.w1(32'h3985e7ea),
	.w2(32'h39b24be7),
	.w3(32'h38d55221),
	.w4(32'h3a2789fe),
	.w5(32'h39cb6299),
	.w6(32'h39358491),
	.w7(32'h39988d47),
	.w8(32'hba0724ec),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969834c),
	.w1(32'hb863f3cb),
	.w2(32'h3788bae5),
	.w3(32'h38f60559),
	.w4(32'h3911a29a),
	.w5(32'h38746ccf),
	.w6(32'hb8e770e6),
	.w7(32'h38aaa057),
	.w8(32'hb7c69873),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9210977),
	.w1(32'h39575a55),
	.w2(32'hb9908f3e),
	.w3(32'h3ac4bd40),
	.w4(32'h3a3c5c59),
	.w5(32'hbaa8652c),
	.w6(32'h3a8adfa2),
	.w7(32'h3a4cae58),
	.w8(32'hba81bf53),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a118786),
	.w1(32'h381a1a84),
	.w2(32'h39a7ac95),
	.w3(32'h39aa3458),
	.w4(32'h398e640b),
	.w5(32'hb93d20ab),
	.w6(32'h39ec5cd9),
	.w7(32'h390dbef6),
	.w8(32'hba747f53),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd7da3),
	.w1(32'hb94569c3),
	.w2(32'h3a4af203),
	.w3(32'h37bd314d),
	.w4(32'hba061d5b),
	.w5(32'h3a48091b),
	.w6(32'h3a674633),
	.w7(32'h3a2f233e),
	.w8(32'h3b1435a8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac1e50),
	.w1(32'h384b6514),
	.w2(32'h37a1b03e),
	.w3(32'h37d1f061),
	.w4(32'h3861106b),
	.w5(32'h37e98d2e),
	.w6(32'hb6c18f35),
	.w7(32'h3837707a),
	.w8(32'h37e1073f),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b395214),
	.w1(32'h3aedb29d),
	.w2(32'h3a72918f),
	.w3(32'h3b3112c9),
	.w4(32'h3af1f704),
	.w5(32'hb9fcb217),
	.w6(32'h3a7ec84f),
	.w7(32'hba182430),
	.w8(32'hbaca9e3a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a0f13f),
	.w1(32'hb5e931f8),
	.w2(32'hb7655b0e),
	.w3(32'hb7c80334),
	.w4(32'hb7acc568),
	.w5(32'hb80e1f3f),
	.w6(32'hb7a21e6c),
	.w7(32'hb7d14356),
	.w8(32'hb7c2aaac),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371ac92b),
	.w1(32'h37ab949f),
	.w2(32'hb83240ff),
	.w3(32'h37678158),
	.w4(32'h380478a6),
	.w5(32'hb85b3669),
	.w6(32'h37da0484),
	.w7(32'h3809246e),
	.w8(32'hb8ac0e1b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f7f6c9),
	.w1(32'h392b28a5),
	.w2(32'h38d1b80e),
	.w3(32'h39aa8613),
	.w4(32'h3a20ae1a),
	.w5(32'h3a2da999),
	.w6(32'h394620a8),
	.w7(32'h3994f8ad),
	.w8(32'h396a1923),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8ddb1),
	.w1(32'h3af1fdc0),
	.w2(32'h39ff0f16),
	.w3(32'h39ec67f0),
	.w4(32'hb9803377),
	.w5(32'hbb349b0f),
	.w6(32'hba891463),
	.w7(32'h3a4bef86),
	.w8(32'hbb424d1a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39831a5a),
	.w1(32'h3a071278),
	.w2(32'h390f46d2),
	.w3(32'h39971c90),
	.w4(32'h39e6d19c),
	.w5(32'h3932501f),
	.w6(32'h39aab7d7),
	.w7(32'h39d383ff),
	.w8(32'h389ef23b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dc43dd),
	.w1(32'h3a0c26e6),
	.w2(32'h3a7611c6),
	.w3(32'hb88bb306),
	.w4(32'h3986394f),
	.w5(32'h3aa1bac5),
	.w6(32'hb946dc8c),
	.w7(32'h39210ce0),
	.w8(32'h39fcc7a2),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d56aa),
	.w1(32'h3a1d8978),
	.w2(32'h3959da18),
	.w3(32'h39df179a),
	.w4(32'hb9b88f52),
	.w5(32'h3a513d28),
	.w6(32'hba14143a),
	.w7(32'hba880eaa),
	.w8(32'h3a52ffec),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7dabc4),
	.w1(32'h39b83b35),
	.w2(32'hb8a07ee4),
	.w3(32'h3998fa2d),
	.w4(32'hbabbc116),
	.w5(32'hbb2d94c3),
	.w6(32'hbafeac7e),
	.w7(32'hbb31a39a),
	.w8(32'hbb0eaab9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39056672),
	.w1(32'hba7e5fb2),
	.w2(32'hba737dc6),
	.w3(32'hb97a850e),
	.w4(32'hba850a34),
	.w5(32'hba174143),
	.w6(32'hb9776cbe),
	.w7(32'hba0f6c2d),
	.w8(32'hb98b2700),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982ea2f),
	.w1(32'hb90619c9),
	.w2(32'h39a96a1a),
	.w3(32'hb7c0e879),
	.w4(32'hbaae7d3a),
	.w5(32'hbb2aec9f),
	.w6(32'hb9bbb07d),
	.w7(32'hbaf55e99),
	.w8(32'hbb326dca),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bcb045),
	.w1(32'hb72b5910),
	.w2(32'h382bac21),
	.w3(32'h38723636),
	.w4(32'hb7f566bf),
	.w5(32'h37a780ee),
	.w6(32'h382dbd10),
	.w7(32'hb75fde44),
	.w8(32'h3856723f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a681e7),
	.w1(32'hb9d14922),
	.w2(32'hb8373f86),
	.w3(32'h3a1b4039),
	.w4(32'hb9064367),
	.w5(32'hb930452c),
	.w6(32'h3a5d19be),
	.w7(32'h39f52b36),
	.w8(32'h39d3b42e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb543261b),
	.w1(32'hb5f04821),
	.w2(32'hb75185d1),
	.w3(32'h371c740f),
	.w4(32'h364b2215),
	.w5(32'hb55c420e),
	.w6(32'h37872257),
	.w7(32'h37818636),
	.w8(32'h377e812a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919e5fe),
	.w1(32'hb96dd4a3),
	.w2(32'hb92c89a4),
	.w3(32'hb8dfdc64),
	.w4(32'hb958a0cd),
	.w5(32'h39515bf1),
	.w6(32'hb9942faa),
	.w7(32'hb9cb581f),
	.w8(32'hb9200ad1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394dd9c0),
	.w1(32'h38c1b59f),
	.w2(32'h38b35c70),
	.w3(32'h396d9a66),
	.w4(32'h39b874ea),
	.w5(32'h399b0b29),
	.w6(32'h39500086),
	.w7(32'h391b195d),
	.w8(32'h38d95cb0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14b723),
	.w1(32'hba5e2cd4),
	.w2(32'hbaafd932),
	.w3(32'h3937b010),
	.w4(32'hb99444d8),
	.w5(32'hba17d4e2),
	.w6(32'hba470b25),
	.w7(32'hba5f49c4),
	.w8(32'hb8b7b7f4),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb668cc8a),
	.w1(32'hb6b0aca3),
	.w2(32'h36568035),
	.w3(32'hb7397063),
	.w4(32'hb70af598),
	.w5(32'h368c4218),
	.w6(32'hb6d80deb),
	.w7(32'hb4556d22),
	.w8(32'h376f3b2a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c41414),
	.w1(32'hb7f8bab1),
	.w2(32'hb7dd1568),
	.w3(32'h37a813f6),
	.w4(32'hb76f7674),
	.w5(32'hb6feb57d),
	.w6(32'h36e15dc7),
	.w7(32'hb6a24ee4),
	.w8(32'h37509117),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2451b),
	.w1(32'h3a20646d),
	.w2(32'hb812accd),
	.w3(32'h3a1ea1d6),
	.w4(32'h3982ebf8),
	.w5(32'h3a786b1d),
	.w6(32'h3aa0b59e),
	.w7(32'h39fda845),
	.w8(32'h3a625a0b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca0bb3),
	.w1(32'hb96f01e6),
	.w2(32'hbb39876e),
	.w3(32'h3a57cb5e),
	.w4(32'h3a670004),
	.w5(32'hbb0a59f3),
	.w6(32'h3aa3ae9b),
	.w7(32'h3ab7bd34),
	.w8(32'hba843ada),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb866b0b4),
	.w1(32'hba00576e),
	.w2(32'hbae499a4),
	.w3(32'hba9618ba),
	.w4(32'h3b4339a7),
	.w5(32'h3af22111),
	.w6(32'hbac3e90b),
	.w7(32'h3b16f2d1),
	.w8(32'hba8326e6),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b9f802),
	.w1(32'hb8876e87),
	.w2(32'h36b88a90),
	.w3(32'hb7bf2fe2),
	.w4(32'h376ea6ca),
	.w5(32'h38a97567),
	.w6(32'h3793005f),
	.w7(32'hb88d93d4),
	.w8(32'h37da22ce),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba322bac),
	.w1(32'hb9a23afa),
	.w2(32'hb942037b),
	.w3(32'h3a429b88),
	.w4(32'hbb608cf8),
	.w5(32'hbbe0c0b7),
	.w6(32'hba04aeab),
	.w7(32'hbb44dfa7),
	.w8(32'hbbbee7b4),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a128c19),
	.w1(32'h3acd847f),
	.w2(32'h3b0dcbf7),
	.w3(32'h3a3f7fb4),
	.w4(32'h3a951ac9),
	.w5(32'h3bfdc9e3),
	.w6(32'h3a89c1f2),
	.w7(32'hba86be16),
	.w8(32'h3b9673ec),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ce750),
	.w1(32'h3a311d07),
	.w2(32'h38a81242),
	.w3(32'h3a485441),
	.w4(32'h3aa33ec2),
	.w5(32'h390d2700),
	.w6(32'h3a4cb599),
	.w7(32'h3a1e8040),
	.w8(32'hba8516fc),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb768cdd0),
	.w1(32'hb7bd2fde),
	.w2(32'hb81007bf),
	.w3(32'h37fed5b4),
	.w4(32'hb7cf15b2),
	.w5(32'hb8239e91),
	.w6(32'h3818501e),
	.w7(32'h3769a561),
	.w8(32'h3811d00d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80f4451),
	.w1(32'h379ac2cc),
	.w2(32'hb8ca1dbd),
	.w3(32'hb70ac89e),
	.w4(32'h360d53c7),
	.w5(32'hb87df979),
	.w6(32'h3742851a),
	.w7(32'h3864e9a1),
	.w8(32'hb6986cfc),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb612181c),
	.w1(32'h36a0a14a),
	.w2(32'h36d694f0),
	.w3(32'h35725dcb),
	.w4(32'hb61bd932),
	.w5(32'h361ac670),
	.w6(32'h366c3c8e),
	.w7(32'h36b1b970),
	.w8(32'h366a781f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee957b),
	.w1(32'h3b0440c1),
	.w2(32'h3a8c0f9a),
	.w3(32'h3afe6cac),
	.w4(32'h3b2f1ce5),
	.w5(32'hb9f83f19),
	.w6(32'h3ac0e135),
	.w7(32'h3b159158),
	.w8(32'hbad488ab),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1864b1),
	.w1(32'h39a535c7),
	.w2(32'h39b09f14),
	.w3(32'hb7c43b42),
	.w4(32'h3a105603),
	.w5(32'h38a9319e),
	.w6(32'hb980f592),
	.w7(32'hb9951ca6),
	.w8(32'hba88b29f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a84182),
	.w1(32'hb97a4ce9),
	.w2(32'hbaa068d3),
	.w3(32'hb98f3687),
	.w4(32'h3a4b4de5),
	.w5(32'h3a255bd1),
	.w6(32'h3855e892),
	.w7(32'h3ac1e7ef),
	.w8(32'h3a79e3e1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc27e6),
	.w1(32'hb93e10cb),
	.w2(32'hb8dab64f),
	.w3(32'h38959f4e),
	.w4(32'h39008679),
	.w5(32'h392c2a47),
	.w6(32'h39b4f3ae),
	.w7(32'h3a1278b5),
	.w8(32'h39f9c888),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990a3d1),
	.w1(32'h3bedca93),
	.w2(32'h3bed015a),
	.w3(32'h3a2213d7),
	.w4(32'h3abb492a),
	.w5(32'hbb3692f5),
	.w6(32'h38e043da),
	.w7(32'h3b35911e),
	.w8(32'hbaca3223),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba10aff),
	.w1(32'h3ae10860),
	.w2(32'hbadd6d89),
	.w3(32'h3bf94565),
	.w4(32'hbaa28100),
	.w5(32'hbabb9d79),
	.w6(32'h3b57b576),
	.w7(32'hba73df89),
	.w8(32'hbb8409f9),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99bad7),
	.w1(32'hbbca2ed8),
	.w2(32'hbb33a50f),
	.w3(32'h3aade8bf),
	.w4(32'hbbf65c8b),
	.w5(32'hbbe11b48),
	.w6(32'hbb92bd92),
	.w7(32'h3c6af38c),
	.w8(32'h3ce8da66),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5319be),
	.w1(32'hbb274ee6),
	.w2(32'h39eba2aa),
	.w3(32'h3b9019b5),
	.w4(32'hbc4cb790),
	.w5(32'hbc4bcd47),
	.w6(32'h3c1b7b55),
	.w7(32'hbc228f59),
	.w8(32'hbb425b04),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5e9e7),
	.w1(32'h3b774f47),
	.w2(32'h3c4fe28e),
	.w3(32'h39eca41f),
	.w4(32'h3c03cbed),
	.w5(32'h3c1a5eed),
	.w6(32'h3b97580b),
	.w7(32'hbc3f0ab4),
	.w8(32'hbc917020),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d4654),
	.w1(32'hbb129f0b),
	.w2(32'hbc0eae6b),
	.w3(32'hbb7db597),
	.w4(32'hba4cf985),
	.w5(32'hbaa99d0d),
	.w6(32'hbc45156b),
	.w7(32'hbbe0b287),
	.w8(32'hbbec09fb),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb11161),
	.w1(32'hbb809466),
	.w2(32'h3b6fad14),
	.w3(32'h3ba9a781),
	.w4(32'h39c9f20e),
	.w5(32'h3c199151),
	.w6(32'hbbd00817),
	.w7(32'hbb75d5b3),
	.w8(32'hbb6b967b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392624c9),
	.w1(32'h3b0115bc),
	.w2(32'h3aff17ae),
	.w3(32'h3b89ca6c),
	.w4(32'h3ae61190),
	.w5(32'h3bb798ca),
	.w6(32'hbbc2239b),
	.w7(32'h3b8b49a7),
	.w8(32'h3b04bd45),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb712caf9),
	.w1(32'hbaa5e0d2),
	.w2(32'h3b686464),
	.w3(32'hbbb80cf5),
	.w4(32'h39c5e9e1),
	.w5(32'h3a7754d6),
	.w6(32'hba9bb02a),
	.w7(32'hbc287e88),
	.w8(32'hbc331a3a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c46a5),
	.w1(32'hbb76959a),
	.w2(32'hbbd31e7b),
	.w3(32'h3c44bae7),
	.w4(32'hbc177fb0),
	.w5(32'hbad319d9),
	.w6(32'hbbd57df1),
	.w7(32'hbb5a0f6a),
	.w8(32'h3b08525d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ea258),
	.w1(32'h3bcc622e),
	.w2(32'h395ad816),
	.w3(32'h3c2ef6a7),
	.w4(32'h3c0ba8fe),
	.w5(32'hbab59c13),
	.w6(32'hbb1b944a),
	.w7(32'hba3ce747),
	.w8(32'hbb507b71),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc18b41),
	.w1(32'h3c85bdef),
	.w2(32'h3b8b1491),
	.w3(32'hbbf86f39),
	.w4(32'h3c376dd8),
	.w5(32'h3a6786ce),
	.w6(32'h3aa72d47),
	.w7(32'h3c59ca21),
	.w8(32'hbbb873a7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb906a1),
	.w1(32'h3a3d2015),
	.w2(32'h3b1e61af),
	.w3(32'hb9669177),
	.w4(32'h3ab6bc16),
	.w5(32'h3a3dd6d7),
	.w6(32'h3b8c20a6),
	.w7(32'hba139219),
	.w8(32'h39a7a7cc),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fd4cd),
	.w1(32'hbc711f6b),
	.w2(32'hbc6a7a1b),
	.w3(32'hbb299a54),
	.w4(32'hbc856c63),
	.w5(32'hbc71bb86),
	.w6(32'h3b83d0f7),
	.w7(32'h3bea1f8f),
	.w8(32'h3cb5d2e9),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc910b4c),
	.w1(32'hbc02f4ab),
	.w2(32'h3b51c55e),
	.w3(32'hbbeea452),
	.w4(32'hbbe2f61a),
	.w5(32'hbbc856cd),
	.w6(32'h3c3c2384),
	.w7(32'h3b071e7f),
	.w8(32'hbb8492d8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c98d2),
	.w1(32'hbc3caa9e),
	.w2(32'hbc39bf4c),
	.w3(32'hbb568e51),
	.w4(32'h3b5572e5),
	.w5(32'hba5f1d50),
	.w6(32'h3b5aa7be),
	.w7(32'hbb50e934),
	.w8(32'h3bdee4b9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ce42f),
	.w1(32'hbbb0a878),
	.w2(32'h3a2d793c),
	.w3(32'hbc1512ac),
	.w4(32'hbb878d9a),
	.w5(32'hbbc281fc),
	.w6(32'h3c2352aa),
	.w7(32'h3b394cdf),
	.w8(32'hb9238908),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f129d),
	.w1(32'h3baa9b27),
	.w2(32'h3b408037),
	.w3(32'hba8f324f),
	.w4(32'h3bddf733),
	.w5(32'h3bfda85d),
	.w6(32'h3c11dbab),
	.w7(32'h3a1c2b0e),
	.w8(32'hbba4179a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba87ed4),
	.w1(32'hbc6449a5),
	.w2(32'h3bd67dcd),
	.w3(32'h3c800486),
	.w4(32'hbb329c0c),
	.w5(32'h3cb77308),
	.w6(32'hba83ceb7),
	.w7(32'hbc896b85),
	.w8(32'hbbc3b0c4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eeac6),
	.w1(32'hbc2e9a48),
	.w2(32'hbc00da46),
	.w3(32'h3c424fba),
	.w4(32'hbba1584f),
	.w5(32'hbade1470),
	.w6(32'hbbcc7057),
	.w7(32'hbb830d5f),
	.w8(32'hbae6ccce),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b856e39),
	.w1(32'hbb63aa8a),
	.w2(32'hbc089f1d),
	.w3(32'h3b6141f2),
	.w4(32'hbbb1cad9),
	.w5(32'hbc6a5aec),
	.w6(32'hb8ef8322),
	.w7(32'h3b4fdbf4),
	.w8(32'hbad86769),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dc7fe),
	.w1(32'hbc14b4be),
	.w2(32'hba149e0f),
	.w3(32'hbbf47c3d),
	.w4(32'hbbebdd52),
	.w5(32'hbc349211),
	.w6(32'hbab535e4),
	.w7(32'hbc47b5f5),
	.w8(32'hbc0a2df5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a702ea0),
	.w1(32'hbb88bade),
	.w2(32'hbb6f9fba),
	.w3(32'hbc13763c),
	.w4(32'hbb6f43bb),
	.w5(32'hba575f94),
	.w6(32'hbb0cb75e),
	.w7(32'h3b106b70),
	.w8(32'hbc1dca75),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cd9fc),
	.w1(32'hbc9fbfcc),
	.w2(32'hbccf5f6c),
	.w3(32'h3b1adbd5),
	.w4(32'hba9c614d),
	.w5(32'h3afaf2ac),
	.w6(32'hbbe8d508),
	.w7(32'h3c8e876b),
	.w8(32'h3d028f42),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd0c075),
	.w1(32'h3bd25e4b),
	.w2(32'h3beadb71),
	.w3(32'h3bbb406d),
	.w4(32'h3b9d62d0),
	.w5(32'h3b1bc18d),
	.w6(32'h3cc81fba),
	.w7(32'h3b20ee61),
	.w8(32'hbbec8268),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcd872),
	.w1(32'hbbfdb85b),
	.w2(32'h39a26921),
	.w3(32'hbb00745e),
	.w4(32'hbbed11ad),
	.w5(32'hbc02b4d0),
	.w6(32'h3aea3e2e),
	.w7(32'hbbda97cc),
	.w8(32'hbbbb75e8),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33c2c2),
	.w1(32'hbc178ac8),
	.w2(32'h3b12143f),
	.w3(32'hbba80889),
	.w4(32'h3bdd1f0e),
	.w5(32'h3c8e66f8),
	.w6(32'hba82d1e9),
	.w7(32'hbc6276f1),
	.w8(32'hbc36b6c8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d6896),
	.w1(32'hbc8a97de),
	.w2(32'hbb478688),
	.w3(32'hbc441fe9),
	.w4(32'h3c163d2b),
	.w5(32'h3cd3f563),
	.w6(32'hbbd3326e),
	.w7(32'hbc2404d8),
	.w8(32'hbb409026),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d2da2),
	.w1(32'h3bf25679),
	.w2(32'h3b189f41),
	.w3(32'h3c2fbb05),
	.w4(32'h3b35c60f),
	.w5(32'hbc2e42b5),
	.w6(32'h3b80e325),
	.w7(32'h3b1d4e26),
	.w8(32'hba8465e6),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24caec),
	.w1(32'h3ada24f5),
	.w2(32'h3a95a093),
	.w3(32'hbc042c5c),
	.w4(32'hbb3370f4),
	.w5(32'hbc73a990),
	.w6(32'hbb2f7100),
	.w7(32'h3b821512),
	.w8(32'h3c385558),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8721a8),
	.w1(32'h3b974350),
	.w2(32'hbbae5442),
	.w3(32'hbb6ed5e6),
	.w4(32'hb8a1869c),
	.w5(32'hba7b595f),
	.w6(32'h3c2a14c3),
	.w7(32'h3bdc31de),
	.w8(32'h3a82be09),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd66405),
	.w1(32'hbb8b65b6),
	.w2(32'h3bf93ae8),
	.w3(32'h3bc569a4),
	.w4(32'h3a704556),
	.w5(32'h3c3ecadc),
	.w6(32'h3bb90a1b),
	.w7(32'hbb526f84),
	.w8(32'hbbd4b737),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c2902),
	.w1(32'hbb863adc),
	.w2(32'hbbe658fb),
	.w3(32'h3b9794f7),
	.w4(32'h3bed4acc),
	.w5(32'h3c1cb646),
	.w6(32'hbb0e0560),
	.w7(32'hbbf7b60d),
	.w8(32'h3b2ba537),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39806705),
	.w1(32'hbb1cf405),
	.w2(32'h3c99404c),
	.w3(32'h3baf28ed),
	.w4(32'hbb4d66f3),
	.w5(32'h3bc557d2),
	.w6(32'h3befef07),
	.w7(32'h3b8d59ef),
	.w8(32'h3c3ca1f0),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980e381),
	.w1(32'hbb978815),
	.w2(32'hbb4fb34e),
	.w3(32'hb9f050d0),
	.w4(32'h3c645f3c),
	.w5(32'hbb2a0eea),
	.w6(32'h3c18e060),
	.w7(32'h3aa05cdb),
	.w8(32'h3abda58c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8ec31),
	.w1(32'hbc292116),
	.w2(32'hbc6f800e),
	.w3(32'h3b75ca57),
	.w4(32'hbbd2141e),
	.w5(32'hbb4b3c8a),
	.w6(32'h39322567),
	.w7(32'h3a5265ea),
	.w8(32'h3c42430c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c3e7f),
	.w1(32'hbc003996),
	.w2(32'hbc385201),
	.w3(32'h3b89b18a),
	.w4(32'hbb761919),
	.w5(32'hbbc24608),
	.w6(32'h3bcbd92f),
	.w7(32'h3bbe5e78),
	.w8(32'h3c16bbe0),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb18e2),
	.w1(32'h3bfd7bb7),
	.w2(32'h3c12e78e),
	.w3(32'hbad21cd0),
	.w4(32'hba15459d),
	.w5(32'h3bb33993),
	.w6(32'h3bc299c3),
	.w7(32'hb922ae10),
	.w8(32'hbaadba99),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10a405),
	.w1(32'h3aaa9c84),
	.w2(32'hbb744bfb),
	.w3(32'hbc1d6384),
	.w4(32'hbb85e115),
	.w5(32'hbc02f45f),
	.w6(32'hbc67fd0b),
	.w7(32'hbb189a43),
	.w8(32'hba54e2d5),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9043b7),
	.w1(32'hbc06e8f2),
	.w2(32'hbc1ab293),
	.w3(32'hbbcacefa),
	.w4(32'hbb81d353),
	.w5(32'h3bcc61a2),
	.w6(32'h3b08003c),
	.w7(32'hbb4f74d3),
	.w8(32'h3c9360a1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83f7fb),
	.w1(32'hbbc5896e),
	.w2(32'hbc36e588),
	.w3(32'h3be6c91b),
	.w4(32'h3bd629c5),
	.w5(32'h3c4cb131),
	.w6(32'h3c315504),
	.w7(32'hba6ec74f),
	.w8(32'h3ccd4ea4),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaecbb3),
	.w1(32'h3a31f6c6),
	.w2(32'h3bfa5c29),
	.w3(32'h3af743f6),
	.w4(32'hbabf6a21),
	.w5(32'hbbd735d5),
	.w6(32'h3cb2133f),
	.w7(32'hbba314a0),
	.w8(32'h3b1afb91),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0791f9),
	.w1(32'h38d468e8),
	.w2(32'hbb533c9f),
	.w3(32'hbb164df3),
	.w4(32'hbb10c874),
	.w5(32'hbbeba474),
	.w6(32'h3a8e0051),
	.w7(32'hbba96bf0),
	.w8(32'hbc269c0e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f2f8e),
	.w1(32'h3b13a25c),
	.w2(32'h3c1ba8e9),
	.w3(32'h3b167583),
	.w4(32'h3b8ca0a8),
	.w5(32'hbb4e3f43),
	.w6(32'hbb9a8a2b),
	.w7(32'hbc503eff),
	.w8(32'hbcac5186),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd30f33),
	.w1(32'hbaeb804d),
	.w2(32'h3b2241b0),
	.w3(32'hbbf5d0dc),
	.w4(32'hba840a1e),
	.w5(32'h3cfa8dca),
	.w6(32'hbc3d139c),
	.w7(32'hbc456a0d),
	.w8(32'hbca71433),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10a40e),
	.w1(32'hbafa476d),
	.w2(32'hbbfcaae3),
	.w3(32'h3b849a5a),
	.w4(32'hbbdb7e64),
	.w5(32'hbc2af21c),
	.w6(32'hbbf61bc8),
	.w7(32'h3b809007),
	.w8(32'hb9d899ad),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a312f),
	.w1(32'h3a53706b),
	.w2(32'hb9de8c0b),
	.w3(32'h3c5195ad),
	.w4(32'hbb3066c5),
	.w5(32'hba8dc11e),
	.w6(32'h3b507423),
	.w7(32'h3b555388),
	.w8(32'h3b7afcea),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14ed57),
	.w1(32'hbb963091),
	.w2(32'hbb957bfb),
	.w3(32'h3bcb2710),
	.w4(32'h3be67ae6),
	.w5(32'h3c0c31b0),
	.w6(32'h3b9d50ff),
	.w7(32'h3b494f7a),
	.w8(32'h3bb189b1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d87bd),
	.w1(32'hbc8c6ab6),
	.w2(32'hbca81372),
	.w3(32'hba1cea4c),
	.w4(32'hb869d6ad),
	.w5(32'hbc130304),
	.w6(32'hbb13cad7),
	.w7(32'h3cba5081),
	.w8(32'h3ccb2d33),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd9adf1),
	.w1(32'hbbab5775),
	.w2(32'h3b4cb004),
	.w3(32'hbc4a33ab),
	.w4(32'h399120a4),
	.w5(32'h3c86133d),
	.w6(32'h3c8c664b),
	.w7(32'hbca571a5),
	.w8(32'hbc7c604e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa87e5b),
	.w1(32'h3a4c8ca8),
	.w2(32'h3a8d7467),
	.w3(32'h3c2ded66),
	.w4(32'hb9b0ffbb),
	.w5(32'hbbc1d6e9),
	.w6(32'hbc35dbc2),
	.w7(32'h39bbc0de),
	.w8(32'hb99c8089),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e1fce),
	.w1(32'hba957c68),
	.w2(32'hbb574f9e),
	.w3(32'h3c4a1318),
	.w4(32'h3bb0d6f1),
	.w5(32'h3b299aee),
	.w6(32'h3ae98a7c),
	.w7(32'h3b0a84ec),
	.w8(32'hba62d41d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5b981),
	.w1(32'hbbee7f57),
	.w2(32'hbc0639a7),
	.w3(32'h399c4c86),
	.w4(32'hbb459222),
	.w5(32'h3a0e2f24),
	.w6(32'h3a760ec1),
	.w7(32'h3b4239fa),
	.w8(32'h3c03e2b8),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ab0d1),
	.w1(32'hbaf1bd41),
	.w2(32'h3bb67ff7),
	.w3(32'h3b7e45a3),
	.w4(32'hbb3a71b9),
	.w5(32'h3942d0f0),
	.w6(32'h3c21181e),
	.w7(32'hbc33541b),
	.w8(32'hbc0fa007),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a941d5b),
	.w1(32'h3a7aac17),
	.w2(32'hbb329830),
	.w3(32'hbba8478d),
	.w4(32'h3bcaf3c2),
	.w5(32'h3bc609ee),
	.w6(32'hbbf39e10),
	.w7(32'h3b5dabf0),
	.w8(32'h3b32cca1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51ec32),
	.w1(32'hbc525ad3),
	.w2(32'hbbd5d5b3),
	.w3(32'h3a47b459),
	.w4(32'h3b0af7ac),
	.w5(32'h3c3f9449),
	.w6(32'h3bfcd208),
	.w7(32'h3c28796c),
	.w8(32'h3d096429),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc279fcb),
	.w1(32'hbb803d17),
	.w2(32'hbba132cd),
	.w3(32'h3c1e78d3),
	.w4(32'hbb8ced8f),
	.w5(32'hbbe3d804),
	.w6(32'h3ca50eec),
	.w7(32'hbb400487),
	.w8(32'h3b97e423),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb05125),
	.w1(32'hbc324244),
	.w2(32'hbbacc446),
	.w3(32'h3c41fdd4),
	.w4(32'hbc2b320c),
	.w5(32'hbc8dbe28),
	.w6(32'h3c3cb764),
	.w7(32'hbc131827),
	.w8(32'hbb9e82f2),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ec3f1),
	.w1(32'hbc21f9ab),
	.w2(32'h3a9389ec),
	.w3(32'hbbc4235f),
	.w4(32'hbbfbd46c),
	.w5(32'hbb12fef4),
	.w6(32'hbba68130),
	.w7(32'h3ba517d0),
	.w8(32'h3c13c634),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule