module layer_8_featuremap_212(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0b789),
	.w1(32'h3a8c7031),
	.w2(32'hbb861a67),
	.w3(32'h3c0c5c24),
	.w4(32'h3a894f9d),
	.w5(32'hbc1bfdf9),
	.w6(32'h3ba370d5),
	.w7(32'h3c1ab0ea),
	.w8(32'h3c2e7777),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a930714),
	.w1(32'h3b979cb1),
	.w2(32'h3b569410),
	.w3(32'hbb86163a),
	.w4(32'h3b3fbdb7),
	.w5(32'h3b1f9ce0),
	.w6(32'h3b160030),
	.w7(32'hb93641ef),
	.w8(32'hbb07eb9d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf24938),
	.w1(32'h3baa63be),
	.w2(32'hb99b49e4),
	.w3(32'h3b5007a6),
	.w4(32'h3b4d966d),
	.w5(32'hbb0349c1),
	.w6(32'h3c6daebf),
	.w7(32'h3c630d91),
	.w8(32'h3bdfbb00),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385924f8),
	.w1(32'hbca62d54),
	.w2(32'hbc3736c0),
	.w3(32'hbc0e5e05),
	.w4(32'hbb86bc63),
	.w5(32'hbc8586cc),
	.w6(32'hb9a97954),
	.w7(32'hbb78dbf9),
	.w8(32'hbb3ef7d9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5784e),
	.w1(32'h3aafecc7),
	.w2(32'h3bb4d877),
	.w3(32'hbc3b9498),
	.w4(32'h3a3c6301),
	.w5(32'h385ab86d),
	.w6(32'h37cecbdc),
	.w7(32'h3ae82b0c),
	.w8(32'h394b0c08),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad61fe1),
	.w1(32'hbc486247),
	.w2(32'h3b0ca40e),
	.w3(32'h3b2028db),
	.w4(32'h3b7bba6b),
	.w5(32'h3b6d882b),
	.w6(32'hbc7b8b2d),
	.w7(32'hbb892271),
	.w8(32'hbb76edcb),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2aa29),
	.w1(32'hbaa75dca),
	.w2(32'hb977449a),
	.w3(32'h3c029b7e),
	.w4(32'h3ab43ed4),
	.w5(32'hba64448d),
	.w6(32'h3a55847f),
	.w7(32'hbac16b02),
	.w8(32'hbb1d5630),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e6c48),
	.w1(32'h3ba26961),
	.w2(32'h3c339b32),
	.w3(32'h3c1c5307),
	.w4(32'h3bca94f6),
	.w5(32'hb98dfc17),
	.w6(32'h3c6c221b),
	.w7(32'h3cae5a2c),
	.w8(32'h3c258c7e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9635a),
	.w1(32'h3a7d7a0f),
	.w2(32'h3bb38123),
	.w3(32'hbb8a26b2),
	.w4(32'hbb62fc23),
	.w5(32'hbb323ef5),
	.w6(32'h3c6cd94c),
	.w7(32'h3c5abe75),
	.w8(32'h3c2356ea),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca00888),
	.w1(32'h3c5af1eb),
	.w2(32'h3b8fe523),
	.w3(32'h3bf7eaf7),
	.w4(32'hba91eb85),
	.w5(32'hba57aec0),
	.w6(32'h3c6fa206),
	.w7(32'h3c42fbb3),
	.w8(32'hbc26aaff),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c2400),
	.w1(32'h3c8bc7bf),
	.w2(32'hbcd60261),
	.w3(32'hbb74c680),
	.w4(32'h3ccbf2c9),
	.w5(32'hbbf02e6d),
	.w6(32'hbbe37974),
	.w7(32'hbcc36db8),
	.w8(32'hbc295610),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce7b084),
	.w1(32'hbb19a344),
	.w2(32'hbc02aca3),
	.w3(32'hbccab8e9),
	.w4(32'hbbdde58d),
	.w5(32'hbc45b939),
	.w6(32'hba1aa9b2),
	.w7(32'hbaae577e),
	.w8(32'hbb9fed9a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06c699),
	.w1(32'h3c71f526),
	.w2(32'h3b71be9b),
	.w3(32'hbbd068e3),
	.w4(32'hbb65d0c7),
	.w5(32'hbc0a6e24),
	.w6(32'h3c65f8cc),
	.w7(32'h3c5e72cc),
	.w8(32'hbc19213f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc704bbb),
	.w1(32'h3c0f7655),
	.w2(32'h38de1c89),
	.w3(32'hbc5fe2d2),
	.w4(32'h3bb7d219),
	.w5(32'h3c82a259),
	.w6(32'h3b717ba6),
	.w7(32'h3a78741d),
	.w8(32'hbb9b7a17),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be59266),
	.w1(32'hbba5cacb),
	.w2(32'hbb2e0ce1),
	.w3(32'h3bc160c5),
	.w4(32'hbb704853),
	.w5(32'hbb8a2bb0),
	.w6(32'hba217f3e),
	.w7(32'hbb0f05a2),
	.w8(32'h3b20ffc1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eaef6),
	.w1(32'h3bcf3d15),
	.w2(32'hbb92f073),
	.w3(32'h3b8db842),
	.w4(32'h3c001c1b),
	.w5(32'h39eb4d40),
	.w6(32'h38f2f489),
	.w7(32'h3ab2a641),
	.w8(32'hbbe4acb7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4638ae),
	.w1(32'hbc10b93d),
	.w2(32'h3b890a74),
	.w3(32'hbafe3cfe),
	.w4(32'hbadf820f),
	.w5(32'hbac32a60),
	.w6(32'hbb870f7f),
	.w7(32'h3bb695a3),
	.w8(32'h3baaf9ff),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cbf09),
	.w1(32'hbb506b10),
	.w2(32'h3ae44e3f),
	.w3(32'h3c2d1cd0),
	.w4(32'h3c4ff798),
	.w5(32'h3c0e7433),
	.w6(32'hbb9a53f1),
	.w7(32'hbbe5c7f4),
	.w8(32'h3be5a309),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceb9847),
	.w1(32'h3baa5e3d),
	.w2(32'h3c1af39e),
	.w3(32'hb90f236a),
	.w4(32'h3c10157e),
	.w5(32'h3ccb318b),
	.w6(32'hbd4270fd),
	.w7(32'hbc690a38),
	.w8(32'hbc6e014b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9393b),
	.w1(32'h3c6a486c),
	.w2(32'h3c3513d7),
	.w3(32'h3b45217a),
	.w4(32'h3c59476b),
	.w5(32'h3c0d0b2c),
	.w6(32'hbbcb64ec),
	.w7(32'hbbb18373),
	.w8(32'hbba42e1d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ee965),
	.w1(32'h3c24db6f),
	.w2(32'h3b7ab472),
	.w3(32'h3b857156),
	.w4(32'h3c2dcc05),
	.w5(32'h3c3373fc),
	.w6(32'hba8fc994),
	.w7(32'h3aeb41b4),
	.w8(32'h3c028010),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c076c3c),
	.w1(32'h3c6a4e91),
	.w2(32'h3cf00d37),
	.w3(32'h3c16cd87),
	.w4(32'h3c8aa786),
	.w5(32'h3cc536a0),
	.w6(32'h3c969a59),
	.w7(32'h3c8b9ce2),
	.w8(32'h3c19932e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a1369),
	.w1(32'h3caab819),
	.w2(32'hbb716af9),
	.w3(32'h3b8d6062),
	.w4(32'h3cfa378e),
	.w5(32'hbb996a08),
	.w6(32'hbbd49230),
	.w7(32'hbb52b49b),
	.w8(32'hbc75c622),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4d2ca),
	.w1(32'h3c890d03),
	.w2(32'h3c83ac20),
	.w3(32'hbca1c8a9),
	.w4(32'h3c364a59),
	.w5(32'h3c814132),
	.w6(32'h3c052b1b),
	.w7(32'h3c174711),
	.w8(32'h3ba19fba),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c129bb4),
	.w1(32'hbb3d8609),
	.w2(32'hbbfb5594),
	.w3(32'h3c0aae0f),
	.w4(32'h3b0f2cee),
	.w5(32'h3ae85a9c),
	.w6(32'h3abaf84a),
	.w7(32'h3bada571),
	.w8(32'h3b1186bc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb584fd6),
	.w1(32'h3c61ad7f),
	.w2(32'h3a6b9d84),
	.w3(32'hbb657968),
	.w4(32'h3b614bd2),
	.w5(32'h3a563b83),
	.w6(32'hbafe8aba),
	.w7(32'hbad41d28),
	.w8(32'h3b19c576),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4761f7),
	.w1(32'h3afa7812),
	.w2(32'h3ad5ded0),
	.w3(32'h3b6bdd6e),
	.w4(32'h3c21bf47),
	.w5(32'h3aed4bf6),
	.w6(32'h3bb3e34f),
	.w7(32'h3a802f99),
	.w8(32'h3b7f0f8b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c3aab),
	.w1(32'h3cffa1ef),
	.w2(32'h3c38560f),
	.w3(32'hbb8828fd),
	.w4(32'hbcfef90d),
	.w5(32'hbd28dc5a),
	.w6(32'hbdde1288),
	.w7(32'hbdd58596),
	.w8(32'h3c0f9a2e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb882d0b),
	.w1(32'h3c69b36b),
	.w2(32'hbc06f1bb),
	.w3(32'hbc44875b),
	.w4(32'h3c8414e1),
	.w5(32'hbb2e3968),
	.w6(32'h3c1a359a),
	.w7(32'hbb33ca53),
	.w8(32'h3ba612db),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91fff4b),
	.w1(32'hbacb5cc7),
	.w2(32'hbb2cc298),
	.w3(32'h3ba59eef),
	.w4(32'hbbfe6cd4),
	.w5(32'hbc6b7c6d),
	.w6(32'h3a7da96b),
	.w7(32'hbac35e25),
	.w8(32'h3c27e5eb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf3ecf),
	.w1(32'h3c7bbf09),
	.w2(32'h39c3527e),
	.w3(32'hbb71e247),
	.w4(32'hbb89b4a7),
	.w5(32'hbbcac5fe),
	.w6(32'h3c4f8978),
	.w7(32'h3c1f35fc),
	.w8(32'hb8ac243b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08d70a),
	.w1(32'h3cf7840d),
	.w2(32'h3c5cfbe5),
	.w3(32'hba94f894),
	.w4(32'h3c38216a),
	.w5(32'h3b901dcf),
	.w6(32'h3c772855),
	.w7(32'h3c0f9394),
	.w8(32'h3ae786ac),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ac811),
	.w1(32'hbbe54f25),
	.w2(32'h3af1f2f5),
	.w3(32'hbc02c82f),
	.w4(32'h3c2066f8),
	.w5(32'h3bd2d1d9),
	.w6(32'h3acdaea3),
	.w7(32'hbbd7573a),
	.w8(32'hbbc0de50),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb44f9),
	.w1(32'hba614b2a),
	.w2(32'hbb89c81f),
	.w3(32'hbc1e070f),
	.w4(32'h3b846804),
	.w5(32'hb92065d4),
	.w6(32'hbc19166e),
	.w7(32'hbc0401ec),
	.w8(32'hbbc86bae),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71d937),
	.w1(32'hbc2a1e2c),
	.w2(32'hbc5a34a8),
	.w3(32'hb9eddf0f),
	.w4(32'hbc10eb9d),
	.w5(32'hbc3d4595),
	.w6(32'hbb644377),
	.w7(32'hbbd189c8),
	.w8(32'hbbb54994),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c0961),
	.w1(32'h3c76d0cd),
	.w2(32'h3c06f9a0),
	.w3(32'hbbc63687),
	.w4(32'h3ba53e99),
	.w5(32'h3c0e6f25),
	.w6(32'hbc3249d3),
	.w7(32'hba79493d),
	.w8(32'h3bf2ba17),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39b928),
	.w1(32'hbc3ec38c),
	.w2(32'hbc8e11bd),
	.w3(32'h3b98c2a2),
	.w4(32'hbbe31430),
	.w5(32'hbc6887c2),
	.w6(32'hbb59b06c),
	.w7(32'hbb9d77d9),
	.w8(32'h3c3b220b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb911a6),
	.w1(32'hbc48fe02),
	.w2(32'h3abc7b84),
	.w3(32'hbae386ce),
	.w4(32'hbc4d4b1f),
	.w5(32'hbb84ab6e),
	.w6(32'hbbe35bdf),
	.w7(32'hbb489255),
	.w8(32'h3baea9a6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c246a5b),
	.w1(32'h3c45e44c),
	.w2(32'h3bf757e2),
	.w3(32'h3bea811e),
	.w4(32'h3b593cfc),
	.w5(32'hbbc7822a),
	.w6(32'h3c2e8ec2),
	.w7(32'hbb8473ea),
	.w8(32'hbb454f9b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f8ab5),
	.w1(32'hbb18591d),
	.w2(32'hbaa000a9),
	.w3(32'hbbc433fd),
	.w4(32'h3a358dea),
	.w5(32'h3b49a542),
	.w6(32'h3a9b41f7),
	.w7(32'h3a672a32),
	.w8(32'hbb7d8ca5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d1abf),
	.w1(32'hbc448a9b),
	.w2(32'hbc1de85a),
	.w3(32'hbbca51e4),
	.w4(32'hbc5075aa),
	.w5(32'hbbd28291),
	.w6(32'hbc86d345),
	.w7(32'hbc4fb45f),
	.w8(32'hbabd8073),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6be0a),
	.w1(32'h3b9fbd2c),
	.w2(32'h3bc40ddd),
	.w3(32'hbb5e8905),
	.w4(32'h3c04cfae),
	.w5(32'h3c1ae258),
	.w6(32'hbc0c14f5),
	.w7(32'hbb797c76),
	.w8(32'hbc6a18c4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22408a),
	.w1(32'hbc03f00a),
	.w2(32'hbcbe1acb),
	.w3(32'hbc3f1985),
	.w4(32'h3bc695f2),
	.w5(32'hbc8c4781),
	.w6(32'h3a6c0273),
	.w7(32'hbb98beb0),
	.w8(32'h3b982055),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08f9b9),
	.w1(32'h3c8a2bac),
	.w2(32'h3c85303d),
	.w3(32'hbb63b2d8),
	.w4(32'h3c855693),
	.w5(32'h3c8b18ca),
	.w6(32'h3b8b8cf9),
	.w7(32'hbb237491),
	.w8(32'hbaa47613),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d9f2f),
	.w1(32'hbb24837e),
	.w2(32'hbc699212),
	.w3(32'hbaa2691f),
	.w4(32'h3ac8ce5c),
	.w5(32'hbb534034),
	.w6(32'hbc17d674),
	.w7(32'hbb44da51),
	.w8(32'h3a94f2cc),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45f726),
	.w1(32'h3b0a86d0),
	.w2(32'hbb908db3),
	.w3(32'h3c5e4ef9),
	.w4(32'h3b258294),
	.w5(32'hbb2beb99),
	.w6(32'h3bbc42a9),
	.w7(32'hbad54b6f),
	.w8(32'h3a8e1b86),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31f06b),
	.w1(32'h3c44b2d4),
	.w2(32'hba345a3f),
	.w3(32'h3b7f56ab),
	.w4(32'h3c4a4598),
	.w5(32'hba8e5d9f),
	.w6(32'hbab6bdc9),
	.w7(32'hbbfae27d),
	.w8(32'hbc7bbb6c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fd4eb),
	.w1(32'h3c9135c6),
	.w2(32'h3bc8ac41),
	.w3(32'hbb503df1),
	.w4(32'h3c527794),
	.w5(32'h3c46a550),
	.w6(32'hbbb4bb61),
	.w7(32'h3aab47d3),
	.w8(32'h3afdca35),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88bd55),
	.w1(32'h3c41aab4),
	.w2(32'h3c54875f),
	.w3(32'h3c8cf420),
	.w4(32'h3c7904ff),
	.w5(32'hb6f87576),
	.w6(32'h3afa907d),
	.w7(32'h3b3f6cb2),
	.w8(32'h3a67927d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ffcfa),
	.w1(32'hbc13fda1),
	.w2(32'hbca8a1f9),
	.w3(32'hbb9e9702),
	.w4(32'hbb828d7d),
	.w5(32'hbc949f33),
	.w6(32'hbc5acc24),
	.w7(32'hbc364119),
	.w8(32'hbc3c8403),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc061a3b),
	.w1(32'hbbb6dd5a),
	.w2(32'hbc450a37),
	.w3(32'hbbf8ee31),
	.w4(32'hbc1f126e),
	.w5(32'hbc3c10aa),
	.w6(32'h3b61baad),
	.w7(32'hbc02b65c),
	.w8(32'hbc1eea4f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a885dd0),
	.w1(32'h3901af9e),
	.w2(32'hbb8d381c),
	.w3(32'h3c5ba45e),
	.w4(32'h3c5fbdf1),
	.w5(32'h3c40f1aa),
	.w6(32'hbcd6953c),
	.w7(32'hbbb36a9f),
	.w8(32'hbcb44018),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ded8c),
	.w1(32'hbb69687c),
	.w2(32'hbba4f9cb),
	.w3(32'h3c3da0fa),
	.w4(32'h3b1ca9be),
	.w5(32'hbb6ab8a6),
	.w6(32'hbbcdaef4),
	.w7(32'hbbc1ca7e),
	.w8(32'hbb8715cd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccec8f),
	.w1(32'hbbb25267),
	.w2(32'h3b076b94),
	.w3(32'h3b4f54eb),
	.w4(32'hbc0ac5cf),
	.w5(32'h3c68a3d5),
	.w6(32'hbb3daec3),
	.w7(32'h3bb2bb5b),
	.w8(32'h3b090492),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb1d4e),
	.w1(32'hbc8d0f36),
	.w2(32'h3c72e704),
	.w3(32'h3ac25593),
	.w4(32'hbc35b19e),
	.w5(32'h3c923b03),
	.w6(32'hbc75bbe2),
	.w7(32'hbb142717),
	.w8(32'hbb8b3d88),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c2cda),
	.w1(32'h3c755c2e),
	.w2(32'hba0e9738),
	.w3(32'h3b566a5f),
	.w4(32'h3bca79fc),
	.w5(32'hb9d059ef),
	.w6(32'hbc493b03),
	.w7(32'hbbf389b2),
	.w8(32'h3b78a294),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb1c7b),
	.w1(32'hbc0e50be),
	.w2(32'hbc9c0dd7),
	.w3(32'hbb413478),
	.w4(32'h3bc2056b),
	.w5(32'hbc4a0347),
	.w6(32'hbbd02940),
	.w7(32'hbc6f201f),
	.w8(32'hbc044c85),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b5793),
	.w1(32'hbc5bff4b),
	.w2(32'hbcb4990f),
	.w3(32'h3b5a5c5a),
	.w4(32'hbb2c6371),
	.w5(32'hbc818abf),
	.w6(32'hbbf09889),
	.w7(32'hbb42caef),
	.w8(32'h3c734cf1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bade804),
	.w1(32'h3b821b1a),
	.w2(32'h3b074c96),
	.w3(32'h3c1a7a9b),
	.w4(32'h3c00b64b),
	.w5(32'h3b26b95d),
	.w6(32'hbb08ecd5),
	.w7(32'h39c5e1e8),
	.w8(32'h3ae787e9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a2fc5),
	.w1(32'h3bc4d0ff),
	.w2(32'hbb367c83),
	.w3(32'h3b9e0739),
	.w4(32'h3b139515),
	.w5(32'h3ad29688),
	.w6(32'h3aa23c0b),
	.w7(32'hbb63f9c5),
	.w8(32'hbc0eb02a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd6990),
	.w1(32'h3bb8ce6b),
	.w2(32'h3bb9708a),
	.w3(32'h3c21f75a),
	.w4(32'h3bebef7b),
	.w5(32'h3b5122b4),
	.w6(32'h3bca64e4),
	.w7(32'hb9817b1a),
	.w8(32'h39c207b3),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04b15a),
	.w1(32'hbc4deb94),
	.w2(32'hbc2dce1b),
	.w3(32'hbbaa797b),
	.w4(32'hb9eae3bf),
	.w5(32'hbb9ad702),
	.w6(32'hbb1275f1),
	.w7(32'h3a6a2e9a),
	.w8(32'h3c6636e1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c5149),
	.w1(32'hbb23b506),
	.w2(32'hbb95c25a),
	.w3(32'hbc311d00),
	.w4(32'h3b28792c),
	.w5(32'hba3e761c),
	.w6(32'h3b256985),
	.w7(32'h3bca1df8),
	.w8(32'h3c9b6129),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90f50e),
	.w1(32'hbc1a38f6),
	.w2(32'hbbfb4a2c),
	.w3(32'h3c8b77db),
	.w4(32'hbbf67aa0),
	.w5(32'hbbbcd3d0),
	.w6(32'hbbb56865),
	.w7(32'hbb0421b9),
	.w8(32'hbbd8b846),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc569634),
	.w1(32'h3b85e98d),
	.w2(32'h3aacba9a),
	.w3(32'hbc661ada),
	.w4(32'h3bf75b5b),
	.w5(32'h3b721f1c),
	.w6(32'hba8e4d5a),
	.w7(32'hbb3b99ca),
	.w8(32'hbba5cb5b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f93f),
	.w1(32'h3ba551dc),
	.w2(32'h3b30b77e),
	.w3(32'h3ade9c4f),
	.w4(32'h3b7dcdfe),
	.w5(32'h3c3bd175),
	.w6(32'h39e94679),
	.w7(32'h3a3d2b7e),
	.w8(32'h3aa881eb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf80949),
	.w1(32'hbc1783e5),
	.w2(32'hbb04d4a7),
	.w3(32'h3c07a582),
	.w4(32'h3a9c04f3),
	.w5(32'h39d7f751),
	.w6(32'h3b3c716e),
	.w7(32'hbad39d4b),
	.w8(32'h3b1648f6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d82b7),
	.w1(32'h3bbc2c22),
	.w2(32'hbc68a73f),
	.w3(32'hbabb841b),
	.w4(32'hba3a434f),
	.w5(32'hbbf54b8f),
	.w6(32'h3bf0e255),
	.w7(32'hba97b7b7),
	.w8(32'hbb2f8e50),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa55fe),
	.w1(32'hbae183a1),
	.w2(32'h3b0d53db),
	.w3(32'hbad8f3d7),
	.w4(32'h3c6b77c7),
	.w5(32'h3bf8fad3),
	.w6(32'hbb2b30ac),
	.w7(32'hbbe1e1b8),
	.w8(32'hbb9f4995),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63f422),
	.w1(32'h3c650e97),
	.w2(32'hb941e966),
	.w3(32'h3c00ecf5),
	.w4(32'h3c13f4a0),
	.w5(32'hbaf0f575),
	.w6(32'hbcefcddd),
	.w7(32'hbce7a2d7),
	.w8(32'hbc96f596),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d93d1),
	.w1(32'hbc8e38e2),
	.w2(32'h3c7bfc97),
	.w3(32'hbc2dbaad),
	.w4(32'hbcad3a3c),
	.w5(32'h3c5fe6c0),
	.w6(32'hbbcab90c),
	.w7(32'h3c18acd7),
	.w8(32'hbb81d52c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8468ae),
	.w1(32'h3c6c8908),
	.w2(32'h3c55895b),
	.w3(32'h3c631e15),
	.w4(32'h3c3f091b),
	.w5(32'h3bb2eaf5),
	.w6(32'hbb884f3b),
	.w7(32'h3ab126ac),
	.w8(32'hbb8beb58),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98152b),
	.w1(32'h3b03c616),
	.w2(32'h3c1e94fc),
	.w3(32'h3bdf2d71),
	.w4(32'h3b39e88f),
	.w5(32'h3bd69957),
	.w6(32'hbaac82d9),
	.w7(32'hbadf2934),
	.w8(32'hbae9b0ae),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7be2f3),
	.w1(32'h3bf1fa2c),
	.w2(32'hbc0005db),
	.w3(32'hbb2fb8c7),
	.w4(32'hbb11bb57),
	.w5(32'hbb6c44cf),
	.w6(32'h3b844058),
	.w7(32'h3b745dc0),
	.w8(32'h3b2bd420),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8db950),
	.w1(32'hbadd334c),
	.w2(32'h3c242698),
	.w3(32'hb9bddfd1),
	.w4(32'h3a4a3f57),
	.w5(32'h3c65283f),
	.w6(32'hbbfc2900),
	.w7(32'h3afd9b5e),
	.w8(32'hbb2a9b6e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39301f44),
	.w1(32'hbc2ad6be),
	.w2(32'hbc305578),
	.w3(32'h3ba418ff),
	.w4(32'hbc22adca),
	.w5(32'hbc38987f),
	.w6(32'hbc8145ae),
	.w7(32'hbc85df83),
	.w8(32'hbcf8256e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbaa865),
	.w1(32'h3b0a0959),
	.w2(32'hbc338fb1),
	.w3(32'hbc9f8cb8),
	.w4(32'h3b31f24c),
	.w5(32'hbacb99d1),
	.w6(32'h3a4fe8ed),
	.w7(32'hba7fa414),
	.w8(32'hba32e3b7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bca3a),
	.w1(32'h3b4c81f9),
	.w2(32'hbc9c0a2e),
	.w3(32'h3b4ec27a),
	.w4(32'h3bb9ef6f),
	.w5(32'hbc544ef4),
	.w6(32'hbcabbf1b),
	.w7(32'hbc89a803),
	.w8(32'hbc0607ed),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49b776),
	.w1(32'h3b77038e),
	.w2(32'h3c468b88),
	.w3(32'hbc3163b8),
	.w4(32'h3c07503f),
	.w5(32'h3c612198),
	.w6(32'hbaa42132),
	.w7(32'h3c00104e),
	.w8(32'hbb903490),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf01540),
	.w1(32'h3c26fd19),
	.w2(32'h3988ac50),
	.w3(32'hbba17b24),
	.w4(32'h3c633667),
	.w5(32'h3bab42d1),
	.w6(32'h3b83ac31),
	.w7(32'hbbd36abc),
	.w8(32'h3b98a1b7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf27e94),
	.w1(32'hb9930ee8),
	.w2(32'h3bc81cd5),
	.w3(32'hbb0d6da1),
	.w4(32'h3b3e90a7),
	.w5(32'h3b682f66),
	.w6(32'hba31a232),
	.w7(32'h3ad5fd0a),
	.w8(32'hb8007c35),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c277e8a),
	.w1(32'h3c050713),
	.w2(32'h3c1e7a57),
	.w3(32'h3b6ed2cf),
	.w4(32'h3c94bfa8),
	.w5(32'h3ca8e278),
	.w6(32'hb9cac626),
	.w7(32'h3b46e539),
	.w8(32'hbba1f850),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2340c5),
	.w1(32'hb955908d),
	.w2(32'hbb186602),
	.w3(32'h3c57a68e),
	.w4(32'hbaebcea7),
	.w5(32'hbb100bc1),
	.w6(32'hbc3d1e64),
	.w7(32'hbc406b16),
	.w8(32'hbcbb8d1f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ec55a),
	.w1(32'hbcbe8d73),
	.w2(32'hbc9757f7),
	.w3(32'hbd1bc942),
	.w4(32'hbccf471a),
	.w5(32'h3b4ba02b),
	.w6(32'hbc857300),
	.w7(32'hbc81ebf0),
	.w8(32'hbca473f8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8ccdb),
	.w1(32'h3c0b54df),
	.w2(32'h3b6019cc),
	.w3(32'h3c327bd8),
	.w4(32'h3c0fcb63),
	.w5(32'h3b07a118),
	.w6(32'hbcdd7beb),
	.w7(32'hbc3cfc61),
	.w8(32'hbb87824e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3542c1),
	.w1(32'h391b2c55),
	.w2(32'hb692d8dc),
	.w3(32'hbbbaecc1),
	.w4(32'h3ae0b349),
	.w5(32'hbc0959cc),
	.w6(32'hbbf21bde),
	.w7(32'hbb803a2c),
	.w8(32'hba822239),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd13aea),
	.w1(32'h3c2af054),
	.w2(32'h3c00ae8a),
	.w3(32'hbc0583c8),
	.w4(32'h3bab969d),
	.w5(32'h3bde0d64),
	.w6(32'h3c3684ac),
	.w7(32'h3bf4016b),
	.w8(32'hbbf64515),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed8c36),
	.w1(32'h3bab19b9),
	.w2(32'hbbc8b40c),
	.w3(32'h3bf82349),
	.w4(32'h3ca361b6),
	.w5(32'h3b98e888),
	.w6(32'hbb452ce9),
	.w7(32'hbb923015),
	.w8(32'hb93bede8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2cfe5),
	.w1(32'h3bcb3b82),
	.w2(32'hba4d75ad),
	.w3(32'hbb98ba4b),
	.w4(32'h3b067c58),
	.w5(32'hbaef0161),
	.w6(32'h3c382069),
	.w7(32'h3b8712f6),
	.w8(32'hbba45ce4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd209fc),
	.w1(32'h3c4325d1),
	.w2(32'h3b564475),
	.w3(32'hb930da88),
	.w4(32'h3bddf196),
	.w5(32'hbb302de5),
	.w6(32'h3b946529),
	.w7(32'hbb830428),
	.w8(32'hbc1817c6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fd34f),
	.w1(32'hbbbd6a4d),
	.w2(32'hbaeee756),
	.w3(32'hbb25a56c),
	.w4(32'h3ab44a71),
	.w5(32'h3b8b4c16),
	.w6(32'h3a2cbe0a),
	.w7(32'hbba0e810),
	.w8(32'hbbbf6460),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba012dfe),
	.w1(32'hbba0fe74),
	.w2(32'hbbf733de),
	.w3(32'h3b9584a5),
	.w4(32'h3bb23e30),
	.w5(32'h3c1f88f5),
	.w6(32'hbba2c0f1),
	.w7(32'hbb566e5a),
	.w8(32'hbbe992ce),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb919315),
	.w1(32'h3aa76188),
	.w2(32'hb98dbbdd),
	.w3(32'h3c071d15),
	.w4(32'h3b627fa0),
	.w5(32'h3b42c5f2),
	.w6(32'hbada3c57),
	.w7(32'hbbb6022a),
	.w8(32'hbba4e4ea),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f182e),
	.w1(32'h3c756b78),
	.w2(32'h3bdf2cb0),
	.w3(32'h3bbd5072),
	.w4(32'h3c8440fb),
	.w5(32'h3c395d8a),
	.w6(32'h3ba9017b),
	.w7(32'h3aa9d8ac),
	.w8(32'hbb31bf54),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa984a5),
	.w1(32'hbb8ffa5f),
	.w2(32'hbd0353ab),
	.w3(32'hbab64bf8),
	.w4(32'h390c4a41),
	.w5(32'hbc8004ab),
	.w6(32'h3b835f29),
	.w7(32'hbbf89b87),
	.w8(32'hb980b469),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d942f),
	.w1(32'hbb11860e),
	.w2(32'hbc459512),
	.w3(32'hbc04e025),
	.w4(32'hbab902b2),
	.w5(32'hbb5e6d14),
	.w6(32'hba25c05e),
	.w7(32'hbaa9d7e0),
	.w8(32'h3c10dce6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba01921),
	.w1(32'hbb2558bb),
	.w2(32'hbc2d6628),
	.w3(32'h3c07dfc4),
	.w4(32'h3be93522),
	.w5(32'hb85dc36f),
	.w6(32'hbc865c51),
	.w7(32'hbca9ea8d),
	.w8(32'hbcd5bfff),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd62c30),
	.w1(32'h3c80a99a),
	.w2(32'h3c20caa5),
	.w3(32'h3c49d2d1),
	.w4(32'h3c2f0892),
	.w5(32'h3c2bcc2e),
	.w6(32'h3b734cb3),
	.w7(32'h3bda052c),
	.w8(32'hbba515d4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe481c6),
	.w1(32'h3c3b85f5),
	.w2(32'h3b4ea61d),
	.w3(32'hbbc2db68),
	.w4(32'h3c3d5ef8),
	.w5(32'h3ab98300),
	.w6(32'h3b4c0da9),
	.w7(32'hbb77c147),
	.w8(32'hbb5d30c4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf764e1),
	.w1(32'hbbed39d3),
	.w2(32'hbcaa9c68),
	.w3(32'h3b182a8b),
	.w4(32'hbbaaf10a),
	.w5(32'hbc950ad0),
	.w6(32'hbc227a23),
	.w7(32'hbc76e663),
	.w8(32'hbbb1b558),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc901a4e),
	.w1(32'hbc25be34),
	.w2(32'hbc961cb4),
	.w3(32'hbc6c87e0),
	.w4(32'hb62111fa),
	.w5(32'h3a5abbc6),
	.w6(32'hbb0dc46e),
	.w7(32'hbc696f4e),
	.w8(32'hbbf92ca6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca67e7e),
	.w1(32'hbbad1b96),
	.w2(32'h3658336e),
	.w3(32'h3912a4d4),
	.w4(32'h3ad0e1b8),
	.w5(32'hbb8e73ed),
	.w6(32'h3bbb83ff),
	.w7(32'h3b7bc8d4),
	.w8(32'h3bca6458),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b99d9),
	.w1(32'hbb4c401f),
	.w2(32'h3a1c32b4),
	.w3(32'h3b1000bc),
	.w4(32'h3bb8c608),
	.w5(32'h3c00c806),
	.w6(32'h3b26e189),
	.w7(32'hb98e43b1),
	.w8(32'hbba58534),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b885a27),
	.w1(32'h3c3bec62),
	.w2(32'h3a0c3f70),
	.w3(32'h3c9a49e9),
	.w4(32'h3b558816),
	.w5(32'h3bc924ef),
	.w6(32'h3ba1ca17),
	.w7(32'hbb8ee2de),
	.w8(32'hbc1669a0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93dea0),
	.w1(32'h3bafd6f8),
	.w2(32'hba959117),
	.w3(32'h3c28ec61),
	.w4(32'h3b680499),
	.w5(32'hbc161311),
	.w6(32'h3b1cc7d2),
	.w7(32'h3ac67481),
	.w8(32'h3c16208b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf966f2),
	.w1(32'h3b80f754),
	.w2(32'hbbc6aab8),
	.w3(32'h3c2ab381),
	.w4(32'h3bf3b648),
	.w5(32'hbbbd92e3),
	.w6(32'hbc80994d),
	.w7(32'hbc8bd4c6),
	.w8(32'hbc40f786),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21c574),
	.w1(32'h3c81da94),
	.w2(32'h3a1e0eb5),
	.w3(32'h3bc0827e),
	.w4(32'h3bb02f8d),
	.w5(32'h3b107014),
	.w6(32'h3c58c1c6),
	.w7(32'h3bd58a34),
	.w8(32'hbc30c452),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e1984),
	.w1(32'hbc33ab42),
	.w2(32'hbc7c2b70),
	.w3(32'h3bf82517),
	.w4(32'h3ba44887),
	.w5(32'hbc6184b0),
	.w6(32'h39d02540),
	.w7(32'h3a874ca0),
	.w8(32'h3bb9ecab),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0ee21),
	.w1(32'hbbdf99c8),
	.w2(32'hbb4483af),
	.w3(32'hbb7bfb5c),
	.w4(32'hbb5a62e8),
	.w5(32'hbbdaa6d1),
	.w6(32'h3bd5fbbb),
	.w7(32'h3ba4198c),
	.w8(32'h3c03ae50),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc52dc9),
	.w1(32'h3c544919),
	.w2(32'h3c1fae39),
	.w3(32'h3ba5c5b4),
	.w4(32'h3c409fde),
	.w5(32'h3bf9db0d),
	.w6(32'h3bae6658),
	.w7(32'h3bbd1d65),
	.w8(32'h3ab592ed),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b861337),
	.w1(32'h3a81963f),
	.w2(32'h3b4b6f8b),
	.w3(32'hb724fa99),
	.w4(32'hbaa1a012),
	.w5(32'h3bf20de4),
	.w6(32'h38bf22db),
	.w7(32'hbaf4a877),
	.w8(32'hbbd6c29f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8eb1b),
	.w1(32'h3c621fef),
	.w2(32'h3b181946),
	.w3(32'h3c7cc1db),
	.w4(32'h3c09cb3e),
	.w5(32'h3b06f0ba),
	.w6(32'h3b587fe1),
	.w7(32'hbb320b8b),
	.w8(32'hbbefa42f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4d529),
	.w1(32'hbbe19290),
	.w2(32'hbbbdf0ca),
	.w3(32'hba1ef94a),
	.w4(32'h3aefd1cf),
	.w5(32'hb936794a),
	.w6(32'h398e7599),
	.w7(32'h3b2036b4),
	.w8(32'h3a1d5eba),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6be70),
	.w1(32'hb707ec6d),
	.w2(32'h3b6435d7),
	.w3(32'h3b39cec0),
	.w4(32'h395f8b51),
	.w5(32'h3a5cc871),
	.w6(32'h3ac00134),
	.w7(32'h3bc806fa),
	.w8(32'h3b83f8f6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69be58),
	.w1(32'h3b2e812e),
	.w2(32'h3bd9038d),
	.w3(32'h3b81d7f0),
	.w4(32'hbae284ab),
	.w5(32'h3b6ec24c),
	.w6(32'h3b07ab7d),
	.w7(32'h3b9029c5),
	.w8(32'hbbae3a07),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1054a0),
	.w1(32'h3ba6a9ca),
	.w2(32'h3b65e745),
	.w3(32'hbbaf9811),
	.w4(32'h3b9f5f70),
	.w5(32'h3b3c8c8f),
	.w6(32'hba84325c),
	.w7(32'hb91d0def),
	.w8(32'h3a13d34c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2c84d),
	.w1(32'hbbe2d753),
	.w2(32'h3b05614d),
	.w3(32'h3b2560c7),
	.w4(32'hbc77248c),
	.w5(32'hb9db4211),
	.w6(32'hbbb0c269),
	.w7(32'h3af6c1c1),
	.w8(32'h3c04bd68),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed8345),
	.w1(32'hbc2c2e2d),
	.w2(32'hbc539ba8),
	.w3(32'h3b2af441),
	.w4(32'hbb03ef2d),
	.w5(32'hbbe6e0fa),
	.w6(32'h39d3b514),
	.w7(32'hbc48ad08),
	.w8(32'hbb1bad0b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9de7aa),
	.w1(32'hbc393e7a),
	.w2(32'hbc0509b2),
	.w3(32'hbb31b028),
	.w4(32'h3b88b0f6),
	.w5(32'h3b3450e2),
	.w6(32'hbc6c685a),
	.w7(32'hbc9ce621),
	.w8(32'hbcc3ccf8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83f7c2),
	.w1(32'h3b05d7f8),
	.w2(32'h3c096e7a),
	.w3(32'h39964ad1),
	.w4(32'h3b11567c),
	.w5(32'h3c254dfa),
	.w6(32'hbb70518b),
	.w7(32'h3b160fe2),
	.w8(32'h3982ecd6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae16930),
	.w1(32'h3ac66dbc),
	.w2(32'hbb1b07ac),
	.w3(32'h3c3880bf),
	.w4(32'h3c5a5c6a),
	.w5(32'h3c27cbda),
	.w6(32'h3b466ca5),
	.w7(32'hbbd7fb88),
	.w8(32'h3a95ed0b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b78dd),
	.w1(32'h3c36e875),
	.w2(32'h3a37e224),
	.w3(32'hbb8fff84),
	.w4(32'h3a3fe470),
	.w5(32'h3ae4ecf0),
	.w6(32'hbc03f8bc),
	.w7(32'hbc20cb34),
	.w8(32'hbc550284),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc171be2),
	.w1(32'h3b0defcc),
	.w2(32'hbb79321e),
	.w3(32'hbab3c730),
	.w4(32'hba65de15),
	.w5(32'hbba4ee82),
	.w6(32'h3ab48d45),
	.w7(32'hbb32ae70),
	.w8(32'hbb970864),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cb8c5),
	.w1(32'hbb97eb7a),
	.w2(32'hba5ca4e1),
	.w3(32'hbbb0cf45),
	.w4(32'hbba15084),
	.w5(32'hb9e6de30),
	.w6(32'h3b8a5d4f),
	.w7(32'hbb3d975d),
	.w8(32'h3bba7e81),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1fb28),
	.w1(32'hbade56d5),
	.w2(32'h3be02eef),
	.w3(32'h3ad12b9c),
	.w4(32'h3b23a36e),
	.w5(32'hb9390d45),
	.w6(32'h3ab0122d),
	.w7(32'h39d5bbb0),
	.w8(32'h3b03e6b2),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37df09),
	.w1(32'h3b4fa7d0),
	.w2(32'h3c1616bf),
	.w3(32'h3c19a358),
	.w4(32'h3c21c2a8),
	.w5(32'h3c4e357e),
	.w6(32'h3b7528b6),
	.w7(32'h3bfaa0a5),
	.w8(32'h3b239fcb),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c487921),
	.w1(32'h3b051601),
	.w2(32'hbb253b93),
	.w3(32'h3bfdab0e),
	.w4(32'h3b0b7f5c),
	.w5(32'h39016959),
	.w6(32'h3a2efe0a),
	.w7(32'hbaa1d9f1),
	.w8(32'h3ac0595d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba53c42),
	.w1(32'hbc0b1f8f),
	.w2(32'hbcecb8cb),
	.w3(32'h3b9afc7d),
	.w4(32'hbbd718a6),
	.w5(32'hbca0541a),
	.w6(32'hbb0cce3b),
	.w7(32'hbc955f3c),
	.w8(32'hbad97263),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule