module layer_8_featuremap_20(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51ad8b),
	.w1(32'hbc3a2b24),
	.w2(32'hbc96bf73),
	.w3(32'hbcd34509),
	.w4(32'hbc8c237f),
	.w5(32'h3b5bbc97),
	.w6(32'h3bf39071),
	.w7(32'hba63d290),
	.w8(32'h3c5f7c27),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c424b),
	.w1(32'hbc35d228),
	.w2(32'hbc221a30),
	.w3(32'h3c30a51d),
	.w4(32'h3b7d37ca),
	.w5(32'hbc6461a3),
	.w6(32'h3d929f1d),
	.w7(32'hbb82805a),
	.w8(32'h3c556cb8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd08b76b),
	.w1(32'hbbdca598),
	.w2(32'h3a18be22),
	.w3(32'hb9a7b66e),
	.w4(32'h3a17cd27),
	.w5(32'h3bcd320d),
	.w6(32'hbbd79418),
	.w7(32'h38d8160f),
	.w8(32'hb8496ad9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80e8a6),
	.w1(32'h3b1e7a4d),
	.w2(32'h3c04da69),
	.w3(32'h3b05da1a),
	.w4(32'hbc1970c9),
	.w5(32'h3c8322e3),
	.w6(32'hbc087cc6),
	.w7(32'hbc570315),
	.w8(32'h3c6a9fe0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25f13a),
	.w1(32'hbabd210a),
	.w2(32'hbc177307),
	.w3(32'hbbccbd25),
	.w4(32'hbc190ce7),
	.w5(32'h3a5cb787),
	.w6(32'hbc2f6ab2),
	.w7(32'hbba0336c),
	.w8(32'h3b90c1e1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf548eb),
	.w1(32'hba974025),
	.w2(32'h3c2a4e06),
	.w3(32'hbc27d70c),
	.w4(32'hbc212c21),
	.w5(32'hbc4adf7c),
	.w6(32'h3c41e598),
	.w7(32'h3bc289aa),
	.w8(32'h3c35b5ed),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30f140),
	.w1(32'h3c522ee8),
	.w2(32'h391689dd),
	.w3(32'hbc7ad06e),
	.w4(32'hba5de3ac),
	.w5(32'hbc1d1693),
	.w6(32'hbb496d77),
	.w7(32'hbbaef2f7),
	.w8(32'hbafd78a5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0178f),
	.w1(32'h3b3e946f),
	.w2(32'h3c6876a4),
	.w3(32'hbb4351b6),
	.w4(32'h3b95823b),
	.w5(32'hbc85c8e2),
	.w6(32'hbc11cc12),
	.w7(32'hbcaea0c7),
	.w8(32'hba9e94d8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32c2c9),
	.w1(32'hbb37409e),
	.w2(32'h3b534d7b),
	.w3(32'h3c89c475),
	.w4(32'hbca77f3e),
	.w5(32'h3a49b2e6),
	.w6(32'hba529472),
	.w7(32'h3b94ddc4),
	.w8(32'hbcb746cf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a33c0),
	.w1(32'hbc29d64a),
	.w2(32'hbbc46da3),
	.w3(32'h3c833668),
	.w4(32'hbc7fb329),
	.w5(32'hbab80ba5),
	.w6(32'hbb6d1db0),
	.w7(32'hbc29a560),
	.w8(32'h3b62de97),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81705d),
	.w1(32'h3b2a523d),
	.w2(32'hbc27505d),
	.w3(32'hbbdfada8),
	.w4(32'h39fa3da6),
	.w5(32'h3bdd78b1),
	.w6(32'h3acce77d),
	.w7(32'hbb69f75b),
	.w8(32'h3c74b906),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7ed4df),
	.w1(32'hbc97f861),
	.w2(32'h37388f19),
	.w3(32'hbb31bc8e),
	.w4(32'h3c62e889),
	.w5(32'hbad02348),
	.w6(32'h3a18a17f),
	.w7(32'hbcbbe052),
	.w8(32'hbcc8dc1e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb97c2),
	.w1(32'h3bc59aba),
	.w2(32'h3abf64e9),
	.w3(32'h3c1d8981),
	.w4(32'hbb544031),
	.w5(32'h3b9a0b1e),
	.w6(32'h3cbc6d8f),
	.w7(32'h3d5ee922),
	.w8(32'h3c0645ee),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc846d18),
	.w1(32'h3c362e52),
	.w2(32'hbba27331),
	.w3(32'h3c7b160f),
	.w4(32'h3af47678),
	.w5(32'hbcb4d8fb),
	.w6(32'h3c7524db),
	.w7(32'h3da0f350),
	.w8(32'h3ba74a72),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4874a6),
	.w1(32'h3b0c9a68),
	.w2(32'h3bd7a635),
	.w3(32'h3b030d4d),
	.w4(32'hbaad08cd),
	.w5(32'h3cf336fc),
	.w6(32'h3d2ac81e),
	.w7(32'h3c16a26a),
	.w8(32'hb9cdbf03),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4643c6),
	.w1(32'hbc342381),
	.w2(32'hbbb7b4d5),
	.w3(32'h3c0ce3dc),
	.w4(32'h3b265fa7),
	.w5(32'hbd8c3d2c),
	.w6(32'h3a303795),
	.w7(32'h3ae2dc32),
	.w8(32'h3c0dda04),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1e111b),
	.w1(32'h3baa6108),
	.w2(32'h3b3c28ad),
	.w3(32'hbcbf6fa4),
	.w4(32'h3cb6a3c2),
	.w5(32'h3d0273d9),
	.w6(32'hbc025045),
	.w7(32'h3b1ec2cf),
	.w8(32'h3b5beb7d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd19b2f),
	.w1(32'hbc6dc999),
	.w2(32'h39860da1),
	.w3(32'hbc068a8e),
	.w4(32'h3ba0cc47),
	.w5(32'hbc91c147),
	.w6(32'hbd74b35c),
	.w7(32'hba17c012),
	.w8(32'hba5d127e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb273e0b),
	.w1(32'h3884fe77),
	.w2(32'hbbb47d34),
	.w3(32'h39edf535),
	.w4(32'h3c29ed8c),
	.w5(32'hbba685a3),
	.w6(32'hbc450f93),
	.w7(32'h3b1c7b79),
	.w8(32'h3aed51c2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26c565),
	.w1(32'h3b3d1eaa),
	.w2(32'hbc56882f),
	.w3(32'hbc230f75),
	.w4(32'h3d657b1d),
	.w5(32'hbd0b3a43),
	.w6(32'hbaba3ffe),
	.w7(32'hbcb7b5c3),
	.w8(32'h3b2f54bd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b2666),
	.w1(32'hbc4ee1a8),
	.w2(32'hba80df41),
	.w3(32'hbc4822a9),
	.w4(32'h3d7fba9f),
	.w5(32'h3c9215ab),
	.w6(32'h3b04f576),
	.w7(32'hbb6eb191),
	.w8(32'h3be09924),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cc7a0),
	.w1(32'h3bff4d41),
	.w2(32'hbb8747a7),
	.w3(32'h3b4d048a),
	.w4(32'hbb20d623),
	.w5(32'h3a6cd51f),
	.w6(32'h3b57f889),
	.w7(32'hbc050ea1),
	.w8(32'hbb9ddedb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe54806),
	.w1(32'hbd88ab5e),
	.w2(32'hbb9388f0),
	.w3(32'h3b37ecaf),
	.w4(32'h3b70a65b),
	.w5(32'h3b4d6c91),
	.w6(32'h3b6b5545),
	.w7(32'h3b56087b),
	.w8(32'hbc7b0922),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98c87b),
	.w1(32'h3c253b4f),
	.w2(32'h3c00c2db),
	.w3(32'hbb8fd540),
	.w4(32'hbbcd152f),
	.w5(32'h3b121bbf),
	.w6(32'h3b510725),
	.w7(32'h3b297edd),
	.w8(32'h3c1e267d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba548cce),
	.w1(32'hbc25fb8d),
	.w2(32'hbbca3670),
	.w3(32'hbb3794cc),
	.w4(32'h3c2f38dd),
	.w5(32'hbc7912a8),
	.w6(32'h3af5739e),
	.w7(32'h3c2b29c6),
	.w8(32'hbaee2348),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae0f80),
	.w1(32'hbc394e25),
	.w2(32'h3bbd7109),
	.w3(32'h3c056853),
	.w4(32'hbc59b3de),
	.w5(32'h3b46650d),
	.w6(32'h3bdbe53f),
	.w7(32'h3c672187),
	.w8(32'h3b40dca0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82361b),
	.w1(32'h3ba245b6),
	.w2(32'h3bb65920),
	.w3(32'h3aaacde5),
	.w4(32'hbbfeb336),
	.w5(32'h3a7a01d3),
	.w6(32'hbc3fab44),
	.w7(32'hbb6c9874),
	.w8(32'hbb027236),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbda97b),
	.w1(32'h3bcea7d4),
	.w2(32'h3b44d42a),
	.w3(32'hbba0b7ce),
	.w4(32'hbc1433fc),
	.w5(32'h3ca690aa),
	.w6(32'hba0298a4),
	.w7(32'h3bbd12d9),
	.w8(32'hbab6a73f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8686e0),
	.w1(32'hbb36f64f),
	.w2(32'hbb2b950a),
	.w3(32'hba30f560),
	.w4(32'h3c4d694d),
	.w5(32'hbb503d29),
	.w6(32'hba114bfd),
	.w7(32'hba88061d),
	.w8(32'hb91619bf),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87e80f),
	.w1(32'hb8cb57c6),
	.w2(32'hbbd066d7),
	.w3(32'hbc3cee06),
	.w4(32'h3b3f58de),
	.w5(32'hba397e20),
	.w6(32'hbb092a35),
	.w7(32'h3b2ced98),
	.w8(32'hbadf5fb2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3d30e),
	.w1(32'h3b853ef3),
	.w2(32'h3b4eb99b),
	.w3(32'h3bed9b69),
	.w4(32'h3ba2edfe),
	.w5(32'hbbbd56ab),
	.w6(32'hbb14f845),
	.w7(32'hbbdc096a),
	.w8(32'h3a152f62),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13e604),
	.w1(32'hbadcfbe0),
	.w2(32'hbb100288),
	.w3(32'hba4444cb),
	.w4(32'hbb495b83),
	.w5(32'hbacaca7f),
	.w6(32'hbb2c59cb),
	.w7(32'h3ae4ae6d),
	.w8(32'h3b498b6f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6614c1),
	.w1(32'hbc2bd348),
	.w2(32'h3b03c413),
	.w3(32'h3aa71eb1),
	.w4(32'h3a92de5f),
	.w5(32'h3aa7554e),
	.w6(32'hbb6a2dbf),
	.w7(32'h3ada8e93),
	.w8(32'h3bdb54ce),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae923d),
	.w1(32'h3b4b5049),
	.w2(32'h3bac4156),
	.w3(32'h3bc04102),
	.w4(32'h3acc2ddc),
	.w5(32'hbbf76be5),
	.w6(32'h3b42e3a4),
	.w7(32'h3c8ad215),
	.w8(32'h3b8c3928),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59e4f7),
	.w1(32'hbbf5064e),
	.w2(32'h3c3d9df4),
	.w3(32'h3ab0d90c),
	.w4(32'hbbde6dac),
	.w5(32'hbb92aa1a),
	.w6(32'h3918fa60),
	.w7(32'h3bd4679b),
	.w8(32'hbb293328),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d1c73),
	.w1(32'h3a719781),
	.w2(32'hbbd6b24f),
	.w3(32'h3b3965ac),
	.w4(32'h3c318ec6),
	.w5(32'hbba5cbf1),
	.w6(32'h3c5e05e4),
	.w7(32'h3c87c347),
	.w8(32'hbbc44e9d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30f74a),
	.w1(32'hbadd284c),
	.w2(32'h377e745e),
	.w3(32'h3c057a9d),
	.w4(32'h3962a622),
	.w5(32'hbbb5f6f8),
	.w6(32'hbb892b05),
	.w7(32'hbb7c5006),
	.w8(32'hbbc54767),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb938776),
	.w1(32'h3b954f4f),
	.w2(32'h3c3add47),
	.w3(32'hbb0004de),
	.w4(32'h39a91372),
	.w5(32'h3bef9556),
	.w6(32'h3aac65dc),
	.w7(32'h3b8e0556),
	.w8(32'hbaf377b7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d0ae8),
	.w1(32'h3bcd6a0e),
	.w2(32'h3c862afe),
	.w3(32'hbbc12658),
	.w4(32'hbacf3c99),
	.w5(32'h3c4f757b),
	.w6(32'hbb30ece4),
	.w7(32'h3be2019b),
	.w8(32'hbb9ffac7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbb373),
	.w1(32'h3b86b8d5),
	.w2(32'hbba4f21a),
	.w3(32'hbaf187d8),
	.w4(32'hbac46348),
	.w5(32'h3b3e4c1e),
	.w6(32'h3a840419),
	.w7(32'h3aca8d16),
	.w8(32'hbbd737b9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33c2ac),
	.w1(32'h3ad7e9d4),
	.w2(32'hbb072b46),
	.w3(32'h3a154770),
	.w4(32'h3b767386),
	.w5(32'hb7dd073f),
	.w6(32'hbb758402),
	.w7(32'hbb21066c),
	.w8(32'h3af7ac52),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6b0a8),
	.w1(32'h3c228bbb),
	.w2(32'hbb8ad217),
	.w3(32'hbbfc22de),
	.w4(32'hbbd857ea),
	.w5(32'h38845853),
	.w6(32'h3b990927),
	.w7(32'hbc3b251d),
	.w8(32'hbb4b307a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce8924d),
	.w1(32'h3be1bbd2),
	.w2(32'h3bf1fef2),
	.w3(32'h3c3f2ad7),
	.w4(32'hbb6a9c4b),
	.w5(32'hbc705791),
	.w6(32'h3c8fc38c),
	.w7(32'h3bebe00d),
	.w8(32'hbb0b91cc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce4fae),
	.w1(32'h3c287a8f),
	.w2(32'hbbd376b4),
	.w3(32'hbbb69fd5),
	.w4(32'h3c175161),
	.w5(32'h3c346da7),
	.w6(32'hba236ca3),
	.w7(32'h3a5b4dc5),
	.w8(32'hbb811975),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e5729),
	.w1(32'hbbd6ea20),
	.w2(32'h3c8c111c),
	.w3(32'h3ac6c9a2),
	.w4(32'h3ca3d63f),
	.w5(32'hbc12d014),
	.w6(32'h3c87b9cf),
	.w7(32'h3c219281),
	.w8(32'hbb6168db),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1458a6),
	.w1(32'h3b0f1a2f),
	.w2(32'h3bc75e9a),
	.w3(32'hb97791ae),
	.w4(32'hbbd25753),
	.w5(32'h3c8c6a50),
	.w6(32'hbc628647),
	.w7(32'h3bb92680),
	.w8(32'hba4c5414),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf97841),
	.w1(32'h3a0cba29),
	.w2(32'h3cab1de9),
	.w3(32'hba94e883),
	.w4(32'h3c02fd3e),
	.w5(32'h3c8e50a5),
	.w6(32'h3cae84a8),
	.w7(32'h3b1baaa2),
	.w8(32'hba2a255d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb016fd4),
	.w1(32'h3c6271f8),
	.w2(32'h3c06bcbc),
	.w3(32'hbc29dec6),
	.w4(32'hb9ca11cf),
	.w5(32'hbbcbdbe8),
	.w6(32'h39f8a3ff),
	.w7(32'h3c952905),
	.w8(32'hbc92afc1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d50f3),
	.w1(32'hbc4b8e3f),
	.w2(32'h3bf20479),
	.w3(32'h3c2efad2),
	.w4(32'hbc02d6f8),
	.w5(32'h3ca236ae),
	.w6(32'h3ce26b33),
	.w7(32'hbb5af911),
	.w8(32'hbc9aacf6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89d622),
	.w1(32'hbab1b7c4),
	.w2(32'h3c1fa685),
	.w3(32'h38d14cc7),
	.w4(32'h3b644668),
	.w5(32'h3bf62dd3),
	.w6(32'hbb1d3bbf),
	.w7(32'h3bdc20af),
	.w8(32'hbb34d03c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43c982),
	.w1(32'hb9f63f93),
	.w2(32'hb9dd7db3),
	.w3(32'h3bbe4329),
	.w4(32'h3be61e90),
	.w5(32'h3c6504ea),
	.w6(32'hba79fc61),
	.w7(32'hbc39d551),
	.w8(32'hb9db3578),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97f7e9),
	.w1(32'hbc07c978),
	.w2(32'hb9305fd2),
	.w3(32'h3c62e8c2),
	.w4(32'h3b88f4cb),
	.w5(32'h3cc4ac10),
	.w6(32'hbc372e59),
	.w7(32'h3c89d152),
	.w8(32'h3add7445),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b054c30),
	.w1(32'hbc584f06),
	.w2(32'hbb75d90e),
	.w3(32'h3ce40187),
	.w4(32'hbb83961f),
	.w5(32'h3c08c630),
	.w6(32'hbb8e9f5f),
	.w7(32'hbab46924),
	.w8(32'h3c059273),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2b5d4),
	.w1(32'hbb0ed65c),
	.w2(32'hbbe26e4f),
	.w3(32'hbbc20870),
	.w4(32'h3bfe92c0),
	.w5(32'h3c3b7eae),
	.w6(32'hbbbeb99e),
	.w7(32'hbb8bb24c),
	.w8(32'h3c331d1c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b367bd3),
	.w1(32'hba690f2e),
	.w2(32'h3c5e9f81),
	.w3(32'hbbbf03f5),
	.w4(32'hbaa72cd5),
	.w5(32'hbb80e042),
	.w6(32'hbba1bcbb),
	.w7(32'h3c941b6a),
	.w8(32'h3a1adc87),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65bb2b),
	.w1(32'hba9587e9),
	.w2(32'hbbc9ea14),
	.w3(32'hb9b270ed),
	.w4(32'h3b88ee78),
	.w5(32'h3b10a912),
	.w6(32'h3b9ba2c3),
	.w7(32'hb7901655),
	.w8(32'h3b386b46),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b333174),
	.w1(32'hbb4e9ce6),
	.w2(32'h3c036c3b),
	.w3(32'hbad3fd82),
	.w4(32'h3a8b6b04),
	.w5(32'hba14026b),
	.w6(32'h3c612d35),
	.w7(32'h3aaac5c8),
	.w8(32'h3baff175),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39948cd9),
	.w1(32'h3add4158),
	.w2(32'hbb650d08),
	.w3(32'hbad7d702),
	.w4(32'h3b97a11b),
	.w5(32'hbb686c7d),
	.w6(32'h392a4ea6),
	.w7(32'h3b9a59c6),
	.w8(32'hba8850dd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb818587b),
	.w1(32'hbae6f838),
	.w2(32'hbb668856),
	.w3(32'h3af31d67),
	.w4(32'hbc07386e),
	.w5(32'hbabc88a7),
	.w6(32'hba60d203),
	.w7(32'h3aec42c9),
	.w8(32'hbaa0fb6c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bbf50),
	.w1(32'h3a576fa4),
	.w2(32'hb9dc9883),
	.w3(32'h39bea9ad),
	.w4(32'hbb1b0240),
	.w5(32'hbb624f6e),
	.w6(32'h3acff0c0),
	.w7(32'h3ab15475),
	.w8(32'hbbc66875),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab36e20),
	.w1(32'h3afba6f8),
	.w2(32'hbb853f9a),
	.w3(32'hbaa9d365),
	.w4(32'h3c147fd4),
	.w5(32'h3a99c1aa),
	.w6(32'h3bfb8fd1),
	.w7(32'hbac4a5ba),
	.w8(32'hbb1153ee),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa648e),
	.w1(32'hbb455391),
	.w2(32'h3adc558f),
	.w3(32'hbb24c648),
	.w4(32'hbaa1cd6d),
	.w5(32'h3b6ba44c),
	.w6(32'hbae68915),
	.w7(32'hba0976ab),
	.w8(32'hba6e44a9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa60c9),
	.w1(32'h3a3f70c5),
	.w2(32'hb8a6ce67),
	.w3(32'h3c05a63e),
	.w4(32'hbb486e47),
	.w5(32'h3b785299),
	.w6(32'hbbdac4b4),
	.w7(32'h3a9d51df),
	.w8(32'hb9b99529),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87bd744),
	.w1(32'hb9fe978b),
	.w2(32'hbc3d522e),
	.w3(32'h3c0d3644),
	.w4(32'h3a4d1b19),
	.w5(32'h3995cf8d),
	.w6(32'hbb723f30),
	.w7(32'h3b093a93),
	.w8(32'h3b81722b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b854fe9),
	.w1(32'hbbab0258),
	.w2(32'h3ac76b9c),
	.w3(32'h3b240931),
	.w4(32'hbaac3115),
	.w5(32'hba16833c),
	.w6(32'hbbd8752c),
	.w7(32'hb87b6ace),
	.w8(32'h3a173481),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0a702),
	.w1(32'hbb7f6941),
	.w2(32'h3ad2fe50),
	.w3(32'h3a16417f),
	.w4(32'h3a80d689),
	.w5(32'h39102bed),
	.w6(32'hbb0cd1d3),
	.w7(32'hbb384ed6),
	.w8(32'h3a08fa7b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab91b34),
	.w1(32'hba160b63),
	.w2(32'h3a17aeb6),
	.w3(32'hbb220a90),
	.w4(32'hbad31ab9),
	.w5(32'h37da305c),
	.w6(32'hba8896d8),
	.w7(32'hbba12970),
	.w8(32'h3aa4d193),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94aa18),
	.w1(32'hbb5fcc8f),
	.w2(32'h3a604dbe),
	.w3(32'h3bb0bc98),
	.w4(32'h3a1eb76c),
	.w5(32'hbcb9e18f),
	.w6(32'h3b834297),
	.w7(32'hbb257b31),
	.w8(32'h3af59aef),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cb409),
	.w1(32'hbc667aa9),
	.w2(32'hbae1b151),
	.w3(32'h3b0766fb),
	.w4(32'h3aaaa0be),
	.w5(32'h3ba8c413),
	.w6(32'hbb556dba),
	.w7(32'h3a082631),
	.w8(32'h3a7d8585),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a784d),
	.w1(32'hbb3d3f6f),
	.w2(32'h3be5b4ff),
	.w3(32'hb9d1aa7e),
	.w4(32'h3d8379ad),
	.w5(32'hbc79118c),
	.w6(32'hbaae8784),
	.w7(32'hb9b7bcdb),
	.w8(32'hbc0c30f9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad8f5f),
	.w1(32'hbb02aa1d),
	.w2(32'hbcdf6250),
	.w3(32'hbba9ba18),
	.w4(32'h3d9305a0),
	.w5(32'h3c49bf5a),
	.w6(32'h3c7d2112),
	.w7(32'h3c2646dc),
	.w8(32'hbc9ff673),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc860fed),
	.w1(32'hb90db340),
	.w2(32'h3c9174c4),
	.w3(32'h3d51d8aa),
	.w4(32'hbc19272c),
	.w5(32'h3c564e0d),
	.w6(32'h3b35e375),
	.w7(32'hbd074b2d),
	.w8(32'hbba463ce),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a3fbd),
	.w1(32'h3b75f3cb),
	.w2(32'hbd784940),
	.w3(32'hbbb33a62),
	.w4(32'hbb3fa83e),
	.w5(32'h3c627906),
	.w6(32'hbb061e32),
	.w7(32'hb8e7daff),
	.w8(32'hbce81181),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7e0990),
	.w1(32'h3cd702d1),
	.w2(32'h3d464d04),
	.w3(32'h3c9cdf31),
	.w4(32'h3b2e5244),
	.w5(32'hbc524006),
	.w6(32'h3c36d686),
	.w7(32'h3b47aa16),
	.w8(32'h3bd4355a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e7711),
	.w1(32'hbc559cd1),
	.w2(32'hbc7f2618),
	.w3(32'hbd673460),
	.w4(32'h3bba18ff),
	.w5(32'hbc222e27),
	.w6(32'hb97667f0),
	.w7(32'hbbbc9d5c),
	.w8(32'hbbad6892),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfd267),
	.w1(32'h3c8a25fd),
	.w2(32'h39ae3fb7),
	.w3(32'hbaecf032),
	.w4(32'h3b29c738),
	.w5(32'hbb3f2127),
	.w6(32'hbbb0c832),
	.w7(32'hbb0d58b9),
	.w8(32'h3b176b71),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0359c1),
	.w1(32'h3d702cfb),
	.w2(32'hbd0dc861),
	.w3(32'hbbc2c617),
	.w4(32'hbc8828cb),
	.w5(32'h3c0fced9),
	.w6(32'hbb42fb6b),
	.w7(32'h3c5a8f2c),
	.w8(32'hbb8cb35d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06d3b0),
	.w1(32'h3d92b25c),
	.w2(32'h3c9ed781),
	.w3(32'hbbc22796),
	.w4(32'h3bab1929),
	.w5(32'h3be4691c),
	.w6(32'h3c16cbbb),
	.w7(32'hbc35bb92),
	.w8(32'h3af96950),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2168b9),
	.w1(32'h3a662ec8),
	.w2(32'h3984a946),
	.w3(32'h3beb39de),
	.w4(32'h3bd37817),
	.w5(32'hbbb1c295),
	.w6(32'h3c5a2bf7),
	.w7(32'h3aff0cc3),
	.w8(32'h3b46557d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3156bb),
	.w1(32'h3b80a9ac),
	.w2(32'h3c00a90c),
	.w3(32'h3b774399),
	.w4(32'hbc565a03),
	.w5(32'hbc8e7267),
	.w6(32'hbd846ece),
	.w7(32'h3ab272be),
	.w8(32'hbcaa0e55),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a69fb),
	.w1(32'hbbe9f92e),
	.w2(32'h3c0c08a3),
	.w3(32'h3b704ea9),
	.w4(32'hbc1dd483),
	.w5(32'h3c828bc8),
	.w6(32'hbafca59a),
	.w7(32'hbd14c8de),
	.w8(32'h3ba20a4b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bea1e),
	.w1(32'h3c7ed84d),
	.w2(32'hbc5e6a3b),
	.w3(32'h3b9c4089),
	.w4(32'h3c4e60c3),
	.w5(32'hbb971d43),
	.w6(32'hbbaf27cd),
	.w7(32'h3cabc987),
	.w8(32'hbcd89908),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd31199),
	.w1(32'hbc86e8d1),
	.w2(32'h3a184ec4),
	.w3(32'h3a1d3085),
	.w4(32'h3bbfd3f9),
	.w5(32'h3b4ecc5f),
	.w6(32'hbac37d44),
	.w7(32'h3c9c5149),
	.w8(32'h3b4d8e7e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2671d),
	.w1(32'hbb9affab),
	.w2(32'hbc916fe9),
	.w3(32'hbbcc0760),
	.w4(32'hb9ceb029),
	.w5(32'hbba8cf2f),
	.w6(32'h3cbcd7cd),
	.w7(32'hb962b66b),
	.w8(32'h3c23c6fe),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb880eca),
	.w1(32'hbba6d8f7),
	.w2(32'hbcdb7ce4),
	.w3(32'h3b3e04e7),
	.w4(32'hbb2e84fb),
	.w5(32'h3bea79d7),
	.w6(32'hbb72be7b),
	.w7(32'hbbbfcb89),
	.w8(32'h3c0bcc90),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22e5d9),
	.w1(32'hbb9059d4),
	.w2(32'hba0e5bb0),
	.w3(32'h3a8ed1a9),
	.w4(32'hbadc65f9),
	.w5(32'hbbb5d959),
	.w6(32'h3b77c11d),
	.w7(32'h3b214c91),
	.w8(32'hbbf30c37),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ba8d8),
	.w1(32'h3bb9a972),
	.w2(32'h3b0ccec2),
	.w3(32'h3b50b512),
	.w4(32'h3c965020),
	.w5(32'h3bd261a4),
	.w6(32'hbbf6bdc8),
	.w7(32'h3c0dae0e),
	.w8(32'h3ceadeb7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ca1fe),
	.w1(32'h3b9fdc49),
	.w2(32'hbb58781f),
	.w3(32'h3c89b688),
	.w4(32'h3b3c2ff6),
	.w5(32'hba099239),
	.w6(32'h3c1f19ab),
	.w7(32'hbb0beb65),
	.w8(32'hbc8e84c5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2acae3),
	.w1(32'h3c98810d),
	.w2(32'hbc2f7db5),
	.w3(32'hbad6bc91),
	.w4(32'h3c9354d7),
	.w5(32'hbc08fcf0),
	.w6(32'h3c680f68),
	.w7(32'h3a4c6e1b),
	.w8(32'h3c6bce4f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa4e3d),
	.w1(32'h3cc25778),
	.w2(32'hba523ec6),
	.w3(32'h39b6b795),
	.w4(32'h3bcb0106),
	.w5(32'hbbb4c7fd),
	.w6(32'hbbd33be6),
	.w7(32'hbb335c13),
	.w8(32'hb84d3e65),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8978f),
	.w1(32'h3aeeabc1),
	.w2(32'h3b46ca45),
	.w3(32'hba3b9d67),
	.w4(32'h3ba67659),
	.w5(32'h3cc86094),
	.w6(32'h3c93a466),
	.w7(32'hbc82d8e2),
	.w8(32'h3ccb6b1f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97fc5c),
	.w1(32'h3bca7e46),
	.w2(32'h3b8fd0ca),
	.w3(32'hbadd767d),
	.w4(32'h3c26f0dc),
	.w5(32'h3b62c711),
	.w6(32'hba33fa3d),
	.w7(32'hbc6f5afc),
	.w8(32'hbb85f576),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8832ce),
	.w1(32'h3be9cb57),
	.w2(32'h3b62a135),
	.w3(32'h3bf9d603),
	.w4(32'h3c090df5),
	.w5(32'h3b1d1d8f),
	.w6(32'h3bf4186b),
	.w7(32'hb98baca7),
	.w8(32'h3bedae0f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69d1d1),
	.w1(32'hba755836),
	.w2(32'h391575d6),
	.w3(32'h3ae31af4),
	.w4(32'h3cd024e6),
	.w5(32'h3b837e29),
	.w6(32'hbb0e5c01),
	.w7(32'hbaa9cd80),
	.w8(32'h3b4ac41f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0af875),
	.w1(32'hba619eb3),
	.w2(32'h3beb566b),
	.w3(32'h3c11b31e),
	.w4(32'h3ade4eac),
	.w5(32'hbc0a6627),
	.w6(32'h3c359ba1),
	.w7(32'hbb43ba62),
	.w8(32'hbb6b1f8f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb370137),
	.w1(32'h3abd681b),
	.w2(32'h3bc5ce00),
	.w3(32'h3b9210c8),
	.w4(32'hbb081258),
	.w5(32'h3c15746a),
	.w6(32'h3ac4cb1d),
	.w7(32'h3bf48b2d),
	.w8(32'h39d2f366),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ebb5f),
	.w1(32'h3a81548c),
	.w2(32'h3b8a9efd),
	.w3(32'h3c86c5a6),
	.w4(32'h3c8cd65b),
	.w5(32'h3c2f765d),
	.w6(32'h3c7caa23),
	.w7(32'h3c09501e),
	.w8(32'hbbab0272),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bd07f),
	.w1(32'h3cd61520),
	.w2(32'h3a0231ce),
	.w3(32'h3b09850b),
	.w4(32'h3bd453e4),
	.w5(32'h3b1f246d),
	.w6(32'hb9ed22cb),
	.w7(32'h3a33172e),
	.w8(32'hbc9963b7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac01a9),
	.w1(32'h3b83cf79),
	.w2(32'hbb6ce060),
	.w3(32'hbae6eefe),
	.w4(32'hbb9705c7),
	.w5(32'hba968493),
	.w6(32'hbae1a001),
	.w7(32'hba3be5e4),
	.w8(32'hbccc2853),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eb39aa),
	.w1(32'hbab709ca),
	.w2(32'h3b69cc7e),
	.w3(32'h3bddbcb1),
	.w4(32'hbbb10ecc),
	.w5(32'h3b05f42b),
	.w6(32'hba506503),
	.w7(32'hbca57bc3),
	.w8(32'hbaf1ed1c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e502a2),
	.w1(32'hbad88510),
	.w2(32'h3b644814),
	.w3(32'hbc0cc687),
	.w4(32'hba102a9e),
	.w5(32'hba602f56),
	.w6(32'h3b40353e),
	.w7(32'h3a9b0fc6),
	.w8(32'h3b33b38a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b315e59),
	.w1(32'h3c47063a),
	.w2(32'h3b392048),
	.w3(32'h3cd4861a),
	.w4(32'h3c4f5730),
	.w5(32'hbb8b4342),
	.w6(32'hbb05ee98),
	.w7(32'h3b8ec2f6),
	.w8(32'hba1e5a93),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba836160),
	.w1(32'h3b19196a),
	.w2(32'h3b994ba4),
	.w3(32'hbc6858ec),
	.w4(32'h3b879317),
	.w5(32'hbb37a82b),
	.w6(32'hbae67df0),
	.w7(32'h3ca7faf7),
	.w8(32'h3b1a8798),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c99e2),
	.w1(32'hbb02ba26),
	.w2(32'hbb134f30),
	.w3(32'hbb3469aa),
	.w4(32'h39c0f90d),
	.w5(32'hbb9a6d6a),
	.w6(32'hbac8de40),
	.w7(32'h3bb834ef),
	.w8(32'h3aa67a9c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8629ff),
	.w1(32'hba35c8a1),
	.w2(32'h3b3ef06e),
	.w3(32'hba72953f),
	.w4(32'h3b479f2f),
	.w5(32'hbc97898c),
	.w6(32'hbaa06ef7),
	.w7(32'hbaceba1a),
	.w8(32'h3cb6f3be),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b587281),
	.w1(32'h3b957aac),
	.w2(32'h3ab527b1),
	.w3(32'h3be3d359),
	.w4(32'h3ab5c8ad),
	.w5(32'hbcb77624),
	.w6(32'h3b0938ca),
	.w7(32'hbabd5d07),
	.w8(32'hbab6f4c0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcfc8a),
	.w1(32'h3bef5a22),
	.w2(32'hbb75c2fc),
	.w3(32'hbb8724a6),
	.w4(32'hbb093277),
	.w5(32'hba57a5e5),
	.w6(32'hbb15de3d),
	.w7(32'hbb2adec5),
	.w8(32'h3a12a149),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b363d),
	.w1(32'hba02bac0),
	.w2(32'h3cc77a73),
	.w3(32'h3a929a96),
	.w4(32'hb9cd9d21),
	.w5(32'hbabafca1),
	.w6(32'h3b5e11e4),
	.w7(32'hbaac1c06),
	.w8(32'hbb437bb8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ac914),
	.w1(32'h3ba85ec4),
	.w2(32'hba9c9168),
	.w3(32'h3b0b4abb),
	.w4(32'hba1d0f85),
	.w5(32'hbac22a70),
	.w6(32'h3bead709),
	.w7(32'hba9ed063),
	.w8(32'hbab6b6bf),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdbc0f),
	.w1(32'hbabe52db),
	.w2(32'h3b02cb9e),
	.w3(32'hbb11f2b4),
	.w4(32'h3a60ab3e),
	.w5(32'hbb9da257),
	.w6(32'h3b913326),
	.w7(32'h3b11660f),
	.w8(32'hbb82504f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba69233),
	.w1(32'h3b85bd8d),
	.w2(32'h3b285445),
	.w3(32'h3bc275e2),
	.w4(32'h3be2f407),
	.w5(32'h3aef83d4),
	.w6(32'hbb3f127b),
	.w7(32'hba84ee93),
	.w8(32'h3b38fddd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74fc1e),
	.w1(32'hbad5789a),
	.w2(32'h3bb19268),
	.w3(32'h3a9e78a7),
	.w4(32'hbb602122),
	.w5(32'h3a867105),
	.w6(32'hba7bac48),
	.w7(32'h3b8258ed),
	.w8(32'hbb2177d3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbed34d20),
	.w1(32'hbf5d874a),
	.w2(32'hbf738070),
	.w3(32'h3f5638d6),
	.w4(32'hbf529526),
	.w5(32'hbf2c66d1),
	.w6(32'hbf454214),
	.w7(32'hbf737740),
	.w8(32'hbf5013e9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf2b7a53),
	.w1(32'h3f7f90bc),
	.w2(32'hbf34e67c),
	.w3(32'h3f991894),
	.w4(32'hbf02924c),
	.w5(32'hbfebe823),
	.w6(32'hbf0feb3b),
	.w7(32'hbf1382b2),
	.w8(32'hbf0ac835),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf179824),
	.w1(32'hbf2f6b85),
	.w2(32'hbf351b08),
	.w3(32'hbf3ee617),
	.w4(32'hbf1936a5),
	.w5(32'hbeefd547),
	.w6(32'hbed1e5a2),
	.w7(32'hbec9f6a5),
	.w8(32'hbe06e030),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf21a77f),
	.w1(32'h3f86a0fd),
	.w2(32'h3fca9961),
	.w3(32'hbf0231c2),
	.w4(32'hbf86834d),
	.w5(32'hbf3eabea),
	.w6(32'hbf1c7798),
	.w7(32'h3e9e063c),
	.w8(32'hbf2ceb58),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf35b1c2),
	.w1(32'h3f469a6b),
	.w2(32'hbf065205),
	.w3(32'hbf0f4197),
	.w4(32'hbf2183be),
	.w5(32'h3f402aa8),
	.w6(32'h3e0da163),
	.w7(32'hbef2cce1),
	.w8(32'hbe200eb2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbebf2b97),
	.w1(32'h3f00117c),
	.w2(32'hbed4e846),
	.w3(32'hbf34f44d),
	.w4(32'hbf1bc337),
	.w5(32'hbf27fc45),
	.w6(32'hbf19c8e9),
	.w7(32'hbf142ca8),
	.w8(32'hbdc5c85e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf4d7b38),
	.w1(32'hbec1cd3c),
	.w2(32'hbf31b718),
	.w3(32'hbf2b5546),
	.w4(32'hbf23011f),
	.w5(32'hbf0a6233),
	.w6(32'hbf251489),
	.w7(32'h3ea437ea),
	.w8(32'hbef5b8d2),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f2898e8),
	.w1(32'h3dc97259),
	.w2(32'hbee8169f),
	.w3(32'h3f989c7e),
	.w4(32'hbe986eb8),
	.w5(32'hbee93307),
	.w6(32'hbea907f3),
	.w7(32'hbf24a0e0),
	.w8(32'hbf541df6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f244616),
	.w1(32'hbe89f1cf),
	.w2(32'hbe097f75),
	.w3(32'hbf13af9a),
	.w4(32'h3e1062e8),
	.w5(32'h3da214c7),
	.w6(32'hbefabbc3),
	.w7(32'hbf00764c),
	.w8(32'hbd8f630f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf21f1a5),
	.w1(32'hbf27e261),
	.w2(32'hbf2cf0f2),
	.w3(32'hbf1555d2),
	.w4(32'hbf0066c2),
	.w5(32'h3e23224a),
	.w6(32'hbf16e3ce),
	.w7(32'hbea51dcc),
	.w8(32'h3f8ac6af),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e84d34b),
	.w1(32'hbefd02b2),
	.w2(32'hbec43d30),
	.w3(32'hbf19f805),
	.w4(32'hbf30f712),
	.w5(32'h3e2d3a9f),
	.w6(32'hbefdd6a0),
	.w7(32'hbf89e5e9),
	.w8(32'hbf067622),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf1d08b2),
	.w1(32'hbf1f9095),
	.w2(32'hbf1e9bc1),
	.w3(32'hbf23e64c),
	.w4(32'hbf480d09),
	.w5(32'hbf08ef2e),
	.w6(32'hbf3c5edc),
	.w7(32'hbf0db20d),
	.w8(32'hbf04dd21),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38cbd3),
	.w1(32'hbf1a6c40),
	.w2(32'hbefd05ff),
	.w3(32'hbb1f431b),
	.w4(32'hbf0f52f6),
	.w5(32'hbf56ca76),
	.w6(32'hbed9c80f),
	.w7(32'hbd1cd132),
	.w8(32'h3e853fee),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf38173c),
	.w1(32'hbf0bd1ca),
	.w2(32'h3f4fac65),
	.w3(32'hbebdc6a0),
	.w4(32'hbe267b56),
	.w5(32'h3da84027),
	.w6(32'hbf0e4566),
	.w7(32'hbf209644),
	.w8(32'hbee66c4d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf102dbc),
	.w1(32'h3fbb7279),
	.w2(32'h3eb1d919),
	.w3(32'hbf1ae13c),
	.w4(32'h3e5c2c26),
	.w5(32'h3e4c871f),
	.w6(32'hb75fee0a),
	.w7(32'h3eb67605),
	.w8(32'h3e99363b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e6a5ab4),
	.w1(32'h3f36de02),
	.w2(32'h3e905a03),
	.w3(32'hbeb88b37),
	.w4(32'h3f65588b),
	.w5(32'h3f634ce3),
	.w6(32'h3e53cfc0),
	.w7(32'h3f6e089a),
	.w8(32'h371d0351),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule