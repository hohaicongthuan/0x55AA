module layer_10_featuremap_89(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e3654),
	.w1(32'hbb105e50),
	.w2(32'h3aa22127),
	.w3(32'hbab3be72),
	.w4(32'hbb6762ef),
	.w5(32'hbb192d9d),
	.w6(32'h3c5fc63f),
	.w7(32'h37c5a155),
	.w8(32'h3b0f7336),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc5997),
	.w1(32'h3b28356f),
	.w2(32'hba1203e5),
	.w3(32'hbaf0f394),
	.w4(32'hb9db1f03),
	.w5(32'h3a44f412),
	.w6(32'h39f340fb),
	.w7(32'hbb539300),
	.w8(32'hb81dca74),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7aa7d),
	.w1(32'h3b209413),
	.w2(32'h3b4c8a25),
	.w3(32'hba8e1b3c),
	.w4(32'h3c06bd95),
	.w5(32'hbbc9eba9),
	.w6(32'h3aed6128),
	.w7(32'h396fc82f),
	.w8(32'hbb4aa6d3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b586934),
	.w1(32'hbb57c542),
	.w2(32'hb9d5e1d2),
	.w3(32'h3b21cd59),
	.w4(32'h39dce3a3),
	.w5(32'hbb1f22d7),
	.w6(32'h3a8ea965),
	.w7(32'h3adb07ed),
	.w8(32'h38c6aac0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adaa560),
	.w1(32'h3a3e9439),
	.w2(32'h3b5e7584),
	.w3(32'hbb836398),
	.w4(32'h3b14d9ef),
	.w5(32'h38a16839),
	.w6(32'hbb033349),
	.w7(32'h3b292352),
	.w8(32'h39817e61),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadda726),
	.w1(32'h3a673303),
	.w2(32'hbab7b41a),
	.w3(32'hbb471ce2),
	.w4(32'h39522dde),
	.w5(32'hbafff0cb),
	.w6(32'h3bfa0f98),
	.w7(32'h3a956592),
	.w8(32'hbb4eec47),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb364e27),
	.w1(32'h3969c00b),
	.w2(32'hbaa01fde),
	.w3(32'hbbfb1eab),
	.w4(32'h3aac861d),
	.w5(32'hb94fa4be),
	.w6(32'hbb77e9bf),
	.w7(32'h3b69bda5),
	.w8(32'h3b861574),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1eef2f),
	.w1(32'h3c346bb5),
	.w2(32'h3baef10f),
	.w3(32'h3be96baf),
	.w4(32'h3bf92507),
	.w5(32'h3b8e2e62),
	.w6(32'h3c258040),
	.w7(32'hbaec62e1),
	.w8(32'h3b32fb45),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc40c5d),
	.w1(32'hbb5909fa),
	.w2(32'h3b870ff2),
	.w3(32'h3afbf142),
	.w4(32'h3b35619e),
	.w5(32'h3ac96919),
	.w6(32'hbad43baa),
	.w7(32'hba5a99cb),
	.w8(32'hb9ab7810),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37e688),
	.w1(32'h3badd9b1),
	.w2(32'h3c15e8f2),
	.w3(32'h39bc7ee1),
	.w4(32'hba19db8d),
	.w5(32'h3ae23952),
	.w6(32'hba8b7270),
	.w7(32'h3acf9560),
	.w8(32'hbb279174),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4630b6),
	.w1(32'hbabe40ed),
	.w2(32'h3925755c),
	.w3(32'h3c08788a),
	.w4(32'hbb64fd05),
	.w5(32'h3c4d6ad3),
	.w6(32'hbae4f910),
	.w7(32'hbb117fd5),
	.w8(32'h3a78a182),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c069bd3),
	.w1(32'hbb05877f),
	.w2(32'h3baba656),
	.w3(32'hbbb118fa),
	.w4(32'h3c0843e0),
	.w5(32'hba9aa27c),
	.w6(32'h3a7fbc7a),
	.w7(32'h39c70939),
	.w8(32'hbb28ff3f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd17e2),
	.w1(32'h3bac3b98),
	.w2(32'hb9896a94),
	.w3(32'h3b3ec16f),
	.w4(32'h3be1c38e),
	.w5(32'hbb69d27b),
	.w6(32'hba9b99f5),
	.w7(32'h3bb3bb54),
	.w8(32'hbb4cde13),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20c1ea),
	.w1(32'hbb6b3e5f),
	.w2(32'hbb2b6327),
	.w3(32'h3bbe2f15),
	.w4(32'h3c505d03),
	.w5(32'h3af1205e),
	.w6(32'hbb1272a2),
	.w7(32'hbc06f68f),
	.w8(32'h3b1b02ae),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15c954),
	.w1(32'h3c17ae8e),
	.w2(32'h3bee9b64),
	.w3(32'hbb6a2aca),
	.w4(32'h3a90a5c5),
	.w5(32'h3ae01bf5),
	.w6(32'hba74517b),
	.w7(32'h3bd82c01),
	.w8(32'h3a682d4b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa508e2),
	.w1(32'h3ab65527),
	.w2(32'hbb3dcbc2),
	.w3(32'hbbdbbff9),
	.w4(32'h3a806ebe),
	.w5(32'hba48aa83),
	.w6(32'h3a077f82),
	.w7(32'h3b9b5209),
	.w8(32'hbc2b36c0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82edcd),
	.w1(32'hbbabc97e),
	.w2(32'hb9bb60c4),
	.w3(32'hbb4037f0),
	.w4(32'hb6d0e213),
	.w5(32'h3b24a46a),
	.w6(32'hbb3762b2),
	.w7(32'hbabc7507),
	.w8(32'hb9cce3c3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04ad56),
	.w1(32'h3ca14898),
	.w2(32'h3c933052),
	.w3(32'h3c3dea87),
	.w4(32'h3c5366b6),
	.w5(32'h3aa95ed8),
	.w6(32'h3c1c0635),
	.w7(32'h3c0240d8),
	.w8(32'hbbf6fb82),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab214a3),
	.w1(32'h3c36fab2),
	.w2(32'hbb2b348d),
	.w3(32'h3b8bf7ce),
	.w4(32'h3a913953),
	.w5(32'h3be6151c),
	.w6(32'h3c26143a),
	.w7(32'h3bcd8e49),
	.w8(32'hbb83d980),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37a655),
	.w1(32'h3b824375),
	.w2(32'hbb01d0c3),
	.w3(32'h3a10c88e),
	.w4(32'hbb470dd3),
	.w5(32'h3b18c84a),
	.w6(32'h39708ed2),
	.w7(32'h3b5eddbd),
	.w8(32'hba7e1021),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1e72e),
	.w1(32'h3b34bb71),
	.w2(32'h3a9b173b),
	.w3(32'h3a8e186c),
	.w4(32'h3adf9c23),
	.w5(32'hbb07c505),
	.w6(32'hbbdf55fc),
	.w7(32'h3aea3eb2),
	.w8(32'h3afc4dc0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8580da),
	.w1(32'hb88c8879),
	.w2(32'h3b4e92d4),
	.w3(32'h398c6e4e),
	.w4(32'hb96e4cc2),
	.w5(32'h38e74707),
	.w6(32'hba7ed8bb),
	.w7(32'hb9c74131),
	.w8(32'h3b0d4f79),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0e457),
	.w1(32'h3b81b524),
	.w2(32'h3c2ea91f),
	.w3(32'h3b9d03e6),
	.w4(32'h3c03f337),
	.w5(32'h3b0ac69f),
	.w6(32'h3c13f400),
	.w7(32'h3c18db63),
	.w8(32'h3c0ae28f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b081d72),
	.w1(32'h3bc0a8ed),
	.w2(32'h3b404e63),
	.w3(32'hba8c88ce),
	.w4(32'h3b6a282c),
	.w5(32'h3be2807b),
	.w6(32'hbb3ed968),
	.w7(32'h3c114f9f),
	.w8(32'h3aa05ff6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf6648),
	.w1(32'hbb9ac547),
	.w2(32'h3b8677c1),
	.w3(32'hbbacfa4d),
	.w4(32'hb9d2fce5),
	.w5(32'hba2ef904),
	.w6(32'h3ab64e2f),
	.w7(32'h3b8060f7),
	.w8(32'hbb34f228),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af47863),
	.w1(32'hbbbbebc6),
	.w2(32'hba4156ed),
	.w3(32'hbab78a86),
	.w4(32'hbbf2d977),
	.w5(32'hbb5e1835),
	.w6(32'hbb9bcb9a),
	.w7(32'hb9e4c326),
	.w8(32'hbb0fdaaa),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2df42a),
	.w1(32'hbaa244e5),
	.w2(32'hbb8a0434),
	.w3(32'h3a99114a),
	.w4(32'h3aec15e0),
	.w5(32'h3ba2ed28),
	.w6(32'hba9fa2a9),
	.w7(32'hbb7ff23d),
	.w8(32'hbc0fbcd4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a118c),
	.w1(32'hbbc7d31d),
	.w2(32'h3b8d5b00),
	.w3(32'hbbad6124),
	.w4(32'hbbc95982),
	.w5(32'hbc1b10f3),
	.w6(32'h3abacb80),
	.w7(32'hbd0a47a1),
	.w8(32'hb7b43096),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba358057),
	.w1(32'h3b95da0e),
	.w2(32'h3bc49546),
	.w3(32'hbb971b21),
	.w4(32'hbb75e9d4),
	.w5(32'hbb82b626),
	.w6(32'h3ab403af),
	.w7(32'hbb3a073b),
	.w8(32'h3b820257),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc171df0),
	.w1(32'hba8f5d92),
	.w2(32'h3bffa83c),
	.w3(32'h3a59b7ef),
	.w4(32'hbafb9fe0),
	.w5(32'hbb7c61d7),
	.w6(32'hbbd6a1c4),
	.w7(32'h3b65170f),
	.w8(32'h3b98dee8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecb6b5),
	.w1(32'hb9e9f6ea),
	.w2(32'h3d185664),
	.w3(32'h3abe55d3),
	.w4(32'h3b9b2ccb),
	.w5(32'h3ac33839),
	.w6(32'hbac1a046),
	.w7(32'hba956d74),
	.w8(32'hbccee7ff),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8494e8),
	.w1(32'h3b3a62a2),
	.w2(32'h3a97448e),
	.w3(32'hbb418e67),
	.w4(32'h3a2a1f4d),
	.w5(32'h3a86c100),
	.w6(32'hbbd08945),
	.w7(32'h3b8db61b),
	.w8(32'h3bee5a8e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ab4d9),
	.w1(32'h3a63e1f0),
	.w2(32'hbab0337d),
	.w3(32'h3b2a8a36),
	.w4(32'h3c3a0abc),
	.w5(32'h3a6f1c90),
	.w6(32'h3a068b07),
	.w7(32'hbb61594b),
	.w8(32'hbb66448f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b66d9),
	.w1(32'hbc83a283),
	.w2(32'h3ae74da5),
	.w3(32'hbbbf6cfa),
	.w4(32'h3bbad528),
	.w5(32'hbb8d93a8),
	.w6(32'hba69dbd8),
	.w7(32'h3a677d68),
	.w8(32'h3b610d2c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a0d6b),
	.w1(32'hba6d92f9),
	.w2(32'hb9d3c244),
	.w3(32'h3ad0cae4),
	.w4(32'hba35c21d),
	.w5(32'h3b056c7f),
	.w6(32'h3ae7c58c),
	.w7(32'hbb8bc481),
	.w8(32'hbac5cb8f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c585f),
	.w1(32'hbc17f083),
	.w2(32'h3b51c961),
	.w3(32'h3b4b62a0),
	.w4(32'h3b8dfd79),
	.w5(32'h3abf8d8e),
	.w6(32'h3d32eae0),
	.w7(32'h3b83943e),
	.w8(32'h3ac3b7e2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb966bbf),
	.w1(32'h3beecdec),
	.w2(32'h3c13e887),
	.w3(32'hbc2992d5),
	.w4(32'hbafbe6f5),
	.w5(32'h3c6b09e0),
	.w6(32'h3ac13574),
	.w7(32'h3af669e3),
	.w8(32'h3c00caba),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b7fa9),
	.w1(32'hbb20f228),
	.w2(32'h3b239b3e),
	.w3(32'hbb21d747),
	.w4(32'hbd73889a),
	.w5(32'hbb76b9fa),
	.w6(32'h3bbb681f),
	.w7(32'hbbde8426),
	.w8(32'h3b91e5f2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1a588),
	.w1(32'hbc2b03f8),
	.w2(32'h3a4268bd),
	.w3(32'hbb043d67),
	.w4(32'hbc385620),
	.w5(32'h3b058956),
	.w6(32'h3bf18083),
	.w7(32'h3841c068),
	.w8(32'hbc83a23b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c6788),
	.w1(32'h3bb573af),
	.w2(32'h3b93294c),
	.w3(32'h3a0dd038),
	.w4(32'h3b9208f0),
	.w5(32'h39013107),
	.w6(32'h3c2d8ea1),
	.w7(32'hba8be1a6),
	.w8(32'hbce9e4d9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8845436),
	.w1(32'h3b231c1e),
	.w2(32'h39d2e432),
	.w3(32'hbd21313a),
	.w4(32'hbad4b774),
	.w5(32'hbb968cfe),
	.w6(32'h39c2ba0a),
	.w7(32'hbbd19dad),
	.w8(32'h3b98a19c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25096c),
	.w1(32'hb959c39f),
	.w2(32'h3bd56e53),
	.w3(32'hba9a499e),
	.w4(32'h3b9aaacc),
	.w5(32'hbc61b615),
	.w6(32'h3bd8e21a),
	.w7(32'hbb9c5e80),
	.w8(32'h3c55829f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee33e0),
	.w1(32'hbb28f621),
	.w2(32'hbbe292d2),
	.w3(32'hbb7b6a50),
	.w4(32'h3a4f567f),
	.w5(32'hba4de9ab),
	.w6(32'h3aa95615),
	.w7(32'h3bf15861),
	.w8(32'hbc06d603),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3f7cf),
	.w1(32'h3c3ea78d),
	.w2(32'h39d4e3f2),
	.w3(32'h3bb491dc),
	.w4(32'h3b36fe17),
	.w5(32'hbadee1f0),
	.w6(32'h3c01fc5d),
	.w7(32'h3d304f36),
	.w8(32'h3b0beef7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda9cf6),
	.w1(32'h3c03abe0),
	.w2(32'h3954d131),
	.w3(32'hbbd0cea6),
	.w4(32'hbb034490),
	.w5(32'h3b921f05),
	.w6(32'hbaa9b3c9),
	.w7(32'h3b4846d2),
	.w8(32'h3b076b65),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf22543),
	.w1(32'h3b6acb3c),
	.w2(32'h3bc957fe),
	.w3(32'h3b1a3694),
	.w4(32'hbab8a7c8),
	.w5(32'h3b6ae1a7),
	.w6(32'hbc591a73),
	.w7(32'h3b6ab861),
	.w8(32'h3a3a4230),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc2853c),
	.w1(32'h3ba2dcff),
	.w2(32'hba9425fc),
	.w3(32'hbb296e1a),
	.w4(32'h3bd7e17f),
	.w5(32'h3c855311),
	.w6(32'h3b35ea8e),
	.w7(32'h3b0ccff6),
	.w8(32'hbb0ae525),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befc09e),
	.w1(32'hb9f36217),
	.w2(32'h3bea3dd4),
	.w3(32'h3b6adae4),
	.w4(32'h3d0232ff),
	.w5(32'hbb8e29dc),
	.w6(32'h3c43ca22),
	.w7(32'h3c0670ac),
	.w8(32'h3bb5f3c7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c29d6),
	.w1(32'hbb45a0f4),
	.w2(32'h3cb64914),
	.w3(32'hbb532a6d),
	.w4(32'hbbe0cc09),
	.w5(32'h3b0a78d2),
	.w6(32'hbb186a7b),
	.w7(32'hbb99fa7e),
	.w8(32'hb9e52f11),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b937b46),
	.w1(32'h3854804e),
	.w2(32'h39177863),
	.w3(32'h3c81ca6c),
	.w4(32'hbcabbf0d),
	.w5(32'h3b9d46d5),
	.w6(32'hbaa3601d),
	.w7(32'h3899f3b4),
	.w8(32'hb79837be),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e40f98),
	.w1(32'h3ab24079),
	.w2(32'hba43b649),
	.w3(32'hbb344f45),
	.w4(32'h3aef3989),
	.w5(32'hb89250f3),
	.w6(32'hb9d422bd),
	.w7(32'h3b8b05d9),
	.w8(32'hba62ce1b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacc1a0),
	.w1(32'hbbc7f7b2),
	.w2(32'h3c1d3ab3),
	.w3(32'hbb992aed),
	.w4(32'hbaa67996),
	.w5(32'hb879d064),
	.w6(32'h3c724571),
	.w7(32'h3b260069),
	.w8(32'hbadf8c6d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf43648),
	.w1(32'hba380a69),
	.w2(32'h3ba6934c),
	.w3(32'hbbb57c5d),
	.w4(32'hb910adc6),
	.w5(32'hbbe5c74e),
	.w6(32'h3b44212b),
	.w7(32'hbb305464),
	.w8(32'hbb80c2d5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18ed8a),
	.w1(32'h3bf6be0d),
	.w2(32'hbc817f81),
	.w3(32'h3c4d7fdf),
	.w4(32'h3c3e12d8),
	.w5(32'hb9e533ec),
	.w6(32'h3c335008),
	.w7(32'h3b28dd98),
	.w8(32'h3bb98081),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e8a845),
	.w1(32'h39b08a7b),
	.w2(32'hba3aab62),
	.w3(32'h3aa9345d),
	.w4(32'hb9fbaf71),
	.w5(32'h3b080916),
	.w6(32'hba99b14c),
	.w7(32'hbbab8b62),
	.w8(32'h3a813f5d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba175981),
	.w1(32'hbb48e789),
	.w2(32'h3acd751a),
	.w3(32'hbbd9943e),
	.w4(32'h3b689907),
	.w5(32'hbb3d80e2),
	.w6(32'hba50e218),
	.w7(32'h3c0d99d1),
	.w8(32'h3b03c502),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8637e),
	.w1(32'hba91b0f3),
	.w2(32'h3c6fa78a),
	.w3(32'hbbf66e31),
	.w4(32'hbc24a485),
	.w5(32'hbbd79592),
	.w6(32'h3a0cbc9e),
	.w7(32'h3b375304),
	.w8(32'hba218e3a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93a269),
	.w1(32'hbbc4d23b),
	.w2(32'h3aef2285),
	.w3(32'h3b2b29bf),
	.w4(32'hbc0efc2f),
	.w5(32'hbc282f4f),
	.w6(32'hbb47dffc),
	.w7(32'hbb7276e5),
	.w8(32'h3b9642e9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d913c),
	.w1(32'h3c1144ae),
	.w2(32'h3b7117f5),
	.w3(32'hbb35a05c),
	.w4(32'hbb3b5220),
	.w5(32'hb9423d2c),
	.w6(32'hbaf48c98),
	.w7(32'hba03c7eb),
	.w8(32'hbb66aee0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cec7927),
	.w1(32'hbba01d19),
	.w2(32'hb90b61d8),
	.w3(32'h3c19ae94),
	.w4(32'hba768cac),
	.w5(32'hbbdcfeca),
	.w6(32'hbb13784a),
	.w7(32'hb997dd52),
	.w8(32'h3c2890db),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb990097),
	.w1(32'hbc14d632),
	.w2(32'hb7a60bdc),
	.w3(32'hbac995ed),
	.w4(32'h3af1cdb7),
	.w5(32'h3b25a15d),
	.w6(32'hbb6c4590),
	.w7(32'hbbb13e41),
	.w8(32'hbc06d4e2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4941ae),
	.w1(32'h3b55e542),
	.w2(32'h39950b42),
	.w3(32'h3bf53b9d),
	.w4(32'h3b4875b4),
	.w5(32'h3a218c4b),
	.w6(32'h3bb2df8b),
	.w7(32'hbbec866a),
	.w8(32'hb9911305),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb468ad2),
	.w1(32'hbae061a1),
	.w2(32'h3b8bcd4d),
	.w3(32'h3c164a30),
	.w4(32'h3b89eaac),
	.w5(32'h3c7e75b0),
	.w6(32'h390c0b76),
	.w7(32'hb9dbe818),
	.w8(32'hb8e6bd8c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abab34e),
	.w1(32'h3aa98eed),
	.w2(32'hbaebb3f7),
	.w3(32'hbb7dbbe6),
	.w4(32'hbc179406),
	.w5(32'hbbe9a322),
	.w6(32'hbb23d4c4),
	.w7(32'h3b297b07),
	.w8(32'hbacb5085),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4e2ff),
	.w1(32'hbb7ec35a),
	.w2(32'hba8f824b),
	.w3(32'h395e8851),
	.w4(32'h3b0af217),
	.w5(32'hbb49d0d3),
	.w6(32'hbc0a8a0a),
	.w7(32'h3bf3a0ce),
	.w8(32'h3be53370),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6daedf),
	.w1(32'h3a41fe10),
	.w2(32'hb9e8ed74),
	.w3(32'hbc436836),
	.w4(32'hbac1a83f),
	.w5(32'hb7c094dc),
	.w6(32'hbb9602a9),
	.w7(32'h3c1fc3f2),
	.w8(32'h3c5255d7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c274b55),
	.w1(32'hbc4d5a60),
	.w2(32'hbc15065e),
	.w3(32'h3b86c9a9),
	.w4(32'hbb494d9d),
	.w5(32'hbbcaaf6c),
	.w6(32'h3b62fc45),
	.w7(32'hbb9f71c5),
	.w8(32'hbb11d220),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8caa33),
	.w1(32'h3b8138b8),
	.w2(32'h3ac36fb9),
	.w3(32'h3bd66f5a),
	.w4(32'h3bb033fe),
	.w5(32'h3bae3041),
	.w6(32'h3b8c2921),
	.w7(32'hbbfae8ba),
	.w8(32'hba9e9fbe),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb177d4c),
	.w1(32'h3b83cb87),
	.w2(32'h3a198bb4),
	.w3(32'hba1b9203),
	.w4(32'h3b417990),
	.w5(32'h3b967d83),
	.w6(32'hbb66c5b2),
	.w7(32'hbb5c8fe9),
	.w8(32'hbb817cc9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a285cc9),
	.w1(32'hbc4ad5a4),
	.w2(32'h3c784fda),
	.w3(32'h3b1cad53),
	.w4(32'hbba704bd),
	.w5(32'hbbc209fa),
	.w6(32'hbb9ea9a7),
	.w7(32'h3c2ab075),
	.w8(32'hba82935d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b0e92),
	.w1(32'hbbeec36b),
	.w2(32'hbab39bb2),
	.w3(32'hbb3bb635),
	.w4(32'h39ccb046),
	.w5(32'hb92dd07f),
	.w6(32'hbb700517),
	.w7(32'h3bee37f3),
	.w8(32'hbbf5e6ed),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09a3f2),
	.w1(32'hbbe79de4),
	.w2(32'h3a51f6f2),
	.w3(32'h3b5b5e7c),
	.w4(32'h3aca307f),
	.w5(32'hbb0024d9),
	.w6(32'hba93a9fc),
	.w7(32'hba369fb7),
	.w8(32'h3d0b4ce4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdc2fd),
	.w1(32'h3b97b334),
	.w2(32'hbb171659),
	.w3(32'hbb572007),
	.w4(32'hba2a4f2a),
	.w5(32'h3c0b7047),
	.w6(32'h39de480b),
	.w7(32'hbbab81de),
	.w8(32'h3caadb40),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccef3c),
	.w1(32'h39e06b3a),
	.w2(32'h3a90253d),
	.w3(32'h3b9c1c86),
	.w4(32'h3bdb863b),
	.w5(32'h3b2615bb),
	.w6(32'h3b70f33a),
	.w7(32'hbb56dde8),
	.w8(32'hbaf00ae0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6287be),
	.w1(32'hbb848dd7),
	.w2(32'h386ec568),
	.w3(32'hbba47897),
	.w4(32'h3be4c199),
	.w5(32'hbb0b1a6b),
	.w6(32'hbbccff93),
	.w7(32'hbb7f3f6a),
	.w8(32'h3baff708),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b382951),
	.w1(32'h3cc06818),
	.w2(32'hbc499e54),
	.w3(32'h3a1ac01b),
	.w4(32'h3a84d432),
	.w5(32'hbbaf8f8f),
	.w6(32'hbb2ae03a),
	.w7(32'h3b991e3a),
	.w8(32'hbb294ad0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e97c9),
	.w1(32'h3bf49d56),
	.w2(32'h3c4be269),
	.w3(32'h3c41fe89),
	.w4(32'h3c18ae4d),
	.w5(32'h3a9fa998),
	.w6(32'h3c7ee4d4),
	.w7(32'h3b1e7ae1),
	.w8(32'h3bdab9f9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b992a),
	.w1(32'hbaaec327),
	.w2(32'h3a03cbce),
	.w3(32'hbba44ad4),
	.w4(32'h3b5d7197),
	.w5(32'h3aaf916e),
	.w6(32'h3c50890d),
	.w7(32'h3bd5bcde),
	.w8(32'hbab6f245),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373b95e5),
	.w1(32'h3a5bffa6),
	.w2(32'hbb7b6a02),
	.w3(32'hbaf450f5),
	.w4(32'h3ae0b5db),
	.w5(32'hbb898186),
	.w6(32'h3bc825c1),
	.w7(32'hbbb7894a),
	.w8(32'hbbca529d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a8790),
	.w1(32'hba6e6a03),
	.w2(32'hbc2987ad),
	.w3(32'h3a8e5fdd),
	.w4(32'h3abd0304),
	.w5(32'hb9f9f5ca),
	.w6(32'h3a8ec120),
	.w7(32'h3ca4d483),
	.w8(32'h3bb32d3b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c706f3),
	.w1(32'hbc5b9d5b),
	.w2(32'h3992c9f1),
	.w3(32'hbbe679b1),
	.w4(32'h3c73cbaa),
	.w5(32'h3a4f96e5),
	.w6(32'hba6f1bf7),
	.w7(32'hbc605ab0),
	.w8(32'hbc5612dc),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf6fce),
	.w1(32'h3a519cc1),
	.w2(32'hb9cdcced),
	.w3(32'h39f35b00),
	.w4(32'h3c94544e),
	.w5(32'hbbcb473f),
	.w6(32'hbbe0882e),
	.w7(32'h3cd91d6c),
	.w8(32'hb97588fb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfa3c8),
	.w1(32'h3b7f5618),
	.w2(32'hbb1de013),
	.w3(32'h3a05c01a),
	.w4(32'hbb987752),
	.w5(32'hbaf0f896),
	.w6(32'h3c0ac741),
	.w7(32'h3b012707),
	.w8(32'h3bc85eec),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbba1b1),
	.w1(32'hbb55f2c2),
	.w2(32'h3ba0bdf4),
	.w3(32'hbb2822bd),
	.w4(32'hbb9ced54),
	.w5(32'h3b57951c),
	.w6(32'h3bb9326c),
	.w7(32'hbb548ea2),
	.w8(32'h3b74a062),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2aa595),
	.w1(32'hbc00b637),
	.w2(32'h3c27a8aa),
	.w3(32'h3ab79351),
	.w4(32'hbc195585),
	.w5(32'h3b2ff1b5),
	.w6(32'hbb1dd323),
	.w7(32'hbc08f0d8),
	.w8(32'hb96cc9fd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07f7b2),
	.w1(32'hbbae071a),
	.w2(32'hbb916361),
	.w3(32'hbb0733be),
	.w4(32'h39f11e84),
	.w5(32'hb9af03a5),
	.w6(32'h3b85f846),
	.w7(32'hbc2402b2),
	.w8(32'h3ae1d992),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f91f6),
	.w1(32'h3a11bea4),
	.w2(32'h3b8c86c6),
	.w3(32'h3b6897a6),
	.w4(32'h3ada731b),
	.w5(32'hbbadf090),
	.w6(32'h3bb06d77),
	.w7(32'h3c8636ab),
	.w8(32'h3b80453e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a26efe),
	.w1(32'h3c070c37),
	.w2(32'h3b98b597),
	.w3(32'hbb6d799d),
	.w4(32'hbc1e7668),
	.w5(32'h3c9cc513),
	.w6(32'h3bcf1863),
	.w7(32'hbad6e275),
	.w8(32'hba66cbf9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb877108),
	.w1(32'hbb1110f8),
	.w2(32'h3c8f66ff),
	.w3(32'hbb5816d4),
	.w4(32'hbbb61b95),
	.w5(32'h3c4862fc),
	.w6(32'h3be82008),
	.w7(32'h3c1ed6b8),
	.w8(32'h3c3715e3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2900d),
	.w1(32'h3bbc2058),
	.w2(32'hbbf2fb2e),
	.w3(32'h3c3526df),
	.w4(32'h3c9cb6a1),
	.w5(32'hb97a6751),
	.w6(32'h3c0336b0),
	.w7(32'h3b215ab1),
	.w8(32'hba372e7d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51b405),
	.w1(32'hbb9f61c2),
	.w2(32'h3a21782c),
	.w3(32'h3a2e9e27),
	.w4(32'hbb76f4b8),
	.w5(32'h3a80ffb1),
	.w6(32'h3d5090c7),
	.w7(32'h3c8a509d),
	.w8(32'h39d8125a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03126a),
	.w1(32'hbb4932e1),
	.w2(32'h3a824df4),
	.w3(32'h3bdeea65),
	.w4(32'hbb91efec),
	.w5(32'h3c34d8f5),
	.w6(32'h3c145b9f),
	.w7(32'h3ba975af),
	.w8(32'hbb6c2ede),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a78ad),
	.w1(32'hbc0a49e0),
	.w2(32'h3be47473),
	.w3(32'h3c4d4cdf),
	.w4(32'hbbc2c578),
	.w5(32'hbb1a636b),
	.w6(32'hbacf4c21),
	.w7(32'hbb88b29e),
	.w8(32'hb9b7911a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0eac66),
	.w1(32'h3c6a5e95),
	.w2(32'hbc8aaffd),
	.w3(32'hb9e8758e),
	.w4(32'h3c0d441a),
	.w5(32'hbb2605cb),
	.w6(32'hbbf9823b),
	.w7(32'h3c083235),
	.w8(32'hbb43b5d7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9be2a),
	.w1(32'hbc52f0ed),
	.w2(32'h3b01e1f6),
	.w3(32'hbb4d9c86),
	.w4(32'hbb885fe7),
	.w5(32'hbb3241ca),
	.w6(32'h3a37ebbb),
	.w7(32'h3ca89e92),
	.w8(32'hbb6f50ca),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfc2e21),
	.w1(32'h3a31baeb),
	.w2(32'h3b42138c),
	.w3(32'hbbbc88a2),
	.w4(32'hbbbc4654),
	.w5(32'hbaef5b44),
	.w6(32'h3c169db0),
	.w7(32'h3ba2fba4),
	.w8(32'h3b3e8b20),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae6a63),
	.w1(32'hb9d74f5f),
	.w2(32'h3b96bbbd),
	.w3(32'hbc33c20d),
	.w4(32'h3a18fdf3),
	.w5(32'hbad08459),
	.w6(32'hbbbea8c0),
	.w7(32'hbbd3d750),
	.w8(32'hb7c8471e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d837b),
	.w1(32'hbbd621b3),
	.w2(32'hbb76f031),
	.w3(32'h3ae7e2b4),
	.w4(32'h3b23fac6),
	.w5(32'h3b81d11d),
	.w6(32'h3bc8d1e9),
	.w7(32'hbc17c230),
	.w8(32'h3b89ffd9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25fcb3),
	.w1(32'hbb8a18be),
	.w2(32'h3a845d13),
	.w3(32'h3b9758f2),
	.w4(32'hbb634c92),
	.w5(32'hbb9c9497),
	.w6(32'hba1d9105),
	.w7(32'hbc669a36),
	.w8(32'hbb208fcf),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0ce4b),
	.w1(32'h3c0206cf),
	.w2(32'h3c015149),
	.w3(32'h3b1e8c1c),
	.w4(32'h3c173911),
	.w5(32'h3c1c98bf),
	.w6(32'h3c02ca25),
	.w7(32'hbb8bf5e4),
	.w8(32'hbb58d6db),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e711a),
	.w1(32'h3977c46d),
	.w2(32'h38ec6c7c),
	.w3(32'hbbb54982),
	.w4(32'hbbb598c5),
	.w5(32'h3ba05ec8),
	.w6(32'h3baedc0d),
	.w7(32'h3c726628),
	.w8(32'h3b355ccc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb96e3),
	.w1(32'h3a7bd509),
	.w2(32'h3c156526),
	.w3(32'h3a225020),
	.w4(32'hb8d80a4c),
	.w5(32'h3b0fd28f),
	.w6(32'hbae5f04f),
	.w7(32'h3aeeadb7),
	.w8(32'h3b33daba),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ca9b4),
	.w1(32'hbaa51274),
	.w2(32'h3cae1488),
	.w3(32'hbc1b8e77),
	.w4(32'hb9f7eaa6),
	.w5(32'h3c2c45f0),
	.w6(32'hbace2db0),
	.w7(32'h3c07671a),
	.w8(32'h3d37059d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11fe04),
	.w1(32'hbc1e91b2),
	.w2(32'h3b659185),
	.w3(32'hb89751cc),
	.w4(32'h3b46ae64),
	.w5(32'hbac65cef),
	.w6(32'hbba7ba70),
	.w7(32'h3ae2acd5),
	.w8(32'h3bf3804d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47e130),
	.w1(32'h3c9f9baf),
	.w2(32'h3ca0892a),
	.w3(32'hbc08f0d4),
	.w4(32'h3b5d81ba),
	.w5(32'hbbd17d89),
	.w6(32'h3cac914f),
	.w7(32'h3c02e5e1),
	.w8(32'h3b3e012c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac15d88),
	.w1(32'hbb283b25),
	.w2(32'hbaeae080),
	.w3(32'hbb30178d),
	.w4(32'hbb2b2732),
	.w5(32'h3b1c68c6),
	.w6(32'h3b049705),
	.w7(32'h3c0fa5ad),
	.w8(32'h3bb25bd2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7dd45d),
	.w1(32'h3a15947f),
	.w2(32'hba5c7593),
	.w3(32'hbb979b47),
	.w4(32'h3b0d5bd0),
	.w5(32'h3a352ea5),
	.w6(32'h3ae3aa96),
	.w7(32'hba529bce),
	.w8(32'hb9aaaa3a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babc55f),
	.w1(32'hbb557223),
	.w2(32'h3a7ef813),
	.w3(32'hba4e8911),
	.w4(32'hbbdd9d5d),
	.w5(32'hbad32663),
	.w6(32'h3b6e0897),
	.w7(32'hba060a0f),
	.w8(32'h39abe315),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc274276),
	.w1(32'h3be5af1c),
	.w2(32'hbac00543),
	.w3(32'h3c67d99e),
	.w4(32'h3a19138a),
	.w5(32'h3bd16d05),
	.w6(32'h3c827b01),
	.w7(32'h3c0c03bb),
	.w8(32'hbbb7a98f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b784b),
	.w1(32'hb8f4d438),
	.w2(32'h38f994b2),
	.w3(32'h3b8f84b4),
	.w4(32'hbc3f0f8a),
	.w5(32'h3c6ae36f),
	.w6(32'h3a08e6c8),
	.w7(32'hbbd09dab),
	.w8(32'hba6a1be0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38dada),
	.w1(32'hbbd7aa42),
	.w2(32'h3b45fe07),
	.w3(32'h3c041344),
	.w4(32'h3c519544),
	.w5(32'h3a80175c),
	.w6(32'h3cf38399),
	.w7(32'hba0f2c04),
	.w8(32'hbad345e9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9d8fc),
	.w1(32'hbb8d5e49),
	.w2(32'h3b373865),
	.w3(32'hbb90a895),
	.w4(32'hbb27ac91),
	.w5(32'h3aae1782),
	.w6(32'hbb2dca63),
	.w7(32'h3b422a29),
	.w8(32'h3af9c216),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a659b97),
	.w1(32'hba09d867),
	.w2(32'hbb926a91),
	.w3(32'h3bcddfe1),
	.w4(32'hba88b5e7),
	.w5(32'h39e3cd7f),
	.w6(32'hbbabf326),
	.w7(32'hbba08832),
	.w8(32'h3bda5f49),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff23ad),
	.w1(32'hbaccd491),
	.w2(32'hba957f79),
	.w3(32'hbc90165d),
	.w4(32'h39778649),
	.w5(32'h3ac2875d),
	.w6(32'hb9dc6208),
	.w7(32'h3bdc9dfd),
	.w8(32'hba00eb98),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0845c7),
	.w1(32'hbb6b2225),
	.w2(32'hb9ba7be3),
	.w3(32'hbb342bc9),
	.w4(32'hbb381156),
	.w5(32'h3d12ef8b),
	.w6(32'h3a91b99d),
	.w7(32'h3b2285c9),
	.w8(32'h3baa9db0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b585197),
	.w1(32'h3b2509b6),
	.w2(32'h3a91e193),
	.w3(32'hbb5334ce),
	.w4(32'h3a4b49f8),
	.w5(32'hba1b02eb),
	.w6(32'h3ba8544b),
	.w7(32'hbb8578f8),
	.w8(32'h3934d70e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc389ac7),
	.w1(32'h3ac1fa7e),
	.w2(32'hbb57f073),
	.w3(32'hbb3f1789),
	.w4(32'h3b85d88c),
	.w5(32'hba816c37),
	.w6(32'h39493d8a),
	.w7(32'h3b92ac26),
	.w8(32'hba193990),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa176ad),
	.w1(32'h3b7cea9c),
	.w2(32'hbb2fd644),
	.w3(32'hbb009583),
	.w4(32'hba2f0c53),
	.w5(32'hba868b99),
	.w6(32'hb9ed2f2b),
	.w7(32'hba94b364),
	.w8(32'hb8bd0c2d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79938f),
	.w1(32'h3a811a81),
	.w2(32'hbc07873e),
	.w3(32'h3b2cba72),
	.w4(32'h3b821cb9),
	.w5(32'hbb3f157c),
	.w6(32'hbbbb234c),
	.w7(32'h39d1f921),
	.w8(32'hb9813358),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6526d),
	.w1(32'hbad7d26b),
	.w2(32'h3bd84240),
	.w3(32'hbb0336b9),
	.w4(32'h3b08dc9e),
	.w5(32'h3a702594),
	.w6(32'h3b8da3b2),
	.w7(32'h3bc1a4fa),
	.w8(32'h3ba4b7ac),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5b530),
	.w1(32'hbbf3c2ae),
	.w2(32'h3b50882e),
	.w3(32'hba3c2fea),
	.w4(32'hbb12baa3),
	.w5(32'h3a00a62e),
	.w6(32'h3b19a99a),
	.w7(32'h3b0e7e15),
	.w8(32'hbb6b7236),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cea16),
	.w1(32'hbb8ee8b4),
	.w2(32'h3c0c46e1),
	.w3(32'hbae61040),
	.w4(32'h3b77368d),
	.w5(32'h3be02860),
	.w6(32'hba36bc37),
	.w7(32'hb986c1cb),
	.w8(32'hb6e538a1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc029577),
	.w1(32'hbace06d1),
	.w2(32'h3ab9b10d),
	.w3(32'h3a0a29a9),
	.w4(32'hbbc7bdcc),
	.w5(32'hbb70e7b1),
	.w6(32'h3b41e8d6),
	.w7(32'hbaf23800),
	.w8(32'h3ba32ff8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8db48),
	.w1(32'h3c3f2639),
	.w2(32'hbbd02699),
	.w3(32'h38586b73),
	.w4(32'h3abe48c3),
	.w5(32'h3b975cc7),
	.w6(32'h3a5c9819),
	.w7(32'hbbe9837f),
	.w8(32'hbc272378),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc97345),
	.w1(32'h3a8edfeb),
	.w2(32'hbad14fe4),
	.w3(32'h39bd7fdd),
	.w4(32'h3b74af69),
	.w5(32'h3cbc65fc),
	.w6(32'hbbe31059),
	.w7(32'h3cd8969e),
	.w8(32'h3afe2e37),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb036e61),
	.w1(32'hb787e73c),
	.w2(32'h3b967c27),
	.w3(32'h3b1a6648),
	.w4(32'hba088f87),
	.w5(32'hbb3d8e46),
	.w6(32'hb9f61ebd),
	.w7(32'h382d388e),
	.w8(32'hbb40d283),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91b2a8),
	.w1(32'h3b42000b),
	.w2(32'hbb04ddb1),
	.w3(32'hb99811be),
	.w4(32'h3b7e17b7),
	.w5(32'hbbbce0c0),
	.w6(32'h3b2dda1c),
	.w7(32'h3b202b0d),
	.w8(32'h3959cf51),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc90899),
	.w1(32'hbcb70f80),
	.w2(32'h3ae1e7bc),
	.w3(32'hbbdb8683),
	.w4(32'hbad3c462),
	.w5(32'hbb0d1d94),
	.w6(32'h3a355e02),
	.w7(32'hbb173cf7),
	.w8(32'h3b4dd97a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b9cda),
	.w1(32'hbbfba9e8),
	.w2(32'hba951e25),
	.w3(32'h3b4575e6),
	.w4(32'hbacfe197),
	.w5(32'hb9c17f60),
	.w6(32'h3b189767),
	.w7(32'h3b9efe5c),
	.w8(32'h3bae8b8e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb19fb1),
	.w1(32'h3a805333),
	.w2(32'hbc174164),
	.w3(32'h3b8f9705),
	.w4(32'h3c1b53e3),
	.w5(32'h3b0c9a9d),
	.w6(32'hbacd3f78),
	.w7(32'h3bbd7cba),
	.w8(32'hbb28bec7),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb577d),
	.w1(32'h39e02a1a),
	.w2(32'hbab62911),
	.w3(32'hba531780),
	.w4(32'h3b648911),
	.w5(32'hba8ce251),
	.w6(32'h3a40bfcb),
	.w7(32'hbaf25753),
	.w8(32'hbb550ae5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf7e08),
	.w1(32'hbb75d050),
	.w2(32'h396cdf22),
	.w3(32'h3cd335ea),
	.w4(32'h3ccf9fa9),
	.w5(32'hbb87dba4),
	.w6(32'hba5592a5),
	.w7(32'h39b4b3eb),
	.w8(32'h3aa03d5e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb309afa),
	.w1(32'hbb64beba),
	.w2(32'hb9e5afa1),
	.w3(32'h3ce208f9),
	.w4(32'hbbb927b7),
	.w5(32'h3cc54f40),
	.w6(32'h3b01f698),
	.w7(32'hbbb9fc9a),
	.w8(32'hbb1df8d9),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ce64c),
	.w1(32'hbb8548ad),
	.w2(32'hbbb788ba),
	.w3(32'h39f3d19a),
	.w4(32'hbc20f441),
	.w5(32'hbbe648cc),
	.w6(32'h3c090f36),
	.w7(32'h3ad95e4b),
	.w8(32'h3b2032c3),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6c5fc),
	.w1(32'hbaf9ea26),
	.w2(32'hbbb1b05e),
	.w3(32'h3ae47e81),
	.w4(32'h3bbd93ea),
	.w5(32'h3c00fe92),
	.w6(32'h3ba401d3),
	.w7(32'h3a318512),
	.w8(32'h3b28903b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad0885),
	.w1(32'hb918eb63),
	.w2(32'h3bbb6a8d),
	.w3(32'hbaa99006),
	.w4(32'h3b5e042e),
	.w5(32'hb99ef7ff),
	.w6(32'h36af536e),
	.w7(32'h3ae969d0),
	.w8(32'hb9042dce),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64189f),
	.w1(32'h3b9bdc3c),
	.w2(32'hba13ec92),
	.w3(32'hb923d395),
	.w4(32'h3b303b8e),
	.w5(32'hbb11ef7d),
	.w6(32'h3b20f95b),
	.w7(32'hbc1b30f1),
	.w8(32'h3bb88946),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb78737),
	.w1(32'h3aae7e61),
	.w2(32'h3b1d6d30),
	.w3(32'h3c051f7e),
	.w4(32'h3a97bc22),
	.w5(32'h3aebda8c),
	.w6(32'h3bab27d2),
	.w7(32'h3b913cc3),
	.w8(32'h3b5b3eed),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4906c),
	.w1(32'hbb390a70),
	.w2(32'hbbbcbb34),
	.w3(32'h3b3f6a3f),
	.w4(32'hbb32eb40),
	.w5(32'hbc18a5ba),
	.w6(32'hbbbe54db),
	.w7(32'h3a19efe7),
	.w8(32'h3b568456),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2cffe),
	.w1(32'hbadad84d),
	.w2(32'hbbd2b1b4),
	.w3(32'h3ad478a8),
	.w4(32'h3bb6b750),
	.w5(32'h3c0ceb28),
	.w6(32'hbb852123),
	.w7(32'h3a7a21be),
	.w8(32'h3b1d5bad),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f9e9d),
	.w1(32'hbad7e731),
	.w2(32'h3b8b564e),
	.w3(32'hb9d47835),
	.w4(32'h3b46b89a),
	.w5(32'hbc064329),
	.w6(32'h3b6cb4ed),
	.w7(32'h3b9726ea),
	.w8(32'h3a9e0632),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79f2a4),
	.w1(32'hbcde9c8f),
	.w2(32'h3b1c18fb),
	.w3(32'hbbb106b7),
	.w4(32'hbc20a00a),
	.w5(32'h3b8f042e),
	.w6(32'hba5a7029),
	.w7(32'hbb68e1db),
	.w8(32'h3bf8eab4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe26ea),
	.w1(32'h3b2cc776),
	.w2(32'h3ac803f6),
	.w3(32'h3b8a66cd),
	.w4(32'h3c566b67),
	.w5(32'hbb2233bf),
	.w6(32'h37f5627f),
	.w7(32'h3ac124ab),
	.w8(32'hbb545a8e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b988f06),
	.w1(32'h3bd06bd8),
	.w2(32'hbacb3d17),
	.w3(32'hb8f9b51e),
	.w4(32'hbbe1413e),
	.w5(32'h3b1c8e98),
	.w6(32'h3c9148f6),
	.w7(32'hbb4ac48e),
	.w8(32'h386d080e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93a5b4),
	.w1(32'h3ae3d6af),
	.w2(32'h3c080dee),
	.w3(32'h38105573),
	.w4(32'hbc94ea2e),
	.w5(32'h3b70e5a1),
	.w6(32'hbbfc4ada),
	.w7(32'h3b45c37a),
	.w8(32'hbc10fa5d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a656a42),
	.w1(32'hbbcb6eec),
	.w2(32'hbbd972f8),
	.w3(32'hbb79974b),
	.w4(32'h3a59308c),
	.w5(32'hbac76d15),
	.w6(32'h3bf91b9d),
	.w7(32'hbb5fa437),
	.w8(32'hbb26806a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cb31f),
	.w1(32'hbba49061),
	.w2(32'h3b86d7e7),
	.w3(32'hbbbb1709),
	.w4(32'hbbf496ee),
	.w5(32'h3b49a133),
	.w6(32'h3a8bbc63),
	.w7(32'h3b089a51),
	.w8(32'h3beb3e74),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc36c1a),
	.w1(32'h3bbc3e16),
	.w2(32'h3a6ae665),
	.w3(32'hbb597acc),
	.w4(32'h3cb4714b),
	.w5(32'hbbed2bf2),
	.w6(32'hbbb39675),
	.w7(32'hbaf4cec1),
	.w8(32'hbb7a5465),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387d02b9),
	.w1(32'hbbef557e),
	.w2(32'hbc3c718f),
	.w3(32'h3a823b84),
	.w4(32'hba7c6358),
	.w5(32'h3b0f3d7c),
	.w6(32'hbb2b2c85),
	.w7(32'hbb395fd9),
	.w8(32'h3b873de8),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1d9a47),
	.w1(32'hbb3c8e32),
	.w2(32'h3a6becbf),
	.w3(32'hbc0c6b3d),
	.w4(32'hbb59df02),
	.w5(32'hbb64e02d),
	.w6(32'h3bea5ded),
	.w7(32'h3c32b8cb),
	.w8(32'h3c2a89f0),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc1982),
	.w1(32'h39aebc63),
	.w2(32'hbb9936b4),
	.w3(32'hbb53dadc),
	.w4(32'hba8e1640),
	.w5(32'h3b4b7e6c),
	.w6(32'h3b784399),
	.w7(32'h3b81d433),
	.w8(32'h3ca82c68),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10e0a2),
	.w1(32'h3bd9cf20),
	.w2(32'h3acece5d),
	.w3(32'hbaa26eb6),
	.w4(32'hbb0f912f),
	.w5(32'hbc401df8),
	.w6(32'h3c11120b),
	.w7(32'h3add19ae),
	.w8(32'hbb9a0028),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8fefb),
	.w1(32'h3b385535),
	.w2(32'hbcc03138),
	.w3(32'h3bfdd037),
	.w4(32'h3b2357ac),
	.w5(32'h3b082de4),
	.w6(32'hbbe9175c),
	.w7(32'hba97f0ab),
	.w8(32'hba25dfce),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fa8a5),
	.w1(32'hbb40fcb8),
	.w2(32'hbc20e09a),
	.w3(32'h3a309773),
	.w4(32'h3a25425d),
	.w5(32'h3a682169),
	.w6(32'h3c70c45d),
	.w7(32'hbba35f9d),
	.w8(32'h3ba71e5b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e2d40),
	.w1(32'h3b88b37d),
	.w2(32'h3a53f138),
	.w3(32'h3b3e63e2),
	.w4(32'hbb8b8898),
	.w5(32'hbb6b7f21),
	.w6(32'hba5aceca),
	.w7(32'h3ab1f950),
	.w8(32'h3b590772),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c397),
	.w1(32'hbb3701c6),
	.w2(32'hbc8b3eda),
	.w3(32'hbb32e096),
	.w4(32'hbc590505),
	.w5(32'hbc47a316),
	.w6(32'h3b5d48a6),
	.w7(32'hba639ce0),
	.w8(32'h3a12be0b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966e7fa),
	.w1(32'hbbb2225f),
	.w2(32'hb9b64a21),
	.w3(32'h3a98a2ea),
	.w4(32'h3aec0b90),
	.w5(32'hbb7ca2eb),
	.w6(32'hbc3c3a8c),
	.w7(32'h3b29b185),
	.w8(32'hbad1c0cb),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b514256),
	.w1(32'h3cbee5bf),
	.w2(32'hbb267579),
	.w3(32'h3b97800f),
	.w4(32'h3abb5e83),
	.w5(32'hba44ef0d),
	.w6(32'hbbd72477),
	.w7(32'h3a9d1694),
	.w8(32'h3b7c8d50),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb8a1b),
	.w1(32'h3b890344),
	.w2(32'hb97560d7),
	.w3(32'h38dfbe0b),
	.w4(32'h3a8067b3),
	.w5(32'h3a119394),
	.w6(32'h3bec2448),
	.w7(32'h3baae86d),
	.w8(32'hbbd0c147),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e5072),
	.w1(32'hbaf8746a),
	.w2(32'h3a880c22),
	.w3(32'hbb2679bb),
	.w4(32'h3a4c3f9e),
	.w5(32'h3b6cc163),
	.w6(32'hb9e2bb91),
	.w7(32'h3c2c150c),
	.w8(32'h3bdbd213),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01640f),
	.w1(32'h3b6ef783),
	.w2(32'hbac73ef6),
	.w3(32'hbb714e51),
	.w4(32'hbbbbd17b),
	.w5(32'h3bbbc1b7),
	.w6(32'h3c759555),
	.w7(32'h3d344ffe),
	.w8(32'hbc3176cb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a35c5),
	.w1(32'h39d86a07),
	.w2(32'hbc9dae74),
	.w3(32'h3bc84ebf),
	.w4(32'h3b6db349),
	.w5(32'hbaab41c9),
	.w6(32'h3c96acf4),
	.w7(32'h3b0d94ab),
	.w8(32'hbc00022a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab17527),
	.w1(32'hbb99e707),
	.w2(32'hba2162a5),
	.w3(32'hbc20c9d1),
	.w4(32'h3cd53c70),
	.w5(32'hb83382a1),
	.w6(32'hbacf4266),
	.w7(32'hbb51222a),
	.w8(32'hbca38775),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40f949),
	.w1(32'hbab32148),
	.w2(32'h39764da2),
	.w3(32'hbbe66984),
	.w4(32'h39e93c46),
	.w5(32'hb9c5438c),
	.w6(32'hbb54a4c3),
	.w7(32'h3b79c785),
	.w8(32'h3aae6cb1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5f436),
	.w1(32'h3a711342),
	.w2(32'hba1b295b),
	.w3(32'hbbd02c35),
	.w4(32'h3a4b4b5c),
	.w5(32'hbc184086),
	.w6(32'h3a9c708a),
	.w7(32'h3aa72c04),
	.w8(32'hbc1edc70),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49db9c),
	.w1(32'h3b6f124e),
	.w2(32'hbb429013),
	.w3(32'hba5c4ed7),
	.w4(32'hbb14d9b3),
	.w5(32'hbb9dc177),
	.w6(32'hbb8e4bab),
	.w7(32'hba26bb12),
	.w8(32'hb9bfa7e1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae85e3b),
	.w1(32'h3b642124),
	.w2(32'hbaa25a5f),
	.w3(32'hbaef2992),
	.w4(32'h3b6a7a21),
	.w5(32'hbb2716e0),
	.w6(32'h3914b00f),
	.w7(32'h3b323e6e),
	.w8(32'h3b9fc017),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadacd0),
	.w1(32'hbb3e941c),
	.w2(32'h3d25341b),
	.w3(32'hbbe420ed),
	.w4(32'hbcd1034d),
	.w5(32'h3c165b4d),
	.w6(32'h3c2140d6),
	.w7(32'hbae78b59),
	.w8(32'h3c42e0eb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39f151),
	.w1(32'h3b17e30e),
	.w2(32'hbad3aa2b),
	.w3(32'hbab6ea74),
	.w4(32'h3c3ddca7),
	.w5(32'h3c0b7bec),
	.w6(32'h3ad30542),
	.w7(32'h3b81781a),
	.w8(32'hbb11c8e6),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b2d2c),
	.w1(32'h3aa19e08),
	.w2(32'hbbddcf16),
	.w3(32'hbc107250),
	.w4(32'hbb8a7dec),
	.w5(32'h3c61e920),
	.w6(32'h3aa67fa0),
	.w7(32'h3b759812),
	.w8(32'h3cce06fe),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc458e3),
	.w1(32'hb790ef2f),
	.w2(32'hbabad6b6),
	.w3(32'h3a4b377e),
	.w4(32'hbae7a1c8),
	.w5(32'hbb81b8f2),
	.w6(32'hbaa17254),
	.w7(32'h3b1a4b57),
	.w8(32'h3c6bd76a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5859d),
	.w1(32'h398ff88e),
	.w2(32'h3b972794),
	.w3(32'hbac3066f),
	.w4(32'h3c04bd56),
	.w5(32'h3b5c1210),
	.w6(32'hbc6d39e6),
	.w7(32'h39e229b1),
	.w8(32'h3b1e0c2b),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07dd17),
	.w1(32'h3bd864f7),
	.w2(32'hbab46b41),
	.w3(32'h3c249686),
	.w4(32'h3b784c8f),
	.w5(32'h387c8972),
	.w6(32'h3a9a1a7f),
	.w7(32'hbbb26039),
	.w8(32'hbc127e1d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5083ff),
	.w1(32'hbbdbf42d),
	.w2(32'hbb6ef0dd),
	.w3(32'h3c39a232),
	.w4(32'hbac5b164),
	.w5(32'hbc2f37c2),
	.w6(32'h3b35375b),
	.w7(32'h3c070191),
	.w8(32'hba79726c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8667ff),
	.w1(32'hbbbf917f),
	.w2(32'hbc03c2e2),
	.w3(32'h3c23f368),
	.w4(32'h3aa3728c),
	.w5(32'hbbfd0b22),
	.w6(32'h3bffe105),
	.w7(32'h3bad178c),
	.w8(32'hbba635df),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58b3ef),
	.w1(32'h3b07c754),
	.w2(32'hbb5e72ad),
	.w3(32'hbb8a7bd9),
	.w4(32'h3a086de9),
	.w5(32'hbc3ce5ca),
	.w6(32'h3c00a303),
	.w7(32'hbcc97848),
	.w8(32'h3c60aa43),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9626d2a),
	.w1(32'hbb720e48),
	.w2(32'hbb062be0),
	.w3(32'hba4d708a),
	.w4(32'h3c48807f),
	.w5(32'hbc4c7437),
	.w6(32'hbbcdb8bb),
	.w7(32'h3b55b2d9),
	.w8(32'hbbb28cde),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe209b),
	.w1(32'hbba484ab),
	.w2(32'hbb51d74d),
	.w3(32'h3d90c6f2),
	.w4(32'h3c0107d8),
	.w5(32'hbb9a2c92),
	.w6(32'hbbd40b9d),
	.w7(32'hbab6b0fb),
	.w8(32'hb8635d56),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fc071),
	.w1(32'h3c620e9e),
	.w2(32'h3be60b4a),
	.w3(32'h3b5df570),
	.w4(32'hbba1a494),
	.w5(32'hbbdba70a),
	.w6(32'h3b3b5c68),
	.w7(32'h3b75cd5f),
	.w8(32'h3c44cacb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b314295),
	.w1(32'hbaf5dfbd),
	.w2(32'hbb5a22f8),
	.w3(32'h3b49dc88),
	.w4(32'hbbe0ba37),
	.w5(32'hbad77ecf),
	.w6(32'hbc3589c3),
	.w7(32'h370b9348),
	.w8(32'h3d0a4bc7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e5351),
	.w1(32'h3c5444c4),
	.w2(32'h3b02aff9),
	.w3(32'hbb66ee6f),
	.w4(32'hbb585ae9),
	.w5(32'hbbc35ec2),
	.w6(32'h3bb8e868),
	.w7(32'h3bb24a35),
	.w8(32'hba58c34d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abda526),
	.w1(32'hbc26ec6e),
	.w2(32'h3bcd79be),
	.w3(32'h3ba3c276),
	.w4(32'hbbb689ca),
	.w5(32'h3b06a5e4),
	.w6(32'hbb86466e),
	.w7(32'hbbf8528c),
	.w8(32'hbb83ccf9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94f028),
	.w1(32'hbc08ec39),
	.w2(32'hbb86c605),
	.w3(32'h3ceb4590),
	.w4(32'h3720d96d),
	.w5(32'hb7e6a6b4),
	.w6(32'h37d25ed3),
	.w7(32'h3b646ea2),
	.w8(32'hbb0eb5bb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea863d),
	.w1(32'h3bbca425),
	.w2(32'hbb6d2ce5),
	.w3(32'hb9ffb37a),
	.w4(32'h3b7be97c),
	.w5(32'hbc27ca2e),
	.w6(32'hbbb8d4c1),
	.w7(32'hbbaede3a),
	.w8(32'hbc7c7941),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddbc6b),
	.w1(32'h3ad7095b),
	.w2(32'h39503c25),
	.w3(32'hbb8a7c3e),
	.w4(32'h3a2cc11f),
	.w5(32'hbbb90061),
	.w6(32'hbc09ac69),
	.w7(32'h3a865a09),
	.w8(32'hbc854138),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48c99c),
	.w1(32'hba2b3d01),
	.w2(32'h3c65cf27),
	.w3(32'h3b25a526),
	.w4(32'h3a4f30e0),
	.w5(32'hbb921ac2),
	.w6(32'hbb9c8d41),
	.w7(32'hbb88ecef),
	.w8(32'h3b984ce2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8af320),
	.w1(32'h3c54d49b),
	.w2(32'hbbc03c23),
	.w3(32'h3a370976),
	.w4(32'hbb8c2a36),
	.w5(32'h3aecfa86),
	.w6(32'h3b2bd219),
	.w7(32'hbb9e0249),
	.w8(32'h3bb85a9c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0df28),
	.w1(32'h3bc70c27),
	.w2(32'hba10a021),
	.w3(32'h3c153b7f),
	.w4(32'h3befe2d2),
	.w5(32'hbb5ab45d),
	.w6(32'hb996883d),
	.w7(32'hbba594ba),
	.w8(32'h3ac56169),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdb8c79),
	.w1(32'h3be78457),
	.w2(32'hba3c14dc),
	.w3(32'hbc3fec76),
	.w4(32'hbc1d3e9c),
	.w5(32'h3a91d967),
	.w6(32'hbd2df664),
	.w7(32'hba63f8dd),
	.w8(32'h3a6fe3d9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc102b9f),
	.w1(32'hbbdf17ce),
	.w2(32'h3bf1e6b6),
	.w3(32'hbc69337b),
	.w4(32'hbc6e4619),
	.w5(32'hba2a2128),
	.w6(32'hbbea19ed),
	.w7(32'hbb5d4c0e),
	.w8(32'hbaad79ce),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaffe2e),
	.w1(32'h3a89be5a),
	.w2(32'h39af62d3),
	.w3(32'h3d818cfd),
	.w4(32'hbc34f867),
	.w5(32'hbb8b7ae6),
	.w6(32'h3c342cbb),
	.w7(32'hbba8bc7a),
	.w8(32'hbc0587aa),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8493a),
	.w1(32'h3d4d8696),
	.w2(32'h3ceada17),
	.w3(32'hbbc0687e),
	.w4(32'h3afe8603),
	.w5(32'h3b2b2c11),
	.w6(32'h3b6745cf),
	.w7(32'h39ec0ab7),
	.w8(32'h3aa316d7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0587a),
	.w1(32'hbb282ba3),
	.w2(32'h3ad41f1b),
	.w3(32'hba044075),
	.w4(32'h398effb0),
	.w5(32'hbc02810e),
	.w6(32'hb8fd7d17),
	.w7(32'h3acd53cb),
	.w8(32'h3a033c9d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb274713),
	.w1(32'hbd017f92),
	.w2(32'h3bf9dbc8),
	.w3(32'hbb13bb94),
	.w4(32'hbc8fc7c1),
	.w5(32'hbaa9f342),
	.w6(32'hba159bd9),
	.w7(32'h3badd887),
	.w8(32'hbbd5fd45),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfab425),
	.w1(32'hbc000391),
	.w2(32'hbaee710a),
	.w3(32'hbc126317),
	.w4(32'hba9418a3),
	.w5(32'hbb440c4b),
	.w6(32'h3c2c3863),
	.w7(32'h3752a2e7),
	.w8(32'hbb84fc9c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1377f6),
	.w1(32'h3b19aa9a),
	.w2(32'hbbb59cad),
	.w3(32'h3aa5f97a),
	.w4(32'h3b9e0cf6),
	.w5(32'h3b5a4c87),
	.w6(32'h3a7e95fe),
	.w7(32'h3cee234e),
	.w8(32'hbbec1b00),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11bf51),
	.w1(32'hb8fd7e44),
	.w2(32'hbba26cc7),
	.w3(32'hbc137114),
	.w4(32'h3a964a65),
	.w5(32'h3b3de953),
	.w6(32'h390c6f27),
	.w7(32'hb7f642aa),
	.w8(32'hbbefae78),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cb83e),
	.w1(32'hba3c6387),
	.w2(32'hbb17e8e5),
	.w3(32'hbb389250),
	.w4(32'h3b95b5cf),
	.w5(32'hbb6d0d9a),
	.w6(32'hbac28c95),
	.w7(32'hbbfc3c63),
	.w8(32'hbb8d503e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c20c0),
	.w1(32'hbbe615e0),
	.w2(32'hba4e39fa),
	.w3(32'h3c1bc4c3),
	.w4(32'hbc548bf9),
	.w5(32'hba9365fc),
	.w6(32'hbc942179),
	.w7(32'h3a16ab5b),
	.w8(32'h3b49720b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee08ba),
	.w1(32'h3c8fbf09),
	.w2(32'hbbbb74e7),
	.w3(32'hb9916f38),
	.w4(32'h389ba8dd),
	.w5(32'h3c150872),
	.w6(32'hbbc20b3b),
	.w7(32'h3aeb96d2),
	.w8(32'h3c159dc9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6c23f),
	.w1(32'hbbedee10),
	.w2(32'h3b921003),
	.w3(32'hb98b9430),
	.w4(32'h3c8f5f7b),
	.w5(32'h3b17b99e),
	.w6(32'h3bd7d47b),
	.w7(32'hbbdcd4a2),
	.w8(32'hba9030e1),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa90242),
	.w1(32'h3cfc71f4),
	.w2(32'h3c43f704),
	.w3(32'h3a3b6c00),
	.w4(32'hbb3b575a),
	.w5(32'hbbca42ec),
	.w6(32'hbb8f11a7),
	.w7(32'hbd094a25),
	.w8(32'h3b8156de),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc794c73),
	.w1(32'h39e56a3a),
	.w2(32'hba9ea064),
	.w3(32'h3b7a7423),
	.w4(32'h3b1a44bd),
	.w5(32'h3c0f3dc4),
	.w6(32'h3c508181),
	.w7(32'h3c12198c),
	.w8(32'hbc28117b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba277d1d),
	.w1(32'hbb10f21d),
	.w2(32'hbab4c48b),
	.w3(32'h3af72330),
	.w4(32'h3b392282),
	.w5(32'hba9410b9),
	.w6(32'hbb8c7331),
	.w7(32'hbbdd784a),
	.w8(32'h3b03d14d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd97b5f8),
	.w1(32'hbcc0105b),
	.w2(32'hbb98e724),
	.w3(32'h3b8b59d7),
	.w4(32'hbbd88a70),
	.w5(32'hbb4da396),
	.w6(32'hbb8670fc),
	.w7(32'h3b1351b5),
	.w8(32'h3b8bddfc),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f662b),
	.w1(32'hba4e53fc),
	.w2(32'hbc4be313),
	.w3(32'hbaec6ea2),
	.w4(32'hb9d78f42),
	.w5(32'hbaade8a1),
	.w6(32'h3c211bae),
	.w7(32'h3bf88177),
	.w8(32'h3b277da2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9389a9),
	.w1(32'h3b8e8b28),
	.w2(32'h3b80ebf7),
	.w3(32'hbac1a147),
	.w4(32'hbb3b1ba0),
	.w5(32'hba05bb01),
	.w6(32'h3ae03642),
	.w7(32'h3b174346),
	.w8(32'hba26bccb),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a67e2),
	.w1(32'hbc458715),
	.w2(32'h3a59e546),
	.w3(32'hbb1df06a),
	.w4(32'h3bb09bbb),
	.w5(32'hbabdc261),
	.w6(32'h3bfc1671),
	.w7(32'h3b81ca95),
	.w8(32'h39e30471),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be871f6),
	.w1(32'hbb20bdb2),
	.w2(32'h3b8ef383),
	.w3(32'hbc77d41e),
	.w4(32'h3b9147ac),
	.w5(32'hbcd7e2e7),
	.w6(32'h3bf753b5),
	.w7(32'h3b99c3ce),
	.w8(32'hbb6a1232),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66a7eb),
	.w1(32'hbb622977),
	.w2(32'h3a61c854),
	.w3(32'h3ae81aa1),
	.w4(32'h3b824057),
	.w5(32'hb89872dc),
	.w6(32'hbbc4c6fd),
	.w7(32'h3a8bebbd),
	.w8(32'h3bf1be43),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c166d5d),
	.w1(32'hbbe787e5),
	.w2(32'hb8c678c0),
	.w3(32'h3b447846),
	.w4(32'hbad29b07),
	.w5(32'hbd6631b0),
	.w6(32'h3b93e9ed),
	.w7(32'hbcb715c4),
	.w8(32'hb6da39ff),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00eb3f),
	.w1(32'h3c0f6983),
	.w2(32'h3a211698),
	.w3(32'h3a9a4e6f),
	.w4(32'hbb30c812),
	.w5(32'h3b880d5f),
	.w6(32'hbbbe5b09),
	.w7(32'hba90768a),
	.w8(32'hbb83a1df),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade9984),
	.w1(32'h3a46d59e),
	.w2(32'h3b378588),
	.w3(32'h3c4d3992),
	.w4(32'hbc37548b),
	.w5(32'h3ad33834),
	.w6(32'hbc63e366),
	.w7(32'h3b0a8fc4),
	.w8(32'h3b33a861),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53fae7),
	.w1(32'h3b8463d5),
	.w2(32'h3c0a81f6),
	.w3(32'h3b35322e),
	.w4(32'h3bd228df),
	.w5(32'hbbc39680),
	.w6(32'h3aecf196),
	.w7(32'hbc80fb27),
	.w8(32'hbb685e07),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c0c41),
	.w1(32'hbbad0496),
	.w2(32'hbb7e7b23),
	.w3(32'hbbc01ecd),
	.w4(32'hbc7a3cc2),
	.w5(32'hbc383834),
	.w6(32'hbb4b81d5),
	.w7(32'h3aace125),
	.w8(32'h3bab9ba6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd6ff75),
	.w1(32'h3ba3e295),
	.w2(32'hbbf3e768),
	.w3(32'hbac88832),
	.w4(32'hb9a9eb29),
	.w5(32'hbab9132a),
	.w6(32'h3885668c),
	.w7(32'h3965ea4d),
	.w8(32'hb74fd83e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b87c2),
	.w1(32'hbc61d024),
	.w2(32'hbd31c963),
	.w3(32'hbb4445ce),
	.w4(32'hbcc4eaf5),
	.w5(32'hbc4c5b01),
	.w6(32'h3b8c2567),
	.w7(32'hbb96b155),
	.w8(32'hb9cc23be),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaced9),
	.w1(32'hbb82edf6),
	.w2(32'h3aea9aac),
	.w3(32'hbb68d4e8),
	.w4(32'hbc1924cc),
	.w5(32'h3c6e3e90),
	.w6(32'hba51ee41),
	.w7(32'hbb45d84c),
	.w8(32'h3c85fb62),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15483b),
	.w1(32'h3a829014),
	.w2(32'hba8cb955),
	.w3(32'h3c88dc23),
	.w4(32'h3b8d3d55),
	.w5(32'h3a8140f4),
	.w6(32'hbaceb9d9),
	.w7(32'h3d2fea7b),
	.w8(32'hbc46b4cf),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba52efb),
	.w1(32'hbbefc695),
	.w2(32'hb9a12bca),
	.w3(32'hbc52357c),
	.w4(32'h3c0d2d0c),
	.w5(32'h3cdcbc30),
	.w6(32'h3bb4be52),
	.w7(32'h3b4d8b37),
	.w8(32'h3b6a037d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9394fd),
	.w1(32'hbafe4bef),
	.w2(32'h3a20bff7),
	.w3(32'hbc472d9c),
	.w4(32'h3ba14618),
	.w5(32'hba2c2a31),
	.w6(32'hbadbd710),
	.w7(32'hbb4c5acd),
	.w8(32'h3b2d1512),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91adca),
	.w1(32'hba045da6),
	.w2(32'hba50d86e),
	.w3(32'hbbd32557),
	.w4(32'hbb1b7ab3),
	.w5(32'h3cfb1295),
	.w6(32'h3a8b6886),
	.w7(32'h3bb11fce),
	.w8(32'hbc54097c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82dd25),
	.w1(32'hbb6874c7),
	.w2(32'hbb68c7d0),
	.w3(32'h3b71affa),
	.w4(32'hbc594a9b),
	.w5(32'h3bde2a5d),
	.w6(32'hbb69a199),
	.w7(32'hbb0af90b),
	.w8(32'h3bb28a1a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac85a0c),
	.w1(32'h3b7afef5),
	.w2(32'hba45679e),
	.w3(32'hbb933290),
	.w4(32'h3bc4fc98),
	.w5(32'hbac62757),
	.w6(32'h3bcff758),
	.w7(32'hbd187c61),
	.w8(32'hbc2897b3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3593d),
	.w1(32'h3b684f20),
	.w2(32'hbb60a378),
	.w3(32'hbc5e9585),
	.w4(32'hbbe35a46),
	.w5(32'h3c901538),
	.w6(32'hbc186a7b),
	.w7(32'hbbf28608),
	.w8(32'hbb033aee),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17aa5e),
	.w1(32'h3bdbfd1f),
	.w2(32'h3b3f3385),
	.w3(32'hbbc5f410),
	.w4(32'h3aa58d81),
	.w5(32'h3aea400f),
	.w6(32'hbb84de54),
	.w7(32'hbbb62ee6),
	.w8(32'hb9ea2d28),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64e5a0),
	.w1(32'h3a263280),
	.w2(32'h3a8d5217),
	.w3(32'hbb84d983),
	.w4(32'hbb6a698a),
	.w5(32'h39ff8f97),
	.w6(32'h3af65cef),
	.w7(32'h3b82ea6a),
	.w8(32'h3d506a31),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaecb86),
	.w1(32'hba462afd),
	.w2(32'h3b5cea71),
	.w3(32'hbbb4da39),
	.w4(32'h3b546e04),
	.w5(32'hbd37ff87),
	.w6(32'hbb667cc1),
	.w7(32'h3ae1e891),
	.w8(32'h3c05286c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57b326),
	.w1(32'h3b876a2a),
	.w2(32'h3aa349bc),
	.w3(32'hbb609ea9),
	.w4(32'h3b1dd5c5),
	.w5(32'h3a2f79cb),
	.w6(32'h37385746),
	.w7(32'hbd3cfec6),
	.w8(32'h3bcba780),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb861e36),
	.w1(32'h398d015e),
	.w2(32'h3b704c58),
	.w3(32'hbb4bffbb),
	.w4(32'h3b7932fd),
	.w5(32'h3b0998ec),
	.w6(32'h3b1966e7),
	.w7(32'h3b1a1081),
	.w8(32'hbb385f61),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae8e0f),
	.w1(32'h3bad1eb2),
	.w2(32'hbabd9684),
	.w3(32'h3a8bf060),
	.w4(32'h3bc6159e),
	.w5(32'h3ad1f8cc),
	.w6(32'h3b1db1b6),
	.w7(32'h3bbfb7fb),
	.w8(32'h3a609758),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3aa4f5),
	.w1(32'h3aa6fa75),
	.w2(32'hbba2aa3a),
	.w3(32'hbb15f161),
	.w4(32'h3b98b645),
	.w5(32'hbb10fb11),
	.w6(32'h3b2e9331),
	.w7(32'h3bc9cefd),
	.w8(32'hbb97f4ee),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74d9c8),
	.w1(32'h388c456c),
	.w2(32'hbabe5342),
	.w3(32'h39a71130),
	.w4(32'hbc9a717f),
	.w5(32'hbc804931),
	.w6(32'hb934300c),
	.w7(32'h3abc3183),
	.w8(32'hba602214),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b1c4c),
	.w1(32'h3b63ba50),
	.w2(32'h3ba41b0b),
	.w3(32'h3b32d6f8),
	.w4(32'h3b56683c),
	.w5(32'hbb2018e6),
	.w6(32'h3b0687aa),
	.w7(32'h3b9585a9),
	.w8(32'h3b11f1dd),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25ed0f),
	.w1(32'h3b99160f),
	.w2(32'hbbb789f6),
	.w3(32'hba148ea4),
	.w4(32'h3cb23c3c),
	.w5(32'hbbcbbb85),
	.w6(32'hba79cae7),
	.w7(32'h3b839c4a),
	.w8(32'h3bfdd7ad),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f27ae),
	.w1(32'h3ab2f2c6),
	.w2(32'h3bd85b0c),
	.w3(32'h3bb3cbdb),
	.w4(32'hba971af7),
	.w5(32'h3b515750),
	.w6(32'hbbc88175),
	.w7(32'hbc7c4f87),
	.w8(32'h3c86134f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd135e),
	.w1(32'h3b53aec4),
	.w2(32'h3b0575bc),
	.w3(32'hb9c16185),
	.w4(32'hb4fdfbd0),
	.w5(32'h3a018749),
	.w6(32'hbba4fea7),
	.w7(32'hbbd2fd0e),
	.w8(32'hb94b4df7),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39d912),
	.w1(32'h3946308a),
	.w2(32'h3b657da6),
	.w3(32'hbb8e1024),
	.w4(32'h3bd6d312),
	.w5(32'h3bd330e7),
	.w6(32'hba8d91b2),
	.w7(32'hb8f116df),
	.w8(32'hbaddedf5),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba49f5),
	.w1(32'hbd833894),
	.w2(32'h3b4f9b50),
	.w3(32'hba4683a7),
	.w4(32'hbb0860cd),
	.w5(32'h3a0fc53e),
	.w6(32'h3ac78c43),
	.w7(32'hbd341016),
	.w8(32'h3afba302),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba61181),
	.w1(32'h3b1cffc4),
	.w2(32'h3b932a80),
	.w3(32'hba09e4f1),
	.w4(32'h3b3b0be1),
	.w5(32'h3a44345b),
	.w6(32'hbc205313),
	.w7(32'h3ba823f0),
	.w8(32'h3987c140),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f4afe),
	.w1(32'h3af92f17),
	.w2(32'h3b8741e6),
	.w3(32'h3bf1818d),
	.w4(32'h3b1960ab),
	.w5(32'h39bb0e63),
	.w6(32'h3a9e7a4b),
	.w7(32'h3d3a96d8),
	.w8(32'hbbfe8304),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6fc9bd),
	.w1(32'h3b535af4),
	.w2(32'hbb155b3c),
	.w3(32'h3d6d2f95),
	.w4(32'h3b38862b),
	.w5(32'h3a30bb6c),
	.w6(32'h3af94b7f),
	.w7(32'h3b1c03cc),
	.w8(32'hba4e721d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a418d),
	.w1(32'h3a473668),
	.w2(32'hbbefaf12),
	.w3(32'h3b181060),
	.w4(32'hbb667a67),
	.w5(32'hbb6b5fec),
	.w6(32'hbad6d6e9),
	.w7(32'hbba5d03f),
	.w8(32'hbb33ea8d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ef22e),
	.w1(32'h3b6ed52c),
	.w2(32'hbac5182a),
	.w3(32'hbb1cec8d),
	.w4(32'h3d013a38),
	.w5(32'hbac4e68d),
	.w6(32'hb9e2c97c),
	.w7(32'h3ade6787),
	.w8(32'h3d453227),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7583d94),
	.w1(32'hbc7fb3db),
	.w2(32'hbb0da139),
	.w3(32'hba03dac7),
	.w4(32'h3b1312d5),
	.w5(32'h3b2693cd),
	.w6(32'h3b0a32bf),
	.w7(32'hbb627eb7),
	.w8(32'hbd5d0b6e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab47d0f),
	.w1(32'hb8008ee3),
	.w2(32'h39f906ad),
	.w3(32'hbc8b59da),
	.w4(32'hbac1f753),
	.w5(32'hbaf31636),
	.w6(32'hbcf8791e),
	.w7(32'h3c1cdf06),
	.w8(32'hbd033e3b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41c260),
	.w1(32'h3bfb0bac),
	.w2(32'h3b2c5348),
	.w3(32'h3bcc451e),
	.w4(32'h3b5916f0),
	.w5(32'h3abb3fb6),
	.w6(32'hbb3e2310),
	.w7(32'hbd3e2df1),
	.w8(32'hba8791ad),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc4b13),
	.w1(32'h3b39a037),
	.w2(32'hb9bf5035),
	.w3(32'hbb4996dd),
	.w4(32'hb9aa8cc7),
	.w5(32'hbc4f4c2c),
	.w6(32'h3bd03bd4),
	.w7(32'h3b9318c1),
	.w8(32'hba0b223c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b510aee),
	.w1(32'h3b3d296c),
	.w2(32'hba918692),
	.w3(32'h3abb4ca3),
	.w4(32'h3bc5719a),
	.w5(32'hbb3a97fe),
	.w6(32'h3c268995),
	.w7(32'h3c8452d4),
	.w8(32'h3b474dcd),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bc905),
	.w1(32'hb91ddb1d),
	.w2(32'h3b668b63),
	.w3(32'h3a066f0d),
	.w4(32'h3a032cef),
	.w5(32'hb9cd3e1a),
	.w6(32'h3b080be9),
	.w7(32'hba6884ff),
	.w8(32'hb8743e6b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19f23e),
	.w1(32'hbc8b77aa),
	.w2(32'hba898569),
	.w3(32'h3b0cfdea),
	.w4(32'h3aedf72b),
	.w5(32'hbb672e24),
	.w6(32'hbab774c3),
	.w7(32'hbaeadd8f),
	.w8(32'h3ab7bd34),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09f4a9),
	.w1(32'hba1eed8a),
	.w2(32'h3ae2393f),
	.w3(32'hbb1c118c),
	.w4(32'hb7463cda),
	.w5(32'hb8ac8f55),
	.w6(32'hbb2f5d11),
	.w7(32'hb9781d53),
	.w8(32'hbb5ad721),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c163ef4),
	.w1(32'h3ae0332f),
	.w2(32'hbbbcf6f2),
	.w3(32'h3af5f697),
	.w4(32'h3b57485c),
	.w5(32'h3c4157af),
	.w6(32'h3a977a7a),
	.w7(32'h3badcb68),
	.w8(32'h3b6cba1e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c498cb5),
	.w1(32'h3a673216),
	.w2(32'hbbcb0eed),
	.w3(32'h3b69b7f5),
	.w4(32'hba1dbf71),
	.w5(32'hb929545d),
	.w6(32'h3c22c89c),
	.w7(32'h3b896c16),
	.w8(32'h3b3965b9),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e5ce5),
	.w1(32'h3b7ecfbe),
	.w2(32'h3a63b130),
	.w3(32'h3b186974),
	.w4(32'hbb3a891d),
	.w5(32'h3ad11f9c),
	.w6(32'h3b4e0f94),
	.w7(32'h3b7b429d),
	.w8(32'hbb8e4f22),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23e624),
	.w1(32'h3c87ff1c),
	.w2(32'hbb1cdf54),
	.w3(32'hbc1e925a),
	.w4(32'hbb3f4ff6),
	.w5(32'h37602898),
	.w6(32'h3b860616),
	.w7(32'h3abc7674),
	.w8(32'hbb237bd5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule