module layer_10_featuremap_159(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37857c8d),
	.w1(32'hbb6192d1),
	.w2(32'hbbc04ae6),
	.w3(32'hba2b5c35),
	.w4(32'h3b43a433),
	.w5(32'h3c81f53d),
	.w6(32'hbb205ada),
	.w7(32'h3c280d18),
	.w8(32'h3c4095b0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ba311),
	.w1(32'h3a8ee14c),
	.w2(32'h3adced61),
	.w3(32'hb8f2f1ad),
	.w4(32'hba4de6c2),
	.w5(32'hbaf545cb),
	.w6(32'hbb0d7f6b),
	.w7(32'hbad0d845),
	.w8(32'hba5dae1f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a243f19),
	.w1(32'hbaf36884),
	.w2(32'hbb124be0),
	.w3(32'hba4b965b),
	.w4(32'hbb3bdf45),
	.w5(32'hbb1a5c53),
	.w6(32'h3a2a9ba1),
	.w7(32'h3b69f1e8),
	.w8(32'h390f0611),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2acbe6),
	.w1(32'hbb8dd7b7),
	.w2(32'h3cd2a10b),
	.w3(32'hbb412ac0),
	.w4(32'h3c11175a),
	.w5(32'hbac15d2b),
	.w6(32'hb9624b0e),
	.w7(32'hbc2d942d),
	.w8(32'hbb6803e1),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16354d),
	.w1(32'h3a4cc899),
	.w2(32'h3bfce562),
	.w3(32'h3b5e3fca),
	.w4(32'h390cbd0f),
	.w5(32'hbb9b5049),
	.w6(32'h3b5477a0),
	.w7(32'h3a917b89),
	.w8(32'hbc27a97a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ba435),
	.w1(32'h3a5a818a),
	.w2(32'h3a605391),
	.w3(32'h3b2c6798),
	.w4(32'hb8c00ae9),
	.w5(32'h399eaebc),
	.w6(32'h3b1f23e8),
	.w7(32'h3bd97bed),
	.w8(32'h3b5fdae2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc2cb7),
	.w1(32'h3b17d5ba),
	.w2(32'hbacddbf9),
	.w3(32'h3bb64e3c),
	.w4(32'hbb0ebeed),
	.w5(32'hbbcf7a3f),
	.w6(32'h3becdf1c),
	.w7(32'h3b34d402),
	.w8(32'hbc226120),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23be95),
	.w1(32'hbbe2240e),
	.w2(32'hbb9b72b8),
	.w3(32'hbbcc78f8),
	.w4(32'hbc398d38),
	.w5(32'hbb835521),
	.w6(32'hba05a12d),
	.w7(32'hbb6267b5),
	.w8(32'hba19c2e7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d19c7),
	.w1(32'hba7c614c),
	.w2(32'hbb9c4145),
	.w3(32'h3aed7739),
	.w4(32'h3a93b497),
	.w5(32'hbac19597),
	.w6(32'h3b178e0b),
	.w7(32'h39d389dc),
	.w8(32'hba11ab2a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57a2cb),
	.w1(32'h3b664be2),
	.w2(32'h3abcfcd5),
	.w3(32'h3ab50e72),
	.w4(32'h3ae3824a),
	.w5(32'hbb3e1446),
	.w6(32'h3b298e9d),
	.w7(32'hbbbad5dc),
	.w8(32'hbbbf51b1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90e312),
	.w1(32'hbc8a2771),
	.w2(32'hbbd8aa07),
	.w3(32'h3a987242),
	.w4(32'hba34cfd9),
	.w5(32'h3ad4d2c6),
	.w6(32'hbb4039c2),
	.w7(32'hbaa54a65),
	.w8(32'hba738d52),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b0377),
	.w1(32'h3c1f249a),
	.w2(32'h3d115699),
	.w3(32'h3c236f75),
	.w4(32'h3c28760c),
	.w5(32'hbc6860d4),
	.w6(32'h3c76a01f),
	.w7(32'hb8aee743),
	.w8(32'h3b90d23d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c191a60),
	.w1(32'hbb5f8a93),
	.w2(32'hbbc8a425),
	.w3(32'h3bb8b401),
	.w4(32'hb9d290da),
	.w5(32'hbab60da7),
	.w6(32'h3b43861f),
	.w7(32'hbb7b515e),
	.w8(32'hbbd9ce65),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b28a4c),
	.w1(32'h39d8a9ab),
	.w2(32'hbb954afb),
	.w3(32'h3abc9376),
	.w4(32'h3ab7bd2b),
	.w5(32'h3aa01553),
	.w6(32'h3bc23fc5),
	.w7(32'hbb4ab368),
	.w8(32'h3b6efe4e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c6738),
	.w1(32'h3b52660f),
	.w2(32'h3d5cdb87),
	.w3(32'h3bb5fc22),
	.w4(32'h3bf4b238),
	.w5(32'hbcbef244),
	.w6(32'h3c0b9166),
	.w7(32'hbc1e3ad5),
	.w8(32'hbbbd79e2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b9aa2),
	.w1(32'hbad905c1),
	.w2(32'hbb82cf23),
	.w3(32'hbacfe645),
	.w4(32'hbae9f08e),
	.w5(32'hbb3c3422),
	.w6(32'hbb782a19),
	.w7(32'hbbbe33a5),
	.w8(32'hbb90b2e4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40de2e),
	.w1(32'h3b14a47c),
	.w2(32'hba984aa3),
	.w3(32'hbb0d1d43),
	.w4(32'h3b5ed4de),
	.w5(32'h3bdd3bed),
	.w6(32'h3ba9f0f4),
	.w7(32'h3bf3a4a0),
	.w8(32'hbb2b7958),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee1f4d),
	.w1(32'hbaa55601),
	.w2(32'h3ac4c4b2),
	.w3(32'h3b1ac4fc),
	.w4(32'hbc05f31b),
	.w5(32'hbb172c3c),
	.w6(32'h3a96d04d),
	.w7(32'hbc0bd83a),
	.w8(32'hbc0f4578),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38660a),
	.w1(32'h37937852),
	.w2(32'h3a101648),
	.w3(32'hba8c7fdd),
	.w4(32'hbb073211),
	.w5(32'hbad298ed),
	.w6(32'h3b9caf16),
	.w7(32'hbace5b9f),
	.w8(32'hbb93e66a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7337552),
	.w1(32'hba9d63ad),
	.w2(32'hbb4a5120),
	.w3(32'h3969f043),
	.w4(32'h39c934cc),
	.w5(32'hba08df93),
	.w6(32'hba0d2d64),
	.w7(32'hba41e67a),
	.w8(32'hba143178),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb699e41),
	.w1(32'h3a062341),
	.w2(32'hb949fd99),
	.w3(32'hba4a131e),
	.w4(32'h3a0d9251),
	.w5(32'hbae4eabd),
	.w6(32'h3b75ef23),
	.w7(32'h3ba176ac),
	.w8(32'h3b3bdbf1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39372890),
	.w1(32'h3939d51d),
	.w2(32'h3b94e577),
	.w3(32'h3aa1c1b7),
	.w4(32'hbc3a9119),
	.w5(32'h3b141c84),
	.w6(32'hbc1721cc),
	.w7(32'h3b91be31),
	.w8(32'hbc3acd82),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bf7b4),
	.w1(32'hbbb1b6c5),
	.w2(32'hbc3b910a),
	.w3(32'hbca7f8c2),
	.w4(32'hbbb5f557),
	.w5(32'hbc5df050),
	.w6(32'hbbbbb242),
	.w7(32'hbc7f66f8),
	.w8(32'hbc9be93b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd57bab),
	.w1(32'hbaece13a),
	.w2(32'hbb3696ba),
	.w3(32'h3a0fa202),
	.w4(32'h3a1b0ec2),
	.w5(32'hbb0a5d01),
	.w6(32'h3b774d55),
	.w7(32'h3b0470ff),
	.w8(32'hbb13ad43),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace8db0),
	.w1(32'hb9ea63dc),
	.w2(32'h3b95ca89),
	.w3(32'h3a9d13a6),
	.w4(32'h3b8c8957),
	.w5(32'hb7a15c98),
	.w6(32'hbc0fb974),
	.w7(32'hbbf806b9),
	.w8(32'hbb053c9e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b392a2f),
	.w1(32'hbc0ba1e4),
	.w2(32'hbb420056),
	.w3(32'h3b47eaf3),
	.w4(32'hbb78d01b),
	.w5(32'hbc2a0ff0),
	.w6(32'hbb113112),
	.w7(32'hbb9c4e6a),
	.w8(32'hbb339a6e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc438f21),
	.w1(32'hb8d9cff3),
	.w2(32'hba5a3fad),
	.w3(32'h3a8ff97f),
	.w4(32'h396c7ff4),
	.w5(32'h39d8686c),
	.w6(32'h393ae2bf),
	.w7(32'h3ad24f56),
	.w8(32'h3afd80f8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc42af),
	.w1(32'hbbcb5e05),
	.w2(32'h3af62773),
	.w3(32'h3a62c7c0),
	.w4(32'h3b3f2648),
	.w5(32'hba0f0d55),
	.w6(32'hbbb2a4fa),
	.w7(32'hbc21067f),
	.w8(32'h3b69a0ac),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad4e3f),
	.w1(32'h3a277a15),
	.w2(32'hbb195f2f),
	.w3(32'h36e2a61d),
	.w4(32'h3b38d781),
	.w5(32'h3a4ed124),
	.w6(32'h3b1fde43),
	.w7(32'h3ada7a21),
	.w8(32'h3b048172),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c19b79),
	.w1(32'h3b33d9de),
	.w2(32'h3a9a9d94),
	.w3(32'h3b73d324),
	.w4(32'h3b9fa5f7),
	.w5(32'hba265582),
	.w6(32'h3b22c5cd),
	.w7(32'h3a2e6410),
	.w8(32'hbb704625),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f48da),
	.w1(32'hba3fd06f),
	.w2(32'hbb1fa437),
	.w3(32'h3a8a63be),
	.w4(32'h3a1b5b65),
	.w5(32'hb89529bb),
	.w6(32'h3a367c59),
	.w7(32'h3b3523a7),
	.w8(32'h3a528cba),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac249a2),
	.w1(32'hbac8c553),
	.w2(32'hbb385d0e),
	.w3(32'h3a3cc2de),
	.w4(32'hba48684c),
	.w5(32'hbadc368f),
	.w6(32'h37bab209),
	.w7(32'h3aa4ac0a),
	.w8(32'h39809ab3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395143f9),
	.w1(32'h3a5cafb0),
	.w2(32'hbbdc7898),
	.w3(32'h3b0346ef),
	.w4(32'h3a4435fe),
	.w5(32'h3a8ba509),
	.w6(32'h3b77f514),
	.w7(32'hbb22c58c),
	.w8(32'hbbf05348),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf91c13),
	.w1(32'hbb686543),
	.w2(32'hbbb284ab),
	.w3(32'h3a42d144),
	.w4(32'h3835b454),
	.w5(32'hbb93ce01),
	.w6(32'hbb9ecbaa),
	.w7(32'hbb3c3f6d),
	.w8(32'hbb4943b0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb940451),
	.w1(32'h3ab60171),
	.w2(32'h3b40448f),
	.w3(32'hbbf23ebc),
	.w4(32'h3b30f4f6),
	.w5(32'h3a5dc48e),
	.w6(32'h3a66b75a),
	.w7(32'h3a2515f6),
	.w8(32'h3b905dea),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd006c),
	.w1(32'hbbabc010),
	.w2(32'hbb347f9e),
	.w3(32'h3ba016cd),
	.w4(32'hbb0a2898),
	.w5(32'hbbc079dd),
	.w6(32'hb9b84276),
	.w7(32'hbb08bd44),
	.w8(32'hbb9f81d4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c76e8),
	.w1(32'h3b20a2c9),
	.w2(32'h3be0ceba),
	.w3(32'h3ab0c1b9),
	.w4(32'h3b97787e),
	.w5(32'hbb840539),
	.w6(32'h3a4e7b8e),
	.w7(32'hbb6bf2d7),
	.w8(32'hbc7ec336),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a88c0),
	.w1(32'h3bf7a43d),
	.w2(32'h3b1a66ef),
	.w3(32'h3b1f93ef),
	.w4(32'h3c187a86),
	.w5(32'h3b05f657),
	.w6(32'hbb6cc23b),
	.w7(32'h3be72718),
	.w8(32'h3a286d4b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa9944),
	.w1(32'h3b66a0c5),
	.w2(32'hbb49e676),
	.w3(32'h3b42ca5a),
	.w4(32'h3bd9eac4),
	.w5(32'hb9ead246),
	.w6(32'h3adfb2c3),
	.w7(32'h3afbd3b1),
	.w8(32'hba0cf6b5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0aa5b),
	.w1(32'h3a8c116e),
	.w2(32'h3b8421c9),
	.w3(32'hb9988f63),
	.w4(32'hb7b60874),
	.w5(32'hba557ec8),
	.w6(32'hbab66b86),
	.w7(32'hba9ba277),
	.w8(32'hbb873cd8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebeda4),
	.w1(32'hba691e5f),
	.w2(32'hba9e48ad),
	.w3(32'hb9703f3c),
	.w4(32'h3a8028c5),
	.w5(32'h3ada4048),
	.w6(32'hb9ef2941),
	.w7(32'h3a999ecf),
	.w8(32'hbaaed785),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97c5f7),
	.w1(32'hbc1e1777),
	.w2(32'h3b749c31),
	.w3(32'h3a14b342),
	.w4(32'hba704916),
	.w5(32'hbbd9c0aa),
	.w6(32'hbb94266a),
	.w7(32'hbc09bc48),
	.w8(32'hbb5b794c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabf3e6),
	.w1(32'hba142b6a),
	.w2(32'hbb24cc75),
	.w3(32'h3a81c915),
	.w4(32'h3ac641b3),
	.w5(32'hba407fff),
	.w6(32'hbad4c9cd),
	.w7(32'h39d1b177),
	.w8(32'hb919922b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f8ca),
	.w1(32'h3b8306bc),
	.w2(32'h3aa31499),
	.w3(32'hba9121ef),
	.w4(32'hbac87e9b),
	.w5(32'hb935b330),
	.w6(32'hb96938f2),
	.w7(32'hbc1039d5),
	.w8(32'hbbec146f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8da7c3),
	.w1(32'hbb3cdab3),
	.w2(32'hbc4b4e82),
	.w3(32'h3b876d31),
	.w4(32'h3bdcf501),
	.w5(32'h3c062c84),
	.w6(32'hbab5d75b),
	.w7(32'hbb9c42f8),
	.w8(32'hbbc41d6c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9390d0),
	.w1(32'hbb487c95),
	.w2(32'hbbd6660b),
	.w3(32'h3ba6cf7c),
	.w4(32'h3ad4fa58),
	.w5(32'h3c0c4d1b),
	.w6(32'hbbad1c1e),
	.w7(32'hbb507738),
	.w8(32'hbc2196e4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf898ca),
	.w1(32'h3bfe9623),
	.w2(32'h3d639dd5),
	.w3(32'h3af2756a),
	.w4(32'h3c0a9bd7),
	.w5(32'hbc732bcd),
	.w6(32'h3b04e88b),
	.w7(32'hbc465741),
	.w8(32'hbb9cc1bd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bb03b),
	.w1(32'hbb67b941),
	.w2(32'hbc1af22c),
	.w3(32'hba1d846a),
	.w4(32'hbbbd72cc),
	.w5(32'hbbeb1f07),
	.w6(32'h3b312880),
	.w7(32'hbc142da2),
	.w8(32'hbc478635),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbceccc0),
	.w1(32'hbaa5effb),
	.w2(32'hbb0d7aad),
	.w3(32'hbab397da),
	.w4(32'hba22d9cd),
	.w5(32'h39f17c6a),
	.w6(32'hba776412),
	.w7(32'h39452184),
	.w8(32'h3af10d94),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad29af9),
	.w1(32'hba21ad32),
	.w2(32'hbade6c9f),
	.w3(32'hb84b7811),
	.w4(32'hba38af6d),
	.w5(32'h399f0b49),
	.w6(32'h3acc5452),
	.w7(32'h3a9b6f81),
	.w8(32'h3a92f930),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f8ae5),
	.w1(32'h3b24af19),
	.w2(32'hbb9dc867),
	.w3(32'h3a9bb3c6),
	.w4(32'hba81fee6),
	.w5(32'hbb9c1bc3),
	.w6(32'h3b0f483d),
	.w7(32'hbb9e9d94),
	.w8(32'hba86eb8b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60fd03),
	.w1(32'hb96a2ed2),
	.w2(32'h3c781488),
	.w3(32'hbb08da5d),
	.w4(32'hbae10a39),
	.w5(32'hbc706a43),
	.w6(32'hbbc91533),
	.w7(32'hbbedae0f),
	.w8(32'h3c307f76),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a3437),
	.w1(32'hbb4713c3),
	.w2(32'hbba5393c),
	.w3(32'hbbb1cb43),
	.w4(32'hbb0a1944),
	.w5(32'hbb7a247f),
	.w6(32'hba2060e1),
	.w7(32'hbaf437f9),
	.w8(32'hbaaa034e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadcb7b),
	.w1(32'hba1fb506),
	.w2(32'hbb97f645),
	.w3(32'hbb2b022d),
	.w4(32'hbb7b00e4),
	.w5(32'hbb51a452),
	.w6(32'h3af5b00a),
	.w7(32'hba617e94),
	.w8(32'hbc53a24c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb888a3f),
	.w1(32'h3a44aaf9),
	.w2(32'hb9e53c73),
	.w3(32'h3b0e47e1),
	.w4(32'h391f077d),
	.w5(32'h3a064af0),
	.w6(32'h3b4e07c1),
	.w7(32'h3aa51111),
	.w8(32'h3a665ae5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab909a6),
	.w1(32'hbb07db9f),
	.w2(32'hba76da05),
	.w3(32'h3b90c832),
	.w4(32'h3a7a8515),
	.w5(32'hb95a08bb),
	.w6(32'hba84938f),
	.w7(32'h3abd8a2f),
	.w8(32'hbaeca55b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f78b3),
	.w1(32'h3ae32506),
	.w2(32'hb9809ca1),
	.w3(32'h3ac1446e),
	.w4(32'h3b8c7834),
	.w5(32'h3bcef120),
	.w6(32'h3b736a45),
	.w7(32'h3b0ca59d),
	.w8(32'h3b4a6377),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cfeb5),
	.w1(32'hb8ee8e99),
	.w2(32'hbb007ff2),
	.w3(32'h3b9a3c70),
	.w4(32'hbb0f9faf),
	.w5(32'hbae169cd),
	.w6(32'h3b87475d),
	.w7(32'h3b27c120),
	.w8(32'hbb9075bf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee0e1f),
	.w1(32'h3a1fda1b),
	.w2(32'h3a9d83c8),
	.w3(32'h3b942f4b),
	.w4(32'hbaf448fc),
	.w5(32'hbb34fdb1),
	.w6(32'h3aa4dd30),
	.w7(32'h3b3fd49a),
	.w8(32'h3b0818e6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15045f),
	.w1(32'hba83bb54),
	.w2(32'hbaea42fe),
	.w3(32'hbb8152a4),
	.w4(32'h38c75d04),
	.w5(32'hba3df1fc),
	.w6(32'h3b02ffe5),
	.w7(32'h3b2541a2),
	.w8(32'h3a468d6c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3af352),
	.w1(32'hb9063e29),
	.w2(32'h3ae68458),
	.w3(32'hba63d6b0),
	.w4(32'hbb578c73),
	.w5(32'hbb16c95f),
	.w6(32'hb8895615),
	.w7(32'hba9bcf43),
	.w8(32'h3a524e44),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfc066),
	.w1(32'hbbe08c7f),
	.w2(32'hbc02c94c),
	.w3(32'hbbc10ab0),
	.w4(32'h36c3b0f8),
	.w5(32'h3bd3b2a5),
	.w6(32'hbbf52371),
	.w7(32'hbb87a266),
	.w8(32'hbb482f38),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f7584),
	.w1(32'h3ae4499f),
	.w2(32'hbbdf1679),
	.w3(32'h3b1b7b3c),
	.w4(32'h3a950d04),
	.w5(32'h3b2e103b),
	.w6(32'h3b18cbb3),
	.w7(32'h3b0e2d4c),
	.w8(32'h3a83aab0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04c2d1),
	.w1(32'h3b4ef8ee),
	.w2(32'h3b7bade1),
	.w3(32'hbb4a045f),
	.w4(32'h3a7b6e54),
	.w5(32'h3a7cc831),
	.w6(32'hb9fd3880),
	.w7(32'hbafc7023),
	.w8(32'hba592dca),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e61c0),
	.w1(32'h38c83843),
	.w2(32'hb9bf3876),
	.w3(32'h3ab55552),
	.w4(32'hb94599ba),
	.w5(32'hbacbe2ce),
	.w6(32'hba248162),
	.w7(32'hbab5e036),
	.w8(32'h38b19365),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acce311),
	.w1(32'hbb03f4a4),
	.w2(32'hbc157d88),
	.w3(32'h3a0529af),
	.w4(32'h39942de2),
	.w5(32'h3bda7578),
	.w6(32'hb84d5784),
	.w7(32'h3b402c12),
	.w8(32'hbbb9482d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf18e06),
	.w1(32'hba996dba),
	.w2(32'hb9036e3b),
	.w3(32'h393ff316),
	.w4(32'h3b001aaa),
	.w5(32'h3bd13150),
	.w6(32'h36d273ca),
	.w7(32'hbb98bb7c),
	.w8(32'hbb3c64f4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cdabd),
	.w1(32'h3ae93962),
	.w2(32'hbac9c743),
	.w3(32'h3bd342cb),
	.w4(32'h39f5df7b),
	.w5(32'hbc0273c0),
	.w6(32'h3a6aaebb),
	.w7(32'hbb1a340b),
	.w8(32'hbbcd0452),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba23bdd),
	.w1(32'hbc065f80),
	.w2(32'hbbbcaf61),
	.w3(32'hbb5b8949),
	.w4(32'hbbc4d187),
	.w5(32'hbbfbec34),
	.w6(32'hbbbc9e6e),
	.w7(32'hbbc68f83),
	.w8(32'hbc01d8cf),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aade0e),
	.w1(32'h3aa05b55),
	.w2(32'hbb543b26),
	.w3(32'h3b048d55),
	.w4(32'h3c0e24fc),
	.w5(32'h3babfe61),
	.w6(32'hbacba789),
	.w7(32'hbbeaf8c7),
	.w8(32'hbc0582b5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b8ff5),
	.w1(32'h3ab04345),
	.w2(32'h3b5fd076),
	.w3(32'h3baa03bf),
	.w4(32'h39e2a595),
	.w5(32'h3a3c0bdf),
	.w6(32'h3aaa8db1),
	.w7(32'h3b199128),
	.w8(32'h3acbb625),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af92306),
	.w1(32'hbb065b02),
	.w2(32'hbaba6226),
	.w3(32'hba53e752),
	.w4(32'hbaa4fd93),
	.w5(32'hb9ec2561),
	.w6(32'h3addc85f),
	.w7(32'h3b6d1976),
	.w8(32'hba995b4d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba296c95),
	.w1(32'hba4dfa82),
	.w2(32'hba1c5501),
	.w3(32'h3a918ae7),
	.w4(32'hb898dcdd),
	.w5(32'hbab08617),
	.w6(32'h3ae9b3aa),
	.w7(32'h3b480ebb),
	.w8(32'h3aaf17a4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc5c2c),
	.w1(32'hbb6e57ac),
	.w2(32'hbb52d2fb),
	.w3(32'hba74d499),
	.w4(32'hbaf6482f),
	.w5(32'hbb679963),
	.w6(32'hbb19bcb4),
	.w7(32'hbb149617),
	.w8(32'hba98ab43),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ec21e),
	.w1(32'hbb2434b2),
	.w2(32'h3b223d74),
	.w3(32'hba986987),
	.w4(32'hbb5cf4fb),
	.w5(32'hbba23a98),
	.w6(32'hbb9cde4d),
	.w7(32'hbbb55c0b),
	.w8(32'h3a495276),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379bcc86),
	.w1(32'hbc3c859d),
	.w2(32'h3c725bdd),
	.w3(32'hbb455c25),
	.w4(32'h3a6fe750),
	.w5(32'hbca93e42),
	.w6(32'h3c025052),
	.w7(32'hbc60ef80),
	.w8(32'hba9e448d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47fcce),
	.w1(32'hbb7134bd),
	.w2(32'hbc0d239c),
	.w3(32'h3b916d4f),
	.w4(32'hbb91a976),
	.w5(32'hbb45bc22),
	.w6(32'h3ae8f509),
	.w7(32'hbb83f69b),
	.w8(32'hbbc1c15a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94a9c6),
	.w1(32'h3b8fc370),
	.w2(32'h3b142286),
	.w3(32'h3b580115),
	.w4(32'h3b85d74f),
	.w5(32'hba0d3d39),
	.w6(32'h3a98f064),
	.w7(32'h3b510dca),
	.w8(32'h3b5d40d1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07c053),
	.w1(32'hbb2ff77a),
	.w2(32'hbba62c09),
	.w3(32'hbb2da952),
	.w4(32'hbb7edf19),
	.w5(32'hbb76f8c6),
	.w6(32'h3b07c685),
	.w7(32'hba1edc66),
	.w8(32'hbb3b15f7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb204de7),
	.w1(32'hb99f8df3),
	.w2(32'hbb344903),
	.w3(32'h3b992cc4),
	.w4(32'h3b207fe6),
	.w5(32'hb9deadaa),
	.w6(32'h3bdc5c58),
	.w7(32'h3b2da900),
	.w8(32'hbb5adaaf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306e69),
	.w1(32'hba566db8),
	.w2(32'hbba12586),
	.w3(32'h3a61f0b3),
	.w4(32'h391facd3),
	.w5(32'hbb39aea7),
	.w6(32'h3a9428cf),
	.w7(32'hbacf8f79),
	.w8(32'hbac73cf9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b7263),
	.w1(32'hbbacb320),
	.w2(32'hbb94725c),
	.w3(32'hbaa18bd5),
	.w4(32'hbc011eda),
	.w5(32'hbb9be529),
	.w6(32'hba9a4cea),
	.w7(32'hbb55e47e),
	.w8(32'hbb8dea00),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a592bf3),
	.w1(32'hbaed579a),
	.w2(32'hba98dab9),
	.w3(32'hba990367),
	.w4(32'hb9efb2d6),
	.w5(32'hba7a4e85),
	.w6(32'hbaffa5e5),
	.w7(32'hbb6e59b5),
	.w8(32'hbb7002ca),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a297e),
	.w1(32'hbb26efd0),
	.w2(32'hbb3a0430),
	.w3(32'hba01c54c),
	.w4(32'hbb72dfca),
	.w5(32'hb949a0cd),
	.w6(32'h398efd6b),
	.w7(32'h3b4e4f87),
	.w8(32'h3b3aeada),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9297ef2),
	.w1(32'h3ad38b1e),
	.w2(32'hb9e8ba92),
	.w3(32'hbb676718),
	.w4(32'h39b2d695),
	.w5(32'hbaa80c5f),
	.w6(32'h3b7c1f75),
	.w7(32'h3b1ae3a9),
	.w8(32'h3b920ec5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcc65d),
	.w1(32'h3b34d4bf),
	.w2(32'h3b57704e),
	.w3(32'hbb286598),
	.w4(32'h3a3baae8),
	.w5(32'h3b332777),
	.w6(32'h3b88f81a),
	.w7(32'h3bf0ec65),
	.w8(32'h3b608d39),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0582ae),
	.w1(32'h3b295463),
	.w2(32'h3bb38638),
	.w3(32'h3aa40322),
	.w4(32'h3bd562f8),
	.w5(32'hba7158e2),
	.w6(32'hb8811fd1),
	.w7(32'hbbe64ba1),
	.w8(32'hbb2089d8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20c93f),
	.w1(32'hba0aaab9),
	.w2(32'hbaf280fc),
	.w3(32'h3992c9f4),
	.w4(32'h3a03b802),
	.w5(32'hba803053),
	.w6(32'h3a0841a4),
	.w7(32'h3b320b8f),
	.w8(32'h3a9bb632),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23ae32),
	.w1(32'h3a90a367),
	.w2(32'h3b131bd2),
	.w3(32'h3a6c578d),
	.w4(32'h3b360450),
	.w5(32'h3a8480b7),
	.w6(32'h3b66e166),
	.w7(32'h3ae0723c),
	.w8(32'hb8cc868b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82e9c3),
	.w1(32'hbbe73634),
	.w2(32'hbc020ea1),
	.w3(32'hb9ae6468),
	.w4(32'hbbe894c7),
	.w5(32'hbbd74ca9),
	.w6(32'hbaa3c172),
	.w7(32'hbba71fda),
	.w8(32'hbbc6cefc),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b28d4),
	.w1(32'hbaac2b5c),
	.w2(32'hbb90bef6),
	.w3(32'h3a10fefb),
	.w4(32'h3b12a334),
	.w5(32'h39af88ce),
	.w6(32'hbadb074e),
	.w7(32'h3b1b3065),
	.w8(32'hb999cf96),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48d352),
	.w1(32'h3b5af0a4),
	.w2(32'hba93876b),
	.w3(32'h3b02e4b9),
	.w4(32'h3ba0fa5e),
	.w5(32'h3b0aab00),
	.w6(32'h3ba18f01),
	.w7(32'h3b2a0197),
	.w8(32'hbb94e548),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18a3e3),
	.w1(32'hbb526161),
	.w2(32'hbb38229b),
	.w3(32'h3b2fc1cc),
	.w4(32'hbb230b7f),
	.w5(32'hbb06bf8f),
	.w6(32'hbb0658dd),
	.w7(32'hbaa51156),
	.w8(32'h3ad54fd4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac85a2d),
	.w1(32'hbb60730b),
	.w2(32'hbb8146a6),
	.w3(32'hb815c9e0),
	.w4(32'hbb1232ac),
	.w5(32'hba061208),
	.w6(32'h392d1b5c),
	.w7(32'hbb948f76),
	.w8(32'hbb7525c3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aa342),
	.w1(32'hbb355d52),
	.w2(32'hbaff2ae4),
	.w3(32'hb9bde10c),
	.w4(32'hbb2ab13a),
	.w5(32'hbb5745ec),
	.w6(32'hba8579bb),
	.w7(32'hbb3ccc09),
	.w8(32'hbb1ebf81),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba727f03),
	.w1(32'hba084e34),
	.w2(32'hbb7f5124),
	.w3(32'hbb027158),
	.w4(32'hba74b9fb),
	.w5(32'h3bad9fa4),
	.w6(32'hbaa9bc79),
	.w7(32'h3c1af858),
	.w8(32'hbbb30dae),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b146e),
	.w1(32'hb963c5d5),
	.w2(32'h3b43779c),
	.w3(32'hbabb4c08),
	.w4(32'hbb90d404),
	.w5(32'hbb9c43ba),
	.w6(32'hbb209782),
	.w7(32'hbadbdd49),
	.w8(32'hba8b5640),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af67bf2),
	.w1(32'hbba2d3ab),
	.w2(32'hbc10e4d7),
	.w3(32'hba843371),
	.w4(32'hba85a6c9),
	.w5(32'hbbc090e8),
	.w6(32'hb9e5497f),
	.w7(32'hbb0faf96),
	.w8(32'hb980a6e8),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbc198),
	.w1(32'hbba22482),
	.w2(32'hbb7288ee),
	.w3(32'h39ce8ba6),
	.w4(32'h3a95195b),
	.w5(32'h3b0020ac),
	.w6(32'h3b01265a),
	.w7(32'hbad29393),
	.w8(32'hbbb1ebe8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c79fa),
	.w1(32'hbb3bc928),
	.w2(32'hbb9fd9fc),
	.w3(32'hba9c9551),
	.w4(32'h3a4857bd),
	.w5(32'hbbb40513),
	.w6(32'hbb823e65),
	.w7(32'hbb027198),
	.w8(32'hbbaa0b17),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6be835),
	.w1(32'hbb695b08),
	.w2(32'hbc2f642d),
	.w3(32'h3bca5701),
	.w4(32'h3c3b0998),
	.w5(32'hbbfce6bc),
	.w6(32'hbc584aba),
	.w7(32'h3b1f9216),
	.w8(32'hbc1e720e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa526ac),
	.w1(32'h3bd78084),
	.w2(32'hbbaca9b3),
	.w3(32'h3bf3769e),
	.w4(32'h38c5e550),
	.w5(32'h3c58395a),
	.w6(32'hb9ae6414),
	.w7(32'h3c979d1d),
	.w8(32'hbc7d94ca),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4e21b),
	.w1(32'hbbc5bf45),
	.w2(32'hbc1bfe3e),
	.w3(32'h3c4fddab),
	.w4(32'h3b720fbc),
	.w5(32'h39faf905),
	.w6(32'h3bc50cda),
	.w7(32'h3b4d1fb9),
	.w8(32'hbbf9c3b5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae828da),
	.w1(32'hba71019d),
	.w2(32'hb9242e40),
	.w3(32'h3b807182),
	.w4(32'hbaa2a633),
	.w5(32'hba69b553),
	.w6(32'h3a8c0e0d),
	.w7(32'h3b8942b3),
	.w8(32'hba3db07b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07db12),
	.w1(32'hbc39e5f3),
	.w2(32'hbc3de757),
	.w3(32'hbbe74a41),
	.w4(32'hbad90914),
	.w5(32'hbb1c2234),
	.w6(32'hbb638151),
	.w7(32'h3a5cf267),
	.w8(32'hbbe59be6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66f9e7),
	.w1(32'hbb20b5f1),
	.w2(32'hbb9ebe45),
	.w3(32'h3b925296),
	.w4(32'h3b13788c),
	.w5(32'hbbb41904),
	.w6(32'h3b21d33a),
	.w7(32'h3b3a3de4),
	.w8(32'hbb4aaaf9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bc134),
	.w1(32'hbb4ccf67),
	.w2(32'hbb02c8d6),
	.w3(32'hba5ac1a8),
	.w4(32'hbb9af0a7),
	.w5(32'hbb907ce3),
	.w6(32'hb97365a2),
	.w7(32'h3b0783c6),
	.w8(32'h3b2878f5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cee90),
	.w1(32'hbae79caa),
	.w2(32'hbb79a0b7),
	.w3(32'hbbcef20f),
	.w4(32'h3a9574a0),
	.w5(32'hba036fe4),
	.w6(32'hbb26d590),
	.w7(32'h3ae207ab),
	.w8(32'h3abb828c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa37eee),
	.w1(32'h3a00085d),
	.w2(32'hbb898506),
	.w3(32'h3b8de3da),
	.w4(32'h3a614123),
	.w5(32'hba7284f0),
	.w6(32'h3ba06a53),
	.w7(32'hb9232151),
	.w8(32'hbb886634),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a119d9c),
	.w1(32'h3b5176a2),
	.w2(32'hbabae078),
	.w3(32'h3b993986),
	.w4(32'hb9a2b243),
	.w5(32'hbb13f4f4),
	.w6(32'h3b125376),
	.w7(32'hbb7239bc),
	.w8(32'hbb5c2f04),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf791b2),
	.w1(32'hbb39804e),
	.w2(32'hbb902974),
	.w3(32'hbb43c8ef),
	.w4(32'hbace36d5),
	.w5(32'hbbb5a9e4),
	.w6(32'hbb12d4e5),
	.w7(32'hbb7e8f25),
	.w8(32'h39bf025a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a6b48),
	.w1(32'hbb452393),
	.w2(32'hbc4b6bc6),
	.w3(32'hbb7561ec),
	.w4(32'h3bab146b),
	.w5(32'h3b1f043e),
	.w6(32'hb93a49c7),
	.w7(32'hbbcea452),
	.w8(32'h3a9776d6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e3224),
	.w1(32'h3b8de7df),
	.w2(32'h3bc2ace3),
	.w3(32'h3b57b4c4),
	.w4(32'h3b6c14f2),
	.w5(32'hbba41cc1),
	.w6(32'hbb53d5c9),
	.w7(32'h3b1eece0),
	.w8(32'h3a920eee),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab68dde),
	.w1(32'hbb227652),
	.w2(32'h3b840d28),
	.w3(32'hbbd11704),
	.w4(32'hbb1e2e05),
	.w5(32'hbb979675),
	.w6(32'hbb405cdf),
	.w7(32'hbbf1cdda),
	.w8(32'hbb35b35a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2c2b8),
	.w1(32'hbb806970),
	.w2(32'hbbe8867f),
	.w3(32'hbb3bdf4d),
	.w4(32'h3b7e8a68),
	.w5(32'h3b5bdc3a),
	.w6(32'hbb37ea17),
	.w7(32'hbbbde149),
	.w8(32'hb80b3e94),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb799932),
	.w1(32'hbadf0575),
	.w2(32'hbbb2e4fe),
	.w3(32'h3b4fdb90),
	.w4(32'h3a943e68),
	.w5(32'h3acb376c),
	.w6(32'h3b192646),
	.w7(32'h3ac05021),
	.w8(32'h3999c799),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfbec5),
	.w1(32'hbac4b7a7),
	.w2(32'hba98e129),
	.w3(32'h3b1abe93),
	.w4(32'h39aa45a8),
	.w5(32'h39fcc9e9),
	.w6(32'h3b040d96),
	.w7(32'h3b837aaf),
	.w8(32'h3b00a1cf),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4cc5b6),
	.w1(32'hbacf3169),
	.w2(32'hbb0289e9),
	.w3(32'h3acfa126),
	.w4(32'h39b7aa3c),
	.w5(32'h399c6aca),
	.w6(32'h3b0210ec),
	.w7(32'h3b6dc8fb),
	.w8(32'h3ab3bdb2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378f9797),
	.w1(32'hbb15bfec),
	.w2(32'hba8fba2e),
	.w3(32'h3ad31c33),
	.w4(32'h3c037af0),
	.w5(32'h3cb6955d),
	.w6(32'hbbe2aea7),
	.w7(32'hbaa93cb2),
	.w8(32'hbc166078),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecbb02),
	.w1(32'h3bb680a1),
	.w2(32'hbaeb04d0),
	.w3(32'h3c0e6b78),
	.w4(32'h3ae2e602),
	.w5(32'hbab5497d),
	.w6(32'h3bb39a32),
	.w7(32'h3ac208e8),
	.w8(32'hbbde1d7d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb050009),
	.w1(32'hbbc3fb40),
	.w2(32'hbbdb8935),
	.w3(32'hbabcc43d),
	.w4(32'hba9b80d7),
	.w5(32'hbb3231f7),
	.w6(32'hbb631db2),
	.w7(32'hbb98049a),
	.w8(32'hbb7047a8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7699d),
	.w1(32'hbbd2579c),
	.w2(32'hbc040a32),
	.w3(32'hba8af64d),
	.w4(32'hba859b9b),
	.w5(32'hbab7abd0),
	.w6(32'hba4cd885),
	.w7(32'hbb705649),
	.w8(32'hbad0afb0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaa720),
	.w1(32'h3b1418a5),
	.w2(32'hb9bb3ea4),
	.w3(32'h3943e802),
	.w4(32'h3b5a5cba),
	.w5(32'h3a2d2dde),
	.w6(32'hba927ed7),
	.w7(32'h3b2f591c),
	.w8(32'h39883d73),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaceebda),
	.w1(32'h3b7e1da6),
	.w2(32'h3b79f059),
	.w3(32'h3a46b4c1),
	.w4(32'h3b940644),
	.w5(32'h3cbcd4fe),
	.w6(32'hbb269ff9),
	.w7(32'h3ca6c3d6),
	.w8(32'h3ab477e0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc15f82),
	.w1(32'h39c0df1f),
	.w2(32'hbb8be895),
	.w3(32'h3b8727e4),
	.w4(32'hba03477a),
	.w5(32'hb9ca8d4e),
	.w6(32'h3b8bae81),
	.w7(32'h3b8f080d),
	.w8(32'hbad75e3f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb677cae),
	.w1(32'hbabd57f9),
	.w2(32'hbb80711e),
	.w3(32'hba2cce13),
	.w4(32'hb989d141),
	.w5(32'hbb327f56),
	.w6(32'hb8d9a101),
	.w7(32'h3a0bf394),
	.w8(32'hba3f643a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b1277),
	.w1(32'h390394a9),
	.w2(32'h3bd1de4b),
	.w3(32'h39401a8e),
	.w4(32'h3b6d4fef),
	.w5(32'hba45c65f),
	.w6(32'hbb2a31c5),
	.w7(32'hbcbb1f8c),
	.w8(32'hbb018b9b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c7915),
	.w1(32'hbb55b179),
	.w2(32'h3cbe946c),
	.w3(32'h3c11a942),
	.w4(32'hbb0f662c),
	.w5(32'hb9d86ec2),
	.w6(32'h3bfd2f9a),
	.w7(32'hbc53bcb3),
	.w8(32'hbaffc62f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06140a),
	.w1(32'h3c7282bc),
	.w2(32'h3bb35011),
	.w3(32'hbbdcc7fc),
	.w4(32'h3bae4c4f),
	.w5(32'hbc18e61f),
	.w6(32'h3bcb596f),
	.w7(32'hbb898765),
	.w8(32'hbc785ce0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63001c),
	.w1(32'h3c29b8c7),
	.w2(32'hbcf33468),
	.w3(32'hbbbea3a0),
	.w4(32'hbb4a5e6c),
	.w5(32'hbcf5b16a),
	.w6(32'h3c6d8180),
	.w7(32'h3d32edda),
	.w8(32'h3c4b4cba),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34f821),
	.w1(32'hbba3e30c),
	.w2(32'hbcf69a5a),
	.w3(32'hbbc22651),
	.w4(32'hbb384d9a),
	.w5(32'hbbeec888),
	.w6(32'h3bbf24c0),
	.w7(32'h3cb5b218),
	.w8(32'h3bf38241),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03f276),
	.w1(32'hbc0d94be),
	.w2(32'hbab55102),
	.w3(32'hb8be53ab),
	.w4(32'h3986bf4c),
	.w5(32'h3c35eb1f),
	.w6(32'h3b9baf9e),
	.w7(32'hbbc3df67),
	.w8(32'h3ac74ac9),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb580775),
	.w1(32'hbb189a64),
	.w2(32'h3c4c3c08),
	.w3(32'h3c55ea46),
	.w4(32'hb9c9d046),
	.w5(32'h3bb17919),
	.w6(32'hbb96807e),
	.w7(32'hbba99ec5),
	.w8(32'h3b35a2c7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf179e2),
	.w1(32'hbbf4a20a),
	.w2(32'h3c791606),
	.w3(32'hbb7a9701),
	.w4(32'hbaa466c7),
	.w5(32'h3bf8cd13),
	.w6(32'h3bac9ebb),
	.w7(32'hbc0e15c1),
	.w8(32'h3c2405c0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb2886),
	.w1(32'h3c0fda12),
	.w2(32'hbcec9964),
	.w3(32'hbb81a61c),
	.w4(32'hbbb8a1b5),
	.w5(32'hbcdec078),
	.w6(32'h3c66d63c),
	.w7(32'h3d2e7d4e),
	.w8(32'h3b882aa9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0aea8),
	.w1(32'hbc1599ef),
	.w2(32'h3cdad245),
	.w3(32'hbc1ea922),
	.w4(32'hbb8e997d),
	.w5(32'h3b94bd72),
	.w6(32'hbb1b5351),
	.w7(32'hbcc9caf0),
	.w8(32'hbbaad96c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdeea6b),
	.w1(32'h3c13b1a1),
	.w2(32'h3c6a1bfc),
	.w3(32'hbc7bf9b2),
	.w4(32'h3b04d2b9),
	.w5(32'hba651f42),
	.w6(32'h3af5d15c),
	.w7(32'hbbb91a95),
	.w8(32'h3b2733ee),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80a01c),
	.w1(32'h3b6f3372),
	.w2(32'hbd76e506),
	.w3(32'hbbe537ea),
	.w4(32'hbb70023a),
	.w5(32'hbcbd54c7),
	.w6(32'h3cba7cc0),
	.w7(32'h3d7a531f),
	.w8(32'h3c1d7734),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12aa01),
	.w1(32'hbc67a561),
	.w2(32'hbc9058fc),
	.w3(32'h3b65a5f4),
	.w4(32'h3a3b5332),
	.w5(32'hbb98630b),
	.w6(32'hbb94c524),
	.w7(32'hbc18e9e6),
	.w8(32'hba1718ed),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81f545),
	.w1(32'hb98c822a),
	.w2(32'hbaacd2bc),
	.w3(32'h3bb4b576),
	.w4(32'h392f0b29),
	.w5(32'hbaacf5d4),
	.w6(32'h3b01e40b),
	.w7(32'hba88654e),
	.w8(32'hbb22bb6b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ab54c),
	.w1(32'hbc1e2d09),
	.w2(32'hbc3b733d),
	.w3(32'hbb46a36c),
	.w4(32'hbb9204fc),
	.w5(32'hbb96d782),
	.w6(32'h3aa42a66),
	.w7(32'hbc52ff08),
	.w8(32'hbb3f535a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe15359),
	.w1(32'hbbafc73f),
	.w2(32'h3d3435e6),
	.w3(32'h3a1bfde8),
	.w4(32'h3b894c9e),
	.w5(32'h3cda145d),
	.w6(32'h3a4a3f97),
	.w7(32'hbcd55b10),
	.w8(32'h3be79ef5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80f5db),
	.w1(32'h3b780804),
	.w2(32'hbb9f5212),
	.w3(32'hbbb54e95),
	.w4(32'h3a093263),
	.w5(32'h39fffa79),
	.w6(32'hbb265213),
	.w7(32'h3ad79ff3),
	.w8(32'hbc154b91),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc412882),
	.w1(32'h3b6532a9),
	.w2(32'h3c8df676),
	.w3(32'hbb900a86),
	.w4(32'hbbf79791),
	.w5(32'hbb96bec1),
	.w6(32'h3b038952),
	.w7(32'hbae0c6db),
	.w8(32'h3bd380e0),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1bf05),
	.w1(32'h3bb260db),
	.w2(32'h3b30a9d4),
	.w3(32'hbc2b2b62),
	.w4(32'hbba6c206),
	.w5(32'hbc055a02),
	.w6(32'hba641172),
	.w7(32'h3b05fa83),
	.w8(32'hbb09120d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26176e),
	.w1(32'h3c033541),
	.w2(32'hbd3772ac),
	.w3(32'hba33b3d2),
	.w4(32'hbbed9950),
	.w5(32'hbd000377),
	.w6(32'h3c6c0b8d),
	.w7(32'h3d6894c1),
	.w8(32'h3bcec70d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79a200),
	.w1(32'h3b7d8d96),
	.w2(32'hbc12e597),
	.w3(32'hbbc10dcd),
	.w4(32'hbc0d0ed3),
	.w5(32'hbc76ed14),
	.w6(32'h3be3af6f),
	.w7(32'h3d00f584),
	.w8(32'h3c255d57),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7da2c),
	.w1(32'h3b5f9dea),
	.w2(32'h3c0429ee),
	.w3(32'hbb89c509),
	.w4(32'hbb0c21f6),
	.w5(32'hbb2eee74),
	.w6(32'h3b41a245),
	.w7(32'hbb2b8536),
	.w8(32'h3b6c01fd),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39f90c),
	.w1(32'hbc5bc0ce),
	.w2(32'h3c21ceb4),
	.w3(32'hbbacafb0),
	.w4(32'hbbee8e51),
	.w5(32'h3af466c4),
	.w6(32'hbc72fa5b),
	.w7(32'hbcd4e042),
	.w8(32'hbc0bddad),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96db6e),
	.w1(32'hbc0aa507),
	.w2(32'hbc98b694),
	.w3(32'hbaebfc25),
	.w4(32'hbb6a4500),
	.w5(32'hbaa0cc84),
	.w6(32'hbb509305),
	.w7(32'hbb4e07a7),
	.w8(32'hbc41e8dd),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbd308),
	.w1(32'hbb8950dd),
	.w2(32'hbc1d9506),
	.w3(32'h39dda44c),
	.w4(32'h3a7cd2a9),
	.w5(32'hbba08166),
	.w6(32'hbad8da0f),
	.w7(32'hbc8603a6),
	.w8(32'hbb65b566),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55b5ad),
	.w1(32'hbc1b4d1b),
	.w2(32'h3cba3180),
	.w3(32'h3b8e5ed2),
	.w4(32'hbba978b1),
	.w5(32'hb9bf8cba),
	.w6(32'h3ab52a2d),
	.w7(32'hbcc60d77),
	.w8(32'hbc18cdb8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba27457),
	.w1(32'hbbe43381),
	.w2(32'hbc852673),
	.w3(32'hbc6e791b),
	.w4(32'h39de1dd2),
	.w5(32'hbb25e9af),
	.w6(32'h3b77347f),
	.w7(32'h3b27ef3b),
	.w8(32'h3b4c1b32),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a680965),
	.w1(32'hbc2db9bd),
	.w2(32'hbc79c8fb),
	.w3(32'h38943b6a),
	.w4(32'hbc1b045f),
	.w5(32'h3a931702),
	.w6(32'hb86b4e24),
	.w7(32'hba88e1ce),
	.w8(32'hbaeda87d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbb2b7),
	.w1(32'hbb01c958),
	.w2(32'h3bddade9),
	.w3(32'hbbf02411),
	.w4(32'hbbe1ab6f),
	.w5(32'hbbdae0e2),
	.w6(32'h3b153b4d),
	.w7(32'hbb8ca7ab),
	.w8(32'h3ae48d63),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8914b07),
	.w1(32'hbb54798b),
	.w2(32'hbc65b309),
	.w3(32'hbbda9625),
	.w4(32'hbbb1e4f6),
	.w5(32'hbace44aa),
	.w6(32'h3c1e7b42),
	.w7(32'h3b0d3c71),
	.w8(32'hbb4d7bff),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55318e),
	.w1(32'hbb45842b),
	.w2(32'hbc69d9c7),
	.w3(32'h3a7f63bb),
	.w4(32'h3c0ddc0b),
	.w5(32'hbc080eb4),
	.w6(32'h3b19ce3d),
	.w7(32'hbc6b9cb2),
	.w8(32'hbb01d5b9),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6a2f8),
	.w1(32'h3bee445a),
	.w2(32'h3c0f69e6),
	.w3(32'hb8aa18f9),
	.w4(32'h3bbf3baa),
	.w5(32'h3bedbbe0),
	.w6(32'hbb2de1cb),
	.w7(32'h3b67b725),
	.w8(32'h3aa7d3bb),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d67c4),
	.w1(32'hbc32a683),
	.w2(32'h3a991fed),
	.w3(32'h3b8ed5a6),
	.w4(32'hbbe6942c),
	.w5(32'hbb632cdf),
	.w6(32'hbc0df7b4),
	.w7(32'hbc6848fb),
	.w8(32'hbbca9571),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae6275),
	.w1(32'hbc30f0d6),
	.w2(32'hba9058d2),
	.w3(32'hbbadfcf3),
	.w4(32'hbc032281),
	.w5(32'hbc04bb9e),
	.w6(32'hbb118062),
	.w7(32'hbc2fcacb),
	.w8(32'hbb4b944e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85f261),
	.w1(32'hb964f44e),
	.w2(32'h3bbb0dff),
	.w3(32'hbbcf5b87),
	.w4(32'hbc09efdd),
	.w5(32'h3a195cca),
	.w6(32'h3be89b0d),
	.w7(32'h3a856415),
	.w8(32'h3ac8b901),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffeae6),
	.w1(32'h3c0a492d),
	.w2(32'hbb5d3df6),
	.w3(32'hbc14ed4c),
	.w4(32'h3b93f5dc),
	.w5(32'hb9a80031),
	.w6(32'h3c6c1526),
	.w7(32'hbb799bcd),
	.w8(32'hbb5a1263),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7897f),
	.w1(32'h3bb1d5f7),
	.w2(32'hbd48794c),
	.w3(32'hbc5332ed),
	.w4(32'hbc14e233),
	.w5(32'hbd0cabc0),
	.w6(32'h3c7224dc),
	.w7(32'h3d3c5a75),
	.w8(32'h3baa2b87),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc632bb7),
	.w1(32'hbc101bb7),
	.w2(32'hbbc24b77),
	.w3(32'hbc3cae7c),
	.w4(32'hbc317ae7),
	.w5(32'hbc98a805),
	.w6(32'hbac57ec8),
	.w7(32'hbbb88123),
	.w8(32'hba979e3e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8723f3),
	.w1(32'h3bdbaa4d),
	.w2(32'hbd0941f6),
	.w3(32'hbbf640f9),
	.w4(32'h3a561c54),
	.w5(32'hbcbf6adb),
	.w6(32'h3c06392f),
	.w7(32'h3d108ab1),
	.w8(32'h3b0e6427),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc989e0b),
	.w1(32'h3c52d29c),
	.w2(32'hbcc05a98),
	.w3(32'hbc0fbd6f),
	.w4(32'hbb5f800d),
	.w5(32'hbcb61b50),
	.w6(32'h3c8281d6),
	.w7(32'h3d350606),
	.w8(32'h3c647d08),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d504f),
	.w1(32'hbb2d585a),
	.w2(32'h3cda3327),
	.w3(32'hbb96c5f2),
	.w4(32'hbac9d0df),
	.w5(32'h3bb69db4),
	.w6(32'h3b437033),
	.w7(32'hbc6a9463),
	.w8(32'hbaca2e02),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f305a2),
	.w1(32'h3c08776d),
	.w2(32'hbc8fc160),
	.w3(32'hbc139a35),
	.w4(32'hbb2882fd),
	.w5(32'hbc8bb171),
	.w6(32'h3c029812),
	.w7(32'h3d079066),
	.w8(32'h3bef65b9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ee0c4),
	.w1(32'h3bceaee0),
	.w2(32'h3b51d4a7),
	.w3(32'hbbb3276e),
	.w4(32'h3be17ebf),
	.w5(32'hb9ae2711),
	.w6(32'hbb238907),
	.w7(32'hbc2e66aa),
	.w8(32'hbc7f3eed),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e5534),
	.w1(32'h3b5100e2),
	.w2(32'hbc927430),
	.w3(32'h3b7e1444),
	.w4(32'hbb9c9ad2),
	.w5(32'hbc8b1b77),
	.w6(32'h3b3f32f6),
	.w7(32'h3c987565),
	.w8(32'h3bfb0adc),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abee72a),
	.w1(32'hbbbfb3ab),
	.w2(32'h3b22f22d),
	.w3(32'hbaada456),
	.w4(32'hbb37a77b),
	.w5(32'hbb2e1949),
	.w6(32'hbac0054e),
	.w7(32'hbc60923a),
	.w8(32'hbbbd5627),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d757b4),
	.w1(32'h3ca59bde),
	.w2(32'hbd6d0377),
	.w3(32'hbb6b8fce),
	.w4(32'h3bad29c6),
	.w5(32'hbca61042),
	.w6(32'h3d08fd44),
	.w7(32'h3da0667e),
	.w8(32'h3c49d318),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc859436),
	.w1(32'hba090471),
	.w2(32'hbc8ab2a2),
	.w3(32'h3c08d976),
	.w4(32'hbc107afb),
	.w5(32'hbc8f2306),
	.w6(32'h3b4b7454),
	.w7(32'h3cdc74a9),
	.w8(32'h3c78e374),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cd8d0),
	.w1(32'h3b3a83e1),
	.w2(32'hbc435294),
	.w3(32'hbbae4782),
	.w4(32'hbc331c45),
	.w5(32'hbc8c7c42),
	.w6(32'h3bec7445),
	.w7(32'h3cc75f49),
	.w8(32'h3c0ea53e),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937e629),
	.w1(32'hbb5f612f),
	.w2(32'hb9fdf1fe),
	.w3(32'hbb9eb0a3),
	.w4(32'h3b830baf),
	.w5(32'h3bf59ad3),
	.w6(32'hbb156091),
	.w7(32'hbc2f7cfd),
	.w8(32'hbc3b9b0d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcae11),
	.w1(32'hba9ca1bd),
	.w2(32'hbb18427a),
	.w3(32'h3be3baea),
	.w4(32'hbaa5803a),
	.w5(32'hba787f1a),
	.w6(32'hbb16d452),
	.w7(32'h3b45e1f6),
	.w8(32'hbb7a5d8f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce14c7),
	.w1(32'hbbda065e),
	.w2(32'hbb02f3e9),
	.w3(32'h3a031523),
	.w4(32'hbb8bc34f),
	.w5(32'hbb676c92),
	.w6(32'h3b3af455),
	.w7(32'hbc19f490),
	.w8(32'hba423c6f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb153679),
	.w1(32'hbbea75a8),
	.w2(32'h3cf6a867),
	.w3(32'hbb87c5d7),
	.w4(32'hbbb6d56d),
	.w5(32'h3be01525),
	.w6(32'h39eee83c),
	.w7(32'hbc86ff4b),
	.w8(32'h3b31569d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e7d5a),
	.w1(32'h3b258f5b),
	.w2(32'hbcdbed75),
	.w3(32'hbc39302b),
	.w4(32'hbc064806),
	.w5(32'hbc7b05ac),
	.w6(32'h3c29e6eb),
	.w7(32'h3cf48103),
	.w8(32'h3c2458ed),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9940df),
	.w1(32'hba338e27),
	.w2(32'hbb9119c3),
	.w3(32'h3a754fb4),
	.w4(32'hbc098e1d),
	.w5(32'hbb8963db),
	.w6(32'hba366d4f),
	.w7(32'hbbaf4ccf),
	.w8(32'hbba26c7e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fb664),
	.w1(32'hbb9d4c9c),
	.w2(32'h3c083150),
	.w3(32'hba9dbdb6),
	.w4(32'hbc01b40c),
	.w5(32'hbc23e3cd),
	.w6(32'h3b338137),
	.w7(32'h3ad5835f),
	.w8(32'h3c25a489),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e21d0),
	.w1(32'hbc36a623),
	.w2(32'hbb147ec3),
	.w3(32'hbc3e7870),
	.w4(32'hbb9a4819),
	.w5(32'hbb9deae7),
	.w6(32'hbb9f6430),
	.w7(32'h3b8bb737),
	.w8(32'h3b994f3d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef96d1),
	.w1(32'hbaf2ff05),
	.w2(32'hbc48fa01),
	.w3(32'hbbdd0c05),
	.w4(32'hba8db428),
	.w5(32'hbc1f1d9c),
	.w6(32'h3c11b8cf),
	.w7(32'h3c9526ec),
	.w8(32'h3bd7e94e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09b7bc),
	.w1(32'hbb27fdea),
	.w2(32'hbad14cdf),
	.w3(32'h3b7c74fe),
	.w4(32'h3b061b20),
	.w5(32'hbb8d5bf4),
	.w6(32'hbb955301),
	.w7(32'hbc727c99),
	.w8(32'hbbd259e0),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a032fdd),
	.w1(32'hbbcdbdf5),
	.w2(32'hbc4bfe5c),
	.w3(32'h3b3865ae),
	.w4(32'hbb2a7b7c),
	.w5(32'hbc62e0bd),
	.w6(32'h3a5214df),
	.w7(32'h3c636288),
	.w8(32'h3be3d889),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71e1a9),
	.w1(32'h3ac834fa),
	.w2(32'h3c0a59a0),
	.w3(32'h3af64bc8),
	.w4(32'hbc22490e),
	.w5(32'hbc267448),
	.w6(32'h3c2c58fd),
	.w7(32'hbb776c80),
	.w8(32'hbb837a5b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c613f60),
	.w1(32'h3b63c909),
	.w2(32'hbd016174),
	.w3(32'h3b664cd7),
	.w4(32'hbbce9033),
	.w5(32'hbcd5cfff),
	.w6(32'h3c9d6b59),
	.w7(32'h3d2fbca9),
	.w8(32'h3b485f5a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80eb1b),
	.w1(32'hbc202a3e),
	.w2(32'h3cbddade),
	.w3(32'h3b62b0d6),
	.w4(32'hbbd2b23d),
	.w5(32'h398ce10e),
	.w6(32'h3ba84d59),
	.w7(32'hbcbe58f9),
	.w8(32'hbc1ca4c3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc38e8c),
	.w1(32'h3ac6b0d6),
	.w2(32'hbce07f4a),
	.w3(32'hbc62bd34),
	.w4(32'hbb209c47),
	.w5(32'hbc958826),
	.w6(32'h3bd6ac82),
	.w7(32'h3d2d5a67),
	.w8(32'h3ca152b9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11e591),
	.w1(32'hbbef45db),
	.w2(32'h3c3e6c87),
	.w3(32'hbbaf226e),
	.w4(32'hb9fbaf8b),
	.w5(32'h3beea1c2),
	.w6(32'hbb0e145b),
	.w7(32'hbc678e7b),
	.w8(32'hbbf4f361),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8af882),
	.w1(32'hbbf7ffbc),
	.w2(32'h3c211d8b),
	.w3(32'hbc79cafa),
	.w4(32'hbc502441),
	.w5(32'hbc0acf66),
	.w6(32'h3b2598fb),
	.w7(32'h3c53f75c),
	.w8(32'h3c57dcc8),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d9610),
	.w1(32'h3c6281bf),
	.w2(32'hbd2b17ca),
	.w3(32'hbbab8961),
	.w4(32'h3b24cb39),
	.w5(32'hbc8c1d9e),
	.w6(32'h3cc2e3af),
	.w7(32'h3d6a06c1),
	.w8(32'h3c25e06e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc096d54),
	.w1(32'hbaaf39d6),
	.w2(32'hbc1068ac),
	.w3(32'h3bb979b5),
	.w4(32'hbb6df710),
	.w5(32'hbbfa4ebe),
	.w6(32'h3ba52bee),
	.w7(32'h3cc75e19),
	.w8(32'h3c0880de),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef645b),
	.w1(32'hbae32349),
	.w2(32'h3ab8d6f8),
	.w3(32'hbb4c473c),
	.w4(32'hba26baf1),
	.w5(32'h3b97535a),
	.w6(32'h3c3bcf7a),
	.w7(32'hbc1befc1),
	.w8(32'hbbcab3a1),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a9740),
	.w1(32'h3b5e0e9f),
	.w2(32'hbb4726af),
	.w3(32'h3c623f8b),
	.w4(32'h3b3daee2),
	.w5(32'h3a39162b),
	.w6(32'h3b32c3bd),
	.w7(32'h3ad92b74),
	.w8(32'hb8d0e930),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe7a72),
	.w1(32'hbb5d5b48),
	.w2(32'hbb843155),
	.w3(32'h3bd54483),
	.w4(32'h39a627b9),
	.w5(32'hbb8e426e),
	.w6(32'hbbb3adfc),
	.w7(32'hbc2bd4dd),
	.w8(32'hbbed0931),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba923f26),
	.w1(32'hbb4b7271),
	.w2(32'h3cd13d80),
	.w3(32'h3b9abab3),
	.w4(32'hbc28a1e6),
	.w5(32'hbc2b28c9),
	.w6(32'h3b1c52de),
	.w7(32'hb9edcfee),
	.w8(32'h3b242a61),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99386b),
	.w1(32'hbbd8f857),
	.w2(32'hbc487bed),
	.w3(32'hbc81e3d0),
	.w4(32'hbbab4d22),
	.w5(32'hbc396e5a),
	.w6(32'h3bc11985),
	.w7(32'h3b8eb91b),
	.w8(32'hba39e31f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44115b),
	.w1(32'h3bedb4b3),
	.w2(32'hbd08e220),
	.w3(32'h3bc1975c),
	.w4(32'hbb9b6c9a),
	.w5(32'hbcee1653),
	.w6(32'h3c3ff871),
	.w7(32'h3d28b5ad),
	.w8(32'h3b62c6d1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbef149),
	.w1(32'hbb4e174d),
	.w2(32'h3ca8d5aa),
	.w3(32'hbb48e596),
	.w4(32'hbbd54ae7),
	.w5(32'hbbaf5ec4),
	.w6(32'h3b9ec75c),
	.w7(32'hbc1f8604),
	.w8(32'hbac9190b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a4f51),
	.w1(32'hbb4739b8),
	.w2(32'h3cc500b7),
	.w3(32'hbc80074a),
	.w4(32'hbb28297c),
	.w5(32'h3b121236),
	.w6(32'h3aa5b26a),
	.w7(32'hbc4c6f61),
	.w8(32'hbb24bdae),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e43a8),
	.w1(32'hbc7d9e14),
	.w2(32'hbaaadc5e),
	.w3(32'hbc3a6472),
	.w4(32'hbc47ef9e),
	.w5(32'hbc7157eb),
	.w6(32'hbb4f54cf),
	.w7(32'hbc2fabe0),
	.w8(32'hba8382a4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bf9b8),
	.w1(32'hba26587a),
	.w2(32'hbceea4d5),
	.w3(32'hbc662475),
	.w4(32'hbbcbf608),
	.w5(32'hbca03d43),
	.w6(32'h3c627105),
	.w7(32'h3d143b56),
	.w8(32'h3ba8d688),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b5fa2),
	.w1(32'hbc0f8b8c),
	.w2(32'hbcb73e05),
	.w3(32'h3b6faea4),
	.w4(32'hbadc1b86),
	.w5(32'h3b4e380e),
	.w6(32'hbc0e479f),
	.w7(32'h3aa0f762),
	.w8(32'hba6fdc73),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a3047),
	.w1(32'hbc4e385f),
	.w2(32'h3d0ca5ec),
	.w3(32'h3b346875),
	.w4(32'hb8c859ff),
	.w5(32'h3c9df3a1),
	.w6(32'hbb79b26c),
	.w7(32'hbd13f04a),
	.w8(32'hbbb8993a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3a0b9),
	.w1(32'hbb9b907f),
	.w2(32'hbcbca1bf),
	.w3(32'hbc173c50),
	.w4(32'hbc970a21),
	.w5(32'hbcd61263),
	.w6(32'h3bd0d8b4),
	.w7(32'h3d2b4c62),
	.w8(32'h3c855087),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0d69e),
	.w1(32'hb986d307),
	.w2(32'hbae9a32f),
	.w3(32'hbc10929b),
	.w4(32'h3b3a4ef7),
	.w5(32'h3a672b71),
	.w6(32'h3ad2ce33),
	.w7(32'hbb008878),
	.w8(32'hbb438b22),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3794a7),
	.w1(32'hbc2073e0),
	.w2(32'h3be041a7),
	.w3(32'h3adbf9c9),
	.w4(32'hbba6c536),
	.w5(32'hbbbac878),
	.w6(32'hbc521360),
	.w7(32'hbcdbdd27),
	.w8(32'hbc09e031),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9344f7),
	.w1(32'hbb88ce2e),
	.w2(32'hbba658c2),
	.w3(32'hbb1b86ec),
	.w4(32'h3b1ec702),
	.w5(32'hbbf2171a),
	.w6(32'hbb66d61e),
	.w7(32'hbc2cfd92),
	.w8(32'hbc0b71c2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8c9ed),
	.w1(32'h3ba0c5ba),
	.w2(32'hbca7f84e),
	.w3(32'h3b2b313a),
	.w4(32'hbb822b4d),
	.w5(32'hbce64039),
	.w6(32'h3bcad351),
	.w7(32'h3d16b370),
	.w8(32'h3c6fa7fc),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb916fb8d),
	.w1(32'hbba2a7de),
	.w2(32'hbbda7feb),
	.w3(32'hbc37e069),
	.w4(32'hbbe1129b),
	.w5(32'hbb9ff0cf),
	.w6(32'hbb2ec636),
	.w7(32'h3b35c8ab),
	.w8(32'h39585a21),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05f56c),
	.w1(32'h3ba625d5),
	.w2(32'hbcabf4b8),
	.w3(32'h3bee5d1d),
	.w4(32'hbbe4c375),
	.w5(32'hbce8809b),
	.w6(32'h3c3b1e12),
	.w7(32'h3d10281d),
	.w8(32'h3b7a96b2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a3ca6),
	.w1(32'hbaed5bcb),
	.w2(32'hbb1c9f22),
	.w3(32'hbbfd0a88),
	.w4(32'hbaf41eb4),
	.w5(32'hbc18bbb7),
	.w6(32'h39902647),
	.w7(32'hbb6d64d9),
	.w8(32'hbc8324fa),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16bbf5),
	.w1(32'h395d3516),
	.w2(32'hbc826775),
	.w3(32'hbb2b00fb),
	.w4(32'hbba6734c),
	.w5(32'hbc88eb35),
	.w6(32'h3b849be7),
	.w7(32'h3c6c122a),
	.w8(32'h3b33137e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06eae6),
	.w1(32'hbb61c639),
	.w2(32'hbb8a2608),
	.w3(32'h3baf2c37),
	.w4(32'hbc0cd0b0),
	.w5(32'hbc0207aa),
	.w6(32'hba3d6bd6),
	.w7(32'h3b5769cf),
	.w8(32'hbc421024),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e1faf),
	.w1(32'hbc2ec243),
	.w2(32'h3b57b571),
	.w3(32'hbacc4c83),
	.w4(32'hbbe01209),
	.w5(32'hbb836b15),
	.w6(32'hbc27b6a8),
	.w7(32'hbc6ab02c),
	.w8(32'hbbb5fcfb),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ce3b2),
	.w1(32'h3b143cea),
	.w2(32'hbbf234a7),
	.w3(32'hbbd5d39c),
	.w4(32'hb9ed40e5),
	.w5(32'hbbe85758),
	.w6(32'h3c290858),
	.w7(32'h3cad3e3f),
	.w8(32'h3c08010b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f591b),
	.w1(32'hbbbf4d36),
	.w2(32'h3bcea25f),
	.w3(32'h3c0c7688),
	.w4(32'hbb539742),
	.w5(32'hbc2dce56),
	.w6(32'hbc023977),
	.w7(32'hbc9c57cd),
	.w8(32'hbc5c824b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99664f),
	.w1(32'hbcdc43fc),
	.w2(32'hbbc8fbc7),
	.w3(32'hbbccecfa),
	.w4(32'hbc577698),
	.w5(32'hbbb5ac58),
	.w6(32'hbba2c9c9),
	.w7(32'hbc7fcdd7),
	.w8(32'hbbe1284a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4717ce),
	.w1(32'h3beb29c0),
	.w2(32'hbd0787bf),
	.w3(32'hbb7eca95),
	.w4(32'hbaa90b2a),
	.w5(32'hbcb2ba26),
	.w6(32'h3c7e68df),
	.w7(32'h3d4b232e),
	.w8(32'h3c60b134),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b91d3),
	.w1(32'h3b9e3c67),
	.w2(32'hbc16e80e),
	.w3(32'hb941c95b),
	.w4(32'hbba17b2e),
	.w5(32'hbcc2f8ae),
	.w6(32'h3bf79838),
	.w7(32'h3cf899be),
	.w8(32'h3c351301),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd8587),
	.w1(32'hbc22167a),
	.w2(32'hbc613370),
	.w3(32'hbc06fc49),
	.w4(32'hb9564541),
	.w5(32'hbc5cd768),
	.w6(32'hbc450d09),
	.w7(32'hbca1db0b),
	.w8(32'hbc112696),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb30a85),
	.w1(32'h3b7398d7),
	.w2(32'hbc9379fc),
	.w3(32'h3a865218),
	.w4(32'hbb0c5186),
	.w5(32'hbc42e5bb),
	.w6(32'h3b2bddab),
	.w7(32'h3c798119),
	.w8(32'h3a4fb214),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb205a63),
	.w1(32'hbc0ae9fc),
	.w2(32'h3b6deea4),
	.w3(32'hbae7a082),
	.w4(32'hbb4df767),
	.w5(32'hbad64594),
	.w6(32'h3b89c9b1),
	.w7(32'hb9f7c855),
	.w8(32'hbb27afb1),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6944a0),
	.w1(32'h3ac4d7cd),
	.w2(32'h3bd14d05),
	.w3(32'hbab2bb81),
	.w4(32'h3ac24c1d),
	.w5(32'h3bfb5aa4),
	.w6(32'hba3df618),
	.w7(32'h3b637251),
	.w8(32'h3b1ce35f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae42d17),
	.w1(32'hba36a54c),
	.w2(32'h3b190c87),
	.w3(32'h3b814274),
	.w4(32'h3abeedd5),
	.w5(32'h3c310437),
	.w6(32'h3c39260b),
	.w7(32'h3bde7f33),
	.w8(32'hbae07cc9),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79353d),
	.w1(32'h3b98f953),
	.w2(32'hbcb745df),
	.w3(32'h38a412e3),
	.w4(32'hbc25d3ff),
	.w5(32'hbcf262ee),
	.w6(32'h3c65b3cd),
	.w7(32'h3d4a46d2),
	.w8(32'h3c934762),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02123c),
	.w1(32'hbb721710),
	.w2(32'hbc55cfa6),
	.w3(32'hbc801bb1),
	.w4(32'hbb936c3c),
	.w5(32'hbc786c44),
	.w6(32'h3b241e5c),
	.w7(32'h3bd71613),
	.w8(32'hba83386a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb401d68),
	.w1(32'h3b0fe745),
	.w2(32'h3be1a3a9),
	.w3(32'hbb9dc8c7),
	.w4(32'h3809bb49),
	.w5(32'hbba789bc),
	.w6(32'h3b9948eb),
	.w7(32'h3b89f879),
	.w8(32'h3c17745d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ca3e1),
	.w1(32'hbc031d60),
	.w2(32'hba9a74da),
	.w3(32'hbc44aaf5),
	.w4(32'hbbeb6b95),
	.w5(32'hbc3d6164),
	.w6(32'hbb06b8fd),
	.w7(32'h3b04731d),
	.w8(32'h3bd56b40),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b9585),
	.w1(32'hbcb51bf6),
	.w2(32'h3d51fedd),
	.w3(32'h3ba687df),
	.w4(32'hbb8fbcdb),
	.w5(32'h3ce525bb),
	.w6(32'hba26f146),
	.w7(32'hbd5a8168),
	.w8(32'hbc55e922),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9c3a4),
	.w1(32'hbb4750ce),
	.w2(32'h3cc74815),
	.w3(32'hbc5319da),
	.w4(32'hbbdec1b5),
	.w5(32'hbb9778b5),
	.w6(32'h3be94ca0),
	.w7(32'hbc67c395),
	.w8(32'hbac2a7f7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71fa1d),
	.w1(32'hbc1d5d47),
	.w2(32'h3cda2a5e),
	.w3(32'hbc45cfd9),
	.w4(32'hba445161),
	.w5(32'h3c700a7b),
	.w6(32'hbb269f9b),
	.w7(32'hbcd9e243),
	.w8(32'hbb2de6ef),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92fa10),
	.w1(32'h3a6b1a5b),
	.w2(32'h3b93d640),
	.w3(32'hbbe3f23b),
	.w4(32'hbb5c9ecc),
	.w5(32'hbb54e8cf),
	.w6(32'h3b918c98),
	.w7(32'hbbedc90a),
	.w8(32'hbb3a2712),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa57d96),
	.w1(32'h3a2fb300),
	.w2(32'hbca042e8),
	.w3(32'hbb762226),
	.w4(32'hba166377),
	.w5(32'hbc3e82d0),
	.w6(32'h3c5477cc),
	.w7(32'h3cda33cd),
	.w8(32'h36bf2a22),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2d037),
	.w1(32'hbcabf212),
	.w2(32'hba30632f),
	.w3(32'hbb00abfc),
	.w4(32'hbc20df90),
	.w5(32'hbac1952d),
	.w6(32'hbc519879),
	.w7(32'hbc8e566b),
	.w8(32'hbbd6ee13),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc199c13),
	.w1(32'hbc2976b3),
	.w2(32'h3ce61bea),
	.w3(32'hbb8daf77),
	.w4(32'hba8bcbc0),
	.w5(32'h3c85d898),
	.w6(32'hbaeb5712),
	.w7(32'hbce34f8e),
	.w8(32'hbb0df9fc),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98f600),
	.w1(32'hba5c3a70),
	.w2(32'hbce96101),
	.w3(32'hbbfe6a92),
	.w4(32'hbb77acb3),
	.w5(32'hbc936b6d),
	.w6(32'h3c1fc106),
	.w7(32'h3d06c742),
	.w8(32'h3c220f57),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b215519),
	.w1(32'h3ac08a32),
	.w2(32'h3cc21508),
	.w3(32'hbb915154),
	.w4(32'hbb71cc56),
	.w5(32'h3b1867ce),
	.w6(32'h3bc11705),
	.w7(32'hba835521),
	.w8(32'h3bd83bf2),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb92e24),
	.w1(32'hbb11e511),
	.w2(32'h3bb175c6),
	.w3(32'hbc1a9aaa),
	.w4(32'h3c06c7cc),
	.w5(32'h3bdb9508),
	.w6(32'hbc538fc3),
	.w7(32'hbc17360a),
	.w8(32'hbb4bbccb),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc120227),
	.w1(32'hb990c557),
	.w2(32'h3caa7ae4),
	.w3(32'hbc54d299),
	.w4(32'hbc261ebb),
	.w5(32'hbbd901b2),
	.w6(32'h3c13d0ce),
	.w7(32'hba572c60),
	.w8(32'h3b7c6683),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b4aec),
	.w1(32'h3a9c4e10),
	.w2(32'hbd12f448),
	.w3(32'hbc2edf14),
	.w4(32'h3a9bc2e7),
	.w5(32'hbc3fead5),
	.w6(32'h3c3aaca0),
	.w7(32'h3c73859d),
	.w8(32'hbc56f755),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf95c12),
	.w1(32'hbbb6bc7b),
	.w2(32'h3c8bb128),
	.w3(32'h3c0ae54b),
	.w4(32'hbbf3b8ad),
	.w5(32'h3c062de2),
	.w6(32'hba148591),
	.w7(32'hbc123ed9),
	.w8(32'h3c43dd48),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc795a),
	.w1(32'hbc6bb787),
	.w2(32'h3d2346d8),
	.w3(32'hbc155e3f),
	.w4(32'hbaa1fb97),
	.w5(32'h3cbc2d4b),
	.w6(32'hbb486039),
	.w7(32'hbd2316d8),
	.w8(32'hbb701569),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2437b),
	.w1(32'hbc333da9),
	.w2(32'h3cb2c4af),
	.w3(32'hbc2c757a),
	.w4(32'hbbb69b3c),
	.w5(32'h3a8f23a4),
	.w6(32'hbb5fe14d),
	.w7(32'hbca971d8),
	.w8(32'hbb56bb94),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58d3a9),
	.w1(32'hbc456a15),
	.w2(32'h3cc22d85),
	.w3(32'hbc5cf093),
	.w4(32'hbbbe0ae9),
	.w5(32'h3b386926),
	.w6(32'hbbb8d30d),
	.w7(32'hbcb52bda),
	.w8(32'hbb40d6ad),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd16b3d),
	.w1(32'hbc5f5428),
	.w2(32'hbc5acfcb),
	.w3(32'hbc792c12),
	.w4(32'hba5fe09b),
	.w5(32'hbaf01ced),
	.w6(32'hbb9c8c5b),
	.w7(32'hbaab2521),
	.w8(32'h3b9fea82),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc578907),
	.w1(32'h3ba1e0fc),
	.w2(32'hbbacb5af),
	.w3(32'hbbd27000),
	.w4(32'hbbab0a15),
	.w5(32'hbb163343),
	.w6(32'h3c3b0c38),
	.w7(32'h3d1fcb0d),
	.w8(32'h3b58430e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc084675),
	.w1(32'hbb804440),
	.w2(32'h3c1ce0d4),
	.w3(32'hbbbbaff7),
	.w4(32'hbc16cb16),
	.w5(32'hbbdeeb9d),
	.w6(32'h3bc8010b),
	.w7(32'h3b5bc948),
	.w8(32'h3c3f6a2f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b964452),
	.w1(32'hbb0e3bd4),
	.w2(32'h3bbfd1ea),
	.w3(32'hbc439f57),
	.w4(32'hbbaa5339),
	.w5(32'hba9701e9),
	.w6(32'h3b3605f8),
	.w7(32'h3b7ac5b8),
	.w8(32'h3c5d6f0e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9613e6),
	.w1(32'hbc0c7570),
	.w2(32'h3cca94f5),
	.w3(32'hb9c1d1fd),
	.w4(32'hbbc6ba55),
	.w5(32'h3aa4bb15),
	.w6(32'hba620e60),
	.w7(32'hbcb61d28),
	.w8(32'hbb7ba435),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb961f73),
	.w1(32'hbc08fa9e),
	.w2(32'hbb987fec),
	.w3(32'hbc8020d6),
	.w4(32'h3baaa1ff),
	.w5(32'h3c0b37db),
	.w6(32'h3a1aa737),
	.w7(32'h3aead060),
	.w8(32'h399a3758),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0c19d),
	.w1(32'hbbfb8b8d),
	.w2(32'h3c5b877b),
	.w3(32'h3bea5a79),
	.w4(32'hbb9ed888),
	.w5(32'hbab9a6d4),
	.w6(32'h3b9a42ed),
	.w7(32'h3b85ec89),
	.w8(32'h3c46e4de),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86994c),
	.w1(32'hbc8e3d31),
	.w2(32'hb9f529c2),
	.w3(32'hbc448e25),
	.w4(32'hbc382de5),
	.w5(32'hbb26cd32),
	.w6(32'hbcaafd12),
	.w7(32'hbcb9a563),
	.w8(32'hbbef324e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc031103),
	.w1(32'hb9b31aca),
	.w2(32'hb9ddd43a),
	.w3(32'hbc05b63f),
	.w4(32'hb9c48e0d),
	.w5(32'hba0a0642),
	.w6(32'hb9372bf9),
	.w7(32'hb9c2ec26),
	.w8(32'hb8b04d4b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30779e),
	.w1(32'h39009a7d),
	.w2(32'h3ae9f483),
	.w3(32'h3aa8c0f4),
	.w4(32'h3b3b17f0),
	.w5(32'h38a23171),
	.w6(32'hbb2e13b6),
	.w7(32'h3a1adbf5),
	.w8(32'hba39e708),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule