module layer_8_featuremap_233(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1db83),
	.w1(32'h3c0d85c5),
	.w2(32'hba974627),
	.w3(32'h3b56b09f),
	.w4(32'h3b980dd1),
	.w5(32'h3c41664a),
	.w6(32'h3bc68fd7),
	.w7(32'h395eb186),
	.w8(32'h3bc6d35e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c9ccf),
	.w1(32'hbb4458be),
	.w2(32'hbb3ecd53),
	.w3(32'h3c18b65a),
	.w4(32'hbb4ae7cd),
	.w5(32'hbbd847f6),
	.w6(32'hbb87f1cc),
	.w7(32'hbb7472dd),
	.w8(32'hbaf249d0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ec5cd),
	.w1(32'h3bc8ab8c),
	.w2(32'h3bf554b2),
	.w3(32'hbb44286b),
	.w4(32'h3bae38be),
	.w5(32'h3bd182c5),
	.w6(32'hbb30ba00),
	.w7(32'h3bd87caa),
	.w8(32'h3a91dc47),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83cf30),
	.w1(32'h3bc6d079),
	.w2(32'h3c31fa9b),
	.w3(32'h3bc02dd7),
	.w4(32'hbc43f3e8),
	.w5(32'h39538cf3),
	.w6(32'h3aa1d1c2),
	.w7(32'h3b4d4a3d),
	.w8(32'h3c36094d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88d828),
	.w1(32'h3bd81623),
	.w2(32'h3bb1e660),
	.w3(32'h3c088ae3),
	.w4(32'h3b70f2f5),
	.w5(32'h3ae1f4b2),
	.w6(32'h3ae6eef8),
	.w7(32'h3abfc2f9),
	.w8(32'h3b15eae4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c667266),
	.w1(32'h3c4fccf9),
	.w2(32'h3c0bf0d9),
	.w3(32'h3c00f21d),
	.w4(32'h3c2a01ce),
	.w5(32'h3bc511fc),
	.w6(32'h3c2f747a),
	.w7(32'h3c24c853),
	.w8(32'hbbdef0c7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa90d90),
	.w1(32'hbab8e6df),
	.w2(32'hbb292919),
	.w3(32'h3b3d882d),
	.w4(32'hba57b2b6),
	.w5(32'h3ab0dd2f),
	.w6(32'hbb08035a),
	.w7(32'hba814367),
	.w8(32'hbb9e7a0c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc85026),
	.w1(32'hbc179375),
	.w2(32'hbb8f8dc1),
	.w3(32'hbacba542),
	.w4(32'hbc519a8d),
	.w5(32'h3b8cf128),
	.w6(32'hbcd5cb17),
	.w7(32'hbc03db6a),
	.w8(32'hbc4a7f80),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3347e),
	.w1(32'hbc233c90),
	.w2(32'hbb51a956),
	.w3(32'hbb7b7bf5),
	.w4(32'hbc4a7a5a),
	.w5(32'hbc294321),
	.w6(32'hbc736487),
	.w7(32'hbc1cc713),
	.w8(32'hbbce8ff2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc05150),
	.w1(32'hbb96edcd),
	.w2(32'h3bd1e1af),
	.w3(32'hbc2451cf),
	.w4(32'h3801411b),
	.w5(32'h3bc82730),
	.w6(32'hbb311aa3),
	.w7(32'hbb1b8e6a),
	.w8(32'h3a8c9ead),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc77445),
	.w1(32'hbc6ebda1),
	.w2(32'h3b6591cd),
	.w3(32'h3b0908a1),
	.w4(32'hbc97784d),
	.w5(32'hbbc35330),
	.w6(32'hbc128b74),
	.w7(32'hbbba1511),
	.w8(32'hbbd1f1a1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b177978),
	.w1(32'h3b36368e),
	.w2(32'h39f05d6e),
	.w3(32'hbacabce1),
	.w4(32'h3b8c29f8),
	.w5(32'h39ed6bd3),
	.w6(32'h3b8c327b),
	.w7(32'h3b52f52e),
	.w8(32'h39449e7c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc9507),
	.w1(32'hbab29073),
	.w2(32'hbba25091),
	.w3(32'h3b8f56cc),
	.w4(32'hbc12fa62),
	.w5(32'hbc43faf3),
	.w6(32'hbb3e1abb),
	.w7(32'hbc0cdc05),
	.w8(32'hbb19f0e5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc539760),
	.w1(32'h3b5f3f71),
	.w2(32'h3bdc7cc5),
	.w3(32'hbc3de815),
	.w4(32'h3c0399d4),
	.w5(32'h3c49b585),
	.w6(32'hb7a4d57e),
	.w7(32'hbaee1e64),
	.w8(32'h3ba1b2ed),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c665f15),
	.w1(32'hba0095e3),
	.w2(32'h3b02b7b2),
	.w3(32'h3c087d97),
	.w4(32'hbae558e8),
	.w5(32'h3b26fc99),
	.w6(32'h396e1510),
	.w7(32'h3ae1e8dc),
	.w8(32'hbb95f1ea),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb927346),
	.w1(32'h3c1558ed),
	.w2(32'h3a7c2119),
	.w3(32'hbb85d529),
	.w4(32'hbaea42ee),
	.w5(32'hbb522891),
	.w6(32'h3be7091e),
	.w7(32'h3b287054),
	.w8(32'h3b293208),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb636da4),
	.w1(32'hbc239484),
	.w2(32'hbc920b8e),
	.w3(32'hb9f40314),
	.w4(32'hbcb37979),
	.w5(32'hbced5e76),
	.w6(32'hbc5503b4),
	.w7(32'hbcb5c30b),
	.w8(32'hbc218597),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd013b4),
	.w1(32'hbd13cde6),
	.w2(32'hbd5996b2),
	.w3(32'hbc7600e6),
	.w4(32'hbcaa5b6f),
	.w5(32'hbd3954c0),
	.w6(32'hbc91801e),
	.w7(32'hbcee5677),
	.w8(32'hbc686674),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd386684),
	.w1(32'hbb9a3345),
	.w2(32'hbb81b128),
	.w3(32'hbca1412b),
	.w4(32'hbb52558e),
	.w5(32'h3c0a3a66),
	.w6(32'hbabc4f14),
	.w7(32'hbc1ee78b),
	.w8(32'h3b9e7e64),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5134d8),
	.w1(32'hbb8beaf4),
	.w2(32'hbb5ad45d),
	.w3(32'hbbcedd3c),
	.w4(32'hba3d1c49),
	.w5(32'h3a4acb6d),
	.w6(32'hba54d37f),
	.w7(32'hbb3c15de),
	.w8(32'hbb7d8c5d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79db6e),
	.w1(32'h3c24823e),
	.w2(32'h3cd87f1d),
	.w3(32'h3c1452cc),
	.w4(32'h3bef95ff),
	.w5(32'h3c607a6e),
	.w6(32'h3bdffdc9),
	.w7(32'h3c9be72b),
	.w8(32'h3bf75d2e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bfeca),
	.w1(32'h3d0d6566),
	.w2(32'h3d427530),
	.w3(32'h3c4266ab),
	.w4(32'h3cf627a0),
	.w5(32'h3d2ccbc0),
	.w6(32'h3c4812b3),
	.w7(32'h3cc909ae),
	.w8(32'h3ca9381d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce3993e),
	.w1(32'h3aa0e2f7),
	.w2(32'h3baace51),
	.w3(32'h3cc92651),
	.w4(32'hbaf67b3d),
	.w5(32'h3b925b56),
	.w6(32'h3c12e581),
	.w7(32'h3b6663cb),
	.w8(32'h3c746435),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac8078),
	.w1(32'h3d2fb4a1),
	.w2(32'h3d80614f),
	.w3(32'hbb7a1dac),
	.w4(32'h3d1dfe36),
	.w5(32'h3d5e4b72),
	.w6(32'h3c703147),
	.w7(32'h3cf80175),
	.w8(32'h3c8beb3b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d16de0b),
	.w1(32'hbb168d7b),
	.w2(32'h3bf47c34),
	.w3(32'h3cd296cf),
	.w4(32'h3b861040),
	.w5(32'h3b9c4084),
	.w6(32'h3bd1a9cc),
	.w7(32'h3bb23dc0),
	.w8(32'h3a23cf2f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1de504),
	.w1(32'h3bb86f27),
	.w2(32'h3c96a0d4),
	.w3(32'h3c2aceb7),
	.w4(32'h3c02f597),
	.w5(32'h3c38071b),
	.w6(32'h3b4bb1d9),
	.w7(32'h3bef4ee5),
	.w8(32'h3ba22385),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2cc5b),
	.w1(32'hbb22efbe),
	.w2(32'h3b24e26c),
	.w3(32'h3af97518),
	.w4(32'hbbacc661),
	.w5(32'h3b1bbcec),
	.w6(32'hb9a34691),
	.w7(32'hbb15af5b),
	.w8(32'h398c8779),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f35e0),
	.w1(32'hbd18f0f2),
	.w2(32'hbc817d3c),
	.w3(32'hbbd4c5e4),
	.w4(32'hbcf1305b),
	.w5(32'hbcf5520f),
	.w6(32'hbcce2bd7),
	.w7(32'hbba7c702),
	.w8(32'h3babe2e5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00894f),
	.w1(32'h39631c72),
	.w2(32'h3bd92251),
	.w3(32'hbc959b9d),
	.w4(32'h39b2dad7),
	.w5(32'h3abb770e),
	.w6(32'hbb90d9a1),
	.w7(32'h3a9bc497),
	.w8(32'hb9e687fd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80a9c7),
	.w1(32'h3bbf1846),
	.w2(32'h3bc02ba9),
	.w3(32'h3bae267e),
	.w4(32'h3b4f246e),
	.w5(32'h3bf1e777),
	.w6(32'hbb3366b4),
	.w7(32'h392ca590),
	.w8(32'h3a4835b8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f78f3),
	.w1(32'h3bd8114b),
	.w2(32'h3c066415),
	.w3(32'h3b7885d1),
	.w4(32'h3b02d438),
	.w5(32'h3c0a0485),
	.w6(32'h3b802710),
	.w7(32'h3b0b2cd7),
	.w8(32'hbbd679ab),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab635aa),
	.w1(32'h3c513bc4),
	.w2(32'h3cac7911),
	.w3(32'h3be3a94d),
	.w4(32'h39a4d15f),
	.w5(32'h3bf2640c),
	.w6(32'hba54ce2a),
	.w7(32'h39ed757b),
	.w8(32'hbc16855d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb9db8),
	.w1(32'hbcdbc9bf),
	.w2(32'hbcfb99bd),
	.w3(32'hb9d5909f),
	.w4(32'hbc43b61d),
	.w5(32'hbc0d0f15),
	.w6(32'hbc2b4903),
	.w7(32'hbc80cfd5),
	.w8(32'hba732c76),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6dde09),
	.w1(32'hbd1d8021),
	.w2(32'hbd78522a),
	.w3(32'hbc22aaf3),
	.w4(32'hbca5a400),
	.w5(32'hbd19191c),
	.w6(32'hbcc6ac45),
	.w7(32'hbd23924a),
	.w8(32'hbcc45e94),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2d1654),
	.w1(32'hb9c7a84a),
	.w2(32'h3a3dd655),
	.w3(32'hbce1437f),
	.w4(32'hbb908d7a),
	.w5(32'h3b7c4be2),
	.w6(32'h3baa9330),
	.w7(32'h3bd45dfd),
	.w8(32'hbad598d3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f6e0f),
	.w1(32'hbbe4c6fa),
	.w2(32'h3c4cca5c),
	.w3(32'hbbe846a8),
	.w4(32'hbbc1eb09),
	.w5(32'h3c971be1),
	.w6(32'hbba48a91),
	.w7(32'h3bc7d323),
	.w8(32'hba83a7f1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e2859),
	.w1(32'h3b96bf0b),
	.w2(32'h3b8715af),
	.w3(32'h3c23e607),
	.w4(32'h3b49b88a),
	.w5(32'h3b746285),
	.w6(32'h3b487c58),
	.w7(32'h3ade9cd2),
	.w8(32'h3bc15228),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ffa45),
	.w1(32'h3bab8ee4),
	.w2(32'h3bed7819),
	.w3(32'h3b57a9df),
	.w4(32'h3946dea6),
	.w5(32'h3ba1c5d1),
	.w6(32'hb9a31633),
	.w7(32'h3b19104c),
	.w8(32'h3b788982),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbee528),
	.w1(32'h3cae6fc1),
	.w2(32'h3d1ec30b),
	.w3(32'h3ae554e5),
	.w4(32'h3ca70eae),
	.w5(32'h3ccfed1e),
	.w6(32'h3c60a860),
	.w7(32'h3c9ac0f8),
	.w8(32'h3c0eb554),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc7c139),
	.w1(32'h3bfaeaf2),
	.w2(32'h3c8c1090),
	.w3(32'h3cc3e10d),
	.w4(32'h3a84b13e),
	.w5(32'h3c64d79f),
	.w6(32'hbb8052b1),
	.w7(32'h39e137ad),
	.w8(32'hbaa188de),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9608cf),
	.w1(32'h3b41a8dc),
	.w2(32'h3c4bef3b),
	.w3(32'h3bb23bc3),
	.w4(32'h3b3dcfd5),
	.w5(32'h3c184834),
	.w6(32'h3be66cfe),
	.w7(32'h3c883d42),
	.w8(32'h3c05d1bb),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2ac8a),
	.w1(32'hbbd0a66c),
	.w2(32'hb98407f2),
	.w3(32'h3ad9a91a),
	.w4(32'hbc023d37),
	.w5(32'h3b94e349),
	.w6(32'hbc23c19d),
	.w7(32'hbc361492),
	.w8(32'hbb6c36d0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6e9c2),
	.w1(32'hba05d1cb),
	.w2(32'h3bfa2839),
	.w3(32'h3b3fb8ad),
	.w4(32'h3a93731c),
	.w5(32'h3a49e639),
	.w6(32'hbb03f0d4),
	.w7(32'h3c45d0b4),
	.w8(32'h3c5061c3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11ca8c),
	.w1(32'hbd014b08),
	.w2(32'hbd9806f9),
	.w3(32'h3ba7f006),
	.w4(32'hbca90b81),
	.w5(32'hbd5ad3fb),
	.w6(32'hbb9c466a),
	.w7(32'hbd0bd618),
	.w8(32'hbcec7bfc),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4fa8f6),
	.w1(32'h3b1ac3da),
	.w2(32'h3d108b71),
	.w3(32'hbca4b03e),
	.w4(32'hbc37f5c5),
	.w5(32'h3c96b921),
	.w6(32'hba3fbf51),
	.w7(32'h3c647c80),
	.w8(32'h3c55b744),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb57a8d),
	.w1(32'hbbd8f485),
	.w2(32'hbbb88ce4),
	.w3(32'h3c360e46),
	.w4(32'hbb29926e),
	.w5(32'hba5971cd),
	.w6(32'h3a9b9b7c),
	.w7(32'hbb449fbd),
	.w8(32'hbb95870e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb44df),
	.w1(32'h3c22bd88),
	.w2(32'h3ca1a4bb),
	.w3(32'hbaddfc44),
	.w4(32'h3c5db6f5),
	.w5(32'h3c52cb2a),
	.w6(32'h3b7ec9d1),
	.w7(32'h3c18fc6c),
	.w8(32'hbb3341a2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf0451),
	.w1(32'hbc932004),
	.w2(32'hbc085447),
	.w3(32'h3ad293f8),
	.w4(32'hbb65f43e),
	.w5(32'hbb94fc59),
	.w6(32'hbbb67a0a),
	.w7(32'hbc53fcd3),
	.w8(32'hbc003219),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7adb15),
	.w1(32'hbc35ee00),
	.w2(32'hbc8b283e),
	.w3(32'h3ba3f9ed),
	.w4(32'hbc176153),
	.w5(32'hbba4ec2b),
	.w6(32'hbc1ccd96),
	.w7(32'hbc57e516),
	.w8(32'hbc1057dd),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e4a68),
	.w1(32'hbb8018c6),
	.w2(32'hbcd4a8a2),
	.w3(32'hbc41800a),
	.w4(32'hbb39c47d),
	.w5(32'hbc6de4d4),
	.w6(32'hbc78f697),
	.w7(32'hbb8a060d),
	.w8(32'hbb5316fd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd29636),
	.w1(32'h3c08d218),
	.w2(32'h3c592ad4),
	.w3(32'hba02f0eb),
	.w4(32'h3c35d99d),
	.w5(32'h3bc6d77d),
	.w6(32'h3bf10eea),
	.w7(32'h3c5f024e),
	.w8(32'h3ba7e355),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76120b),
	.w1(32'h3bec6553),
	.w2(32'h3ca37f91),
	.w3(32'hb93a747d),
	.w4(32'h3ac31a6e),
	.w5(32'h3cba82a4),
	.w6(32'h3a9a15af),
	.w7(32'h3b96fa53),
	.w8(32'h3c47b4cd),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c483f87),
	.w1(32'hbaaccead),
	.w2(32'hb958e33d),
	.w3(32'h3b7ac437),
	.w4(32'hbb89ff23),
	.w5(32'hbb5520b9),
	.w6(32'hbb360c8b),
	.w7(32'hbada0344),
	.w8(32'hbb4ecafb),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68f370),
	.w1(32'h3b3c11b6),
	.w2(32'h3c050e34),
	.w3(32'hbc2a277d),
	.w4(32'h3b8bc561),
	.w5(32'h3b7a3640),
	.w6(32'h3b533e64),
	.w7(32'h3c2011a6),
	.w8(32'h3c10c293),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1103fa),
	.w1(32'hbbdbe412),
	.w2(32'hbcd1bb19),
	.w3(32'hbb9a0eae),
	.w4(32'hbb895236),
	.w5(32'hbc40a2ec),
	.w6(32'hbbc1a31f),
	.w7(32'hbc7a31d2),
	.w8(32'hbc55d5ef),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf776d8),
	.w1(32'hbd26402e),
	.w2(32'hbd7e28a8),
	.w3(32'hbc0cba38),
	.w4(32'hbc904da9),
	.w5(32'hbd3ca58c),
	.w6(32'hbcbab8b6),
	.w7(32'hbd09748b),
	.w8(32'hbc93cfdb),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4e7be6),
	.w1(32'h3c094e74),
	.w2(32'h3c143e1e),
	.w3(32'hbd1a9f0e),
	.w4(32'h3c0c9ea5),
	.w5(32'hbb10cc43),
	.w6(32'h3c1b7689),
	.w7(32'h3beac338),
	.w8(32'h3c373e3a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe5e8a),
	.w1(32'hba28070e),
	.w2(32'h3b7fb3b3),
	.w3(32'hbaa2a851),
	.w4(32'hbb9bb6fd),
	.w5(32'h3b4a2cbd),
	.w6(32'hbb8b7e5d),
	.w7(32'hbb5a1357),
	.w8(32'hbb5db522),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cbd66),
	.w1(32'hbba766e1),
	.w2(32'h3aad4ed2),
	.w3(32'hbbdc8663),
	.w4(32'hbb9f3485),
	.w5(32'hbb2ba1e3),
	.w6(32'hbb4bb72b),
	.w7(32'hbb65fa80),
	.w8(32'hbab20499),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cf3e5),
	.w1(32'h3d06a07e),
	.w2(32'h3d66d7ab),
	.w3(32'hbb343b57),
	.w4(32'h3d054026),
	.w5(32'h3d452093),
	.w6(32'h3c52f6fe),
	.w7(32'h3d01b624),
	.w8(32'h3cd524fb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1c38d4),
	.w1(32'hbc006679),
	.w2(32'hbc4eb258),
	.w3(32'h3cdf35a1),
	.w4(32'h3ac129aa),
	.w5(32'hbc044aff),
	.w6(32'hbb481a21),
	.w7(32'hbb0296f9),
	.w8(32'hbc088930),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0291b3),
	.w1(32'h3b4d02c8),
	.w2(32'h3bd2aa52),
	.w3(32'hbbb1248c),
	.w4(32'h3b8e3aeb),
	.w5(32'h3c488712),
	.w6(32'hbc0b418c),
	.w7(32'hbc3d0370),
	.w8(32'hbc4430f8),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a530c43),
	.w1(32'h3aabaae1),
	.w2(32'h3bf05416),
	.w3(32'h3b91a39c),
	.w4(32'hbbfcd1b2),
	.w5(32'h3be39b9d),
	.w6(32'hbba17b75),
	.w7(32'h3a2630b8),
	.w8(32'h38d26442),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf602bb),
	.w1(32'h3b1bc174),
	.w2(32'h3b2ba150),
	.w3(32'h3c14052c),
	.w4(32'h3b0f9522),
	.w5(32'h3a779f24),
	.w6(32'h3b7eafbd),
	.w7(32'h3b87586f),
	.w8(32'h3bc10fc0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fdaa0),
	.w1(32'hb946570d),
	.w2(32'h3ac2504c),
	.w3(32'h39a48834),
	.w4(32'hbc0d5f41),
	.w5(32'hbacd8b24),
	.w6(32'hbb618bc4),
	.w7(32'hbaccec53),
	.w8(32'hbbacbe07),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31e422),
	.w1(32'h3bb7e7e3),
	.w2(32'h3cb6ca39),
	.w3(32'hbb42a8ba),
	.w4(32'h3b9026f8),
	.w5(32'h3c724d80),
	.w6(32'hbbc498e2),
	.w7(32'hbbe5805a),
	.w8(32'h39ce7c55),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fdaeb),
	.w1(32'hbb496d97),
	.w2(32'h3c3a1792),
	.w3(32'h3c0cfd0b),
	.w4(32'hbb51905a),
	.w5(32'hbb51e7c1),
	.w6(32'h3c3bc422),
	.w7(32'h3c504897),
	.w8(32'h3c389ae0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91c650),
	.w1(32'h3c3314a5),
	.w2(32'h3c187e34),
	.w3(32'h3b0a7f82),
	.w4(32'h3c4a7ca1),
	.w5(32'h3af27b22),
	.w6(32'h3aec7590),
	.w7(32'h3b97d667),
	.w8(32'h3b245212),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19fa22),
	.w1(32'hbcd4d897),
	.w2(32'hbd4d00be),
	.w3(32'hbbcde61a),
	.w4(32'hbbf410ed),
	.w5(32'hbcae880d),
	.w6(32'hbc9a04ab),
	.w7(32'hbcdaf12b),
	.w8(32'hbc565575),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd26b30d),
	.w1(32'h3ba6860a),
	.w2(32'h3c09d8ff),
	.w3(32'hbcb8f949),
	.w4(32'hba9662cb),
	.w5(32'h3c8fea2c),
	.w6(32'h3beed0bf),
	.w7(32'h3bbc9348),
	.w8(32'h3c694897),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfc025),
	.w1(32'hbbb422d8),
	.w2(32'h3b8cbaa2),
	.w3(32'h3b7126a5),
	.w4(32'hbb1e3e66),
	.w5(32'h3b07b07c),
	.w6(32'hbbf81663),
	.w7(32'h3bb2515e),
	.w8(32'h3ba674a1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f5c21),
	.w1(32'h3cf404f0),
	.w2(32'h3d380aac),
	.w3(32'h3bc3945d),
	.w4(32'h3c8c0070),
	.w5(32'h3ce837dc),
	.w6(32'h3c70affe),
	.w7(32'h3cd5388c),
	.w8(32'h3ccb46dd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd1512d),
	.w1(32'h3c2d823e),
	.w2(32'h3d13075b),
	.w3(32'h3c8d8c31),
	.w4(32'h3c638c0d),
	.w5(32'h3cfc7d31),
	.w6(32'h3ae0246a),
	.w7(32'h3c6c897b),
	.w8(32'h3c52bd81),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd0c447),
	.w1(32'hbc2e8b90),
	.w2(32'hbb8a22bf),
	.w3(32'h3c84905d),
	.w4(32'hbc43feff),
	.w5(32'hbc286044),
	.w6(32'hbc2c68ef),
	.w7(32'hbbc3a2b4),
	.w8(32'hbc104704),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc286edc),
	.w1(32'hbb165906),
	.w2(32'h3c121b01),
	.w3(32'hbba5a2fa),
	.w4(32'h3b2d5143),
	.w5(32'h3bd9544a),
	.w6(32'h3c005d3d),
	.w7(32'h3b9976a2),
	.w8(32'h3b17d77f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a88d3),
	.w1(32'hb99e211b),
	.w2(32'h396f9fce),
	.w3(32'h3b6b94c6),
	.w4(32'h3ac59a82),
	.w5(32'hbb52b48a),
	.w6(32'h3be895ad),
	.w7(32'h3aa31b61),
	.w8(32'h3bc73b43),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c078618),
	.w1(32'hbb2d6ce7),
	.w2(32'h3a9d1a11),
	.w3(32'h3b507f9d),
	.w4(32'h3b3c3988),
	.w5(32'h3bb2b7bd),
	.w6(32'hbbf0a6f8),
	.w7(32'h39b1412f),
	.w8(32'h3a67f0fa),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd2607),
	.w1(32'hbb1a8763),
	.w2(32'h3b8f82f2),
	.w3(32'h3c02b22b),
	.w4(32'h38846884),
	.w5(32'h3b1fb1ca),
	.w6(32'hbbe3af32),
	.w7(32'hbb2a31f9),
	.w8(32'h3c156617),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b839bfb),
	.w1(32'hbc7951ef),
	.w2(32'hbbb6d207),
	.w3(32'h3b1fb7e3),
	.w4(32'hbbd46538),
	.w5(32'hbb9cf228),
	.w6(32'hbbf693fa),
	.w7(32'hba0068b2),
	.w8(32'h3bf6eaf0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad250d),
	.w1(32'hbd3e01dc),
	.w2(32'hbd6ce294),
	.w3(32'h3b93d5b4),
	.w4(32'hbd0a8233),
	.w5(32'hbd367300),
	.w6(32'hbcab7f82),
	.w7(32'hbd1bc98b),
	.w8(32'hbc8942b3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0a6132),
	.w1(32'h3b961b9c),
	.w2(32'h3bff5ced),
	.w3(32'hbcd090bc),
	.w4(32'h3b9b3013),
	.w5(32'h3c293755),
	.w6(32'hb8a92ee9),
	.w7(32'h3be60e2a),
	.w8(32'h3c3d14bb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5e10f),
	.w1(32'hbce31689),
	.w2(32'hbd21c839),
	.w3(32'h3b9b1fef),
	.w4(32'hbb920175),
	.w5(32'hbc839e9b),
	.w6(32'hbc718fbf),
	.w7(32'hbcf29c66),
	.w8(32'hbc4a4e1a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcace585),
	.w1(32'h3afa0dbe),
	.w2(32'hbb65c0ec),
	.w3(32'hbc3a5e82),
	.w4(32'hbb583fdc),
	.w5(32'hba20fce0),
	.w6(32'h3b700a40),
	.w7(32'hb9638ee9),
	.w8(32'hbaea6e8d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ca18b),
	.w1(32'h3bcde040),
	.w2(32'h3bb56530),
	.w3(32'hb71fae8c),
	.w4(32'h3ac41f99),
	.w5(32'h394f7f8e),
	.w6(32'hbb912f9f),
	.w7(32'h3bb7f8a6),
	.w8(32'hba355b2d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c0286),
	.w1(32'hbbbfbf00),
	.w2(32'h3a925889),
	.w3(32'hbb32e353),
	.w4(32'hbc2fe0f7),
	.w5(32'h3c0ae3de),
	.w6(32'h3b1630a8),
	.w7(32'h3be8a1fe),
	.w8(32'h3c3dea87),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a8397),
	.w1(32'hbae3a47c),
	.w2(32'hbc76b8fc),
	.w3(32'h3b95d925),
	.w4(32'hbc4941ef),
	.w5(32'hba8892ec),
	.w6(32'h3b882786),
	.w7(32'hbc5ab633),
	.w8(32'hbc08ac0d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1babfa),
	.w1(32'hbbbb967d),
	.w2(32'hbb9935b1),
	.w3(32'h3a9d19a9),
	.w4(32'hbb9975d6),
	.w5(32'hbb956477),
	.w6(32'hbad8c777),
	.w7(32'hbae7e84e),
	.w8(32'hb89dcd4e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a265ddb),
	.w1(32'hbbe65124),
	.w2(32'hb9833929),
	.w3(32'h3ab04178),
	.w4(32'hbc4bbceb),
	.w5(32'hb90a79b4),
	.w6(32'hbbe7ced7),
	.w7(32'hbab614bf),
	.w8(32'hba2ed957),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae025d7),
	.w1(32'hbaa41661),
	.w2(32'h39a7a33c),
	.w3(32'h3aa652f5),
	.w4(32'hb9479e3b),
	.w5(32'h3aa04136),
	.w6(32'hba86544d),
	.w7(32'hbb6cb3ba),
	.w8(32'hbb934f20),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cc8b1),
	.w1(32'hbb3d57b3),
	.w2(32'hbb305bc8),
	.w3(32'h3b865553),
	.w4(32'hb9c857ae),
	.w5(32'h3ba2b793),
	.w6(32'hbb696c3d),
	.w7(32'hbae02447),
	.w8(32'h3c2511e6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc362d),
	.w1(32'h3cafa3ab),
	.w2(32'h3d488669),
	.w3(32'h3c0a094b),
	.w4(32'h3ca1303a),
	.w5(32'h3d093f57),
	.w6(32'h3bca09a6),
	.w7(32'h3cafb8a6),
	.w8(32'h3c94b960),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0ab5b7),
	.w1(32'hbc53fc6b),
	.w2(32'hbd3e7db1),
	.w3(32'h3c966b8e),
	.w4(32'hbc368cab),
	.w5(32'hbd0aeaec),
	.w6(32'hbc0f61d2),
	.w7(32'hbcf566db),
	.w8(32'hbc8c2338),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0fee09),
	.w1(32'h3b4d8517),
	.w2(32'h3af3c377),
	.w3(32'hbd057f32),
	.w4(32'h3a114c6a),
	.w5(32'hba1fa93c),
	.w6(32'h3bd9f715),
	.w7(32'h3b4b974e),
	.w8(32'h3b3edb04),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba657bf1),
	.w1(32'hbb21457b),
	.w2(32'h3a8e12db),
	.w3(32'h3b3282ec),
	.w4(32'h38df8c60),
	.w5(32'hba8b297b),
	.w6(32'hbb027628),
	.w7(32'hbb1aa1fb),
	.w8(32'hbb66e584),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf33b6b),
	.w1(32'hbb004bdc),
	.w2(32'hbbd10134),
	.w3(32'hbb0d5919),
	.w4(32'h3c23f827),
	.w5(32'h3c04195b),
	.w6(32'hbba498ef),
	.w7(32'hbbc464f4),
	.w8(32'hbc31d435),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38fc5e),
	.w1(32'hbbabd39b),
	.w2(32'hbba5455f),
	.w3(32'h39df470d),
	.w4(32'hbb492e05),
	.w5(32'hbb05530e),
	.w6(32'hbb361a22),
	.w7(32'hbbb54173),
	.w8(32'hbbe378d3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83685e),
	.w1(32'h3c61a68e),
	.w2(32'h3ca1966b),
	.w3(32'hbba357f3),
	.w4(32'h3c85f4d6),
	.w5(32'h3ca6280a),
	.w6(32'h3c69b190),
	.w7(32'h3c9e029f),
	.w8(32'h3c0e4894),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84c559),
	.w1(32'h3c313479),
	.w2(32'hbb24064a),
	.w3(32'h3c4abcf7),
	.w4(32'h3b983aff),
	.w5(32'hbb05e1d7),
	.w6(32'h399f98c7),
	.w7(32'h3afb9373),
	.w8(32'hba8481b0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89cc5f),
	.w1(32'hb98eecbc),
	.w2(32'hbc2253e0),
	.w3(32'h38e59991),
	.w4(32'hbb5845b3),
	.w5(32'hbc5883e4),
	.w6(32'h3bac9db5),
	.w7(32'h3b5464e6),
	.w8(32'hbacf4307),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd9af8),
	.w1(32'hbc8229e9),
	.w2(32'hbb748600),
	.w3(32'hbb127e3d),
	.w4(32'h3b1912ad),
	.w5(32'hbb10639e),
	.w6(32'h3b241c6b),
	.w7(32'h3a4fb744),
	.w8(32'h3bdbc783),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07de4),
	.w1(32'hbc3f10a2),
	.w2(32'hba4e7857),
	.w3(32'h3ac660bc),
	.w4(32'hbb4a49db),
	.w5(32'hbad3f079),
	.w6(32'hbba381b1),
	.w7(32'hbbaa50e0),
	.w8(32'h3bac628c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c154541),
	.w1(32'h3aeb52e3),
	.w2(32'h3c0182ce),
	.w3(32'h3c3cf9d6),
	.w4(32'hbbdca3cf),
	.w5(32'hba901d9f),
	.w6(32'hba66966d),
	.w7(32'hbb7114aa),
	.w8(32'hbbcebd20),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee5d14),
	.w1(32'h3bc975fe),
	.w2(32'hbc3adc62),
	.w3(32'hbbc114db),
	.w4(32'h3c0b8c09),
	.w5(32'h3badd6e0),
	.w6(32'h3be7ceb8),
	.w7(32'h3a848724),
	.w8(32'h3b597724),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f35c28),
	.w1(32'hbc3b9d36),
	.w2(32'hbba93e88),
	.w3(32'h3b9b8907),
	.w4(32'hbbacffc8),
	.w5(32'hbae3bef7),
	.w6(32'hbc174e4f),
	.w7(32'hbbddd929),
	.w8(32'h3a6fc969),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba92f5d),
	.w1(32'hb960a8a7),
	.w2(32'h3a9240a9),
	.w3(32'hbbdefcfe),
	.w4(32'h3ae430c8),
	.w5(32'h3b6e6f06),
	.w6(32'h3c8c6bb6),
	.w7(32'h3857040f),
	.w8(32'h3b6d73ef),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b677dfc),
	.w1(32'hbb9416e6),
	.w2(32'h3acf3928),
	.w3(32'h3b559972),
	.w4(32'hbb43417e),
	.w5(32'h3b77e90a),
	.w6(32'h3ae91cb7),
	.w7(32'h3b162e40),
	.w8(32'hbb9055b1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc89936),
	.w1(32'h3b0a5ca9),
	.w2(32'h3c568670),
	.w3(32'hbb4f03a8),
	.w4(32'h398704ac),
	.w5(32'h3b8d5a46),
	.w6(32'h3bc268b3),
	.w7(32'h3bb14375),
	.w8(32'h3bb67dfe),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb8808),
	.w1(32'hbbd0672c),
	.w2(32'hbc0a04ec),
	.w3(32'h3bb63793),
	.w4(32'hb9af3d21),
	.w5(32'hbbca9a99),
	.w6(32'hbb59bacf),
	.w7(32'hbbabae88),
	.w8(32'h3a4eed5e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5bd01),
	.w1(32'h3c0c4117),
	.w2(32'h3c85722c),
	.w3(32'h38f1a13d),
	.w4(32'h3be633ba),
	.w5(32'h3c2c5226),
	.w6(32'h39253e8e),
	.w7(32'h3b498d7f),
	.w8(32'h3abc6934),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b978e4f),
	.w1(32'h3b818718),
	.w2(32'h3bb40f61),
	.w3(32'h3ad59576),
	.w4(32'h3a61acdc),
	.w5(32'h3aa3a36f),
	.w6(32'hbb088aca),
	.w7(32'hbaeb4907),
	.w8(32'h3ad7634a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd609d),
	.w1(32'h3c84fc1c),
	.w2(32'h3c8cce68),
	.w3(32'h3aaee377),
	.w4(32'h3c2961ec),
	.w5(32'h3cba7464),
	.w6(32'h3c85c0f1),
	.w7(32'h3c60e2cd),
	.w8(32'h3c3aa38a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e161d),
	.w1(32'h3a3198b6),
	.w2(32'h3b951488),
	.w3(32'h3cc5a231),
	.w4(32'hbbb82e84),
	.w5(32'hba5e5d61),
	.w6(32'hbab079d6),
	.w7(32'hbae03a9f),
	.w8(32'hbc0da4ce),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28e881),
	.w1(32'hbc6906d0),
	.w2(32'hbcca500e),
	.w3(32'h3a685088),
	.w4(32'hbc2802b7),
	.w5(32'hbcceea08),
	.w6(32'hbc5c6df4),
	.w7(32'hbcdf115d),
	.w8(32'hbbe652ff),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87d46b),
	.w1(32'hbbd08edf),
	.w2(32'h3b8243d8),
	.w3(32'hbbc3533b),
	.w4(32'hbb8b1f66),
	.w5(32'hbbf78879),
	.w6(32'hbc420777),
	.w7(32'hbaa61900),
	.w8(32'h3c189a28),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36de15),
	.w1(32'hbb53ec59),
	.w2(32'hb9bb9287),
	.w3(32'hbc2bac47),
	.w4(32'hbc1ba66a),
	.w5(32'hbb7be603),
	.w6(32'h3856d875),
	.w7(32'h3b831423),
	.w8(32'h3a9d3a47),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82db53),
	.w1(32'h3b4dc53c),
	.w2(32'h3b6cbe1c),
	.w3(32'hb9520510),
	.w4(32'h38f0ea34),
	.w5(32'h3b268d8d),
	.w6(32'hba44e118),
	.w7(32'h3aa1e7d0),
	.w8(32'h3ae5df84),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb62a0a),
	.w1(32'hbb4f589b),
	.w2(32'h3b9406bd),
	.w3(32'h3b05b333),
	.w4(32'hba98733a),
	.w5(32'h3b53c494),
	.w6(32'h3a1a247e),
	.w7(32'h3b7c923d),
	.w8(32'h3b04bd84),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0106c2),
	.w1(32'hbc92a6bb),
	.w2(32'hbce665c2),
	.w3(32'h39e32c81),
	.w4(32'hbc53a0a4),
	.w5(32'hbcc4b71b),
	.w6(32'hbc553ebd),
	.w7(32'hbcc2377d),
	.w8(32'hbc2be50f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97527a),
	.w1(32'hbbd7af2c),
	.w2(32'hbcdb48eb),
	.w3(32'hbc869d5d),
	.w4(32'h3ba2a0f2),
	.w5(32'hbb841fe1),
	.w6(32'hbc848c59),
	.w7(32'hbca5a65f),
	.w8(32'hb982d77d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d0e00),
	.w1(32'hbb84db27),
	.w2(32'h38502af0),
	.w3(32'hbc6b22d9),
	.w4(32'hba529eed),
	.w5(32'hbb891ad9),
	.w6(32'h3a55a8cd),
	.w7(32'hbb12aa20),
	.w8(32'hbb739330),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63c4ef),
	.w1(32'hbce01262),
	.w2(32'hbd33b573),
	.w3(32'hbc4268e9),
	.w4(32'hbbf148cf),
	.w5(32'hbcce7eb4),
	.w6(32'hbcb321ce),
	.w7(32'hbcb6dc0c),
	.w8(32'hbc61c9a1),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1c101b),
	.w1(32'hbbc4fb47),
	.w2(32'hba80eb28),
	.w3(32'hbcf8cd9d),
	.w4(32'h3b1fc901),
	.w5(32'h3bb156dd),
	.w6(32'hb9be4eb5),
	.w7(32'hba6945e6),
	.w8(32'h3adca8f3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87470a),
	.w1(32'h3b8f01b1),
	.w2(32'h3b6baf1c),
	.w3(32'hbb3145ef),
	.w4(32'h3b6d3b77),
	.w5(32'h3a4b2649),
	.w6(32'h3b32cc8f),
	.w7(32'hb9cc534b),
	.w8(32'h3b4b0ed5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a0113),
	.w1(32'hbc295fc1),
	.w2(32'hbc056d98),
	.w3(32'h3ae03395),
	.w4(32'hbc20c22f),
	.w5(32'hbbfa8bab),
	.w6(32'hbbd313bb),
	.w7(32'hbc3cdaf3),
	.w8(32'hbb108fea),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac35899),
	.w1(32'h3c368214),
	.w2(32'h3c014bd4),
	.w3(32'h3a36f162),
	.w4(32'h3c91d9c6),
	.w5(32'h3be8e838),
	.w6(32'hbb5e1ac6),
	.w7(32'hbb0ff98c),
	.w8(32'h3c1bbe30),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d46e6),
	.w1(32'hbca051ed),
	.w2(32'hbc739ca8),
	.w3(32'hbb3ec706),
	.w4(32'hbc4775af),
	.w5(32'hbc373312),
	.w6(32'hbbe7eb99),
	.w7(32'hbc987b84),
	.w8(32'hbc2a1efd),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8156d8),
	.w1(32'h3a8a96d9),
	.w2(32'h3a5f15be),
	.w3(32'hb9006f5e),
	.w4(32'h3a664571),
	.w5(32'hbad531e2),
	.w6(32'hba4ae2b3),
	.w7(32'hbab8771c),
	.w8(32'h3a89ff4e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b690c09),
	.w1(32'hbab7ebc7),
	.w2(32'h3b3e8215),
	.w3(32'h3a8423d6),
	.w4(32'hbaffcae9),
	.w5(32'h3b7f9261),
	.w6(32'h392b2a3e),
	.w7(32'h3b2b935c),
	.w8(32'hba61459a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule