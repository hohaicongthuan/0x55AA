module layer_10_featuremap_392(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74d7265),
	.w1(32'h36026329),
	.w2(32'h37887b4e),
	.w3(32'hb7f49476),
	.w4(32'hb75eea35),
	.w5(32'h37620613),
	.w6(32'hb849ddfc),
	.w7(32'hb7d6a7e9),
	.w8(32'hb6b57f37),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba79a69),
	.w1(32'hbbee8570),
	.w2(32'hbbabab99),
	.w3(32'hbbc3a952),
	.w4(32'hbb76c36f),
	.w5(32'hbae4128a),
	.w6(32'hbae9d53d),
	.w7(32'h3aa06972),
	.w8(32'h3a40116d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71667b2),
	.w1(32'hb6bd50da),
	.w2(32'hb66524dc),
	.w3(32'hb7516c0f),
	.w4(32'hb6eff801),
	.w5(32'h3635afba),
	.w6(32'hb79b8742),
	.w7(32'hb73a451d),
	.w8(32'hb705a3e1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0af344),
	.w1(32'h3a39c71e),
	.w2(32'h3a89ff70),
	.w3(32'h398db56e),
	.w4(32'h3a56d41f),
	.w5(32'h3892799e),
	.w6(32'h38f74398),
	.w7(32'h3985017b),
	.w8(32'hb8a8c818),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ee60b),
	.w1(32'hb8a1dc60),
	.w2(32'h398e39a4),
	.w3(32'hb9ab5ac3),
	.w4(32'hb987090a),
	.w5(32'h37e78300),
	.w6(32'hb98f79af),
	.w7(32'hb96f1b93),
	.w8(32'hb8fc64c4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3790fe31),
	.w1(32'h383f9f40),
	.w2(32'h37d23763),
	.w3(32'hb7cf73d3),
	.w4(32'h37449eb9),
	.w5(32'h37016a3b),
	.w6(32'hb85dd47d),
	.w7(32'hb791fb3f),
	.w8(32'hb7d07d7e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18ac6f),
	.w1(32'hbb1db435),
	.w2(32'hbad50f0d),
	.w3(32'hbb28399e),
	.w4(32'hbaa3a332),
	.w5(32'h3a8efa5a),
	.w6(32'h3a14f836),
	.w7(32'h3b04277b),
	.w8(32'h3ac7b999),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b4009),
	.w1(32'h3c1b9109),
	.w2(32'h3bea0b5f),
	.w3(32'h3c9fc3f3),
	.w4(32'h3c0840a5),
	.w5(32'h3b5e4702),
	.w6(32'h3c1bc09c),
	.w7(32'h3b283941),
	.w8(32'hbaf746c0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c0b89),
	.w1(32'h3a508305),
	.w2(32'h3a451ace),
	.w3(32'h3abfa6b9),
	.w4(32'h3aba6760),
	.w5(32'h3a378a67),
	.w6(32'h39f9a665),
	.w7(32'h39ea60c0),
	.w8(32'h3a2104ac),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ca780),
	.w1(32'hbb843a18),
	.w2(32'hbc30d98e),
	.w3(32'hba28676b),
	.w4(32'hb9379f7b),
	.w5(32'hbb0246f2),
	.w6(32'h3b808ae0),
	.w7(32'h3b92872e),
	.w8(32'h3b015699),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b825c),
	.w1(32'h386ef1f9),
	.w2(32'h3a94b0d6),
	.w3(32'h39ca92de),
	.w4(32'h39e37fb0),
	.w5(32'h3a6eb83a),
	.w6(32'h39e21edf),
	.w7(32'h3a061959),
	.w8(32'h3a7888b2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88cf25),
	.w1(32'hba2d6c58),
	.w2(32'hbaae37fc),
	.w3(32'hba7319c0),
	.w4(32'hbb2bba41),
	.w5(32'hbb317138),
	.w6(32'h3a674f4e),
	.w7(32'h3a997b9b),
	.w8(32'hb9438a82),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5a7be),
	.w1(32'hbb03b4b9),
	.w2(32'hbb8ebcfd),
	.w3(32'hb9728bef),
	.w4(32'h3ad97e68),
	.w5(32'h3a0c5f8e),
	.w6(32'h3af0bb86),
	.w7(32'h3b79d194),
	.w8(32'h3a2a4f62),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa97cd0),
	.w1(32'hb9c506da),
	.w2(32'hb88a8834),
	.w3(32'h3aa42020),
	.w4(32'h39802245),
	.w5(32'h3aa2cd84),
	.w6(32'h3a6dacf1),
	.w7(32'h3a766187),
	.w8(32'h3aefcabf),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58a9ef),
	.w1(32'hbb8d3274),
	.w2(32'hbae18087),
	.w3(32'hbb135d07),
	.w4(32'h39e4b015),
	.w5(32'h392034df),
	.w6(32'h3a3e815a),
	.w7(32'h3b170706),
	.w8(32'h39be4a40),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b0d11),
	.w1(32'hbb02c75b),
	.w2(32'hbabfa237),
	.w3(32'h3afdc41a),
	.w4(32'h3b4cc52e),
	.w5(32'hb90ba07c),
	.w6(32'h3bdda6c5),
	.w7(32'h3bd506fa),
	.w8(32'h3b2aa449),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e9a8b),
	.w1(32'hba3cf297),
	.w2(32'hba1c80ad),
	.w3(32'hb78827de),
	.w4(32'h385cc7e3),
	.w5(32'hb9173bd5),
	.w6(32'h387122ef),
	.w7(32'hb9483fe1),
	.w8(32'hb8ae6d9e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4e966),
	.w1(32'h3cad3ba5),
	.w2(32'h3c8ff3a5),
	.w3(32'h3cef04ae),
	.w4(32'h3ca99a0e),
	.w5(32'h3c155e0e),
	.w6(32'h3c9f89a0),
	.w7(32'h3c0f5145),
	.w8(32'h3aa63696),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be74e1c),
	.w1(32'h3bfe275e),
	.w2(32'h3b614506),
	.w3(32'h3c249039),
	.w4(32'h3c003454),
	.w5(32'h3b093618),
	.w6(32'h3c098a0f),
	.w7(32'h3ba5b5f8),
	.w8(32'h39f02b86),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb895d080),
	.w1(32'hb7824e0f),
	.w2(32'hb781cec7),
	.w3(32'hb868a355),
	.w4(32'hb8049895),
	.w5(32'hb7b0aefc),
	.w6(32'hb88e5553),
	.w7(32'hb8390418),
	.w8(32'hb7ae11ae),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b371b7),
	.w1(32'h393bdec5),
	.w2(32'h39132d0d),
	.w3(32'h37b22c7c),
	.w4(32'h38db774e),
	.w5(32'h38cb0ab5),
	.w6(32'hb87caaf1),
	.w7(32'hb8302edb),
	.w8(32'hb85158b0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad19626),
	.w1(32'hba964565),
	.w2(32'hb966f32b),
	.w3(32'hbaf8fc36),
	.w4(32'hba65f789),
	.w5(32'hb964cb9b),
	.w6(32'hba8afc79),
	.w7(32'hb9b62331),
	.w8(32'hb908e102),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd044b6),
	.w1(32'h3cdf22d4),
	.w2(32'h3c5b82c7),
	.w3(32'h3d0a52cd),
	.w4(32'h3c836b1d),
	.w5(32'h3c448200),
	.w6(32'h3d05f8fc),
	.w7(32'h3c43a482),
	.w8(32'h3b7bb33e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe40e2),
	.w1(32'hbbb1789f),
	.w2(32'hbc3e1668),
	.w3(32'hbb9b2dc1),
	.w4(32'hbb7a7d9b),
	.w5(32'hbb8e8754),
	.w6(32'h3aaf158d),
	.w7(32'h3ab55d5d),
	.w8(32'hba14f55e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8286fe),
	.w1(32'hbbf3c455),
	.w2(32'hbc37e2be),
	.w3(32'hbc06297b),
	.w4(32'hbbfce25d),
	.w5(32'hbb79cd87),
	.w6(32'h3af344a2),
	.w7(32'h3b81c0dc),
	.w8(32'h3b0d8879),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc3725),
	.w1(32'hba280c94),
	.w2(32'hb97d48bf),
	.w3(32'hb90c5814),
	.w4(32'hb8487f03),
	.w5(32'h3980d908),
	.w6(32'hb7f2fb28),
	.w7(32'hb94fbee6),
	.w8(32'hb779b173),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb922c9c1),
	.w1(32'hb886abda),
	.w2(32'hb81563e0),
	.w3(32'hb9733711),
	.w4(32'hb91a5ef4),
	.w5(32'hb85546d4),
	.w6(32'hb9994bda),
	.w7(32'hb90a81fc),
	.w8(32'hb8e0a078),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dafe6),
	.w1(32'hbb999c1c),
	.w2(32'hbad4cd5f),
	.w3(32'hbbbfc9d0),
	.w4(32'hbbd187c1),
	.w5(32'h39d0b516),
	.w6(32'hbabae9e8),
	.w7(32'h3aab8bf1),
	.w8(32'h3ba25866),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85223b),
	.w1(32'hba89a80f),
	.w2(32'h390eda01),
	.w3(32'hbafbc50d),
	.w4(32'hbb195236),
	.w5(32'hbb1b349e),
	.w6(32'hbb12a626),
	.w7(32'hbb1e67a8),
	.w8(32'hbb063643),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65bf99),
	.w1(32'hbbfe1f33),
	.w2(32'hbc08f69a),
	.w3(32'hbbd803ef),
	.w4(32'hbb75f16b),
	.w5(32'hba8e6a05),
	.w6(32'hbac8d375),
	.w7(32'h3aef3a0d),
	.w8(32'h3b366ea9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83de610),
	.w1(32'hb83bb0fb),
	.w2(32'hb8285963),
	.w3(32'hb86922d7),
	.w4(32'hb8288c62),
	.w5(32'hb7eec048),
	.w6(32'hb8a32bc0),
	.w7(32'hb7f25ab4),
	.w8(32'hb7919c8d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5ec67f7),
	.w1(32'hb8684b71),
	.w2(32'hb959c714),
	.w3(32'hb745800a),
	.w4(32'hb813fa43),
	.w5(32'hb987f137),
	.w6(32'hb8074004),
	.w7(32'hb8bd55b1),
	.w8(32'hb99e81f5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a64ee0),
	.w1(32'hbae1dbd7),
	.w2(32'hbb718c50),
	.w3(32'h3a22f9a9),
	.w4(32'hba481ad9),
	.w5(32'hbb0eb0f5),
	.w6(32'h3ae0760c),
	.w7(32'hb95fb1c7),
	.w8(32'hbae93ae1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3879128f),
	.w1(32'hbab7bdc1),
	.w2(32'hbb226b3f),
	.w3(32'hba8dcf66),
	.w4(32'h37fde515),
	.w5(32'hba7f1f9a),
	.w6(32'h3aa1f4a4),
	.w7(32'h3ae464b8),
	.w8(32'hb85626b9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97132a4),
	.w1(32'hb9c4227d),
	.w2(32'hba031dd9),
	.w3(32'hb8c4293f),
	.w4(32'hb94ed157),
	.w5(32'hb9eeb5ad),
	.w6(32'h39ef30a8),
	.w7(32'h3a04066d),
	.w8(32'h39a20e78),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaaabaa),
	.w1(32'hba027ee9),
	.w2(32'hbae43980),
	.w3(32'h3a940193),
	.w4(32'h39d683dd),
	.w5(32'hba498f44),
	.w6(32'h3a9faf0c),
	.w7(32'h38c3c0db),
	.w8(32'hbab09d69),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0912fa),
	.w1(32'h3c0907e9),
	.w2(32'h3b4b2372),
	.w3(32'h3b8141eb),
	.w4(32'h3c0703f0),
	.w5(32'hba0633d9),
	.w6(32'h3c0ba8fe),
	.w7(32'h3c0065f2),
	.w8(32'h3b32a838),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc062273),
	.w1(32'hbc681e99),
	.w2(32'hbc13f163),
	.w3(32'hbcaa9589),
	.w4(32'hbc580663),
	.w5(32'hbb849ce3),
	.w6(32'hbbaec2a4),
	.w7(32'h3a4ee0c0),
	.w8(32'h3b3ab40c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38dfd2),
	.w1(32'hbc73ec4c),
	.w2(32'hbbebe5b8),
	.w3(32'hbcadd2f9),
	.w4(32'hbc551989),
	.w5(32'hbae3453c),
	.w6(32'hbc3edbfa),
	.w7(32'hba703530),
	.w8(32'h3b936f36),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3959d3),
	.w1(32'hbb08b4c4),
	.w2(32'hbab2d805),
	.w3(32'hbb78f6f3),
	.w4(32'hba14fe8f),
	.w5(32'h39adf5ee),
	.w6(32'hba8870c8),
	.w7(32'h3a7c53ab),
	.w8(32'h3aa1ff40),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f0ec02),
	.w1(32'h39e43c9d),
	.w2(32'h38ec1bdf),
	.w3(32'h39ef7a6d),
	.w4(32'h39a9daf3),
	.w5(32'h38b0031d),
	.w6(32'h39790668),
	.w7(32'h3934beba),
	.w8(32'h38501896),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f1b96),
	.w1(32'hb97db93e),
	.w2(32'hb8b0d67f),
	.w3(32'hb9e69a92),
	.w4(32'hb97d8e0e),
	.w5(32'hb881a7fa),
	.w6(32'hb9de09b0),
	.w7(32'hb9569a68),
	.w8(32'hb7c9e147),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25f6d2),
	.w1(32'hba2a9152),
	.w2(32'hbaedd459),
	.w3(32'h3a03e6de),
	.w4(32'hba53b3a8),
	.w5(32'hba5b693d),
	.w6(32'h394f48b5),
	.w7(32'hba4c26cb),
	.w8(32'hba1b312a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9363ff),
	.w1(32'hba29ba2f),
	.w2(32'hbb6c7b8d),
	.w3(32'h3bdd7db5),
	.w4(32'h38a5113b),
	.w5(32'hba8ba539),
	.w6(32'h3bd758e4),
	.w7(32'h3ac6fe3a),
	.w8(32'hba4ade49),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab554b3),
	.w1(32'hbba4c1c5),
	.w2(32'hbbed8902),
	.w3(32'hbb63bdc7),
	.w4(32'hbb3add64),
	.w5(32'hbb39509e),
	.w6(32'h3a24eb48),
	.w7(32'h3ad51c41),
	.w8(32'hb8a87048),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95fa526),
	.w1(32'hbbb5e620),
	.w2(32'hbc5825bb),
	.w3(32'hbb958f6a),
	.w4(32'hbb32e456),
	.w5(32'hbb979592),
	.w6(32'h3b4457f6),
	.w7(32'h3af1d64f),
	.w8(32'hbb258a67),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b680def),
	.w1(32'h3b17ca8d),
	.w2(32'hbb5e4df8),
	.w3(32'h3ba3e7cd),
	.w4(32'h3b813d4c),
	.w5(32'hbaa34d41),
	.w6(32'h3c205455),
	.w7(32'h3b996f7e),
	.w8(32'hb99d0793),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc81714),
	.w1(32'h3cdec3a6),
	.w2(32'h3c9349d5),
	.w3(32'h3d092965),
	.w4(32'h3cc422ab),
	.w5(32'h3c167ac6),
	.w6(32'h3ccfbd29),
	.w7(32'h3c3e5958),
	.w8(32'h3a76e193),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b3459),
	.w1(32'hb996dcbf),
	.w2(32'hb934408f),
	.w3(32'hb8bb3893),
	.w4(32'hba09bf1d),
	.w5(32'hb9503bb4),
	.w6(32'hb996edcf),
	.w7(32'hba01f844),
	.w8(32'hba0c0436),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e9d5e),
	.w1(32'h39f6e233),
	.w2(32'h39c80d83),
	.w3(32'h3a935d9c),
	.w4(32'h3a925adc),
	.w5(32'h3a8833b3),
	.w6(32'h3aa84d4f),
	.w7(32'h3aa18ab7),
	.w8(32'h3aae49f7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0d0d3),
	.w1(32'hba1a060a),
	.w2(32'h3986066a),
	.w3(32'hba26d054),
	.w4(32'hba3fda08),
	.w5(32'hb98a686e),
	.w6(32'hba206449),
	.w7(32'hb9ea7e50),
	.w8(32'hb91cb650),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33a575),
	.w1(32'h3a38ea32),
	.w2(32'hb9a2f9b9),
	.w3(32'h3ae0117f),
	.w4(32'hbaa8de26),
	.w5(32'h38884a3c),
	.w6(32'h3b208aff),
	.w7(32'h3ab70e05),
	.w8(32'h3aa94c65),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bc777),
	.w1(32'h3b0698a2),
	.w2(32'h3abb7b26),
	.w3(32'h3b2c827d),
	.w4(32'h3b0511c6),
	.w5(32'h3a1b78ba),
	.w6(32'h3b2afc8a),
	.w7(32'h3a3b2d3a),
	.w8(32'h39bcb25c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6626ed),
	.w1(32'h3c5838d0),
	.w2(32'h3ba0b4e3),
	.w3(32'h3ca3058c),
	.w4(32'h3c4a4bb6),
	.w5(32'hba40ec2f),
	.w6(32'h3c72f596),
	.w7(32'h3bc7c364),
	.w8(32'hb9eb9c03),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36f762),
	.w1(32'h3b1d1330),
	.w2(32'h3b35536c),
	.w3(32'h3ab71d16),
	.w4(32'h3a7850f7),
	.w5(32'h3a81723a),
	.w6(32'h39a5c2da),
	.w7(32'hba044085),
	.w8(32'h38f0bcbe),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94215ad),
	.w1(32'hb852f31c),
	.w2(32'h386d37c1),
	.w3(32'hb8fa573e),
	.w4(32'h38099438),
	.w5(32'h382c9b8e),
	.w6(32'hb8a552c7),
	.w7(32'h38b9e935),
	.w8(32'h389f5492),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72d9596),
	.w1(32'h3600eb5f),
	.w2(32'hb7227a1f),
	.w3(32'hb8299fb3),
	.w4(32'h36948b9d),
	.w5(32'hb6a330df),
	.w6(32'hb875bc73),
	.w7(32'hb6c133ab),
	.w8(32'hb73832f9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3895ca2c),
	.w1(32'h3917be14),
	.w2(32'hb89d934d),
	.w3(32'hb93dcddc),
	.w4(32'hb987f932),
	.w5(32'hb7874681),
	.w6(32'hb980101f),
	.w7(32'hb89431f3),
	.w8(32'h385a73bc),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27da33),
	.w1(32'hba0066d4),
	.w2(32'hb991dd09),
	.w3(32'hba0a2543),
	.w4(32'hba095d63),
	.w5(32'hb97f230c),
	.w6(32'hb9d1df29),
	.w7(32'hb9c9fb03),
	.w8(32'hb80f6a67),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940bd0b),
	.w1(32'hba01ead1),
	.w2(32'hb9c4d045),
	.w3(32'h393bcb59),
	.w4(32'hb9f52bc4),
	.w5(32'hb8a9f5c0),
	.w6(32'hb906b774),
	.w7(32'hb9ac2fd4),
	.w8(32'h38312424),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7f7ef),
	.w1(32'h3bc1bae7),
	.w2(32'h3b528f8c),
	.w3(32'h3c00fbb8),
	.w4(32'h3b95b587),
	.w5(32'h3ad9ddc9),
	.w6(32'h3baa1d00),
	.w7(32'h3ac8a65f),
	.w8(32'h3a11353a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27f8f3),
	.w1(32'h3be25e99),
	.w2(32'h3b7d00cc),
	.w3(32'h3c3cff8d),
	.w4(32'h3adf17e9),
	.w5(32'h3bada0fc),
	.w6(32'h3bbf973a),
	.w7(32'h3aac1a31),
	.w8(32'h3b44e79a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380f6c55),
	.w1(32'hb8442bae),
	.w2(32'hb8f2db31),
	.w3(32'h3798c5c5),
	.w4(32'hb8dd8b18),
	.w5(32'hb92a3b0a),
	.w6(32'hb853c003),
	.w7(32'hb8f408ca),
	.w8(32'hb958f738),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c19910),
	.w1(32'h37a9375e),
	.w2(32'h37572810),
	.w3(32'h373d197e),
	.w4(32'h37ea3ad4),
	.w5(32'h375f041c),
	.w6(32'hb78cc619),
	.w7(32'hb6ea94fa),
	.w8(32'hb78df88b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e11f87),
	.w1(32'hb951cc0c),
	.w2(32'h37756184),
	.w3(32'hb9b01bd0),
	.w4(32'hb9146a3a),
	.w5(32'hb8052c4d),
	.w6(32'hb9b3d1ac),
	.w7(32'hb96d4c05),
	.w8(32'hb9099b9c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f6a838),
	.w1(32'h382f53cc),
	.w2(32'hb6903493),
	.w3(32'hb870450d),
	.w4(32'hb81e81bd),
	.w5(32'hb8487492),
	.w6(32'hb8f7e264),
	.w7(32'hb8ccd2c7),
	.w8(32'hb8e9ac5d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa01d3f),
	.w1(32'h39b69f35),
	.w2(32'hba39effd),
	.w3(32'h3b4b8278),
	.w4(32'hbada1db6),
	.w5(32'hbb4003f3),
	.w6(32'h3bd5a51c),
	.w7(32'h3b9892bb),
	.w8(32'h3b4d02d8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3506b0),
	.w1(32'hbbabcf1d),
	.w2(32'hbc07e84c),
	.w3(32'hbb9505f9),
	.w4(32'hbac3f752),
	.w5(32'hba965e4e),
	.w6(32'h3b493ce3),
	.w7(32'h3a9784cb),
	.w8(32'hbab6c14c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ed3c8),
	.w1(32'h3c0267ee),
	.w2(32'h3a4f3cd5),
	.w3(32'h3c162ff6),
	.w4(32'hb9043823),
	.w5(32'hbade843f),
	.w6(32'h3c04d72c),
	.w7(32'h3ad1b76b),
	.w8(32'hba7f6126),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc0740),
	.w1(32'hbc375d24),
	.w2(32'hbc059e3f),
	.w3(32'hbc42c4a7),
	.w4(32'hbb668a84),
	.w5(32'h3c76aad0),
	.w6(32'h3a0c55f7),
	.w7(32'h3c095c72),
	.w8(32'h3c797cd8),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e5c76),
	.w1(32'hbb804f8d),
	.w2(32'hbbf101d2),
	.w3(32'hbc15f260),
	.w4(32'hbb40f933),
	.w5(32'hbbce1080),
	.w6(32'hbc98275c),
	.w7(32'hbbce8e09),
	.w8(32'hbb969586),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4844b0),
	.w1(32'hb98b99dd),
	.w2(32'hbb233fa8),
	.w3(32'hbab14ed7),
	.w4(32'hbbc68977),
	.w5(32'hbac6ef03),
	.w6(32'h3bc41b85),
	.w7(32'hba994016),
	.w8(32'h3b950c6e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e20a1),
	.w1(32'h3ac6dc3e),
	.w2(32'h3b81002a),
	.w3(32'hbbc4f689),
	.w4(32'h3b4d5965),
	.w5(32'h3bbf6ff9),
	.w6(32'hbacc384d),
	.w7(32'hba9974be),
	.w8(32'h3b1f103c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7ef7e),
	.w1(32'h3b9819ef),
	.w2(32'h3bd1e669),
	.w3(32'hb9df9259),
	.w4(32'h3b32f2da),
	.w5(32'h3c15a06b),
	.w6(32'h397e5709),
	.w7(32'h39a3570b),
	.w8(32'hbaea1316),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381ea192),
	.w1(32'h3b136ab8),
	.w2(32'hba71f8cd),
	.w3(32'hbb29d08c),
	.w4(32'hbafa0912),
	.w5(32'h3abe2e1e),
	.w6(32'hbb5e2e91),
	.w7(32'hbac17b9a),
	.w8(32'hbb3b0621),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ed218),
	.w1(32'h3c303836),
	.w2(32'h3c1f421b),
	.w3(32'h3c4a7c45),
	.w4(32'h3c129a78),
	.w5(32'hbaa86dd4),
	.w6(32'h3c2b4fb2),
	.w7(32'h3a24f7d4),
	.w8(32'hbb2676c1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b7f1e),
	.w1(32'h3c87f19d),
	.w2(32'h3c72abb3),
	.w3(32'h3cbb9e1e),
	.w4(32'h3d0819e0),
	.w5(32'hbb7ebbd5),
	.w6(32'h3c996359),
	.w7(32'h3c600fa2),
	.w8(32'h3ad20ac3),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a58fb),
	.w1(32'hbc6c908a),
	.w2(32'hbb152acd),
	.w3(32'hbc16e3a9),
	.w4(32'hbb106cc2),
	.w5(32'h3a833d3e),
	.w6(32'h3abbee75),
	.w7(32'hbb4956d4),
	.w8(32'hbbfb42fb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4723e4),
	.w1(32'hbb71c282),
	.w2(32'h3c01c1f5),
	.w3(32'hbaf22daa),
	.w4(32'hbb68070a),
	.w5(32'h3c48e82f),
	.w6(32'hbc1cc90e),
	.w7(32'hbb8faa17),
	.w8(32'h3b184e2d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1dffa0),
	.w1(32'hbb334ad9),
	.w2(32'hbbddf33b),
	.w3(32'hbab690d7),
	.w4(32'hbb81d734),
	.w5(32'hbbdfcdc2),
	.w6(32'h3c0a42f5),
	.w7(32'h3b8175cd),
	.w8(32'h3b56ec00),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ee414a),
	.w1(32'h3c01bba4),
	.w2(32'h3c89a8b8),
	.w3(32'hbb1d893b),
	.w4(32'h3c415a63),
	.w5(32'hbad88a1b),
	.w6(32'hbb3302de),
	.w7(32'h3c6cad78),
	.w8(32'h3caf18d9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c0552),
	.w1(32'h3bd634cf),
	.w2(32'hba2316d4),
	.w3(32'h3c99381e),
	.w4(32'h3a721f53),
	.w5(32'h3ad98f36),
	.w6(32'h3cbfa8be),
	.w7(32'h3a0ec883),
	.w8(32'hbbd32a7f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb896899),
	.w1(32'hb99a3023),
	.w2(32'hba6ff4b7),
	.w3(32'hbbdd58bf),
	.w4(32'hba1f543c),
	.w5(32'hbb517b75),
	.w6(32'hbb07b9eb),
	.w7(32'hb976a992),
	.w8(32'hbb9089fb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e592f),
	.w1(32'h3c393ffa),
	.w2(32'hb8d9fb3d),
	.w3(32'hba108d2b),
	.w4(32'h3c2eb0bf),
	.w5(32'h3c3e793f),
	.w6(32'h3acd0b92),
	.w7(32'h3b8bc311),
	.w8(32'h3b2be824),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab32e21),
	.w1(32'hbbbd01dc),
	.w2(32'hbc286b54),
	.w3(32'h3b97344c),
	.w4(32'hbb3c4685),
	.w5(32'hbc246d9b),
	.w6(32'h3b55878d),
	.w7(32'hbb85152b),
	.w8(32'hbb5a34da),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b572e57),
	.w1(32'hbb826338),
	.w2(32'h3ad67c27),
	.w3(32'hbb630c46),
	.w4(32'hbb41d709),
	.w5(32'hba455e87),
	.w6(32'hbada6fa1),
	.w7(32'hbbfe2724),
	.w8(32'hbba211c4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1254f6),
	.w1(32'hbb96e595),
	.w2(32'hbb928319),
	.w3(32'hbc4ddc4c),
	.w4(32'h39585ce9),
	.w5(32'h3afdf70c),
	.w6(32'hbc14c1cf),
	.w7(32'h3b372b4d),
	.w8(32'h3bf153c0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b109e3b),
	.w1(32'h3aa731d5),
	.w2(32'h3bd50b92),
	.w3(32'h3b5855b7),
	.w4(32'hbb14e3ba),
	.w5(32'h3b01007a),
	.w6(32'hba54c74c),
	.w7(32'hbba0fa5a),
	.w8(32'h3b817101),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae786c7),
	.w1(32'hbb91892e),
	.w2(32'h3a6cae58),
	.w3(32'hbbfadcdc),
	.w4(32'h3c0a7e51),
	.w5(32'h3b69e790),
	.w6(32'h3b61036c),
	.w7(32'hba540af2),
	.w8(32'hbb1bb6f5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb96981),
	.w1(32'h3c7a4213),
	.w2(32'h3ba0ce4a),
	.w3(32'h3d0fb38f),
	.w4(32'h3c8c2b3f),
	.w5(32'h3be8d94f),
	.w6(32'h3cbef9e9),
	.w7(32'h3b1ea100),
	.w8(32'hbb458dc4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e135a),
	.w1(32'hbbb5fab2),
	.w2(32'hbb67a445),
	.w3(32'hbbfcbb11),
	.w4(32'hbbfb09c2),
	.w5(32'hba143862),
	.w6(32'hb95ce206),
	.w7(32'hbbb6faa0),
	.w8(32'h3a32986b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf17e2),
	.w1(32'h3ba87ac9),
	.w2(32'h3c0be348),
	.w3(32'h3c18690b),
	.w4(32'hbb8ffe93),
	.w5(32'hbb0bf434),
	.w6(32'h3be98113),
	.w7(32'h3c639b32),
	.w8(32'h3c11086b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac8d94),
	.w1(32'hbc803317),
	.w2(32'hbbb3d3f5),
	.w3(32'hbbd90b21),
	.w4(32'hbc8a53bb),
	.w5(32'hbb50b57f),
	.w6(32'hbb755aef),
	.w7(32'hbb649877),
	.w8(32'hba9f795b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba37e81),
	.w1(32'hbbc51144),
	.w2(32'hbbe60ded),
	.w3(32'h3b5eadb9),
	.w4(32'hbb31af78),
	.w5(32'hbb27ae85),
	.w6(32'h3b3cfe56),
	.w7(32'hbab96d11),
	.w8(32'h3b382c44),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0896fb),
	.w1(32'hbb97960c),
	.w2(32'hbbdd3460),
	.w3(32'hbb845199),
	.w4(32'hba73a6c8),
	.w5(32'h3b744d82),
	.w6(32'h3a91c20e),
	.w7(32'hba648719),
	.w8(32'hbb6240be),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69e329),
	.w1(32'h3ad5031a),
	.w2(32'hbada8cae),
	.w3(32'h3b20e196),
	.w4(32'hbb67fa60),
	.w5(32'h3a33e5c7),
	.w6(32'hbb464520),
	.w7(32'h39e77250),
	.w8(32'h3a98059a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa9a20),
	.w1(32'h3b7b7c1b),
	.w2(32'hbb818e76),
	.w3(32'hbb31a418),
	.w4(32'h3a71a1e5),
	.w5(32'hb919d748),
	.w6(32'hbb6e2d06),
	.w7(32'hbb8904c4),
	.w8(32'hbc0951fd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb894a2ed),
	.w1(32'h3b8fe0a9),
	.w2(32'hbc15425d),
	.w3(32'h3b52985c),
	.w4(32'h3b34ec27),
	.w5(32'hbbb020d1),
	.w6(32'h3c10f79a),
	.w7(32'h3c0a14bb),
	.w8(32'h396354e2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5e1a5),
	.w1(32'hbb1a8066),
	.w2(32'hbc025131),
	.w3(32'hba9fa1b5),
	.w4(32'hbc0789d5),
	.w5(32'hbbb00c9a),
	.w6(32'h3abf4e8b),
	.w7(32'hba25735e),
	.w8(32'h3b342577),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c570a3a),
	.w1(32'h3cb374e3),
	.w2(32'h3c6c7652),
	.w3(32'h3d073c7e),
	.w4(32'h3c8982dd),
	.w5(32'h3b008ce3),
	.w6(32'h3cc91c26),
	.w7(32'h39a30f10),
	.w8(32'hbc3ec963),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b626c),
	.w1(32'hbc85da8f),
	.w2(32'hbc44664d),
	.w3(32'hbc7a75f6),
	.w4(32'hbc1f9241),
	.w5(32'hbb1fa276),
	.w6(32'hbc65d8bc),
	.w7(32'hbad94c44),
	.w8(32'h3b316614),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8439fa),
	.w1(32'hbc19f687),
	.w2(32'hbc332ac2),
	.w3(32'hbc5e0f5c),
	.w4(32'h3a8647df),
	.w5(32'h3bd186ea),
	.w6(32'h3bca5c69),
	.w7(32'h3bbedbf0),
	.w8(32'h39f1a221),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d168f),
	.w1(32'h3bad85fc),
	.w2(32'hbb53b1e4),
	.w3(32'h3be9d645),
	.w4(32'hba0db4a8),
	.w5(32'hbb8f69e3),
	.w6(32'h3c31d155),
	.w7(32'h3a812bc8),
	.w8(32'h3a31e0c3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa57ae),
	.w1(32'hbb9ac3d8),
	.w2(32'hbb3159c3),
	.w3(32'h3afbb12a),
	.w4(32'hbbbcd48a),
	.w5(32'h3b4e409b),
	.w6(32'hbaef29ba),
	.w7(32'hbbd1f787),
	.w8(32'hbb8169d2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb76b15),
	.w1(32'h3d0a8bea),
	.w2(32'h3cab91aa),
	.w3(32'h3cdefa56),
	.w4(32'h3cd26699),
	.w5(32'h3bced2f2),
	.w6(32'h3ce6039c),
	.w7(32'h3c96912e),
	.w8(32'h3bb08930),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1705a5),
	.w1(32'hbb590310),
	.w2(32'h3ad77339),
	.w3(32'hbbcfaee9),
	.w4(32'h3a9704be),
	.w5(32'h3b9ab547),
	.w6(32'h3ba22a8d),
	.w7(32'h3b3c1e94),
	.w8(32'h3b1c672a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b086d70),
	.w1(32'h3a7faa23),
	.w2(32'h3ab83c11),
	.w3(32'hba9f40d0),
	.w4(32'h3aa860ef),
	.w5(32'h3bcbf2ea),
	.w6(32'h3b0855b4),
	.w7(32'h392ad32e),
	.w8(32'hbb4e099c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25950e),
	.w1(32'h3a8ac82b),
	.w2(32'hbb69c1ae),
	.w3(32'hbab6af65),
	.w4(32'h3b8af6ee),
	.w5(32'hbb9f2f7c),
	.w6(32'h3b152485),
	.w7(32'h3b80ebd6),
	.w8(32'hba84adbf),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b725e96),
	.w1(32'hb820704f),
	.w2(32'h398d09c8),
	.w3(32'hb9bca9be),
	.w4(32'hbb13b863),
	.w5(32'h3b49c4ce),
	.w6(32'hbaf7d912),
	.w7(32'h3b99b3e2),
	.w8(32'h3b4410dc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39976b5b),
	.w1(32'h3a688434),
	.w2(32'h3b4f22e9),
	.w3(32'h3b117896),
	.w4(32'hbb60fbbf),
	.w5(32'hbbb2dca1),
	.w6(32'hbb24a950),
	.w7(32'hbb049698),
	.w8(32'hbb596227),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0073da),
	.w1(32'hbc12ab2c),
	.w2(32'h3b0332b3),
	.w3(32'hbad06a56),
	.w4(32'hbc18e20e),
	.w5(32'hbb3b2c93),
	.w6(32'hbbebd811),
	.w7(32'hbb807904),
	.w8(32'hbb928eba),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49045c),
	.w1(32'hbb174ba2),
	.w2(32'hbb686c33),
	.w3(32'hbb5f9521),
	.w4(32'h3b6bd823),
	.w5(32'h3c891795),
	.w6(32'hb9fbfdcc),
	.w7(32'h3b767c68),
	.w8(32'hbacafac2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beff595),
	.w1(32'h3b80bcde),
	.w2(32'hbb2953b2),
	.w3(32'h3b8217a6),
	.w4(32'hbaaf2d22),
	.w5(32'h3bf74a55),
	.w6(32'h3b58cab9),
	.w7(32'hbb7b41a5),
	.w8(32'hbc0daa06),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dfc36),
	.w1(32'h3a7501bb),
	.w2(32'hba27185b),
	.w3(32'hba95c4c5),
	.w4(32'h3a064b2f),
	.w5(32'hbc2ad8b4),
	.w6(32'h3ba9c001),
	.w7(32'h3b1caaf0),
	.w8(32'h3aeddb05),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb754297),
	.w1(32'hbb00770b),
	.w2(32'hb76de26e),
	.w3(32'h3bbbd3dc),
	.w4(32'hbc047485),
	.w5(32'h3cd5f38d),
	.w6(32'hbbec09b2),
	.w7(32'h3b0f85c0),
	.w8(32'h3c1c0b77),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea0ab7),
	.w1(32'hbaf2b53b),
	.w2(32'h3b2c5b64),
	.w3(32'h3a69093f),
	.w4(32'h3b4bd5b7),
	.w5(32'h3bcf7a89),
	.w6(32'hbba7158a),
	.w7(32'h399144ec),
	.w8(32'hbb34f76c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ae656),
	.w1(32'hbaddadf9),
	.w2(32'h3bae4f7f),
	.w3(32'h3b9d904f),
	.w4(32'hb98c45be),
	.w5(32'h3c5c1db7),
	.w6(32'h3be0449c),
	.w7(32'h39cab176),
	.w8(32'h3be0612f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3620ed),
	.w1(32'hbb3ed8f8),
	.w2(32'hbbf3d26d),
	.w3(32'hbbe61c6b),
	.w4(32'hbb94bc3c),
	.w5(32'hbac54450),
	.w6(32'hbb780d92),
	.w7(32'h3b9fe12b),
	.w8(32'hbb9df160),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba746c5),
	.w1(32'hbb5f5545),
	.w2(32'hbb0d4466),
	.w3(32'h38db783d),
	.w4(32'hbb29e5b3),
	.w5(32'h3b1f03d8),
	.w6(32'hbb46114d),
	.w7(32'h3b39ccf6),
	.w8(32'h3b9c38c8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb07079),
	.w1(32'hbbf85c2c),
	.w2(32'hbc2a856d),
	.w3(32'hbc46e447),
	.w4(32'hbaacfeb0),
	.w5(32'hbb221298),
	.w6(32'hbb00dc4a),
	.w7(32'hba74472d),
	.w8(32'h3a14977d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb840e1b8),
	.w1(32'h3a61a36f),
	.w2(32'hba1c3da7),
	.w3(32'hbbbce230),
	.w4(32'hba8274e8),
	.w5(32'hbb59b10a),
	.w6(32'hbb3e001f),
	.w7(32'hbaa3d914),
	.w8(32'hbaa81467),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba16be1),
	.w1(32'h3bed16ce),
	.w2(32'h3b8bf33c),
	.w3(32'h3b31d73f),
	.w4(32'h3c49513e),
	.w5(32'h3babfdb5),
	.w6(32'h3b9ccd29),
	.w7(32'h3bdb2901),
	.w8(32'h3c4687d7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11f13b),
	.w1(32'hbc1a0849),
	.w2(32'hbc240f5b),
	.w3(32'h3c96c2ff),
	.w4(32'hbb52ea98),
	.w5(32'hbb006f3f),
	.w6(32'hbc49a644),
	.w7(32'hbabf2c2f),
	.w8(32'h3b1903b4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb057a6),
	.w1(32'hbb0f9685),
	.w2(32'hba5fab33),
	.w3(32'hbb2d1e20),
	.w4(32'h3b2586bb),
	.w5(32'h3c061849),
	.w6(32'h3c10442a),
	.w7(32'h3a191515),
	.w8(32'hbabf541a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9a864),
	.w1(32'h3adce7c6),
	.w2(32'h3bf7c509),
	.w3(32'hbc0b1462),
	.w4(32'hbabaeb8d),
	.w5(32'hbab41239),
	.w6(32'hbbd9668e),
	.w7(32'h3b23ea68),
	.w8(32'h3bd5a397),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4afa99),
	.w1(32'h3bc84e11),
	.w2(32'hb99b7e8e),
	.w3(32'hbba629cb),
	.w4(32'hba41aa09),
	.w5(32'hb9fcb572),
	.w6(32'hbb53af14),
	.w7(32'hb996efa4),
	.w8(32'hbbb482b9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2ce19),
	.w1(32'hbba4e0eb),
	.w2(32'hbb80c515),
	.w3(32'hbb8685dc),
	.w4(32'hbbcbd7b3),
	.w5(32'h3afbae45),
	.w6(32'hbb710052),
	.w7(32'hbbb3b62d),
	.w8(32'hbba4ad42),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ea2bb),
	.w1(32'hbad1ec38),
	.w2(32'hbb9dd35d),
	.w3(32'hbbdb61a8),
	.w4(32'h3b84982a),
	.w5(32'h3bb633c7),
	.w6(32'hbb9814b7),
	.w7(32'hbb3e0aa6),
	.w8(32'h3b04c28b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395feb82),
	.w1(32'h3bc80901),
	.w2(32'hbb8875ff),
	.w3(32'h3ac65a63),
	.w4(32'h3c505c79),
	.w5(32'hbcc418ec),
	.w6(32'h3c2311d7),
	.w7(32'h3ba7ba37),
	.w8(32'hbb2a9f50),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4040b),
	.w1(32'h3b67630f),
	.w2(32'hbb6b6f23),
	.w3(32'h3c6c8791),
	.w4(32'h3b793fd0),
	.w5(32'h3b00de47),
	.w6(32'h3c219f68),
	.w7(32'hbb5461d9),
	.w8(32'hbbbe6e17),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef6f98),
	.w1(32'h3b475dd2),
	.w2(32'hba15aaa1),
	.w3(32'hb9b99fa9),
	.w4(32'h3ade899e),
	.w5(32'hbb8c2e3b),
	.w6(32'hbb186b77),
	.w7(32'hbb452bcb),
	.w8(32'h3b12ad14),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd8db6),
	.w1(32'h3a467c3a),
	.w2(32'h3b1f09ea),
	.w3(32'hb9b81a87),
	.w4(32'hbaa93973),
	.w5(32'hbbaca32d),
	.w6(32'hbb300598),
	.w7(32'hba08ed88),
	.w8(32'h3c4eab22),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eaf21),
	.w1(32'h3b7434cf),
	.w2(32'h3aa26f19),
	.w3(32'h3c218fdb),
	.w4(32'h3bd8b3f1),
	.w5(32'h3ad7e4cb),
	.w6(32'h3a8c161f),
	.w7(32'h3ac5c184),
	.w8(32'hb9a84ef9),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e1ab4),
	.w1(32'hbc422927),
	.w2(32'hbbfa7824),
	.w3(32'hbb60c4ae),
	.w4(32'hbc51949e),
	.w5(32'h3c8a2f81),
	.w6(32'hba35361e),
	.w7(32'hb9aa425a),
	.w8(32'hbbaaebf9),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c023c52),
	.w1(32'h3c7558f6),
	.w2(32'h3c19df4a),
	.w3(32'h3c537e24),
	.w4(32'h3c2033ef),
	.w5(32'h3a0c2de4),
	.w6(32'h3bd0e388),
	.w7(32'h3b8c191e),
	.w8(32'hb9541e36),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27be2d),
	.w1(32'hbbc6fdeb),
	.w2(32'hbbad2565),
	.w3(32'hbc3d93a0),
	.w4(32'hbbad62d4),
	.w5(32'hbb12f25d),
	.w6(32'hbb6f3b08),
	.w7(32'hb999479b),
	.w8(32'h3b13a2be),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff6519),
	.w1(32'h3bb14862),
	.w2(32'hbad35de8),
	.w3(32'h3baefe6a),
	.w4(32'hb8e0ed00),
	.w5(32'h3af356d2),
	.w6(32'h3c01bd20),
	.w7(32'h3b1cf721),
	.w8(32'h3b5d29a6),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c382f2c),
	.w1(32'h3c7d6dfc),
	.w2(32'h3c2c55a9),
	.w3(32'h3c63d72d),
	.w4(32'h3c789abe),
	.w5(32'hba1a0e13),
	.w6(32'h3c10b69f),
	.w7(32'h3b641bd0),
	.w8(32'hb9f3d941),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb587d68),
	.w1(32'h3b97706a),
	.w2(32'hbb97f688),
	.w3(32'h3ba984ed),
	.w4(32'h3a812a5c),
	.w5(32'hbb8a87e6),
	.w6(32'hbb5c9c63),
	.w7(32'h3a38cf6c),
	.w8(32'hbafe2875),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86dfe2),
	.w1(32'hbadb8489),
	.w2(32'h3a813e65),
	.w3(32'h3b6b265c),
	.w4(32'h3b800c0a),
	.w5(32'h3c2ec612),
	.w6(32'h3abf6ed5),
	.w7(32'h3a69b8c8),
	.w8(32'h399ca3c7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60a7ee),
	.w1(32'hba5a436b),
	.w2(32'hbbe4b463),
	.w3(32'hbbaf52ad),
	.w4(32'h3aa7ed97),
	.w5(32'h3c4b2bae),
	.w6(32'h3b008617),
	.w7(32'hbb8c206f),
	.w8(32'hbbd4d761),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a486d),
	.w1(32'hbbabe46a),
	.w2(32'hbbbb5171),
	.w3(32'hbc908ade),
	.w4(32'hbc5c05b0),
	.w5(32'hbb4413b3),
	.w6(32'hbb7dba08),
	.w7(32'hb9cdba54),
	.w8(32'h3b9186e1),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacae236),
	.w1(32'hbbd54543),
	.w2(32'hbbce65c8),
	.w3(32'hba630ecd),
	.w4(32'hb9ee6cb7),
	.w5(32'hba849826),
	.w6(32'h3b2a20cc),
	.w7(32'hbb737a6a),
	.w8(32'hbbf97de6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba75b15),
	.w1(32'hbb9b22a8),
	.w2(32'hbb5c1be0),
	.w3(32'h3a84a157),
	.w4(32'hbc004f2c),
	.w5(32'h3ad176b4),
	.w6(32'hb9a1f35d),
	.w7(32'hbc444e77),
	.w8(32'hbb712d75),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaff561),
	.w1(32'hb9d5200b),
	.w2(32'hbab6cb0c),
	.w3(32'h3a20e8ba),
	.w4(32'hba8a94fb),
	.w5(32'hbb82012d),
	.w6(32'h3b0e397d),
	.w7(32'h3b017684),
	.w8(32'h3b60d78d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba25878),
	.w1(32'h3b3c8150),
	.w2(32'hbba241c5),
	.w3(32'hbbc52552),
	.w4(32'hbc0fcf88),
	.w5(32'hbc4d60f4),
	.w6(32'h3b46c9b8),
	.w7(32'h382c0a16),
	.w8(32'hbbd494ca),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9fda0),
	.w1(32'hbb8b50e2),
	.w2(32'hbb8ef993),
	.w3(32'h3aadc556),
	.w4(32'h3b51f125),
	.w5(32'h3b9802a5),
	.w6(32'h3b709816),
	.w7(32'h3b100ee6),
	.w8(32'hbb011e70),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83429e),
	.w1(32'hbbde76b4),
	.w2(32'hbc3d7eb0),
	.w3(32'hba2ee53c),
	.w4(32'hb998b1e2),
	.w5(32'hbc88ba6d),
	.w6(32'h3a290990),
	.w7(32'h3b9b7d1a),
	.w8(32'hbc4e0d3f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa02f34),
	.w1(32'hbb84206b),
	.w2(32'hb986e211),
	.w3(32'hbb252592),
	.w4(32'hbb660654),
	.w5(32'h3c8b3695),
	.w6(32'hbbb4f338),
	.w7(32'hbb10b276),
	.w8(32'hbbb8e85f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb332fba),
	.w1(32'hbac5c6db),
	.w2(32'hbcb564d2),
	.w3(32'hbb1c13c9),
	.w4(32'h3aa51774),
	.w5(32'hbc8710c9),
	.w6(32'hbc35bc19),
	.w7(32'h3abd4237),
	.w8(32'hbc3d71ac),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbd645),
	.w1(32'h3b64c961),
	.w2(32'hbb81dc9a),
	.w3(32'hbc0c678c),
	.w4(32'h3c6b847d),
	.w5(32'h3d529c77),
	.w6(32'hbba1740d),
	.w7(32'h3a566f50),
	.w8(32'hb929db6a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7f2ca),
	.w1(32'h3c2242f3),
	.w2(32'hb9e84c0b),
	.w3(32'h3c932a85),
	.w4(32'h3c0cfeca),
	.w5(32'hbb31536d),
	.w6(32'h3c1b662c),
	.w7(32'h3b76305a),
	.w8(32'hbbfc6f81),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98d2d2),
	.w1(32'hbbccd9e1),
	.w2(32'hbc1e8fa0),
	.w3(32'hbc4f2b27),
	.w4(32'hbc7a314c),
	.w5(32'h3c58d036),
	.w6(32'hbc414940),
	.w7(32'hbc7d357c),
	.w8(32'h3b853262),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe24da5),
	.w1(32'hbb673b4c),
	.w2(32'hbb89f192),
	.w3(32'hbc25e95f),
	.w4(32'hbc153bee),
	.w5(32'hbc2ee45d),
	.w6(32'hbc9aa404),
	.w7(32'hbad67d07),
	.w8(32'hbbd4518a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da57fa),
	.w1(32'h3c36c76a),
	.w2(32'hba59f715),
	.w3(32'hba4d6a50),
	.w4(32'h3bd3cdd6),
	.w5(32'h3aef217e),
	.w6(32'hbc03d2fd),
	.w7(32'hbb4fe37f),
	.w8(32'h3ab437ac),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f3888),
	.w1(32'h3c23d613),
	.w2(32'h3a40f36c),
	.w3(32'h3c1bb875),
	.w4(32'h3b89e548),
	.w5(32'hbbde23d6),
	.w6(32'h3c19f986),
	.w7(32'h3b80f8ef),
	.w8(32'h3bc14562),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a68605),
	.w1(32'h3b83a205),
	.w2(32'h3b8d6864),
	.w3(32'h3afde3dc),
	.w4(32'h3ba269bf),
	.w5(32'h3c1c4aa8),
	.w6(32'hbc4578fb),
	.w7(32'h3bcc493e),
	.w8(32'hba836fbb),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a87a2),
	.w1(32'hbb8c6dc9),
	.w2(32'hba91aa98),
	.w3(32'hbc5c8503),
	.w4(32'h3a0d9b8b),
	.w5(32'h3c0899b6),
	.w6(32'h3a2c407f),
	.w7(32'h3b45f532),
	.w8(32'hbbc2d7ec),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5dad7),
	.w1(32'h3bc4b93a),
	.w2(32'h3c5465dc),
	.w3(32'hbb13da46),
	.w4(32'h3b8f4af6),
	.w5(32'h3b2dfd6e),
	.w6(32'h3aed8cff),
	.w7(32'h3b3004af),
	.w8(32'hbb8844a3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d103f),
	.w1(32'h3bb23c8f),
	.w2(32'h3b6feb85),
	.w3(32'h3a50dd61),
	.w4(32'h3c1ae8a3),
	.w5(32'h3b6f69c0),
	.w6(32'h396652be),
	.w7(32'h3b72c106),
	.w8(32'h3b9c1a42),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9a57b),
	.w1(32'hbae3669a),
	.w2(32'hbaff7241),
	.w3(32'h3b994d07),
	.w4(32'hbb11677f),
	.w5(32'hbbc0ce6e),
	.w6(32'h3b85ce84),
	.w7(32'hbbfc3395),
	.w8(32'h3bbdaa95),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ca979),
	.w1(32'h3b8e5f6f),
	.w2(32'h3b9c4b79),
	.w3(32'hb98ecef2),
	.w4(32'h3aa0967d),
	.w5(32'hbb3bcac9),
	.w6(32'hbac4c2c5),
	.w7(32'h3ad0bf99),
	.w8(32'h3a6cd204),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38d830),
	.w1(32'hb9d65ba7),
	.w2(32'hbbab0dc9),
	.w3(32'h3c0c9c0c),
	.w4(32'hbc6df38e),
	.w5(32'hbc1812e3),
	.w6(32'hbbb1af30),
	.w7(32'hbb94ec87),
	.w8(32'hbb33b4d8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61c45fd),
	.w1(32'hbb3a0aa8),
	.w2(32'h3ba06470),
	.w3(32'h3be061b7),
	.w4(32'hbb593847),
	.w5(32'h3c0a0246),
	.w6(32'h3b49d016),
	.w7(32'hbb642d91),
	.w8(32'h3b55b315),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb484c8),
	.w1(32'hbc32f1e8),
	.w2(32'hbc14a9e0),
	.w3(32'hbbc1f444),
	.w4(32'hbc075795),
	.w5(32'hbb8999d7),
	.w6(32'hbb635564),
	.w7(32'hbbd5e0b5),
	.w8(32'hbb9b702c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb229ed4),
	.w1(32'hbb9b5dd2),
	.w2(32'h3b099266),
	.w3(32'hbaa5a9d9),
	.w4(32'hb8eae5d7),
	.w5(32'h3c05ae3a),
	.w6(32'hbabf6111),
	.w7(32'hbb8cf216),
	.w8(32'hbb326b81),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3759b),
	.w1(32'h3c17338f),
	.w2(32'h3b61c76f),
	.w3(32'hbb5d817e),
	.w4(32'h3c0e6fdd),
	.w5(32'hbc6c9697),
	.w6(32'hbb6041d8),
	.w7(32'h3bbfcdc3),
	.w8(32'hbb7377d8),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a75a3),
	.w1(32'h3ad15ff1),
	.w2(32'hbb8096b9),
	.w3(32'hbb99f6dd),
	.w4(32'h3c23b66c),
	.w5(32'hbc62941f),
	.w6(32'hbc2cf93a),
	.w7(32'hba2a9e7a),
	.w8(32'hbbb08ab9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd05bb0),
	.w1(32'h3b7c15a7),
	.w2(32'hbc3059ef),
	.w3(32'h3c9cac6d),
	.w4(32'h3c850aad),
	.w5(32'hbc23318d),
	.w6(32'h3c3bdc7a),
	.w7(32'h3a10ad66),
	.w8(32'hbb5e1a6b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0c9bd),
	.w1(32'h3982ac36),
	.w2(32'hbbea354d),
	.w3(32'h3a3f953b),
	.w4(32'h3c05acce),
	.w5(32'h3a6e4e45),
	.w6(32'hba836902),
	.w7(32'h3adecba0),
	.w8(32'hbbb2166d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4a49e),
	.w1(32'h3b1cfb55),
	.w2(32'h3a9c755d),
	.w3(32'hbbaf03f8),
	.w4(32'h3bb4fa36),
	.w5(32'h3bf721a8),
	.w6(32'hbb43cd3d),
	.w7(32'h3ac2164b),
	.w8(32'hb91c9c92),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb076eb6),
	.w1(32'h3c26aaf0),
	.w2(32'h3bc576de),
	.w3(32'h3a862d74),
	.w4(32'h3c8fea6d),
	.w5(32'hbc9451f0),
	.w6(32'h3aa87af2),
	.w7(32'h3c0a5d3b),
	.w8(32'h3c1b7550),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89d927),
	.w1(32'hba1fd775),
	.w2(32'hbbac5c20),
	.w3(32'h3c977b86),
	.w4(32'hb94daa52),
	.w5(32'h3a6e92c9),
	.w6(32'h3be488be),
	.w7(32'hbae50f95),
	.w8(32'hbbe0f4ca),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923e7a8),
	.w1(32'h3a4ef834),
	.w2(32'hbb94a306),
	.w3(32'h39a77ac8),
	.w4(32'hbbb8731b),
	.w5(32'hbb91e9a6),
	.w6(32'h3b830f41),
	.w7(32'hbb9e6a8a),
	.w8(32'h3a24181c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87e210),
	.w1(32'hb8c47c57),
	.w2(32'hbad82fc1),
	.w3(32'h3c6ea6ad),
	.w4(32'h38be9638),
	.w5(32'hbbefc1fc),
	.w6(32'h3c3ab5fa),
	.w7(32'hbb8dd53d),
	.w8(32'hbb98f481),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384ab5d2),
	.w1(32'h3b3f4942),
	.w2(32'h38e94f98),
	.w3(32'hbb4d840d),
	.w4(32'hbbc9ba0e),
	.w5(32'h3b3cdae1),
	.w6(32'hbb965d23),
	.w7(32'h3b174441),
	.w8(32'hb87563be),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadab987),
	.w1(32'hbbcb60d3),
	.w2(32'h3acca3d0),
	.w3(32'hbbb4ae2c),
	.w4(32'hbbcb5db7),
	.w5(32'h3b71992f),
	.w6(32'hb9be4989),
	.w7(32'hba229680),
	.w8(32'h3bdea98d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908b6aa),
	.w1(32'hbbc61a0f),
	.w2(32'h3bc2d68a),
	.w3(32'hb9d5580b),
	.w4(32'h39c18c05),
	.w5(32'h3c3ea0f4),
	.w6(32'h3a524dd5),
	.w7(32'hba63d007),
	.w8(32'h3b412cb9),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3347d),
	.w1(32'hbaf08711),
	.w2(32'h3b807a05),
	.w3(32'hbbb3ca26),
	.w4(32'hbc0c99ac),
	.w5(32'h3ce68b4c),
	.w6(32'hbbb5ea5e),
	.w7(32'hba199e1f),
	.w8(32'hbba3ffda),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90af7c),
	.w1(32'h3ae6860c),
	.w2(32'hbbcbb919),
	.w3(32'hbbf9b151),
	.w4(32'hbb078919),
	.w5(32'hbc14c03e),
	.w6(32'hbbea6a52),
	.w7(32'h3b3123be),
	.w8(32'h3a93d917),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb076b56),
	.w1(32'hbb5b0dbb),
	.w2(32'h3a7ba5e8),
	.w3(32'h3af2ead1),
	.w4(32'hbb136302),
	.w5(32'h3c1bf95f),
	.w6(32'h3b16ffa7),
	.w7(32'h3b2fcde6),
	.w8(32'hb8c628df),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af34195),
	.w1(32'h3b9afc61),
	.w2(32'h3bce9ee8),
	.w3(32'h3b6188aa),
	.w4(32'hbb492eca),
	.w5(32'hba13c48c),
	.w6(32'hba566019),
	.w7(32'hbb972a3b),
	.w8(32'h3b613597),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfa351),
	.w1(32'h3b5a028d),
	.w2(32'h3adb1392),
	.w3(32'h3bd2d323),
	.w4(32'h3c3bb384),
	.w5(32'hbb00eb3e),
	.w6(32'h3b5bfa19),
	.w7(32'h3b45b2e5),
	.w8(32'hba609876),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c5025),
	.w1(32'h3b6cc63a),
	.w2(32'h3b80de6e),
	.w3(32'hbae4abdc),
	.w4(32'h3b6e54b6),
	.w5(32'hba080274),
	.w6(32'h39be9669),
	.w7(32'hba0a29bd),
	.w8(32'hb9c55f75),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c3773a),
	.w1(32'h3bb583de),
	.w2(32'h3b3fbf2e),
	.w3(32'hbaa30e77),
	.w4(32'h3ba31889),
	.w5(32'h3c9ffd35),
	.w6(32'h3b0c9996),
	.w7(32'h3b8722ac),
	.w8(32'h3c02073d),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9158c2),
	.w1(32'hbbdb2999),
	.w2(32'hbbcc803f),
	.w3(32'hbc720427),
	.w4(32'hbc4c1b13),
	.w5(32'hbb7c09d4),
	.w6(32'h39f62ba3),
	.w7(32'hbbc453a6),
	.w8(32'hbc30e39c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be2b29),
	.w1(32'h3bc78bbd),
	.w2(32'hba850ed6),
	.w3(32'h3b110b21),
	.w4(32'h3b86c240),
	.w5(32'hbb24c995),
	.w6(32'hbc04af43),
	.w7(32'h3aa57d62),
	.w8(32'h3ad1fcd2),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d233d),
	.w1(32'h3b87cdee),
	.w2(32'hbc01d435),
	.w3(32'h3c0018f8),
	.w4(32'h3c286891),
	.w5(32'h3ae1ad4a),
	.w6(32'h3c2c8d9a),
	.w7(32'h3c127bbc),
	.w8(32'hbc135709),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71da08),
	.w1(32'hbc7e2953),
	.w2(32'hbc835e58),
	.w3(32'hbc882b7b),
	.w4(32'hbc832184),
	.w5(32'hbbc560cd),
	.w6(32'hbc3441f8),
	.w7(32'h3ac57248),
	.w8(32'h3b07664e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a80f),
	.w1(32'h39cb9fab),
	.w2(32'hba7a73bc),
	.w3(32'hbb7c59a6),
	.w4(32'h3b6ffbcd),
	.w5(32'hbc163da4),
	.w6(32'hbba3e542),
	.w7(32'h39a7623c),
	.w8(32'h3ac217d3),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dd287),
	.w1(32'h3b83967d),
	.w2(32'hbc1e7f97),
	.w3(32'h3ad479f7),
	.w4(32'hbb0c5cc4),
	.w5(32'hbc142c22),
	.w6(32'h3b138c90),
	.w7(32'hbaf4eb01),
	.w8(32'hbb6f5f33),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb06e8),
	.w1(32'hb7a08d65),
	.w2(32'h3bf3f806),
	.w3(32'h3bd61f3f),
	.w4(32'h3b19e316),
	.w5(32'h3bf697bc),
	.w6(32'hbb8823e4),
	.w7(32'h3bc647cf),
	.w8(32'hbb47e0ec),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb121e7e),
	.w1(32'h3c2f1042),
	.w2(32'h3bf5eb69),
	.w3(32'hbc1c3ef4),
	.w4(32'h3c14fdb4),
	.w5(32'hbba0e2d1),
	.w6(32'h3b96e667),
	.w7(32'h3c1ff29f),
	.w8(32'h3c011e30),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b517b07),
	.w1(32'h3bc8e846),
	.w2(32'hb814e2a2),
	.w3(32'h3ba83745),
	.w4(32'hbaba55b3),
	.w5(32'hbbff9ea9),
	.w6(32'h3c0fcd3f),
	.w7(32'hba916b1f),
	.w8(32'hbbb2336f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85edb7),
	.w1(32'h3b1e7887),
	.w2(32'hbb8831ae),
	.w3(32'h3af9a362),
	.w4(32'hbba83852),
	.w5(32'hba13b4b2),
	.w6(32'h3ae971d6),
	.w7(32'h3a180226),
	.w8(32'h3b1bd718),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01fa55),
	.w1(32'h3bc8927c),
	.w2(32'hbbbccca1),
	.w3(32'hb80f656d),
	.w4(32'hbb89e5b5),
	.w5(32'hbc0da811),
	.w6(32'h3b2c2d7f),
	.w7(32'h3c2de4b2),
	.w8(32'h3abee7e2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c270715),
	.w1(32'h3a9ff351),
	.w2(32'hbbe2251c),
	.w3(32'h3bb12317),
	.w4(32'hb9236e0e),
	.w5(32'hbb6c7c61),
	.w6(32'h3c3d5930),
	.w7(32'hba113905),
	.w8(32'hbc0c9122),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb55eb8),
	.w1(32'h39d5a9d5),
	.w2(32'hbbc27237),
	.w3(32'hbbdbb10a),
	.w4(32'h3b512f9f),
	.w5(32'hbaca1b05),
	.w6(32'hbbe2d47a),
	.w7(32'h3b94af8f),
	.w8(32'h3a8af65b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b6477),
	.w1(32'h3bbe2bd6),
	.w2(32'h3a25b672),
	.w3(32'h3b87929b),
	.w4(32'h3b851210),
	.w5(32'hbbbb6e5d),
	.w6(32'h3b948996),
	.w7(32'h3c0dd6f0),
	.w8(32'h3b5c0712),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14d150),
	.w1(32'h3a776d0a),
	.w2(32'hba84b826),
	.w3(32'hbb7d193e),
	.w4(32'h3be3cfa4),
	.w5(32'hbc20d1b0),
	.w6(32'hbb8c5476),
	.w7(32'h3ba3f706),
	.w8(32'h3b66a457),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1730b1),
	.w1(32'h3aba0f1f),
	.w2(32'hbab27ef9),
	.w3(32'hba9185e9),
	.w4(32'h3b4e6f17),
	.w5(32'h39541230),
	.w6(32'h3ae15757),
	.w7(32'h3b02d59b),
	.w8(32'hbb58b050),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa72053),
	.w1(32'hbabfd02d),
	.w2(32'hbb340322),
	.w3(32'h385de04c),
	.w4(32'hbba76da6),
	.w5(32'hbb4101cf),
	.w6(32'hbad38e00),
	.w7(32'hbacd3fed),
	.w8(32'hbb8667fe),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2caa7a),
	.w1(32'hb9ad29c6),
	.w2(32'hba313d4b),
	.w3(32'h3a9c8efa),
	.w4(32'hbbafa87d),
	.w5(32'hbb8b87d3),
	.w6(32'hb94c2e10),
	.w7(32'hbb408484),
	.w8(32'hbb835f03),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8051e7),
	.w1(32'hba76f68f),
	.w2(32'h3ac155fc),
	.w3(32'hbc0e84f7),
	.w4(32'hbbcfa919),
	.w5(32'hbb03d164),
	.w6(32'hbb5c7031),
	.w7(32'hbb103f1a),
	.w8(32'h3a010b9f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ca012),
	.w1(32'hbbc7c9a4),
	.w2(32'hbc334871),
	.w3(32'hbb5fe7af),
	.w4(32'hbb2fabea),
	.w5(32'hbaab89b8),
	.w6(32'h3a8a8fba),
	.w7(32'h3b69316d),
	.w8(32'hbad3c1e3),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba18502),
	.w1(32'h3bdb98c7),
	.w2(32'h3c3c6f7b),
	.w3(32'hbbd6e78b),
	.w4(32'h3beacd06),
	.w5(32'h3b20aa43),
	.w6(32'hbbb66153),
	.w7(32'h3af6b633),
	.w8(32'h3aa0c1ca),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8efe8f),
	.w1(32'hbc1a7910),
	.w2(32'hbb66ce94),
	.w3(32'hbb889742),
	.w4(32'hbbc82930),
	.w5(32'hbb76081d),
	.w6(32'hbb7dc228),
	.w7(32'hbb471cf0),
	.w8(32'h39854e92),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbffe29),
	.w1(32'hbb9b6d0e),
	.w2(32'hbbc4264a),
	.w3(32'hbc173999),
	.w4(32'hbbcf35b2),
	.w5(32'hbb8d1a04),
	.w6(32'hbbb2c191),
	.w7(32'hb918b759),
	.w8(32'hbb92596a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ca6da7),
	.w1(32'h3a80f966),
	.w2(32'hbb0ae2c4),
	.w3(32'hb99858c9),
	.w4(32'h3c0bf0be),
	.w5(32'h3bbddc78),
	.w6(32'hbac72391),
	.w7(32'h3b90eebd),
	.w8(32'h3c08038c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb09765),
	.w1(32'h3be182f2),
	.w2(32'h3bc53627),
	.w3(32'h3b30c228),
	.w4(32'h3b96d84a),
	.w5(32'h3b9c6e20),
	.w6(32'h3bd4a27f),
	.w7(32'h3bc7d01f),
	.w8(32'h3c126cce),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b948a90),
	.w1(32'hb93a8129),
	.w2(32'h3b28f96c),
	.w3(32'h3c17fb52),
	.w4(32'hbb726210),
	.w5(32'hbb5742d3),
	.w6(32'h3b897be1),
	.w7(32'hbb8f2736),
	.w8(32'hbb8dc2fc),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeefa5c),
	.w1(32'hbb12083e),
	.w2(32'hbc1505c4),
	.w3(32'hbb52c494),
	.w4(32'hba63a171),
	.w5(32'hbb79b414),
	.w6(32'h3b805edd),
	.w7(32'hba868543),
	.w8(32'hbb8b0a98),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5af134),
	.w1(32'h3c4228e5),
	.w2(32'h3ac1444d),
	.w3(32'h3c24383a),
	.w4(32'h3c5d479b),
	.w5(32'h3bc46c79),
	.w6(32'h3c81e2f6),
	.w7(32'h3c3276f7),
	.w8(32'h3be4416b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdd98a),
	.w1(32'hbbd0da9f),
	.w2(32'hbc2b4e03),
	.w3(32'h3b460950),
	.w4(32'hbab5d1c9),
	.w5(32'hbc1aa4f6),
	.w6(32'h3b9cee29),
	.w7(32'h39ed9dfe),
	.w8(32'hbba287db),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bd956),
	.w1(32'hbafd7f4f),
	.w2(32'hbba5dcf5),
	.w3(32'hbb460d0a),
	.w4(32'hbb023464),
	.w5(32'hba891652),
	.w6(32'h3a6e5181),
	.w7(32'h3c142034),
	.w8(32'h3bc9fb2f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48ba11),
	.w1(32'hbb763880),
	.w2(32'hbb0bdd1d),
	.w3(32'h3ae59033),
	.w4(32'h3a439fe8),
	.w5(32'h3a8ee8bd),
	.w6(32'h3b774c0b),
	.w7(32'h3ba9a6b4),
	.w8(32'h3b90319e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eefe3a),
	.w1(32'hbab02e1e),
	.w2(32'hbbc007fe),
	.w3(32'h3ae11733),
	.w4(32'hbbbec514),
	.w5(32'hbbb01f8e),
	.w6(32'h3b7b6184),
	.w7(32'hbab5e1da),
	.w8(32'hbbdcbd32),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa69cb),
	.w1(32'hbbaea388),
	.w2(32'hbb0ea06e),
	.w3(32'hbb0d89d8),
	.w4(32'hba37bcfc),
	.w5(32'hbc0e1095),
	.w6(32'h3ab527bc),
	.w7(32'h3aaf6ee5),
	.w8(32'hbc0bee89),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e31b6),
	.w1(32'h3c32fd9e),
	.w2(32'hba5be2a2),
	.w3(32'h3c568980),
	.w4(32'h3c03f4a4),
	.w5(32'hbadf6c7a),
	.w6(32'h3bec1d52),
	.w7(32'h3c0891fa),
	.w8(32'hb9254d0d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ac78c),
	.w1(32'h3bbe74db),
	.w2(32'h3bb10018),
	.w3(32'h3c78d3fd),
	.w4(32'h3be689da),
	.w5(32'hbac901ee),
	.w6(32'h3c887668),
	.w7(32'h3ba63ef9),
	.w8(32'h398a18f5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb109c53),
	.w1(32'h3a44f229),
	.w2(32'h3b04aca5),
	.w3(32'hbc0b9d13),
	.w4(32'h3b410ca9),
	.w5(32'h3c01686b),
	.w6(32'hba8a5504),
	.w7(32'hba469ff4),
	.w8(32'h3b0f5cb6),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a98ab),
	.w1(32'hbb999f1b),
	.w2(32'hbb6182c1),
	.w3(32'h3a9ca2bf),
	.w4(32'hbb4face2),
	.w5(32'h3b3b72f1),
	.w6(32'h3b86fc41),
	.w7(32'hbaa1cc12),
	.w8(32'h3b92e272),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75acd6),
	.w1(32'h3ac5de8d),
	.w2(32'h3a173d37),
	.w3(32'h3b73defd),
	.w4(32'hbbfec8c7),
	.w5(32'hbb88b4bb),
	.w6(32'h3b1d4069),
	.w7(32'hbbafa70c),
	.w8(32'hba0846d3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ea4ab),
	.w1(32'hbbc039a0),
	.w2(32'hbbd40ec5),
	.w3(32'hbb94b953),
	.w4(32'hba007648),
	.w5(32'hbb303c7d),
	.w6(32'h395f3075),
	.w7(32'hbbe2d62e),
	.w8(32'hbc160c55),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc9a78),
	.w1(32'h3a614580),
	.w2(32'hb9d7f558),
	.w3(32'hbbfab124),
	.w4(32'h3b6c0187),
	.w5(32'hbaa9a642),
	.w6(32'hbc07a26f),
	.w7(32'h3bf1cee9),
	.w8(32'h3b9042c2),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f6fab),
	.w1(32'hbb5ee871),
	.w2(32'hbb8a8ad8),
	.w3(32'h3b135169),
	.w4(32'hbae5a5db),
	.w5(32'hba2fe1e2),
	.w6(32'hbaacc8cd),
	.w7(32'hba8ed2ab),
	.w8(32'hbb296cb2),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85ce40),
	.w1(32'hbb6f6287),
	.w2(32'hbb1ff350),
	.w3(32'hba00d36b),
	.w4(32'hba58434e),
	.w5(32'hba9af897),
	.w6(32'h3a99f5fd),
	.w7(32'hba5233b2),
	.w8(32'hbb3e1e14),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad51810),
	.w1(32'hbba2a7cc),
	.w2(32'h39861067),
	.w3(32'h3b1d5b24),
	.w4(32'hbb73180d),
	.w5(32'hb97a91f7),
	.w6(32'h3b586ed7),
	.w7(32'hbb5dd4af),
	.w8(32'hbbd2807e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26f15a),
	.w1(32'hbaecf816),
	.w2(32'hbb373001),
	.w3(32'h3a222fd5),
	.w4(32'h3b1cfef9),
	.w5(32'hb97b1d96),
	.w6(32'hbc244278),
	.w7(32'h3b8d9ab6),
	.w8(32'h3bd5171a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d7dc3),
	.w1(32'h38800b0d),
	.w2(32'h395d05db),
	.w3(32'hba4d1765),
	.w4(32'hbaea762d),
	.w5(32'h3be699bc),
	.w6(32'h3a458b3c),
	.w7(32'hbb9fb403),
	.w8(32'hbbeed34b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfed7bc),
	.w1(32'h3c2d8053),
	.w2(32'h3c1f965d),
	.w3(32'h3cba7d29),
	.w4(32'h3c9509cc),
	.w5(32'hba867726),
	.w6(32'h3c7dda90),
	.w7(32'h3c2ad347),
	.w8(32'hbabe331f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f0114),
	.w1(32'h3c1c8f57),
	.w2(32'hb92e08fb),
	.w3(32'h3b71cdc9),
	.w4(32'h3c5a4387),
	.w5(32'h3a934573),
	.w6(32'h3b89f94c),
	.w7(32'h3c2fccb2),
	.w8(32'h3b91f5fa),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba423772),
	.w1(32'h3a67aaf7),
	.w2(32'hb9ac0aec),
	.w3(32'h3a26856f),
	.w4(32'hba212d56),
	.w5(32'hb98f2417),
	.w6(32'hbb1e1e13),
	.w7(32'hbb352336),
	.w8(32'hbb46773b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0a2bf),
	.w1(32'h3ad91948),
	.w2(32'hbb02b372),
	.w3(32'h3b967804),
	.w4(32'h3ba8ad19),
	.w5(32'hbabb829f),
	.w6(32'h3bb1cb4f),
	.w7(32'h3b141b79),
	.w8(32'h3b1e6f33),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6d850),
	.w1(32'h3ad38d5e),
	.w2(32'h3b08cdc4),
	.w3(32'hbb40df70),
	.w4(32'hbb2fece7),
	.w5(32'hba6da428),
	.w6(32'hbb08e82a),
	.w7(32'hba25bbfc),
	.w8(32'h3b966624),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b9c1b),
	.w1(32'h3b1c9b98),
	.w2(32'hb987716d),
	.w3(32'h3b543b57),
	.w4(32'h3bc94812),
	.w5(32'h3b3e7f31),
	.w6(32'h3b9d526c),
	.w7(32'h3ad3d181),
	.w8(32'hbb24853e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0db65),
	.w1(32'h3bf5fe9d),
	.w2(32'h3bd990ea),
	.w3(32'h3b2f7718),
	.w4(32'h3c207e34),
	.w5(32'h3c290821),
	.w6(32'h3b211d38),
	.w7(32'hba98b348),
	.w8(32'h3b0ec229),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4caa69),
	.w1(32'h3ba3e179),
	.w2(32'hbbb24d54),
	.w3(32'h3c07197f),
	.w4(32'h3c1b695c),
	.w5(32'h3c426754),
	.w6(32'h3be70843),
	.w7(32'hbb481f06),
	.w8(32'hbadeff06),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02a842),
	.w1(32'hbb524a4f),
	.w2(32'hbb4ea43b),
	.w3(32'hbab44ac3),
	.w4(32'hbac935e1),
	.w5(32'hbc5125b5),
	.w6(32'hbafa45ee),
	.w7(32'hbc09a46d),
	.w8(32'hbbcdb990),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b095c08),
	.w1(32'hba5e54e0),
	.w2(32'hbb181ec1),
	.w3(32'h3ab47c88),
	.w4(32'hb8befc03),
	.w5(32'hbbe25cf1),
	.w6(32'h3b76f8ef),
	.w7(32'h3b5a5ad4),
	.w8(32'hbb9a0b91),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f7461),
	.w1(32'h3b93d9d5),
	.w2(32'h3b9895db),
	.w3(32'h3bd36a50),
	.w4(32'h3b8f0196),
	.w5(32'h3b397319),
	.w6(32'h3be6313f),
	.w7(32'h3bbeb4b3),
	.w8(32'h3b505cae),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27b260),
	.w1(32'h3bbc6e8b),
	.w2(32'hbc0019c1),
	.w3(32'h3bf4de9f),
	.w4(32'h3c03343a),
	.w5(32'hbb96b681),
	.w6(32'h3c226a20),
	.w7(32'h3b259ba0),
	.w8(32'hb96ec7d5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45e1d5),
	.w1(32'hbbb6fe19),
	.w2(32'hb9e8a8c2),
	.w3(32'hbb921ae4),
	.w4(32'hbb19a388),
	.w5(32'hb9638452),
	.w6(32'hbc0a8b21),
	.w7(32'hbb4f17af),
	.w8(32'h39275725),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae21f8f),
	.w1(32'h3beca16b),
	.w2(32'hbaad5f31),
	.w3(32'h3b5991ca),
	.w4(32'h3c39f77d),
	.w5(32'hba00243f),
	.w6(32'hba2de471),
	.w7(32'h3c33d5e7),
	.w8(32'h3be7b1b0),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d3d8e),
	.w1(32'h3b1026aa),
	.w2(32'h3a2bbe34),
	.w3(32'hba90efb2),
	.w4(32'h3c090ca0),
	.w5(32'h3b7ad104),
	.w6(32'hbb22385d),
	.w7(32'h3c0c2e6c),
	.w8(32'h3b8dae29),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38c17a),
	.w1(32'h3c09651c),
	.w2(32'h3c0f97e9),
	.w3(32'h3c2c7447),
	.w4(32'h3ac78ef2),
	.w5(32'h3b9da28f),
	.w6(32'h3b606df5),
	.w7(32'hbb1928e2),
	.w8(32'h39b7dc97),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e8d90),
	.w1(32'hbb5305a7),
	.w2(32'hbbba2b7e),
	.w3(32'h3c55ebca),
	.w4(32'hbadf2a47),
	.w5(32'hbbdb1f54),
	.w6(32'h3bb07f0c),
	.w7(32'hbb294525),
	.w8(32'hbc1c676a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb89b2e),
	.w1(32'h3b1d407b),
	.w2(32'hb931c824),
	.w3(32'hbb7cc66c),
	.w4(32'h3c2b3e5a),
	.w5(32'hb952ffab),
	.w6(32'hbb981150),
	.w7(32'h3bcaeb3a),
	.w8(32'h3b46ccc9),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28b5eb),
	.w1(32'h3bd17dc2),
	.w2(32'hbbaaa438),
	.w3(32'hbb495383),
	.w4(32'h3bad77c5),
	.w5(32'h3bc29356),
	.w6(32'h3b7c70c9),
	.w7(32'hb8820329),
	.w8(32'hba41c7f6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5cea6),
	.w1(32'hbb1773ab),
	.w2(32'h3b9bd5e3),
	.w3(32'hbb1aa63c),
	.w4(32'h3af6f40f),
	.w5(32'hbb13da10),
	.w6(32'hbac8c5c8),
	.w7(32'hbb20ce66),
	.w8(32'h39b15a44),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0e39a),
	.w1(32'h3a965e48),
	.w2(32'hba679111),
	.w3(32'hbae7152b),
	.w4(32'h3af6b050),
	.w5(32'hbb80908b),
	.w6(32'hba11338e),
	.w7(32'h3a1182f2),
	.w8(32'h3b5ade6b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c95f4),
	.w1(32'h3c2265ba),
	.w2(32'h3c1f7843),
	.w3(32'hbac78f1b),
	.w4(32'h3c1fc93a),
	.w5(32'h3c56ca76),
	.w6(32'h3afa672c),
	.w7(32'h3b9452c3),
	.w8(32'h3bf7338c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39fd1a),
	.w1(32'h3be917f9),
	.w2(32'h3b4d3cd3),
	.w3(32'h3b92c076),
	.w4(32'h3c88df28),
	.w5(32'h3b9e670c),
	.w6(32'h3b8380af),
	.w7(32'h3bd33273),
	.w8(32'h3be1cf92),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ab015),
	.w1(32'h3b1dba1b),
	.w2(32'hba066304),
	.w3(32'h3c16027f),
	.w4(32'h3b96f3d7),
	.w5(32'hbab5d247),
	.w6(32'h3c3a9ea5),
	.w7(32'h3bcd937e),
	.w8(32'h3b3a0719),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ae2482),
	.w1(32'hbb56baee),
	.w2(32'h3aeaa213),
	.w3(32'hbac9f9ce),
	.w4(32'hbbc9b853),
	.w5(32'hba411f15),
	.w6(32'hb9cfc51c),
	.w7(32'hbb530752),
	.w8(32'hbb62c038),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd339c1),
	.w1(32'h3ba1ed63),
	.w2(32'hbb78f7ab),
	.w3(32'h3b63cdba),
	.w4(32'hb966b959),
	.w5(32'hbbe66966),
	.w6(32'hbbc1263f),
	.w7(32'hba2166cf),
	.w8(32'h3a972450),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule