module layer_10_featuremap_118(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ffc045),
	.w1(32'hb9a8f846),
	.w2(32'hba8dfc96),
	.w3(32'h3910bad1),
	.w4(32'hb8244d00),
	.w5(32'hb983421f),
	.w6(32'hb933c486),
	.w7(32'h395b326e),
	.w8(32'h3a14326d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87a2549),
	.w1(32'h3a38bd29),
	.w2(32'hba240371),
	.w3(32'hba32cbc6),
	.w4(32'h393d4de8),
	.w5(32'hbac29b4c),
	.w6(32'h3925a0ae),
	.w7(32'hb9c7360f),
	.w8(32'hbab32394),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a4366a),
	.w1(32'hb9dce44f),
	.w2(32'hba852f2c),
	.w3(32'hb7ea0628),
	.w4(32'hba104cbf),
	.w5(32'hba869acb),
	.w6(32'hb9bdb48b),
	.w7(32'hba549214),
	.w8(32'hba22fb1f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64110b),
	.w1(32'hba96bbd1),
	.w2(32'hbaa1174c),
	.w3(32'hbaa97af0),
	.w4(32'hb92b4258),
	.w5(32'hba8451b6),
	.w6(32'h37e4f816),
	.w7(32'h38cf5ba0),
	.w8(32'h3a456db5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a7abf),
	.w1(32'hb736fe01),
	.w2(32'h3a335a06),
	.w3(32'hba3f7596),
	.w4(32'h3983973c),
	.w5(32'h392feed9),
	.w6(32'h39ac81e3),
	.w7(32'h39535745),
	.w8(32'h3795eae0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91956b9),
	.w1(32'h399a5b94),
	.w2(32'h39f04dd7),
	.w3(32'hb70c8210),
	.w4(32'h39ba9b28),
	.w5(32'h39ea96ee),
	.w6(32'h39c38407),
	.w7(32'h3a10145e),
	.w8(32'h39e82003),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed1f5c),
	.w1(32'hbb85cfad),
	.w2(32'hba4c2280),
	.w3(32'h39a1ae1b),
	.w4(32'hbb107ca4),
	.w5(32'hb98dbba7),
	.w6(32'hbabf1a05),
	.w7(32'hbbaf064c),
	.w8(32'hbb34dd89),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a4c05),
	.w1(32'hbbc5e9c4),
	.w2(32'h3ac0931b),
	.w3(32'hbc6e3c99),
	.w4(32'hbbffced9),
	.w5(32'hbbcb3e36),
	.w6(32'hbc3a4289),
	.w7(32'hbba4b52f),
	.w8(32'hbb77fb0a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e5c1c),
	.w1(32'hb9eb98e6),
	.w2(32'hb9839dd6),
	.w3(32'hba523f5d),
	.w4(32'hb9adf926),
	.w5(32'hb824777d),
	.w6(32'hba38a40b),
	.w7(32'hb9b592d0),
	.w8(32'hb8a93ade),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4ef77),
	.w1(32'hb8f2ac52),
	.w2(32'h3bb5f33a),
	.w3(32'hbb8e7588),
	.w4(32'h3af7ba7f),
	.w5(32'h3bc55892),
	.w6(32'hbb435c13),
	.w7(32'hb904ca86),
	.w8(32'h3b3b3add),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38352f7b),
	.w1(32'hb9923b2a),
	.w2(32'hb9df8d86),
	.w3(32'hb8f300c7),
	.w4(32'h3928a907),
	.w5(32'h39621e72),
	.w6(32'hb97d1756),
	.w7(32'hb9b71abf),
	.w8(32'h39416407),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab85321),
	.w1(32'hbb766edf),
	.w2(32'hbb0124a6),
	.w3(32'h3abec860),
	.w4(32'h3aad4d75),
	.w5(32'h3b0aaf80),
	.w6(32'hba68c5e7),
	.w7(32'hbacdc7d5),
	.w8(32'h37ad9a90),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf10816),
	.w1(32'hbb02d4d1),
	.w2(32'h3b92daf2),
	.w3(32'hbb9da227),
	.w4(32'hba208d8f),
	.w5(32'h3ba28ae2),
	.w6(32'hbb251397),
	.w7(32'hba374ebe),
	.w8(32'h3b175fcf),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d219ed),
	.w1(32'hba407b2c),
	.w2(32'hb9c56965),
	.w3(32'hb966e070),
	.w4(32'h39203afe),
	.w5(32'h3a1fed20),
	.w6(32'h39503817),
	.w7(32'h39771a19),
	.w8(32'hba2d52d1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bd5ca),
	.w1(32'hb8d8a9e1),
	.w2(32'hb9b9cee6),
	.w3(32'hbac162f4),
	.w4(32'hb9fd3291),
	.w5(32'hb933b921),
	.w6(32'hbaf2426c),
	.w7(32'hba08ca8a),
	.w8(32'hba60a793),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba98f1),
	.w1(32'h3a424096),
	.w2(32'h3b4e0f02),
	.w3(32'hbbcc1ecf),
	.w4(32'h3a2b0278),
	.w5(32'h3b907427),
	.w6(32'hbbae1290),
	.w7(32'hb99bcf96),
	.w8(32'h3a9a8e93),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62ae6c3),
	.w1(32'h398f499c),
	.w2(32'h3a9ae5af),
	.w3(32'h38a4897e),
	.w4(32'hb9bd2359),
	.w5(32'h3a38ad47),
	.w6(32'hb9904126),
	.w7(32'h3a86ee94),
	.w8(32'h39f80219),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3f217),
	.w1(32'hbb5d6ec1),
	.w2(32'h3b8244b0),
	.w3(32'hbbc67b65),
	.w4(32'h39061627),
	.w5(32'h3b6fd7b1),
	.w6(32'hbb585964),
	.w7(32'h398fc5ab),
	.w8(32'h3b640ffa),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91ca69),
	.w1(32'hba8c2fec),
	.w2(32'h3b380f6a),
	.w3(32'hbb69b654),
	.w4(32'h38a93240),
	.w5(32'h3b2927ff),
	.w6(32'hbaf4c126),
	.w7(32'hba2c262e),
	.w8(32'h3a9d53a3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ffe1ab),
	.w1(32'hb981dc89),
	.w2(32'h39455dba),
	.w3(32'hb9db8844),
	.w4(32'hb7da9227),
	.w5(32'h37c3205a),
	.w6(32'hb91e9a21),
	.w7(32'h389c4c57),
	.w8(32'hb8920f10),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83490ab),
	.w1(32'hb8ab375f),
	.w2(32'hb9bc024e),
	.w3(32'h381e4b12),
	.w4(32'hb9ba92ae),
	.w5(32'hba0478fd),
	.w6(32'hb936c1db),
	.w7(32'hb985be41),
	.w8(32'hb8f930a6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a033867),
	.w1(32'hb9a9e212),
	.w2(32'hbadad0c4),
	.w3(32'hb8517600),
	.w4(32'h3a14d769),
	.w5(32'hba223490),
	.w6(32'h39cd4300),
	.w7(32'hb9badb30),
	.w8(32'hb9dc8a8a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc371277),
	.w1(32'hbbc5b671),
	.w2(32'h39b51892),
	.w3(32'hbc06e31f),
	.w4(32'hbb8338cd),
	.w5(32'h3ba0ad79),
	.w6(32'hbc25776b),
	.w7(32'hbb887e73),
	.w8(32'h3b0c1150),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a1755),
	.w1(32'h3b0225f0),
	.w2(32'h3ba57eda),
	.w3(32'hbb578714),
	.w4(32'hb836a08d),
	.w5(32'h3b3f9675),
	.w6(32'hbaae3cf8),
	.w7(32'h3adcf8d9),
	.w8(32'h3b432a15),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81bfb4),
	.w1(32'h3b960f31),
	.w2(32'h3aeb2645),
	.w3(32'hba13a0eb),
	.w4(32'hba43bcf0),
	.w5(32'hbababe6b),
	.w6(32'h398bc2d6),
	.w7(32'h3af43050),
	.w8(32'h39c433c2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e21bae),
	.w1(32'h38bb4512),
	.w2(32'h3a9b6e60),
	.w3(32'hb98bbbde),
	.w4(32'hb98712c6),
	.w5(32'h386f7d99),
	.w6(32'hb9e78b27),
	.w7(32'h39a0cb70),
	.w8(32'h39fa34d6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de8289),
	.w1(32'hb956b6f8),
	.w2(32'h3924e5d9),
	.w3(32'hb9b0da77),
	.w4(32'hb9206281),
	.w5(32'hb820fbe2),
	.w6(32'hb8b4f0c9),
	.w7(32'h38f19e37),
	.w8(32'hb6f7e839),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaeb64),
	.w1(32'hbaf7264e),
	.w2(32'h3b05be9d),
	.w3(32'hbbeb8a36),
	.w4(32'h3991d70d),
	.w5(32'h3bab5142),
	.w6(32'hbb8d1647),
	.w7(32'hba8509a4),
	.w8(32'h3b718c4e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e6cb2),
	.w1(32'h392c16de),
	.w2(32'hba017989),
	.w3(32'h3a6b6aca),
	.w4(32'h3a86f5c7),
	.w5(32'hb886cf28),
	.w6(32'h3aa2fda9),
	.w7(32'h3aca437a),
	.w8(32'h3aa258b4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba735e3d),
	.w1(32'h3b1f033a),
	.w2(32'h3babd2e9),
	.w3(32'hbb84c48a),
	.w4(32'h3aa3ae8d),
	.w5(32'h3acee232),
	.w6(32'hba6cfc19),
	.w7(32'h3ad2bbf0),
	.w8(32'h3ac2e6ad),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38acc9fd),
	.w1(32'h387e8b81),
	.w2(32'hb80c78d9),
	.w3(32'hb915cf82),
	.w4(32'hb8ca95db),
	.w5(32'hb8304316),
	.w6(32'h3811b824),
	.w7(32'hb84764f6),
	.w8(32'hb706d925),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38969ffb),
	.w1(32'hb96ce18e),
	.w2(32'hb8b53a07),
	.w3(32'hb71080e2),
	.w4(32'hb9246e92),
	.w5(32'hb7f6e71d),
	.w6(32'hb9902c80),
	.w7(32'hb87c2817),
	.w8(32'h3805594b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf233b4),
	.w1(32'hb9179f8b),
	.w2(32'h3b77bfab),
	.w3(32'hbae5c264),
	.w4(32'h3a2999fb),
	.w5(32'h3b3a05ab),
	.w6(32'hba8a5496),
	.w7(32'h3a0dce76),
	.w8(32'h3a64cd2b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb810d244),
	.w1(32'hb9c1bd58),
	.w2(32'hb9c4f290),
	.w3(32'hba2f397c),
	.w4(32'hba21c807),
	.w5(32'hba8393d6),
	.w6(32'hb6059210),
	.w7(32'h39deb6b7),
	.w8(32'hba9978e4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8876d),
	.w1(32'hb9e9ab23),
	.w2(32'h3976d8f6),
	.w3(32'hba6585c0),
	.w4(32'h37da6f44),
	.w5(32'h3a31dbaa),
	.w6(32'hb9798468),
	.w7(32'hb93b9ba1),
	.w8(32'h3a2359e0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2a43c),
	.w1(32'hbb0819e3),
	.w2(32'hb9ec194e),
	.w3(32'hbaf24df4),
	.w4(32'hbb522cc9),
	.w5(32'hba96201e),
	.w6(32'hbadea820),
	.w7(32'hbab7416c),
	.w8(32'h3abfa0d5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb66ff),
	.w1(32'hbc167c1d),
	.w2(32'hbc09f93f),
	.w3(32'hbc03eba3),
	.w4(32'hbaa8abe0),
	.w5(32'h3b2755a7),
	.w6(32'hbafbea26),
	.w7(32'hbaa3ac36),
	.w8(32'hba1140d4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6093ab),
	.w1(32'h3ae09f27),
	.w2(32'hbaa9d718),
	.w3(32'h3994c5be),
	.w4(32'hb8917056),
	.w5(32'hbb8c8853),
	.w6(32'h3991459a),
	.w7(32'hbabba85d),
	.w8(32'hbb6a2e94),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7030e2),
	.w1(32'h3b8838a2),
	.w2(32'h3ae79dc4),
	.w3(32'h3a445d0c),
	.w4(32'hb9db6b05),
	.w5(32'hbbaa7f29),
	.w6(32'h3a9e25c5),
	.w7(32'hb9a3749f),
	.w8(32'hbb8fa642),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399840da),
	.w1(32'h39730614),
	.w2(32'hb94b92c8),
	.w3(32'hb96ecb43),
	.w4(32'hb9da31a5),
	.w5(32'hba6ea93c),
	.w6(32'hb9f06077),
	.w7(32'hba054966),
	.w8(32'hba6cb979),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba521738),
	.w1(32'hb94d3856),
	.w2(32'h398b92c2),
	.w3(32'hba17f06d),
	.w4(32'hb8901c4f),
	.w5(32'h3994c5c6),
	.w6(32'hb971d5b4),
	.w7(32'h398ef72d),
	.w8(32'hb9847a25),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed4b48),
	.w1(32'hba34469f),
	.w2(32'hba281fd1),
	.w3(32'hb9e09f5b),
	.w4(32'hb9907b61),
	.w5(32'hba08c31c),
	.w6(32'hb9ce7eec),
	.w7(32'hb9f2270c),
	.w8(32'hb9ebd069),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74b71b0),
	.w1(32'hb9c4cdb0),
	.w2(32'h39c45357),
	.w3(32'hb9c5a247),
	.w4(32'hb9496855),
	.w5(32'h39e49466),
	.w6(32'hb9a806fe),
	.w7(32'hb9ac0f33),
	.w8(32'h38511aca),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc219e13),
	.w1(32'h3b6ebe00),
	.w2(32'h3c002643),
	.w3(32'hbbc920ce),
	.w4(32'h3bd946b7),
	.w5(32'h3c2efbbb),
	.w6(32'hbb72fc17),
	.w7(32'h3ba06078),
	.w8(32'h3bd44750),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ffcd1),
	.w1(32'h3b0a2d4d),
	.w2(32'h3b5b0715),
	.w3(32'hbb0693bf),
	.w4(32'h39fd9e10),
	.w5(32'h3b2781ee),
	.w6(32'hbab6a2d3),
	.w7(32'h3a56af51),
	.w8(32'h3a113773),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3329af),
	.w1(32'h3affecaa),
	.w2(32'h3bbe912a),
	.w3(32'hbb76fc94),
	.w4(32'h388a15e7),
	.w5(32'h3b06fa27),
	.w6(32'hbae67cd8),
	.w7(32'h3ab75710),
	.w8(32'h3b4edcff),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba67530),
	.w1(32'hbaa8f345),
	.w2(32'h39bd6429),
	.w3(32'hbb908623),
	.w4(32'hb904c580),
	.w5(32'h3accfe93),
	.w6(32'hbb3996b4),
	.w7(32'hb8d167ef),
	.w8(32'h3999ff5e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc127bb5),
	.w1(32'hbb8f37c6),
	.w2(32'h3b463052),
	.w3(32'hbbc73d80),
	.w4(32'hba80fa60),
	.w5(32'h3ba00410),
	.w6(32'hbb62f5f6),
	.w7(32'hba0a74ea),
	.w8(32'h3b702c4b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aaf23a),
	.w1(32'hb981da9d),
	.w2(32'hb90732dc),
	.w3(32'hb848ef7b),
	.w4(32'h39569185),
	.w5(32'hb98fd22b),
	.w6(32'h391d0888),
	.w7(32'h39a77050),
	.w8(32'hb9bff60c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3757d4),
	.w1(32'hb98973d6),
	.w2(32'hba430edf),
	.w3(32'h38b58b9d),
	.w4(32'hb8255840),
	.w5(32'hb9ea0097),
	.w6(32'hb8058cb0),
	.w7(32'hb9f982c2),
	.w8(32'hba4f1afd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11a38c),
	.w1(32'h384600e3),
	.w2(32'hba8620d8),
	.w3(32'h3ab1080e),
	.w4(32'h399e6264),
	.w5(32'hba5f6e8e),
	.w6(32'h3a389690),
	.w7(32'h398af830),
	.w8(32'hb9cdd9ab),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb804096),
	.w1(32'hbaffc039),
	.w2(32'h3acfc37a),
	.w3(32'hbb78da48),
	.w4(32'hbac43edb),
	.w5(32'h3a9caaf3),
	.w6(32'hbb615d7a),
	.w7(32'hba9352d3),
	.w8(32'h3a26f5c5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b2abe),
	.w1(32'hb63ba6f3),
	.w2(32'h3a990162),
	.w3(32'hba84fbd5),
	.w4(32'h39def12f),
	.w5(32'h3a8bcfdd),
	.w6(32'h36fcc6df),
	.w7(32'h3a51878b),
	.w8(32'h3a61b612),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba910cd),
	.w1(32'hbb0c11a7),
	.w2(32'h3b826418),
	.w3(32'hbb90f6b5),
	.w4(32'h3a7670b1),
	.w5(32'h3b96be69),
	.w6(32'hbb089388),
	.w7(32'h3a741622),
	.w8(32'h3b6f839f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba595973),
	.w1(32'h3a747908),
	.w2(32'h3b1a987b),
	.w3(32'hba7ec031),
	.w4(32'hb7dd13ba),
	.w5(32'h3a0b3f6c),
	.w6(32'h397654e5),
	.w7(32'h3ac55435),
	.w8(32'h3a85b90b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917278a),
	.w1(32'h394dfbc6),
	.w2(32'h386b3a20),
	.w3(32'h3867926e),
	.w4(32'h38e3ef9c),
	.w5(32'h38395b05),
	.w6(32'hb74d9eb4),
	.w7(32'h39ff695b),
	.w8(32'hb881aab4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93cd1b5),
	.w1(32'hb9c36bb3),
	.w2(32'hb9fbad42),
	.w3(32'h39f9df37),
	.w4(32'hb98a79e7),
	.w5(32'hba0672d4),
	.w6(32'hb9d8924f),
	.w7(32'hba7126ae),
	.w8(32'hba85f446),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a50d7),
	.w1(32'hba5a3564),
	.w2(32'h39cb9691),
	.w3(32'hba1d0f02),
	.w4(32'hbaa3304c),
	.w5(32'hbaaf81a3),
	.w6(32'hba3de793),
	.w7(32'hba27fbd3),
	.w8(32'h3a2733c0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b722cd),
	.w1(32'hb7a7965b),
	.w2(32'h3990cf1f),
	.w3(32'hb86d25f8),
	.w4(32'h37ed7ec9),
	.w5(32'h38926ba8),
	.w6(32'hb98e2584),
	.w7(32'hb6ea7c1a),
	.w8(32'h38711b52),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1bc91),
	.w1(32'h39b0aacc),
	.w2(32'h3a5551e5),
	.w3(32'hba36ea60),
	.w4(32'hb95a8ce6),
	.w5(32'h39cbd9cb),
	.w6(32'hb832f19d),
	.w7(32'h39850f5e),
	.w8(32'h3a14482c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51fc83),
	.w1(32'hba5175ae),
	.w2(32'h3aa3576d),
	.w3(32'hbb1fc68f),
	.w4(32'hb91149a1),
	.w5(32'h3a69568e),
	.w6(32'hbadd218a),
	.w7(32'hb80df0ca),
	.w8(32'h3a131d04),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb991047),
	.w1(32'h3b0f1ef7),
	.w2(32'h3b850d75),
	.w3(32'hbb96765a),
	.w4(32'h3afa5116),
	.w5(32'h3b84f779),
	.w6(32'hbb197187),
	.w7(32'h3b0f755b),
	.w8(32'h3a69ceaf),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b79659),
	.w1(32'hba2f3e8b),
	.w2(32'h39f91de1),
	.w3(32'h3906e873),
	.w4(32'hba759739),
	.w5(32'h398c55a6),
	.w6(32'hba621b5d),
	.w7(32'hb9b8c69c),
	.w8(32'hba93d48e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5c4d2),
	.w1(32'h38ccca76),
	.w2(32'h3964da66),
	.w3(32'hbaa936ca),
	.w4(32'h39b71c32),
	.w5(32'h3886797d),
	.w6(32'h39ce1e0f),
	.w7(32'h399228c9),
	.w8(32'h3a31c5c4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efae27),
	.w1(32'h38eca47d),
	.w2(32'hb962e91b),
	.w3(32'h391c05de),
	.w4(32'h37f81982),
	.w5(32'hb932c289),
	.w6(32'h392c6573),
	.w7(32'hb92fc21b),
	.w8(32'hb99e8e40),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f3f59),
	.w1(32'hbaaf2cb1),
	.w2(32'h39f08fd1),
	.w3(32'hb98314e5),
	.w4(32'hba824470),
	.w5(32'hba404f2c),
	.w6(32'hba7a058b),
	.w7(32'hba2a9445),
	.w8(32'hb81ef0d5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc282dc7),
	.w1(32'hbb893b13),
	.w2(32'h3a823274),
	.w3(32'hbbb03f53),
	.w4(32'h3b8fcfd6),
	.w5(32'h3c24cb0d),
	.w6(32'hbbe7a1a8),
	.w7(32'hbb46bdc3),
	.w8(32'hbb09f582),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb317d49),
	.w1(32'h3b0299b8),
	.w2(32'h3bd69001),
	.w3(32'hbbba3956),
	.w4(32'hbb91dc7b),
	.w5(32'hbb417388),
	.w6(32'hbb0d7868),
	.w7(32'h3b503d14),
	.w8(32'h3b5d557e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40c8ed),
	.w1(32'h3ad5ddc3),
	.w2(32'h3b3340b3),
	.w3(32'hbb8df991),
	.w4(32'hb7e9fc57),
	.w5(32'h3ade342e),
	.w6(32'hbae1a79a),
	.w7(32'h3b123ae6),
	.w8(32'h3b6042fe),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afff8d7),
	.w1(32'h3b2afe3f),
	.w2(32'h3ad107e5),
	.w3(32'hbb60c234),
	.w4(32'hbb06d127),
	.w5(32'hbb49a7a3),
	.w6(32'hbb8b964d),
	.w7(32'hba40e72a),
	.w8(32'h39ee3e10),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d53310),
	.w1(32'hba085a90),
	.w2(32'hb8cfc838),
	.w3(32'hb9510129),
	.w4(32'hb980b76b),
	.w5(32'hb969f39c),
	.w6(32'hb9ad362e),
	.w7(32'hb9a2868f),
	.w8(32'hb84b634b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d1ef99),
	.w1(32'hb958c5de),
	.w2(32'hb98a0041),
	.w3(32'hb92502ce),
	.w4(32'hb98bb402),
	.w5(32'hb8c8cff3),
	.w6(32'hb8397a9a),
	.w7(32'hb9650c48),
	.w8(32'hb83dfd52),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fa7657),
	.w1(32'hb786aec1),
	.w2(32'hb8a5273b),
	.w3(32'h38d3dce4),
	.w4(32'hb929a635),
	.w5(32'hb849aaa8),
	.w6(32'hb886fd77),
	.w7(32'hb797bb6f),
	.w8(32'h3856f63f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf559c3),
	.w1(32'hba3a2c3b),
	.w2(32'h392eeb08),
	.w3(32'hbacdb2bd),
	.w4(32'hb9faa151),
	.w5(32'hb8b79336),
	.w6(32'hba85462e),
	.w7(32'hb8e4f57b),
	.w8(32'hb961edfd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9090b68),
	.w1(32'hb9888743),
	.w2(32'hb8dc01a6),
	.w3(32'hb8372896),
	.w4(32'hb66a1623),
	.w5(32'h39027b01),
	.w6(32'h392dc17d),
	.w7(32'h38fbf414),
	.w8(32'h390cb97d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bc0df),
	.w1(32'hbaf8b6bf),
	.w2(32'h38ce949d),
	.w3(32'hbb1ee492),
	.w4(32'hba1b371d),
	.w5(32'h3b2a6ba1),
	.w6(32'hbb3b59a6),
	.w7(32'hbb069767),
	.w8(32'hba15a5a4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9efe30),
	.w1(32'hbb988b98),
	.w2(32'h39c836a9),
	.w3(32'hbbab5c0e),
	.w4(32'hbb88f897),
	.w5(32'h394eacde),
	.w6(32'hbb962d41),
	.w7(32'hbb361600),
	.w8(32'h3a9d448f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94afd9),
	.w1(32'h39be2d3f),
	.w2(32'h3aaab130),
	.w3(32'hbadf205a),
	.w4(32'hb98f4cfe),
	.w5(32'h3a86c677),
	.w6(32'hba4535f6),
	.w7(32'h391d3cea),
	.w8(32'hba0200c3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a642e),
	.w1(32'h3896696a),
	.w2(32'h3b387ea0),
	.w3(32'hbb16ebfa),
	.w4(32'h379456a9),
	.w5(32'h3a96bf91),
	.w6(32'hbab6db0f),
	.w7(32'h391ff162),
	.w8(32'hb9e636da),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7beae8),
	.w1(32'hbb5fe9e1),
	.w2(32'h3a4adf12),
	.w3(32'hbae7551b),
	.w4(32'hba960dfd),
	.w5(32'h3b77bb76),
	.w6(32'hbb18e23e),
	.w7(32'hbb351478),
	.w8(32'hb920c93c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f7ea8),
	.w1(32'h3b0cfbc3),
	.w2(32'h3b1163d4),
	.w3(32'hbab7d18c),
	.w4(32'h3af2dfbb),
	.w5(32'h3b3ca4da),
	.w6(32'hba93a0d6),
	.w7(32'h3b0f5175),
	.w8(32'h3aa0e6e9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ba66e),
	.w1(32'hba7cb940),
	.w2(32'h3ab85354),
	.w3(32'hbb0e4322),
	.w4(32'h3a01241e),
	.w5(32'h3b2f819d),
	.w6(32'hba8ea0ec),
	.w7(32'hb9cbb721),
	.w8(32'h3a93e4cf),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb930529b),
	.w1(32'h384e9988),
	.w2(32'h3949f8d7),
	.w3(32'hb9957905),
	.w4(32'h39337642),
	.w5(32'h38b0fea3),
	.w6(32'h3942a946),
	.w7(32'h399c0447),
	.w8(32'h395a809a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba1d81),
	.w1(32'h38f53475),
	.w2(32'h3868e8fa),
	.w3(32'hb7a4d1db),
	.w4(32'h38ba293c),
	.w5(32'h39a86b8b),
	.w6(32'h38fc9d3e),
	.w7(32'h394961ef),
	.w8(32'hb9113c99),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d5bfe),
	.w1(32'h39e21712),
	.w2(32'h38ff3ab2),
	.w3(32'hb94c2c54),
	.w4(32'h3a58eec2),
	.w5(32'h3a4f55aa),
	.w6(32'h386ffb3f),
	.w7(32'h396d5741),
	.w8(32'h398e0c0e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21cbd9),
	.w1(32'h39993915),
	.w2(32'h388a9793),
	.w3(32'h3a062984),
	.w4(32'h39c04c3f),
	.w5(32'hb98be604),
	.w6(32'h3992942d),
	.w7(32'hb903921f),
	.w8(32'hba0f8906),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c49346),
	.w1(32'h3a35da5e),
	.w2(32'hba9e89bc),
	.w3(32'hbad7a526),
	.w4(32'hba34f12f),
	.w5(32'hbb37657b),
	.w6(32'hb9148739),
	.w7(32'hb68ff92d),
	.w8(32'hbb46bffb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2dc758),
	.w1(32'hb9977c9e),
	.w2(32'hb87fd1eb),
	.w3(32'hba64a324),
	.w4(32'hba1349f8),
	.w5(32'hb9b7f030),
	.w6(32'hb8e8947d),
	.w7(32'hb947a901),
	.w8(32'hb7be3184),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48d96f),
	.w1(32'h3b04d85e),
	.w2(32'h3b30281a),
	.w3(32'hba44cf40),
	.w4(32'hb92610a4),
	.w5(32'h39d4d872),
	.w6(32'hb9096e11),
	.w7(32'h3aca4b2a),
	.w8(32'h3a5f7efb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98cf7e),
	.w1(32'h3b1a6f90),
	.w2(32'h3b70ed7c),
	.w3(32'hb91db0da),
	.w4(32'h39c9a4be),
	.w5(32'h3b221644),
	.w6(32'hb89418cb),
	.w7(32'h39e8c8ad),
	.w8(32'h3b0a2234),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2025d),
	.w1(32'h3a9db69c),
	.w2(32'h38d0d691),
	.w3(32'h3961ff18),
	.w4(32'h39559e44),
	.w5(32'hba876205),
	.w6(32'h3a85bab2),
	.w7(32'hb89a92c0),
	.w8(32'hb84facdd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0da691),
	.w1(32'hbbac78e4),
	.w2(32'h3a6f12d3),
	.w3(32'hbb5ef0b5),
	.w4(32'h3b38b098),
	.w5(32'h3bf58731),
	.w6(32'hbbee2df6),
	.w7(32'hbbb740f9),
	.w8(32'hba03fcd2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca3115),
	.w1(32'h3a12781e),
	.w2(32'h3b27d703),
	.w3(32'hbb0823e9),
	.w4(32'hbb1d7425),
	.w5(32'h3a55b31c),
	.w6(32'hbb0aa93f),
	.w7(32'hbb0f56fb),
	.w8(32'h3a30b325),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb312a51),
	.w1(32'h39c3ab3c),
	.w2(32'h3b4adbf0),
	.w3(32'hbb07deea),
	.w4(32'h3ac22ad6),
	.w5(32'h3b9206ae),
	.w6(32'hbb00f4cc),
	.w7(32'h3a705f44),
	.w8(32'h3996d50c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6999ef),
	.w1(32'h3a2c80b9),
	.w2(32'h3ab0ea67),
	.w3(32'hb9ebaf77),
	.w4(32'h3ae32d15),
	.w5(32'h3b46398a),
	.w6(32'hba094ea4),
	.w7(32'hba5c0b17),
	.w8(32'hbaa5a952),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc19b4),
	.w1(32'h3a22d6e4),
	.w2(32'h3a4beb4b),
	.w3(32'hbb1a89a9),
	.w4(32'hb9adf413),
	.w5(32'hb9767d49),
	.w6(32'h3907728c),
	.w7(32'hb9d8bd08),
	.w8(32'hba8fe0f8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d8af3),
	.w1(32'h3a6255c0),
	.w2(32'hb9f82d2a),
	.w3(32'h3a59c7f0),
	.w4(32'h3a93cc38),
	.w5(32'hb8dedf3a),
	.w6(32'h3a5801fd),
	.w7(32'hba1834b9),
	.w8(32'hb88b1292),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c830d),
	.w1(32'hba859a16),
	.w2(32'h3b428f6b),
	.w3(32'hbb808aa1),
	.w4(32'hb8d21d32),
	.w5(32'h3b228562),
	.w6(32'hbb1f39d7),
	.w7(32'hba87b6c9),
	.w8(32'h3ab38814),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb474c7),
	.w1(32'hbb8493e7),
	.w2(32'h3a0fea2e),
	.w3(32'hbb073baa),
	.w4(32'h3b050f8a),
	.w5(32'h3bd6fc00),
	.w6(32'hbb386854),
	.w7(32'hbb135f9b),
	.w8(32'hbaa48295),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb406fd1),
	.w1(32'hbaf9f041),
	.w2(32'hbb7343c1),
	.w3(32'hbc1b7fa7),
	.w4(32'hbb593c3b),
	.w5(32'h3a86ff8d),
	.w6(32'hbb4d55fb),
	.w7(32'h3ad8d01d),
	.w8(32'h3bf235d4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e7546),
	.w1(32'hbb08d6e4),
	.w2(32'hbabf61d6),
	.w3(32'hba909698),
	.w4(32'hbb619e94),
	.w5(32'hbb7f9e2c),
	.w6(32'hbad3353b),
	.w7(32'hbb14cbe6),
	.w8(32'hbb1c6611),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e6e35),
	.w1(32'h3b897e68),
	.w2(32'h3bd906b7),
	.w3(32'hbafe74f7),
	.w4(32'h3a06f6bd),
	.w5(32'h3af4bda3),
	.w6(32'hb88ad3f8),
	.w7(32'h3b13fd05),
	.w8(32'h3af3d46b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0c7aa),
	.w1(32'hbbd96249),
	.w2(32'hb925f1f8),
	.w3(32'hbb393334),
	.w4(32'h3a925b79),
	.w5(32'h3c026d2c),
	.w6(32'hbb73c20b),
	.w7(32'hbac4d1a7),
	.w8(32'h3b17c46c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0d4d0),
	.w1(32'h3ae60c27),
	.w2(32'hba0f3536),
	.w3(32'h3aea11cc),
	.w4(32'h3b1eaf0f),
	.w5(32'h3ac29bdb),
	.w6(32'h3aa1ef68),
	.w7(32'h3ab9f19a),
	.w8(32'h3a98fbd0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f1fd6),
	.w1(32'hbb14888d),
	.w2(32'hbbe1281b),
	.w3(32'hbc4cbfb4),
	.w4(32'h3af3620e),
	.w5(32'hbae8189a),
	.w6(32'hbb1da04b),
	.w7(32'hbad73ec1),
	.w8(32'hbb0d772d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba813a1b),
	.w1(32'hbb2c19a7),
	.w2(32'h39ebe15b),
	.w3(32'h37b53d34),
	.w4(32'h3a5cad35),
	.w5(32'h3adbaeba),
	.w6(32'hbb0f56ba),
	.w7(32'h38f57ee6),
	.w8(32'h394f2bd8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb932991e),
	.w1(32'hb9afed06),
	.w2(32'hba82a53b),
	.w3(32'hb81c714f),
	.w4(32'hb9c406b7),
	.w5(32'hba0e4946),
	.w6(32'hb8d31f36),
	.w7(32'hba1b3ba7),
	.w8(32'hba3f6ce3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba984a62),
	.w1(32'h3a405b7a),
	.w2(32'hb984ac15),
	.w3(32'hba2da0d2),
	.w4(32'h3a1cd7a8),
	.w5(32'h3a35b06d),
	.w6(32'hb9c90248),
	.w7(32'hb9431810),
	.w8(32'h39a93e43),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dd302),
	.w1(32'h3b0a50bb),
	.w2(32'h3b97a177),
	.w3(32'hbafc641c),
	.w4(32'h3afae5c1),
	.w5(32'h3b80dda9),
	.w6(32'hba02aa44),
	.w7(32'h3aa3f581),
	.w8(32'h3b092ae7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67bcae),
	.w1(32'h3b0d3a50),
	.w2(32'h3aa5d114),
	.w3(32'hb943c559),
	.w4(32'h39f3b226),
	.w5(32'hba4b3233),
	.w6(32'hba0a4662),
	.w7(32'hb96e89ca),
	.w8(32'hbae8b913),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96cbeb),
	.w1(32'hb9e1e300),
	.w2(32'hba22264c),
	.w3(32'hbb8e690c),
	.w4(32'hba2a7985),
	.w5(32'hbb0be8a4),
	.w6(32'hbaa3c15d),
	.w7(32'hb8e3ac68),
	.w8(32'hb9b7dcdc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32b577),
	.w1(32'hba035d41),
	.w2(32'h39cd2148),
	.w3(32'hba7a7fa1),
	.w4(32'h39303e70),
	.w5(32'h3a758e25),
	.w6(32'hb9e7af72),
	.w7(32'h3964445a),
	.w8(32'hba4d361a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae39231),
	.w1(32'h3b3aa91b),
	.w2(32'h3b47be74),
	.w3(32'hbaa99102),
	.w4(32'hba4e858e),
	.w5(32'h3b1c98b5),
	.w6(32'hbafeb7bb),
	.w7(32'h3b09a5a1),
	.w8(32'h3bb7fbe4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0462b8),
	.w1(32'h3aec1bb4),
	.w2(32'h3aedcb33),
	.w3(32'hbb03f24b),
	.w4(32'h3acd750f),
	.w5(32'h3b926e5a),
	.w6(32'hbb28e9d6),
	.w7(32'hba8c592f),
	.w8(32'hb7b5c90d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83feb1),
	.w1(32'h3a928d29),
	.w2(32'h3b21460b),
	.w3(32'hbaf442b2),
	.w4(32'h389638e7),
	.w5(32'h3aa834a8),
	.w6(32'hba29156f),
	.w7(32'h3a8e3540),
	.w8(32'h3a0d1384),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33610e),
	.w1(32'hb92b1859),
	.w2(32'hb9cb82c7),
	.w3(32'hb9a5fe49),
	.w4(32'hb998658c),
	.w5(32'hb90f8a61),
	.w6(32'hb97ad202),
	.w7(32'hb8fb427c),
	.w8(32'h397e9dca),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374563e7),
	.w1(32'h39acd280),
	.w2(32'h395d390d),
	.w3(32'h3839fa7b),
	.w4(32'h37fdbf1f),
	.w5(32'hb8c5d075),
	.w6(32'h396bca39),
	.w7(32'hba30bf8b),
	.w8(32'hb9b47f69),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38343c05),
	.w1(32'h38b4d8d7),
	.w2(32'hb89921b7),
	.w3(32'h398724cf),
	.w4(32'hb7ac0777),
	.w5(32'h3802e4c3),
	.w6(32'h39448578),
	.w7(32'h36e0c3fd),
	.w8(32'h393d169e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945e948),
	.w1(32'hba080731),
	.w2(32'hba6ee22b),
	.w3(32'h39d5f5eb),
	.w4(32'h38e5eb9b),
	.w5(32'h39883e68),
	.w6(32'h3936f7a5),
	.w7(32'hba108d34),
	.w8(32'hba138ce8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6aca0a),
	.w1(32'h3a9a927c),
	.w2(32'h3b4a7736),
	.w3(32'hbad616db),
	.w4(32'hb7cc76c6),
	.w5(32'h3a884b8b),
	.w6(32'hba1f9fb6),
	.w7(32'h3aa00543),
	.w8(32'h3afdce2d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fdb1f),
	.w1(32'h39309622),
	.w2(32'h39e96da8),
	.w3(32'hba642204),
	.w4(32'hb92b2714),
	.w5(32'h39901ebb),
	.w6(32'h388483d5),
	.w7(32'h39c38039),
	.w8(32'h395fd80d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dd94e),
	.w1(32'hbb24db9a),
	.w2(32'h3a238fdc),
	.w3(32'hbb072486),
	.w4(32'hbad1c777),
	.w5(32'h3adfd287),
	.w6(32'hbafbe311),
	.w7(32'hbadff505),
	.w8(32'h3a00ba1e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb871b29b),
	.w1(32'hb894844d),
	.w2(32'hba63cdad),
	.w3(32'hbac64962),
	.w4(32'hbb0693a7),
	.w5(32'hbac3b61d),
	.w6(32'hba445ea3),
	.w7(32'hba28c878),
	.w8(32'hbb00859a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb785721a),
	.w1(32'h390163d1),
	.w2(32'hba51e143),
	.w3(32'h38b9c2f2),
	.w4(32'h3a8dcf2a),
	.w5(32'h38c2778c),
	.w6(32'h399752fa),
	.w7(32'hb98e4956),
	.w8(32'h3930f116),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43b3a2),
	.w1(32'h39bc1227),
	.w2(32'h39ca9444),
	.w3(32'hba02e0f1),
	.w4(32'h3a304ac9),
	.w5(32'h3a43fa2b),
	.w6(32'h3a7d4417),
	.w7(32'h3a80ac9a),
	.w8(32'h3a174432),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdfe24),
	.w1(32'h3909313c),
	.w2(32'h39187801),
	.w3(32'h3a2447db),
	.w4(32'hb909c1cf),
	.w5(32'hb8847815),
	.w6(32'h3965cc59),
	.w7(32'h38507272),
	.w8(32'h376d5f9c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888d4f3),
	.w1(32'hb8effec1),
	.w2(32'hb8af0c92),
	.w3(32'hb91aba53),
	.w4(32'hb93a28ce),
	.w5(32'hb862ecdc),
	.w6(32'hb727d55a),
	.w7(32'hb893c17a),
	.w8(32'hb9059bed),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30b35a),
	.w1(32'hbb186a15),
	.w2(32'h3b223cda),
	.w3(32'hba97df77),
	.w4(32'hbb581b01),
	.w5(32'h3b1f08ea),
	.w6(32'hbac9f7ff),
	.w7(32'h39a57323),
	.w8(32'h3bbabc8a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89ba70),
	.w1(32'hba6e8a42),
	.w2(32'h3b8381ec),
	.w3(32'hbb67880a),
	.w4(32'h3a8be516),
	.w5(32'h3b8aab8f),
	.w6(32'hbae77f60),
	.w7(32'h3a5a5806),
	.w8(32'h3b2872f6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d73906),
	.w1(32'hb90e829e),
	.w2(32'hb9a1d992),
	.w3(32'hb9a54130),
	.w4(32'h39dd27e4),
	.w5(32'h3a1bb03b),
	.w6(32'hb9f0cc58),
	.w7(32'hb8e89960),
	.w8(32'h378ce984),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b46dd),
	.w1(32'h3a17ec7e),
	.w2(32'h3aadd3d1),
	.w3(32'hba82622c),
	.w4(32'hb9db090e),
	.w5(32'hb9f36e32),
	.w6(32'hb8fd655f),
	.w7(32'h3a9ed3b2),
	.w8(32'h39fc73eb),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bae10f),
	.w1(32'hb7bd984e),
	.w2(32'h383d0489),
	.w3(32'hb95a4074),
	.w4(32'hb9877e02),
	.w5(32'h37f64cae),
	.w6(32'h39583115),
	.w7(32'hb83bf1e7),
	.w8(32'hb97ab963),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacef136),
	.w1(32'h3a19d048),
	.w2(32'h3b1794cd),
	.w3(32'hbac5ebfd),
	.w4(32'h39fbbdfd),
	.w5(32'h3ae12c46),
	.w6(32'hba2e2abe),
	.w7(32'h3a06fb28),
	.w8(32'h3aa46c91),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a89f3),
	.w1(32'h3b45983f),
	.w2(32'h3ab94ad6),
	.w3(32'h39eb8870),
	.w4(32'h3b260fd3),
	.w5(32'h3b530fb7),
	.w6(32'h38f80117),
	.w7(32'h3a8744bc),
	.w8(32'h395e3b59),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc013ade),
	.w1(32'hbba12e4f),
	.w2(32'h3a8cdf84),
	.w3(32'hbbc3ad9a),
	.w4(32'hba2ac3ec),
	.w5(32'h3b703005),
	.w6(32'hbb822698),
	.w7(32'hbb064a06),
	.w8(32'h3b054c1e),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8afc91a),
	.w1(32'h3a8350a7),
	.w2(32'h3a84d070),
	.w3(32'hbaa34823),
	.w4(32'h38fa68fe),
	.w5(32'hba0082ec),
	.w6(32'hb981144c),
	.w7(32'hba1fd8b4),
	.w8(32'hba40e479),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39776b),
	.w1(32'hba5be33c),
	.w2(32'h3a320f32),
	.w3(32'hbb4ba0e4),
	.w4(32'hba053547),
	.w5(32'h3b2ec827),
	.w6(32'hbb385bd9),
	.w7(32'hba96f62d),
	.w8(32'h3a1619e7),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88b300),
	.w1(32'hbb4c9c8f),
	.w2(32'h3abc2470),
	.w3(32'hbb58a656),
	.w4(32'hba943edb),
	.w5(32'h3ba4abc0),
	.w6(32'hbb2ec5e5),
	.w7(32'hb89b815c),
	.w8(32'h3b82731c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a913697),
	.w1(32'h3b30e77f),
	.w2(32'h3ab42f50),
	.w3(32'hb9e9c6e5),
	.w4(32'h38b7f7ef),
	.w5(32'hb99906bf),
	.w6(32'hba8ed2fe),
	.w7(32'h39f17d0b),
	.w8(32'h3a574be3),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4124e8),
	.w1(32'hba57781d),
	.w2(32'h3aebf1c2),
	.w3(32'hbac48a80),
	.w4(32'h3a6f216d),
	.w5(32'h3b5ca376),
	.w6(32'hbad8491d),
	.w7(32'hb96e5fb0),
	.w8(32'h3aa3ff7c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc9e02),
	.w1(32'h39fed5de),
	.w2(32'h3a852b5d),
	.w3(32'hb9716277),
	.w4(32'h39a81d8c),
	.w5(32'h3a5aca51),
	.w6(32'hb90c0298),
	.w7(32'h393e9458),
	.w8(32'h39df9386),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9470291),
	.w1(32'hbaa62f53),
	.w2(32'h3b423b82),
	.w3(32'hbb7debf0),
	.w4(32'hbb793bdd),
	.w5(32'hbaff8982),
	.w6(32'hbb2dd21d),
	.w7(32'hbaa0bb3e),
	.w8(32'hb95e262d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd142e),
	.w1(32'h3a0bf339),
	.w2(32'h3aaef08c),
	.w3(32'hb9e3dcdd),
	.w4(32'h39897173),
	.w5(32'h3985ab37),
	.w6(32'hb846452b),
	.w7(32'h394d8c4f),
	.w8(32'hb9bc50a4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bfa14b),
	.w1(32'h3885fd49),
	.w2(32'h392bd36c),
	.w3(32'hb8572ca5),
	.w4(32'h3803633d),
	.w5(32'h38e745a6),
	.w6(32'hb8d4e3c7),
	.w7(32'hb88a5b2d),
	.w8(32'h3786ad20),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d65a53),
	.w1(32'hb873aa1d),
	.w2(32'h37dceb5d),
	.w3(32'h389a8f2f),
	.w4(32'hb7bc45e8),
	.w5(32'h38365b4e),
	.w6(32'h38d50aec),
	.w7(32'hb8f8870c),
	.w8(32'hb894a1be),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87cab5),
	.w1(32'hba650698),
	.w2(32'hb83062db),
	.w3(32'hb9b45671),
	.w4(32'h3964cddc),
	.w5(32'h3a25a656),
	.w6(32'hba64e933),
	.w7(32'h3802d755),
	.w8(32'h378cc4c4),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba948828),
	.w1(32'hb9484fe7),
	.w2(32'hb8df48fb),
	.w3(32'hbb2823ee),
	.w4(32'hba8da3fe),
	.w5(32'hbad2e900),
	.w6(32'hb9e7ad9b),
	.w7(32'hba2572ec),
	.w8(32'hbb1bfc57),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6de360),
	.w1(32'hba30ee48),
	.w2(32'h3b2cdc5b),
	.w3(32'hbb2fba3d),
	.w4(32'hb9bec045),
	.w5(32'h3b03ec5a),
	.w6(32'hbab5cecb),
	.w7(32'h3902b13e),
	.w8(32'h3ab59276),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cb8f5d),
	.w1(32'hb7a67eea),
	.w2(32'h36b31a32),
	.w3(32'hb7956a2c),
	.w4(32'hb7486dc2),
	.w5(32'h37d65f68),
	.w6(32'hb81ae4b7),
	.w7(32'hb8015943),
	.w8(32'h374a7b5e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73633f),
	.w1(32'hb845c9d2),
	.w2(32'h3b767083),
	.w3(32'hbb3bd7d4),
	.w4(32'h3a511e3c),
	.w5(32'h3b78476a),
	.w6(32'hbb00f17a),
	.w7(32'hb9bbbb1f),
	.w8(32'h3aa1833e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9e0c6),
	.w1(32'h3a66588a),
	.w2(32'h3ad19dea),
	.w3(32'hb9e6f0e4),
	.w4(32'hb950b274),
	.w5(32'h3931a95c),
	.w6(32'h39ac3c7a),
	.w7(32'hb8155a2f),
	.w8(32'hb9b2de41),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7e919),
	.w1(32'hbbbc83fa),
	.w2(32'hba4cb32a),
	.w3(32'hbb7a9434),
	.w4(32'hbae9c280),
	.w5(32'h3b77c4df),
	.w6(32'hbba10033),
	.w7(32'hbb93f337),
	.w8(32'h3a31846c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc69944),
	.w1(32'hb9a83c63),
	.w2(32'h3aba3dc8),
	.w3(32'hbbc9eb1b),
	.w4(32'hbac54343),
	.w5(32'h3b56ab62),
	.w6(32'hbb96aad7),
	.w7(32'hba853e6f),
	.w8(32'h3ab0ed14),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc13e5),
	.w1(32'h39ceaa08),
	.w2(32'hbabf4f96),
	.w3(32'h3aa0a7f6),
	.w4(32'h3974b5a1),
	.w5(32'hbb0405cc),
	.w6(32'h3a70792f),
	.w7(32'h3966acd1),
	.w8(32'hbaba28c9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a664764),
	.w1(32'h3a776ee5),
	.w2(32'h389e0ff8),
	.w3(32'h3b1693b7),
	.w4(32'h3b1de771),
	.w5(32'h3ac0cef8),
	.w6(32'h3ae93a17),
	.w7(32'h3ace35ce),
	.w8(32'h3a87c4a9),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab15c51),
	.w1(32'h3a7231a1),
	.w2(32'h3b0128c9),
	.w3(32'hbb0c72ed),
	.w4(32'hb9406013),
	.w5(32'h3a5cb1da),
	.w6(32'hbabd3f6a),
	.w7(32'h3a454704),
	.w8(32'h3a8ba94f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab04e00),
	.w1(32'h3a8dd2ed),
	.w2(32'hb9be1f4b),
	.w3(32'h39d43d2b),
	.w4(32'h3a5ea6e1),
	.w5(32'hba418972),
	.w6(32'h3a6d269d),
	.w7(32'h3a5ce450),
	.w8(32'hbab1eab5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9a505),
	.w1(32'h3a34746c),
	.w2(32'hb994679c),
	.w3(32'h39dc512f),
	.w4(32'h39a25ef6),
	.w5(32'hba8904f1),
	.w6(32'h39ee36ed),
	.w7(32'h38e1384a),
	.w8(32'hba59066f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48ce39),
	.w1(32'hb9fcda84),
	.w2(32'h39c3837c),
	.w3(32'hb961a86f),
	.w4(32'h3a2015fc),
	.w5(32'h3aa58456),
	.w6(32'hba20d7c2),
	.w7(32'hb80bbf9f),
	.w8(32'h3a6c8af8),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f80776),
	.w1(32'hb980bd59),
	.w2(32'hb9340193),
	.w3(32'h395c41f9),
	.w4(32'h3959102b),
	.w5(32'h3967642e),
	.w6(32'h392a0576),
	.w7(32'h3921fcd3),
	.w8(32'h399040ac),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68ee3a),
	.w1(32'hbb0966aa),
	.w2(32'h3aa22d16),
	.w3(32'hbb2afbfa),
	.w4(32'hb909bcda),
	.w5(32'h3b628611),
	.w6(32'hbacaea89),
	.w7(32'h38381480),
	.w8(32'h3b06d3e2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d9d0b),
	.w1(32'hb9abe5fa),
	.w2(32'h39902e38),
	.w3(32'hb903d5f1),
	.w4(32'h3a3f3d2e),
	.w5(32'h3a892bfc),
	.w6(32'hb9892a7c),
	.w7(32'hb91ed910),
	.w8(32'h39e85f95),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f7ee7),
	.w1(32'h3b3f31a7),
	.w2(32'h3b6abaaf),
	.w3(32'hbad913b4),
	.w4(32'hba6d1e41),
	.w5(32'h3a16f5cf),
	.w6(32'hb9cb0a88),
	.w7(32'h3ac1b4da),
	.w8(32'h3ae14673),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80cd7f6),
	.w1(32'hb8ed50ea),
	.w2(32'hb982aa26),
	.w3(32'hb98d485e),
	.w4(32'hb5a2c206),
	.w5(32'hb90b59a7),
	.w6(32'hb931665d),
	.w7(32'h39ac78f0),
	.w8(32'h3950fe2e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb114efa),
	.w1(32'hbad2eca2),
	.w2(32'h39116e64),
	.w3(32'hba8cbcb1),
	.w4(32'hbb14bd70),
	.w5(32'hba428dfe),
	.w6(32'hba8c7413),
	.w7(32'hbb01cf9d),
	.w8(32'h394386d4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eb5cfa),
	.w1(32'h3906e6c5),
	.w2(32'h39408975),
	.w3(32'h3903adb4),
	.w4(32'h398512fc),
	.w5(32'h3999f30d),
	.w6(32'h394e70d9),
	.w7(32'h39a4d866),
	.w8(32'h3998023d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394dc4c1),
	.w1(32'hb928a6bf),
	.w2(32'hb9c81604),
	.w3(32'h3993d47e),
	.w4(32'h3658ad7a),
	.w5(32'hb955f5d4),
	.w6(32'h39489589),
	.w7(32'h383d29c9),
	.w8(32'hb82e963d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab80c98),
	.w1(32'h3a325175),
	.w2(32'h3961a68c),
	.w3(32'hbad4207a),
	.w4(32'h39398f2b),
	.w5(32'hb9a4da36),
	.w6(32'hba3d8f5c),
	.w7(32'h38c93f6d),
	.w8(32'hbab6baa2),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96ca10),
	.w1(32'hba4ea392),
	.w2(32'h3b7dd6cf),
	.w3(32'hbbcb6b3d),
	.w4(32'hbb6fc293),
	.w5(32'h3a28cf06),
	.w6(32'hbb8b2852),
	.w7(32'h3a23da4c),
	.w8(32'h3b6a1f73),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6005fe),
	.w1(32'h39eb902a),
	.w2(32'hb849142a),
	.w3(32'h3a27683f),
	.w4(32'h39d47d54),
	.w5(32'h3892e165),
	.w6(32'h3a32fd96),
	.w7(32'h3a298417),
	.w8(32'h3a4667c6),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4711dc),
	.w1(32'h3b2b11e8),
	.w2(32'h3b4a8c34),
	.w3(32'hba512f5c),
	.w4(32'h3aa3acb0),
	.w5(32'h3abc6e58),
	.w6(32'hb845cad5),
	.w7(32'h3afe9e95),
	.w8(32'h3aa8d553),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba556759),
	.w1(32'h3ae87a88),
	.w2(32'h3aee3650),
	.w3(32'hba4b367c),
	.w4(32'h3ad2db2d),
	.w5(32'h3b00ac96),
	.w6(32'hb99e5e66),
	.w7(32'h3a859fb0),
	.w8(32'h39b2dfb2),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee39dc),
	.w1(32'h3ab5f2ac),
	.w2(32'h3b6b8e5a),
	.w3(32'hbbb00f0f),
	.w4(32'h3b058881),
	.w5(32'h3b8e2119),
	.w6(32'hbb971c18),
	.w7(32'h39d808c4),
	.w8(32'h3a8ea3a2),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8ca15),
	.w1(32'hba125dfb),
	.w2(32'h3927a60c),
	.w3(32'hbac7a0ba),
	.w4(32'hb883608e),
	.w5(32'h3af19ea0),
	.w6(32'hba82686c),
	.w7(32'hba206cce),
	.w8(32'hb925a676),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f1a07),
	.w1(32'h3a0f32f4),
	.w2(32'h3b9021e9),
	.w3(32'hbb2d8239),
	.w4(32'h3b13e784),
	.w5(32'h3b92a194),
	.w6(32'hbac0608c),
	.w7(32'h3a9d3e17),
	.w8(32'h3b092e50),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a030cc2),
	.w1(32'h3a2b89e9),
	.w2(32'h3a2379e4),
	.w3(32'h3a112e2c),
	.w4(32'h3a7ff0a0),
	.w5(32'h3a306c08),
	.w6(32'h3a080f6e),
	.w7(32'h3a9a7e4e),
	.w8(32'h3a8105b2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb410258),
	.w1(32'hba3fe402),
	.w2(32'h3a9edfa8),
	.w3(32'hbb0af38b),
	.w4(32'h3a2cb6c9),
	.w5(32'h3b319518),
	.w6(32'hbb03cf3c),
	.w7(32'hb9ab9e22),
	.w8(32'hb8bcc0e0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e969df),
	.w1(32'h378f20ef),
	.w2(32'h376b69db),
	.w3(32'h380e7a77),
	.w4(32'h37197c42),
	.w5(32'h377f9099),
	.w6(32'h37cd87ae),
	.w7(32'h3635229d),
	.w8(32'h3725888e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c778f),
	.w1(32'hb92f497f),
	.w2(32'h3a79cb4b),
	.w3(32'hba517264),
	.w4(32'h3904cced),
	.w5(32'h3a3604db),
	.w6(32'hba89bcec),
	.w7(32'h3845cfe8),
	.w8(32'h3a0ac691),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38db53eb),
	.w1(32'h398abeac),
	.w2(32'h38cd6752),
	.w3(32'hb945f8ad),
	.w4(32'h398e99bf),
	.w5(32'h374a6f50),
	.w6(32'hb8bc2fda),
	.w7(32'h391522f3),
	.w8(32'hb93e48d8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23a9f1),
	.w1(32'h393d128d),
	.w2(32'h3ad0a7b0),
	.w3(32'hbb3ff6e5),
	.w4(32'h3a05c122),
	.w5(32'h3b191786),
	.w6(32'hbb1b7631),
	.w7(32'h39331f26),
	.w8(32'h38d21a39),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36916bc5),
	.w1(32'h361a8ed3),
	.w2(32'h36c11e03),
	.w3(32'h3538df10),
	.w4(32'h36a81d2a),
	.w5(32'h375b771b),
	.w6(32'h36b4a48f),
	.w7(32'h3782e635),
	.w8(32'h37665248),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86f357c),
	.w1(32'h378375ca),
	.w2(32'hb87693f4),
	.w3(32'h38884dc3),
	.w4(32'h38c862f9),
	.w5(32'hb81ca68a),
	.w6(32'h388c14ef),
	.w7(32'h383a4393),
	.w8(32'hb884665f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c604fd),
	.w1(32'h3aad2d27),
	.w2(32'h3a87562a),
	.w3(32'hba933856),
	.w4(32'hba9052a6),
	.w5(32'hb83b1aff),
	.w6(32'hb9d8ff4a),
	.w7(32'h3a67b3f9),
	.w8(32'h3a57547f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb143d6b),
	.w1(32'hba841143),
	.w2(32'h37dd3f20),
	.w3(32'hba32f2d3),
	.w4(32'h3888c03d),
	.w5(32'hb9f041b7),
	.w6(32'hbaec1271),
	.w7(32'hba573ac8),
	.w8(32'hb9281ae5),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb365265),
	.w1(32'hbb459df2),
	.w2(32'hbb4e067f),
	.w3(32'hbb8267a0),
	.w4(32'hbac331e6),
	.w5(32'hbaf16879),
	.w6(32'hbacb9865),
	.w7(32'hb96f71db),
	.w8(32'hbb127110),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc7e9c),
	.w1(32'h398093a9),
	.w2(32'hb92701b8),
	.w3(32'h39863545),
	.w4(32'h39276b7b),
	.w5(32'hb8e98b43),
	.w6(32'h399f6e90),
	.w7(32'h38b401f0),
	.w8(32'h385cdaec),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ac677),
	.w1(32'hbb4d117f),
	.w2(32'h3bce97c2),
	.w3(32'hbbf8cb83),
	.w4(32'hba600351),
	.w5(32'h3b9108ec),
	.w6(32'hbbac74a3),
	.w7(32'h3a13d6b9),
	.w8(32'h3b9f6e6d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba931a2),
	.w1(32'h3b98d829),
	.w2(32'h38ae2729),
	.w3(32'hbb49198d),
	.w4(32'h3bcb9a5e),
	.w5(32'h3ba28eac),
	.w6(32'hbb676a66),
	.w7(32'h3adf891f),
	.w8(32'hba7ed6f1),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dbb0e),
	.w1(32'hbae491a5),
	.w2(32'hba714aa0),
	.w3(32'hba2f9332),
	.w4(32'hb9bcf21f),
	.w5(32'h3a40211e),
	.w6(32'hba95b1e4),
	.w7(32'hba999d67),
	.w8(32'hbac7d347),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85ff860),
	.w1(32'hb7abb4fa),
	.w2(32'h374e297e),
	.w3(32'hb7ab96ab),
	.w4(32'h37f2d27d),
	.w5(32'h382a643b),
	.w6(32'hb668a207),
	.w7(32'hb768b9bb),
	.w8(32'h36bd77ca),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d59b2),
	.w1(32'hb7ed2e5c),
	.w2(32'hb9987039),
	.w3(32'h38b92c33),
	.w4(32'h38733279),
	.w5(32'hb9197ca6),
	.w6(32'h38474296),
	.w7(32'hb93f5742),
	.w8(32'hb99ca82a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383af34f),
	.w1(32'h3739e2f9),
	.w2(32'hb616e7eb),
	.w3(32'h380fda9e),
	.w4(32'h337be86c),
	.w5(32'hb770c804),
	.w6(32'h37419042),
	.w7(32'hb73cfb35),
	.w8(32'hb6a70a2d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc2bb8),
	.w1(32'hbb104f6f),
	.w2(32'hba0d4487),
	.w3(32'hba872748),
	.w4(32'hbb06b4bf),
	.w5(32'hba8618a1),
	.w6(32'hba57ffa6),
	.w7(32'hbb2aabbb),
	.w8(32'hba8c9e6f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7adaa7),
	.w1(32'hba0a07e8),
	.w2(32'h3a0e9fb3),
	.w3(32'hba9abdaf),
	.w4(32'hb9f20314),
	.w5(32'h395df50a),
	.w6(32'h39bcf272),
	.w7(32'h3a8c9a33),
	.w8(32'h3a8ebcde),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b83de),
	.w1(32'h3a798f58),
	.w2(32'h3a7f1f64),
	.w3(32'hbad82f1a),
	.w4(32'h38be1935),
	.w5(32'hb85c87d4),
	.w6(32'h34dace68),
	.w7(32'h3908968a),
	.w8(32'hba44b83b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e56e97),
	.w1(32'h3a241d38),
	.w2(32'h3aa0857a),
	.w3(32'hb95a8887),
	.w4(32'hb8ca87a1),
	.w5(32'h398710d4),
	.w6(32'h38953b59),
	.w7(32'h39ffd5b5),
	.w8(32'h3a618fa7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a143e),
	.w1(32'hbb095043),
	.w2(32'h3ab86031),
	.w3(32'hbb7db306),
	.w4(32'hba9aa99f),
	.w5(32'h3ab3a3e9),
	.w6(32'hbb3afea7),
	.w7(32'hba1ed813),
	.w8(32'h3a606cc4),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bc87c),
	.w1(32'hbaa11934),
	.w2(32'hb9f87400),
	.w3(32'hba04fd96),
	.w4(32'hba4cb1a5),
	.w5(32'hb99feaa7),
	.w6(32'h393f85dc),
	.w7(32'h3a1ca8c6),
	.w8(32'h3ab8480b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373118b5),
	.w1(32'hb663c277),
	.w2(32'h363b22a8),
	.w3(32'h3703e443),
	.w4(32'h3658cdb5),
	.w5(32'h3719b752),
	.w6(32'h3759ace9),
	.w7(32'h3792ff8e),
	.w8(32'h37436fed),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9183cb3),
	.w1(32'h3ad86467),
	.w2(32'hbb3c051b),
	.w3(32'hbaa5a97f),
	.w4(32'h3a67f752),
	.w5(32'h3a28329e),
	.w6(32'hb990ca3c),
	.w7(32'hba1faba0),
	.w8(32'h3a0a7d93),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384b3f0b),
	.w1(32'h36cb68f0),
	.w2(32'hb710179a),
	.w3(32'h384fcc6b),
	.w4(32'h36b6cb9f),
	.w5(32'h3611cdf6),
	.w6(32'h38425cb1),
	.w7(32'h3780c14e),
	.w8(32'hb77e430a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb478154),
	.w1(32'hbae0cbb7),
	.w2(32'h3a872f1f),
	.w3(32'hbb27f4fb),
	.w4(32'hbb18ebe9),
	.w5(32'h39f0ad0d),
	.w6(32'hbadf6a4d),
	.w7(32'hba83c52a),
	.w8(32'h39255efa),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef6e98),
	.w1(32'h3aa7e02b),
	.w2(32'hbaa1dd58),
	.w3(32'h3918fc1a),
	.w4(32'h391bc9d8),
	.w5(32'hbacd0ae3),
	.w6(32'h3a104a1c),
	.w7(32'h39d22e73),
	.w8(32'hbaa5a7df),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f98258),
	.w1(32'h3ab5e8c1),
	.w2(32'h3acc78fc),
	.w3(32'hba0caf20),
	.w4(32'h3954c7df),
	.w5(32'h3a04debc),
	.w6(32'h37b90a99),
	.w7(32'h3a222d48),
	.w8(32'h3898e9e9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3909af04),
	.w1(32'h3940b555),
	.w2(32'h38dddb85),
	.w3(32'h38359feb),
	.w4(32'h38deec0e),
	.w5(32'h38c49bb2),
	.w6(32'hb7918098),
	.w7(32'h38132e6b),
	.w8(32'h38a346f0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02e5d2),
	.w1(32'h3b1285bc),
	.w2(32'h3b1a35b9),
	.w3(32'hbab3229c),
	.w4(32'h3a81fa3a),
	.w5(32'h3a00a5f8),
	.w6(32'h3a17bb30),
	.w7(32'h3ab6ef69),
	.w8(32'h392bb8cc),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb120ca4),
	.w1(32'hb66af2b2),
	.w2(32'h3b2fc329),
	.w3(32'hbaddf09c),
	.w4(32'h39fc49c1),
	.w5(32'h3b35bb98),
	.w6(32'hbaa6bd04),
	.w7(32'h3a055044),
	.w8(32'h3adf72fe),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fe8c8),
	.w1(32'hbae5ed9f),
	.w2(32'h3ae0c17a),
	.w3(32'hbb802c26),
	.w4(32'hbaaa3b0a),
	.w5(32'h3ab72782),
	.w6(32'hbb43c6b1),
	.w7(32'hba0f67d3),
	.w8(32'h3aa3d856),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387f00b3),
	.w1(32'h372dffda),
	.w2(32'hb783e5c3),
	.w3(32'h38299a95),
	.w4(32'h379b0b33),
	.w5(32'h3715fd02),
	.w6(32'h37fa1522),
	.w7(32'hb718b52b),
	.w8(32'hb7c87b8f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b956bb),
	.w1(32'h3882ae38),
	.w2(32'h38862332),
	.w3(32'h380a79a9),
	.w4(32'hb7d437c5),
	.w5(32'h3817d5d0),
	.w6(32'h3913e0dd),
	.w7(32'h389c5fa5),
	.w8(32'h38d51d84),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2c238),
	.w1(32'h38dbfcd2),
	.w2(32'h3af88e9d),
	.w3(32'hbb15cdf9),
	.w4(32'hbb0e7880),
	.w5(32'hba74d324),
	.w6(32'hbb18a8f6),
	.w7(32'h3b16f1c1),
	.w8(32'h3b9230e8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f6d0d),
	.w1(32'h39d18361),
	.w2(32'h3b76ffc5),
	.w3(32'hbb99472d),
	.w4(32'hbb3bc7ed),
	.w5(32'h36adefd5),
	.w6(32'hbb1fbc83),
	.w7(32'h3a87a92d),
	.w8(32'h3b75c71e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a499c8),
	.w1(32'h3b1a1e7a),
	.w2(32'h3b64b160),
	.w3(32'hbaf72282),
	.w4(32'hb9b01dd2),
	.w5(32'h3a6a70d0),
	.w6(32'hba3413cc),
	.w7(32'h3ac34b6b),
	.w8(32'h3ae07fab),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba59b02),
	.w1(32'hbb564858),
	.w2(32'h3af91dd2),
	.w3(32'hba618cd0),
	.w4(32'h3afbf819),
	.w5(32'h3bca4c55),
	.w6(32'hbb044852),
	.w7(32'hbb1fb5d1),
	.w8(32'hba548e59),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c28c8),
	.w1(32'hb999bd30),
	.w2(32'h3996408e),
	.w3(32'hb93c26af),
	.w4(32'hb90f72bc),
	.w5(32'h381a722c),
	.w6(32'hb9978f24),
	.w7(32'hb9418e48),
	.w8(32'hb963b0f8),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3868fbf5),
	.w1(32'hb98d3706),
	.w2(32'h398d0df2),
	.w3(32'hb9cfc970),
	.w4(32'hb99825a0),
	.w5(32'h386d8f32),
	.w6(32'h39ae02dd),
	.w7(32'h37f352b8),
	.w8(32'h3895ca73),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac6f83),
	.w1(32'hbadc4831),
	.w2(32'hbb0c8ef0),
	.w3(32'hbb741d5c),
	.w4(32'hbb258b49),
	.w5(32'hbb61d1ab),
	.w6(32'hbb768f10),
	.w7(32'hbb3b4f83),
	.w8(32'h3a6fa5bf),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd15ffb),
	.w1(32'hbb403b26),
	.w2(32'h3b84cf33),
	.w3(32'hbb990dcc),
	.w4(32'hbab1802f),
	.w5(32'h3b860ee1),
	.w6(32'hbb69eb7f),
	.w7(32'hb944fdac),
	.w8(32'h3b894654),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba523e9),
	.w1(32'hbb962996),
	.w2(32'hba6baa8b),
	.w3(32'hbb7ca4c4),
	.w4(32'hbaed905a),
	.w5(32'h3ae883c5),
	.w6(32'hbb54df73),
	.w7(32'hba7931da),
	.w8(32'h3a3c122b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff2598),
	.w1(32'h3abf0d69),
	.w2(32'h389df969),
	.w3(32'h39cee416),
	.w4(32'hb98131ef),
	.w5(32'hbac06120),
	.w6(32'h39c5d378),
	.w7(32'hb9fdbb6a),
	.w8(32'hba893a2a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7eff7d),
	.w1(32'h3ad02c3e),
	.w2(32'h3a67c026),
	.w3(32'hba01b1c2),
	.w4(32'h3a0ad7da),
	.w5(32'hb7cb8548),
	.w6(32'hb8280af4),
	.w7(32'hb9e7f2b4),
	.w8(32'hbacf16e4),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bc641b),
	.w1(32'h37899e93),
	.w2(32'h3777d3b6),
	.w3(32'h3789fd76),
	.w4(32'h37436216),
	.w5(32'h37188fc5),
	.w6(32'h378ea02e),
	.w7(32'h3793cadd),
	.w8(32'h37934776),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369474e1),
	.w1(32'hb71c6e26),
	.w2(32'hb6ed4cbd),
	.w3(32'h365edb95),
	.w4(32'hb6fa5769),
	.w5(32'hb696f88c),
	.w6(32'hb62f2c0c),
	.w7(32'h362beb06),
	.w8(32'h35bdd9ae),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a16ff),
	.w1(32'h39b82a8c),
	.w2(32'h3a5d5bea),
	.w3(32'hb90ec3c3),
	.w4(32'hb999f4d7),
	.w5(32'h39e4b6ea),
	.w6(32'h396a10e0),
	.w7(32'h3a96fb1c),
	.w8(32'h3a67a224),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36101845),
	.w1(32'hb697bc3c),
	.w2(32'h35b0b81f),
	.w3(32'hb6275ad8),
	.w4(32'h35bff682),
	.w5(32'h374aa72c),
	.w6(32'h3788ac24),
	.w7(32'h3759cf59),
	.w8(32'h37b96c28),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba836612),
	.w1(32'hbaeaa367),
	.w2(32'hbaad7dc1),
	.w3(32'hba689704),
	.w4(32'hbaf21fdc),
	.w5(32'hbac969e4),
	.w6(32'hba932ed4),
	.w7(32'hba2753d1),
	.w8(32'hba25ae0c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a5ffd),
	.w1(32'hbab2b923),
	.w2(32'h3b0ee5a2),
	.w3(32'hbb1e1dc5),
	.w4(32'hbb41b688),
	.w5(32'h3a4c2c5e),
	.w6(32'hbb3c710d),
	.w7(32'hba1fd05f),
	.w8(32'h3b298892),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdb979),
	.w1(32'h3a14283f),
	.w2(32'h3aa8e6a4),
	.w3(32'hbada352f),
	.w4(32'hb999d1eb),
	.w5(32'h3a341c8b),
	.w6(32'hba07854a),
	.w7(32'h3a2ea288),
	.w8(32'h3a728d95),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83d1a35),
	.w1(32'hb79ad248),
	.w2(32'h37102c69),
	.w3(32'hb7abe50d),
	.w4(32'h37938e29),
	.w5(32'h381b72aa),
	.w6(32'hb839881a),
	.w7(32'h36d14d66),
	.w8(32'h374305bd),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e7863),
	.w1(32'hbc031f8f),
	.w2(32'hbb0e83ca),
	.w3(32'hbbe0ed13),
	.w4(32'hbb7c286f),
	.w5(32'h3b773399),
	.w6(32'hbbc2b8ef),
	.w7(32'hbab69c6e),
	.w8(32'h3b98e034),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13b81c),
	.w1(32'hba8f883b),
	.w2(32'h3a86a9ae),
	.w3(32'hbae19c6a),
	.w4(32'hba037437),
	.w5(32'h3aa8f009),
	.w6(32'hbaa91f58),
	.w7(32'hb9bf3e19),
	.w8(32'h39f29089),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ad7505),
	.w1(32'hb8a6148f),
	.w2(32'hb8f208fe),
	.w3(32'hb80a4007),
	.w4(32'hb87a5a02),
	.w5(32'hb876af43),
	.w6(32'hb86e6f1f),
	.w7(32'hb8313a7c),
	.w8(32'hb81f3769),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb558266),
	.w1(32'hbb2f1c30),
	.w2(32'h3a7ed822),
	.w3(32'hbb151417),
	.w4(32'hba4bb55e),
	.w5(32'h3b127554),
	.w6(32'hbb11d624),
	.w7(32'hba86442f),
	.w8(32'h3aa2e92c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39614e0f),
	.w1(32'h395d4c68),
	.w2(32'h38fbc24c),
	.w3(32'h398ce4c8),
	.w4(32'h3984d317),
	.w5(32'h39170149),
	.w6(32'h39398d6d),
	.w7(32'h392d8a63),
	.w8(32'h38240fc4),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a1c94),
	.w1(32'hb8226f89),
	.w2(32'h3816f294),
	.w3(32'hb8f05c26),
	.w4(32'h38ee69c8),
	.w5(32'h396682ac),
	.w6(32'hb8f33f11),
	.w7(32'h3880a25a),
	.w8(32'h396b499d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75dfe7c),
	.w1(32'hb7495a45),
	.w2(32'h3806bf20),
	.w3(32'hb6a09e58),
	.w4(32'hb6c696dd),
	.w5(32'h37c1eff1),
	.w6(32'hb5cb653a),
	.w7(32'h3775f6a7),
	.w8(32'h37db37d0),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388aaeba),
	.w1(32'h37a28367),
	.w2(32'hb74fe54a),
	.w3(32'h385094e1),
	.w4(32'h379341ab),
	.w5(32'hb6310b09),
	.w6(32'h380c0cfa),
	.w7(32'h37d6f773),
	.w8(32'h382c11aa),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f03c2),
	.w1(32'h38b2fa84),
	.w2(32'hb9ae272c),
	.w3(32'hb9e703c9),
	.w4(32'hba1fa835),
	.w5(32'hbaa7af47),
	.w6(32'hb806f88b),
	.w7(32'hb904cc02),
	.w8(32'hb97686dd),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba93f15),
	.w1(32'h3a493d58),
	.w2(32'h3b8a8965),
	.w3(32'hbb59f7c5),
	.w4(32'h3b4d6515),
	.w5(32'h3c04c4ba),
	.w6(32'hbba17d14),
	.w7(32'hb9f1e6ed),
	.w8(32'h3ab6f664),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb671d34),
	.w1(32'hbab5d9b2),
	.w2(32'h3b36154f),
	.w3(32'hbb377668),
	.w4(32'h39d491b3),
	.w5(32'h3b7c8521),
	.w6(32'hbaece35f),
	.w7(32'h39aa49d2),
	.w8(32'h3b287005),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3fca8),
	.w1(32'hbabc4c10),
	.w2(32'h3b125db5),
	.w3(32'hbb8c2acf),
	.w4(32'h3ad1e8e9),
	.w5(32'h3b89b8c2),
	.w6(32'hbb5830e7),
	.w7(32'hba208f67),
	.w8(32'h3abbc60a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39039bfa),
	.w1(32'h391b8099),
	.w2(32'h38ca3143),
	.w3(32'h38f51651),
	.w4(32'h390f7bef),
	.w5(32'h3894ed90),
	.w6(32'h38eb8476),
	.w7(32'h38fe981b),
	.w8(32'h385e9277),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8f162),
	.w1(32'hb97035ac),
	.w2(32'h3985a187),
	.w3(32'hb99f41c5),
	.w4(32'hb8935d9e),
	.w5(32'h38f53707),
	.w6(32'h391bf9a0),
	.w7(32'hb912c902),
	.w8(32'hb9a2e7a8),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b5007c),
	.w1(32'h350accc6),
	.w2(32'h3886177a),
	.w3(32'hb7fd6d37),
	.w4(32'hb708c091),
	.w5(32'h383bd6c1),
	.w6(32'h369ede58),
	.w7(32'h3747f20d),
	.w8(32'h3873d4a8),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34ad55a1),
	.w1(32'hb687cb69),
	.w2(32'hb56fe265),
	.w3(32'h376faea1),
	.w4(32'hb7368b9f),
	.w5(32'hb717da7e),
	.w6(32'h370fe409),
	.w7(32'hb6bd0efc),
	.w8(32'hb7333d2f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a2ae4),
	.w1(32'hba477cbb),
	.w2(32'h3ac1a25a),
	.w3(32'hbb7d334b),
	.w4(32'hb6ffb83e),
	.w5(32'h3aaee38c),
	.w6(32'hbafe30e7),
	.w7(32'h38239d9c),
	.w8(32'hb97765f4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34b164),
	.w1(32'hb9cfa8b5),
	.w2(32'hb9a4cfc1),
	.w3(32'hb9bd630a),
	.w4(32'hb9806edd),
	.w5(32'hb9be747f),
	.w6(32'hb9e43ce2),
	.w7(32'hb9f5a0ef),
	.w8(32'hba14c53f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398490da),
	.w1(32'h38e9bf94),
	.w2(32'hb9292fba),
	.w3(32'h39a011d0),
	.w4(32'h394019c9),
	.w5(32'hb6be1e87),
	.w6(32'h399082ad),
	.w7(32'h3945ae84),
	.w8(32'h39217374),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17e1de),
	.w1(32'h3a10a142),
	.w2(32'h3a17cfe9),
	.w3(32'hba3eafde),
	.w4(32'h3a6a03fb),
	.w5(32'h3a53695c),
	.w6(32'hb90751eb),
	.w7(32'h3a448983),
	.w8(32'h3a1ead47),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cdc0d7),
	.w1(32'hb84061b1),
	.w2(32'hb728065d),
	.w3(32'h38912995),
	.w4(32'h37588c87),
	.w5(32'h374fd93c),
	.w6(32'h38a6b145),
	.w7(32'hb7d70e5a),
	.w8(32'hb8057e2d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a5184),
	.w1(32'hbaba26b5),
	.w2(32'h38130898),
	.w3(32'hbad4bdbe),
	.w4(32'hba4715b0),
	.w5(32'h395dbec6),
	.w6(32'hbab84832),
	.w7(32'hb9e32e0e),
	.w8(32'h39065b76),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8688ae2),
	.w1(32'hb94b67b9),
	.w2(32'hb906b6fa),
	.w3(32'hb61ae36f),
	.w4(32'hb810f586),
	.w5(32'hb75875e0),
	.w6(32'h391e98e8),
	.w7(32'h38553e51),
	.w8(32'hb9a0a5d3),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf918e),
	.w1(32'h3aa84705),
	.w2(32'h3aa48d3a),
	.w3(32'hbbba8763),
	.w4(32'h3b750691),
	.w5(32'h3bfefa45),
	.w6(32'hbbca6646),
	.w7(32'h3a5fc8c1),
	.w8(32'h39f76c29),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8133605),
	.w1(32'hb991205e),
	.w2(32'hb9a8605d),
	.w3(32'h385e6792),
	.w4(32'h379eea31),
	.w5(32'hba03621c),
	.w6(32'hb849326f),
	.w7(32'hb9852a82),
	.w8(32'hb9ce8ac3),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb91de),
	.w1(32'h3b69cf14),
	.w2(32'h3b94c43d),
	.w3(32'hba408bde),
	.w4(32'hbb45918c),
	.w5(32'hbb863709),
	.w6(32'h39a8615c),
	.w7(32'h3b3a4eb9),
	.w8(32'h3ab99d5f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule