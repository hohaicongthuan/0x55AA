module layer_10_featuremap_457(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dca31),
	.w1(32'h3b2e42bb),
	.w2(32'hbb9c190b),
	.w3(32'hbb064990),
	.w4(32'h3c6a86db),
	.w5(32'h3c04a74d),
	.w6(32'hbb02f44d),
	.w7(32'hbb41435a),
	.w8(32'h3be9d45b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19181b),
	.w1(32'hba0ee82c),
	.w2(32'hbbeced1d),
	.w3(32'hbae6476d),
	.w4(32'hbbf0457d),
	.w5(32'h3a6be67c),
	.w6(32'h3a9499e6),
	.w7(32'hbb9c5f73),
	.w8(32'hbba15cfa),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c21b9),
	.w1(32'h3b2b0f84),
	.w2(32'hbadff085),
	.w3(32'hbbded579),
	.w4(32'h3aac9a5a),
	.w5(32'hbb8707f9),
	.w6(32'hbbbd069f),
	.w7(32'hba465144),
	.w8(32'hbbadbf4c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd541d),
	.w1(32'hb9cb6bc4),
	.w2(32'hbba0ab3b),
	.w3(32'hba46b682),
	.w4(32'hba0e3683),
	.w5(32'hbc6bbf98),
	.w6(32'h39af97dd),
	.w7(32'hba9d2107),
	.w8(32'hbb21445a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a70e8),
	.w1(32'hb9330015),
	.w2(32'hbb67a9af),
	.w3(32'h3ac88dba),
	.w4(32'hb8eb8769),
	.w5(32'hba9aaaa8),
	.w6(32'h3b6eda50),
	.w7(32'hbb4c7928),
	.w8(32'h3a762d1b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85e4cf),
	.w1(32'hbc11f261),
	.w2(32'hbc3b98e7),
	.w3(32'hbb4baad0),
	.w4(32'hbbccf1a9),
	.w5(32'hbc083c80),
	.w6(32'hbbafbb64),
	.w7(32'hbb42a909),
	.w8(32'hbc185969),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06b1ca),
	.w1(32'h3be2f9b1),
	.w2(32'h3bc7d10c),
	.w3(32'hbbab94a4),
	.w4(32'h3a5ab0ff),
	.w5(32'hbcabe6fe),
	.w6(32'hbbd6ac21),
	.w7(32'h3abb20c1),
	.w8(32'hbc1bccaa),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06f2d7),
	.w1(32'hbc4c1146),
	.w2(32'hbca826bf),
	.w3(32'hbb9ceaf3),
	.w4(32'hbc66536c),
	.w5(32'hbc97de81),
	.w6(32'hbbcc2c67),
	.w7(32'h3b0dc12b),
	.w8(32'hbc498fab),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb1c98),
	.w1(32'hbad4e66b),
	.w2(32'hbc1d222c),
	.w3(32'hbacd3a9b),
	.w4(32'hbbca75dc),
	.w5(32'hbc21b8a5),
	.w6(32'hbbefbdd2),
	.w7(32'hbb9f78f8),
	.w8(32'h3b75bf5d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc63f0),
	.w1(32'hb9c74a10),
	.w2(32'h3b862bad),
	.w3(32'hbc415fc9),
	.w4(32'hb9342fba),
	.w5(32'h3b8ec00e),
	.w6(32'hbb275928),
	.w7(32'hbb14ea0d),
	.w8(32'hbb09aa52),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b823d91),
	.w1(32'hbab6f2fe),
	.w2(32'hbaba26bd),
	.w3(32'h3b6df1b3),
	.w4(32'hbbfddcc3),
	.w5(32'h3a5e9415),
	.w6(32'h3ab21499),
	.w7(32'hbbfe7a17),
	.w8(32'hbbd660a6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2038d3),
	.w1(32'h3c466ab6),
	.w2(32'h3cbc8d92),
	.w3(32'h3b819594),
	.w4(32'h3c36a5c7),
	.w5(32'h3c3fad4c),
	.w6(32'hbaa72901),
	.w7(32'h3c008a49),
	.w8(32'h3b7d86e4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0424c7),
	.w1(32'hbc290bef),
	.w2(32'hbbca8e9e),
	.w3(32'h3c634668),
	.w4(32'hba87b975),
	.w5(32'hbc512d3b),
	.w6(32'h3bfb9999),
	.w7(32'hbaf10ce8),
	.w8(32'hbcb387cc),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0db7f3),
	.w1(32'hbb6e6298),
	.w2(32'hbc3f82ea),
	.w3(32'h3a2acd54),
	.w4(32'h3a4a9a35),
	.w5(32'hbb72e1c3),
	.w6(32'hbb9c5e68),
	.w7(32'h3bbd342f),
	.w8(32'h3a542a91),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3afdb1),
	.w1(32'h3b3ae912),
	.w2(32'hba8e4516),
	.w3(32'hbbe77a02),
	.w4(32'h3c174b0c),
	.w5(32'hba804165),
	.w6(32'h3a613187),
	.w7(32'h3b0961ec),
	.w8(32'h3b9a2fee),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab20fc5),
	.w1(32'h3c1a97ed),
	.w2(32'h3bfeef33),
	.w3(32'hbc078ae8),
	.w4(32'h3b4c83a1),
	.w5(32'h3c02b489),
	.w6(32'hbb9d1a27),
	.w7(32'hbbfbfc57),
	.w8(32'hbc0c1aad),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b949c01),
	.w1(32'h3a848012),
	.w2(32'hbab0c805),
	.w3(32'h3b0260b3),
	.w4(32'hbb41b26e),
	.w5(32'hbc2ec134),
	.w6(32'h3aa590cc),
	.w7(32'h3b72bc06),
	.w8(32'hbb30381b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69cad9),
	.w1(32'hba9e8b23),
	.w2(32'h3b45ed10),
	.w3(32'hbbe6b2ef),
	.w4(32'hba36c974),
	.w5(32'hbb800023),
	.w6(32'hbbc2c8b5),
	.w7(32'hb9bbd344),
	.w8(32'hba5ac884),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b605d),
	.w1(32'h3ad4a00a),
	.w2(32'h3bd363e7),
	.w3(32'hbaf2a06a),
	.w4(32'h3b03ca5a),
	.w5(32'hbb7d21aa),
	.w6(32'h3bbb0881),
	.w7(32'hbb6af0b7),
	.w8(32'hbbd7bbff),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b948ebb),
	.w1(32'hba2afd62),
	.w2(32'h3aa259db),
	.w3(32'h3aac4fbd),
	.w4(32'h3bccc56d),
	.w5(32'h3afd9d74),
	.w6(32'hbb274862),
	.w7(32'h3b6e1a0d),
	.w8(32'h3c5f37a8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb438cd2),
	.w1(32'hbac1d82d),
	.w2(32'hba8075e8),
	.w3(32'h3bff554d),
	.w4(32'hbb079dbc),
	.w5(32'hbbb6e1ef),
	.w6(32'h3aae5de8),
	.w7(32'hbb40d4ff),
	.w8(32'hbb4e9c2c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe2147),
	.w1(32'hbba8e8bb),
	.w2(32'hbb95a216),
	.w3(32'hbb164b0b),
	.w4(32'h3b40943b),
	.w5(32'hbb15d85d),
	.w6(32'hbb0905cf),
	.w7(32'hb99258b1),
	.w8(32'hbb88de6f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc63f53),
	.w1(32'hbb889d1f),
	.w2(32'hb9ac56d4),
	.w3(32'hbb8ab372),
	.w4(32'hbbd05faf),
	.w5(32'hbc20bf60),
	.w6(32'hbc415679),
	.w7(32'hbbe838b3),
	.w8(32'hbc22f96e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee980c),
	.w1(32'h3bf56603),
	.w2(32'h3bb95733),
	.w3(32'hbbce0ea7),
	.w4(32'h3c0f7a21),
	.w5(32'h3b8e3130),
	.w6(32'hbb07544c),
	.w7(32'h3b5045f0),
	.w8(32'h3b37ac7c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fb90a),
	.w1(32'hbb5a117d),
	.w2(32'hbbffed28),
	.w3(32'h3becab83),
	.w4(32'hbc6b5e7f),
	.w5(32'hbc05bb50),
	.w6(32'h3b97ffd5),
	.w7(32'hbb416e60),
	.w8(32'hbc05a904),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb41a71),
	.w1(32'hb713b9a7),
	.w2(32'hba81b8b5),
	.w3(32'hbb98c201),
	.w4(32'hbbbd52d6),
	.w5(32'hbb9196e0),
	.w6(32'h3bcc9ce9),
	.w7(32'h3a7e46c9),
	.w8(32'hbb3be155),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b48440),
	.w1(32'hbb56e1ff),
	.w2(32'hba0243db),
	.w3(32'h3b78503c),
	.w4(32'hbc096c21),
	.w5(32'hbc21b92f),
	.w6(32'h3b8b5084),
	.w7(32'hbbdeb557),
	.w8(32'hbbac92b4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc0271),
	.w1(32'h3989322d),
	.w2(32'hbb9d1153),
	.w3(32'hbb8226bf),
	.w4(32'hbc2b57e6),
	.w5(32'hb9c7c181),
	.w6(32'h3b86be5b),
	.w7(32'hbc443e46),
	.w8(32'h3b94863b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98f990),
	.w1(32'h3b755ed9),
	.w2(32'hbb3e6c61),
	.w3(32'hb9f0c16a),
	.w4(32'hbbfca86b),
	.w5(32'hbac6cc10),
	.w6(32'h3ad1bbcc),
	.w7(32'h3a8558e9),
	.w8(32'h3c3ce658),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01019a),
	.w1(32'h3c0d2d3a),
	.w2(32'h3c505440),
	.w3(32'hba48ce06),
	.w4(32'hbbee2d0a),
	.w5(32'h3b2f9be6),
	.w6(32'h3c072f5c),
	.w7(32'hbb15e5a4),
	.w8(32'h3b8432fb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cdfac),
	.w1(32'h3b8daa31),
	.w2(32'h3c014494),
	.w3(32'h3b27b6f1),
	.w4(32'h3abf020b),
	.w5(32'hbbe73a4e),
	.w6(32'hbb12d93e),
	.w7(32'h3b052176),
	.w8(32'h3c0ded60),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390dc3ff),
	.w1(32'hbb3a1984),
	.w2(32'h3a478be0),
	.w3(32'h3bb9a29c),
	.w4(32'h3b0f9263),
	.w5(32'hbaa11945),
	.w6(32'h3b8d1d83),
	.w7(32'h3c007663),
	.w8(32'hbb28de80),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d7cc5),
	.w1(32'h3b919cae),
	.w2(32'hba05d89a),
	.w3(32'hbacd5281),
	.w4(32'h3af7b10d),
	.w5(32'h3b8fc3f2),
	.w6(32'hbb547f49),
	.w7(32'h3b06cda9),
	.w8(32'h3b3ec0a5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad51876),
	.w1(32'h3b6017aa),
	.w2(32'hbb0a8415),
	.w3(32'hbbcc8593),
	.w4(32'h39b5c239),
	.w5(32'hbabbc58e),
	.w6(32'hbac33424),
	.w7(32'hbb2a0168),
	.w8(32'hbb7d4331),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d5868b),
	.w1(32'hba809fda),
	.w2(32'hba4bfb70),
	.w3(32'h3ad4831c),
	.w4(32'h3b5c80bc),
	.w5(32'hbbe0842f),
	.w6(32'hb825e94b),
	.w7(32'h3ab35262),
	.w8(32'hbb3cb942),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c3ba8),
	.w1(32'h3bb41cc2),
	.w2(32'h3b99c04f),
	.w3(32'h3b8b204e),
	.w4(32'h3c16bc38),
	.w5(32'h3ade521c),
	.w6(32'h3b282682),
	.w7(32'h3bac9f76),
	.w8(32'hbb0f068c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19d985),
	.w1(32'hbcc3fbcb),
	.w2(32'h3c71004a),
	.w3(32'hbd025eb8),
	.w4(32'h3c33297f),
	.w5(32'h3ce8de56),
	.w6(32'hbc4bdd50),
	.w7(32'h3cbb1fe8),
	.w8(32'h3c91907d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3eb819),
	.w1(32'hba9b5db8),
	.w2(32'hbb919a85),
	.w3(32'hbbae96b0),
	.w4(32'hb9f26478),
	.w5(32'hbb5ad513),
	.w6(32'hbb60124a),
	.w7(32'h3b1662b3),
	.w8(32'hbb24c7aa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cafc0a7),
	.w1(32'h3b81a581),
	.w2(32'hbc0ea5ac),
	.w3(32'h3bcb6a0a),
	.w4(32'h3a6dcf59),
	.w5(32'h3c157418),
	.w6(32'h3c123705),
	.w7(32'hbb6bfbf6),
	.w8(32'hbbc7c30a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c8c49),
	.w1(32'h38452343),
	.w2(32'h3ac08de4),
	.w3(32'h3a6aaabe),
	.w4(32'hba9b97dc),
	.w5(32'hbaff1555),
	.w6(32'h3a8fc2c0),
	.w7(32'h3b920316),
	.w8(32'hbaa3626b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5501a3),
	.w1(32'hbb2d12a4),
	.w2(32'h3b7e6db4),
	.w3(32'hbadfc1f7),
	.w4(32'hbb1ed55b),
	.w5(32'hb9368f6b),
	.w6(32'hbb49d0db),
	.w7(32'h3b191ba3),
	.w8(32'h3b81914f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b390279),
	.w1(32'hbb385d45),
	.w2(32'hbb9e3e96),
	.w3(32'hbb815b66),
	.w4(32'hba11a96d),
	.w5(32'hbb8b60fd),
	.w6(32'h3a0ad5f3),
	.w7(32'hba39ba49),
	.w8(32'h3a2f516f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb233742),
	.w1(32'hba82910c),
	.w2(32'h3b16a05d),
	.w3(32'hbac65b64),
	.w4(32'h3bb65e5f),
	.w5(32'h3a430be6),
	.w6(32'hbb6bf46d),
	.w7(32'h3bdebae3),
	.w8(32'hbac1d44a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc797a93),
	.w1(32'hbb9706b6),
	.w2(32'hbaab1c71),
	.w3(32'h3bc6fae3),
	.w4(32'hbb75f4fc),
	.w5(32'hbc3bf128),
	.w6(32'h3c1ec7cd),
	.w7(32'hbbab9c47),
	.w8(32'hbc3430a6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd56d17),
	.w1(32'h3a18e92f),
	.w2(32'h3ba0e0e5),
	.w3(32'hbc177f50),
	.w4(32'hbb4226f4),
	.w5(32'h3c06365e),
	.w6(32'hbbe41a32),
	.w7(32'h3a8a9ed5),
	.w8(32'h3bfe2acf),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87daac),
	.w1(32'h3b360ecf),
	.w2(32'h3c12d6f9),
	.w3(32'hbb341b86),
	.w4(32'h3c1df749),
	.w5(32'h3c7ea5db),
	.w6(32'hbb47f41b),
	.w7(32'h3bb86f47),
	.w8(32'h3b09a618),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b7c2c),
	.w1(32'hbbf6c240),
	.w2(32'hba92b101),
	.w3(32'hbb0ccd05),
	.w4(32'h3b2b9628),
	.w5(32'h3c05c393),
	.w6(32'hba2ecd58),
	.w7(32'hba8061cf),
	.w8(32'hbb51d384),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6203dc),
	.w1(32'h3c060ddb),
	.w2(32'h3b96be89),
	.w3(32'hbb201218),
	.w4(32'h3b901cfd),
	.w5(32'hba09dc94),
	.w6(32'hbb30616b),
	.w7(32'h3b8d65ef),
	.w8(32'hbc1fec7f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ba0b3),
	.w1(32'hba178eaf),
	.w2(32'hbac5a415),
	.w3(32'hb8c5dbae),
	.w4(32'hba935742),
	.w5(32'h3ae26aab),
	.w6(32'h3a89aac0),
	.w7(32'h3b4e44f1),
	.w8(32'h3c3392dc),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0533f),
	.w1(32'hbb179ece),
	.w2(32'hbaf47cd3),
	.w3(32'hba9061b9),
	.w4(32'h3b4759a2),
	.w5(32'h3b6ab041),
	.w6(32'h3aa06227),
	.w7(32'h3b905317),
	.w8(32'h3b628b4e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a7a49),
	.w1(32'h3c1d6396),
	.w2(32'h3b628ffe),
	.w3(32'h3a9e537a),
	.w4(32'hbb5c7e06),
	.w5(32'h3b7d3571),
	.w6(32'h3b007c37),
	.w7(32'hbbdc5b33),
	.w8(32'h3ba1095b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fd79c),
	.w1(32'h3b94a3d3),
	.w2(32'h3b8d9b8a),
	.w3(32'hbbe1b20a),
	.w4(32'h3b0a90f1),
	.w5(32'h3c82346a),
	.w6(32'hbb3ea219),
	.w7(32'h39f6d8cc),
	.w8(32'hba60575a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd15b0e),
	.w1(32'hbb7f9ddd),
	.w2(32'hbac9a379),
	.w3(32'h3c6de864),
	.w4(32'hbb6298e0),
	.w5(32'hbba5e12f),
	.w6(32'h3aeb467d),
	.w7(32'hbb812887),
	.w8(32'hbbf58953),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef2f37),
	.w1(32'hbb06bc66),
	.w2(32'hbbd689f1),
	.w3(32'hb9c04a95),
	.w4(32'hbb945829),
	.w5(32'hbb1ce2dc),
	.w6(32'h3aa28857),
	.w7(32'h3b869bdc),
	.w8(32'hbc2f0fb5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9e75c),
	.w1(32'hbbd2685b),
	.w2(32'h3a4b5d47),
	.w3(32'h3aad1d17),
	.w4(32'hbb63fc28),
	.w5(32'hbba71218),
	.w6(32'h3b0ebc15),
	.w7(32'h3b9f8f1b),
	.w8(32'hbac5f8a1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7decc),
	.w1(32'hbb4a9f9a),
	.w2(32'hbbf89987),
	.w3(32'h3bc035e3),
	.w4(32'h3b781d20),
	.w5(32'h399a99cc),
	.w6(32'hba387d24),
	.w7(32'h3bf1aa7c),
	.w8(32'h3bc3ba35),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd90fcc),
	.w1(32'h3b23ea03),
	.w2(32'h3b78e338),
	.w3(32'h3a35f440),
	.w4(32'hbb7bcd94),
	.w5(32'hbbb5b366),
	.w6(32'h3b016483),
	.w7(32'hbbb11564),
	.w8(32'hbbc51679),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b618b4f),
	.w1(32'hbbc54672),
	.w2(32'hbb473cc8),
	.w3(32'h3b4bad43),
	.w4(32'hb927e599),
	.w5(32'hbb8672af),
	.w6(32'h3ac177e4),
	.w7(32'hbb18a448),
	.w8(32'hbb84694c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb038ee),
	.w1(32'hbb056de5),
	.w2(32'h3b4b6e54),
	.w3(32'h3b077b8c),
	.w4(32'h3bc48300),
	.w5(32'hba899be8),
	.w6(32'hbbd56535),
	.w7(32'h3be5aa51),
	.w8(32'hbc11c20d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fd8df),
	.w1(32'hbb64ed97),
	.w2(32'h3b0df9db),
	.w3(32'h3b9ee2b5),
	.w4(32'hbb6a3a57),
	.w5(32'h3bdd1dbe),
	.w6(32'h3b1ae87e),
	.w7(32'h3c02a4b7),
	.w8(32'hbbc60560),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a9c74),
	.w1(32'h3ad0239f),
	.w2(32'h3b87ad81),
	.w3(32'h3bb6cd84),
	.w4(32'h3bb60741),
	.w5(32'hbb69ba6f),
	.w6(32'hbb5a241e),
	.w7(32'hb920a942),
	.w8(32'hbb34d6d4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadb1b3),
	.w1(32'hbb200acf),
	.w2(32'h3a92482a),
	.w3(32'hbb9d9c04),
	.w4(32'hbbcef0ca),
	.w5(32'h3a740e26),
	.w6(32'hb8da0703),
	.w7(32'hbc12bda4),
	.w8(32'h3bebac66),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb88b25),
	.w1(32'hba801a40),
	.w2(32'h3afbe768),
	.w3(32'h3b2d799a),
	.w4(32'hba44e5ea),
	.w5(32'h3a9f178f),
	.w6(32'h3991e18d),
	.w7(32'hbb4b0093),
	.w8(32'hbb7a1774),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fdf4f),
	.w1(32'h3af383de),
	.w2(32'h3be21820),
	.w3(32'h3b4ced40),
	.w4(32'h3c13e8c8),
	.w5(32'h3c477ce5),
	.w6(32'h35b54ede),
	.w7(32'hbbbc7b81),
	.w8(32'h3b1bf053),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6344b3),
	.w1(32'h3b5749b9),
	.w2(32'h3b71e6e3),
	.w3(32'h3c290ecf),
	.w4(32'h3bd478e5),
	.w5(32'h3a8d6307),
	.w6(32'h3b8363cb),
	.w7(32'h3b5c26ca),
	.w8(32'h3b3d67ac),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f995f),
	.w1(32'hbadd8a6d),
	.w2(32'hbbd2d7a6),
	.w3(32'h3b92302c),
	.w4(32'h39d06a2d),
	.w5(32'h3c38125b),
	.w6(32'h3ac9668c),
	.w7(32'h3ac5ce8d),
	.w8(32'h3ae0993c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01bda4),
	.w1(32'hbbcfe5e1),
	.w2(32'hba58dc3e),
	.w3(32'h3b0e9376),
	.w4(32'hbc0cf4b9),
	.w5(32'h384415d2),
	.w6(32'h3cb6ba13),
	.w7(32'hbc63b1b9),
	.w8(32'hbc96fc77),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8adeaa),
	.w1(32'h3b8c7a62),
	.w2(32'hbb267276),
	.w3(32'hbbfeb446),
	.w4(32'h3af32944),
	.w5(32'hbb4af835),
	.w6(32'hbc8c7982),
	.w7(32'h3a64dbf7),
	.w8(32'h3c2abf67),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6552),
	.w1(32'hbc21df3b),
	.w2(32'hbc6364cc),
	.w3(32'h3b10a805),
	.w4(32'hbc65ffe9),
	.w5(32'hbbec4974),
	.w6(32'h3a0ca310),
	.w7(32'hbc8e0438),
	.w8(32'hbc5864cc),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88690b),
	.w1(32'h3b688097),
	.w2(32'h3a8bea3d),
	.w3(32'hbc6ef7d9),
	.w4(32'hb8fa7cda),
	.w5(32'h3b8357b1),
	.w6(32'hbc17d716),
	.w7(32'hbb56e46f),
	.w8(32'h3ba240bb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ce0a1),
	.w1(32'h3aeb3301),
	.w2(32'h3acdfd7a),
	.w3(32'hbb048ba8),
	.w4(32'h3b0eba6f),
	.w5(32'h3abe01dd),
	.w6(32'hb9c4f9c0),
	.w7(32'h3ae4e3cf),
	.w8(32'h3af270c3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39647ef0),
	.w1(32'h39ab2da4),
	.w2(32'hbaa6d30d),
	.w3(32'h3ad64830),
	.w4(32'h3a498a96),
	.w5(32'h3a3908e5),
	.w6(32'h39e76d3d),
	.w7(32'h3a0cd88d),
	.w8(32'h3a97b832),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9361917),
	.w1(32'h3a35e4c7),
	.w2(32'h3b62b25a),
	.w3(32'h3a715b84),
	.w4(32'h39ffa21c),
	.w5(32'h3be3b1f5),
	.w6(32'h3a32cba2),
	.w7(32'h3795a0af),
	.w8(32'h3ba88ae2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981e5be),
	.w1(32'hba937d35),
	.w2(32'hba3f1684),
	.w3(32'h3b3bae9b),
	.w4(32'hb82d0d39),
	.w5(32'hba27250a),
	.w6(32'h3ae50151),
	.w7(32'hb6acc1c9),
	.w8(32'hbb1124c8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9abb60),
	.w1(32'hbb77b208),
	.w2(32'hbbac6f6d),
	.w3(32'hba1b5ec4),
	.w4(32'hbad14ea0),
	.w5(32'hbb104299),
	.w6(32'h391b4c4b),
	.w7(32'hbb5ea92a),
	.w8(32'hbbab7b45),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b5178),
	.w1(32'hbbf4b78f),
	.w2(32'hbb573ef4),
	.w3(32'hbb664f43),
	.w4(32'hbb2d4e09),
	.w5(32'hba948abb),
	.w6(32'hba9ed211),
	.w7(32'hbb25a854),
	.w8(32'hbbc2eb2c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba65616),
	.w1(32'hbb095141),
	.w2(32'h3aabdb2c),
	.w3(32'hbb5cb812),
	.w4(32'h3b829308),
	.w5(32'hbb27bec0),
	.w6(32'hbbdc4785),
	.w7(32'h3c11d84a),
	.w8(32'hbb259889),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8291b5a),
	.w1(32'h3abb65de),
	.w2(32'h3b8efe45),
	.w3(32'hbb782781),
	.w4(32'hbab5cd9c),
	.w5(32'h3b9a9020),
	.w6(32'h398fc526),
	.w7(32'hba81d5e0),
	.w8(32'h3b7b46c9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb14e2),
	.w1(32'h3ac80ee9),
	.w2(32'h3a35380b),
	.w3(32'h3b22ae9c),
	.w4(32'hba06e966),
	.w5(32'hba0bba13),
	.w6(32'h3b255572),
	.w7(32'h3a32f606),
	.w8(32'hbb1890e6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb238581),
	.w1(32'hbb7378a5),
	.w2(32'h3b66cb3c),
	.w3(32'hbb20b172),
	.w4(32'h3b01b2cd),
	.w5(32'h3b329180),
	.w6(32'h3bffffae),
	.w7(32'hbb2965e1),
	.w8(32'hbbe905ff),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad66d90),
	.w1(32'h3b0845f3),
	.w2(32'h3b0bca5a),
	.w3(32'hbb0d0089),
	.w4(32'h3a967de5),
	.w5(32'h3b82ae56),
	.w6(32'hb9c05da3),
	.w7(32'h3b154bc0),
	.w8(32'h3b97ffda),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabeb645),
	.w1(32'hba1cc77e),
	.w2(32'h3b28d71e),
	.w3(32'h3a560c8f),
	.w4(32'h38ccca6e),
	.w5(32'h3a221cb4),
	.w6(32'h3b2f7c26),
	.w7(32'h3a9893d1),
	.w8(32'hba76ab38),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac15e06),
	.w1(32'h3a140342),
	.w2(32'hb7a79587),
	.w3(32'h3a885aa1),
	.w4(32'h391f5d02),
	.w5(32'h37261496),
	.w6(32'h3a6428f7),
	.w7(32'hb91dd7e1),
	.w8(32'h366f8195),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68d10e),
	.w1(32'h3adf12a7),
	.w2(32'h3a3913b3),
	.w3(32'h3a4d23f2),
	.w4(32'h3b580ba1),
	.w5(32'hba001da5),
	.w6(32'h3a1523bc),
	.w7(32'h3b0eb523),
	.w8(32'h3afabf5c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370e8264),
	.w1(32'hba815f0e),
	.w2(32'h3ab5b290),
	.w3(32'hbaa19916),
	.w4(32'hba9a2b97),
	.w5(32'h3b15fc1e),
	.w6(32'hbab3ae47),
	.w7(32'hbab357ae),
	.w8(32'h3a88db96),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4ca05),
	.w1(32'hb98f267e),
	.w2(32'hbba4697d),
	.w3(32'h3ad2cc80),
	.w4(32'hbb738cb1),
	.w5(32'hbbe32b01),
	.w6(32'h3a99103c),
	.w7(32'hbb46eea6),
	.w8(32'hbb72b615),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c9782),
	.w1(32'h3acf3190),
	.w2(32'h3b8773e0),
	.w3(32'hbc16ff1e),
	.w4(32'h3b22462d),
	.w5(32'h3baabee6),
	.w6(32'hbbb333eb),
	.w7(32'hbab4eab3),
	.w8(32'h3b8af011),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e5034),
	.w1(32'hba1106cf),
	.w2(32'h3982cdd9),
	.w3(32'hba13dd4e),
	.w4(32'hbb1058f1),
	.w5(32'hbb0b349a),
	.w6(32'h3a23d41b),
	.w7(32'hba916158),
	.w8(32'h3abef5c6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b50d4),
	.w1(32'h39b602ed),
	.w2(32'h3b31a2fd),
	.w3(32'hbbfb617a),
	.w4(32'h3b6e0e13),
	.w5(32'h3b0c062e),
	.w6(32'hbba987fb),
	.w7(32'h3b51276b),
	.w8(32'h3b04eb53),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfeb59),
	.w1(32'h3b13c42d),
	.w2(32'hb92d87ce),
	.w3(32'h3a61102a),
	.w4(32'hbb01e6ab),
	.w5(32'hbbe6b1b9),
	.w6(32'hba7c1b0d),
	.w7(32'h3a3ddbbe),
	.w8(32'hbc25fbae),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cee41),
	.w1(32'hba27e456),
	.w2(32'h38f6720a),
	.w3(32'hba89e8e6),
	.w4(32'hba4d3bfc),
	.w5(32'h3afc0fcb),
	.w6(32'h3b7692eb),
	.w7(32'hba96d49c),
	.w8(32'h3904533c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc923f0a),
	.w1(32'h3b0812e9),
	.w2(32'h3c07128f),
	.w3(32'hbc553e3c),
	.w4(32'h3c5692d1),
	.w5(32'h3c505f84),
	.w6(32'hb949f929),
	.w7(32'h3b744072),
	.w8(32'hbbcd11e1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a5491),
	.w1(32'h3b4632a8),
	.w2(32'h3b2492b4),
	.w3(32'h3c041dd8),
	.w4(32'h3ac0e011),
	.w5(32'h39b4b84e),
	.w6(32'h3b13d70d),
	.w7(32'hb989e744),
	.w8(32'h3abea95e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dc8c3),
	.w1(32'h3abc4f58),
	.w2(32'hbb89a797),
	.w3(32'h3bb558c0),
	.w4(32'h39b5e380),
	.w5(32'hba793da2),
	.w6(32'h3bbe8bc8),
	.w7(32'h3b3643c8),
	.w8(32'hbb4b8704),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49ce01),
	.w1(32'hba63d779),
	.w2(32'hbb465810),
	.w3(32'hba9a4f07),
	.w4(32'h3b68db50),
	.w5(32'h3b96e8ed),
	.w6(32'h3c059a43),
	.w7(32'hbafcb020),
	.w8(32'hbb4651d9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b217ec4),
	.w1(32'hbb195ae4),
	.w2(32'hbb65cc24),
	.w3(32'hba22b4ce),
	.w4(32'hba6a74bc),
	.w5(32'h3a7eb348),
	.w6(32'h3b251bee),
	.w7(32'hba75911d),
	.w8(32'h3a2e293b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ff3dc6),
	.w1(32'hba155cb4),
	.w2(32'hb9486d10),
	.w3(32'h3b22d70f),
	.w4(32'h3a28317a),
	.w5(32'h3a328795),
	.w6(32'h3af0e203),
	.w7(32'h39f4596e),
	.w8(32'hb957383d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f3a82),
	.w1(32'hb9315a10),
	.w2(32'hba8964c4),
	.w3(32'h3b57f016),
	.w4(32'hbac45741),
	.w5(32'hbb8edc29),
	.w6(32'h3b7b3095),
	.w7(32'h3a7f546a),
	.w8(32'hbc365e57),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12bf1e),
	.w1(32'hbbd263e2),
	.w2(32'h3c10a335),
	.w3(32'hbacd57a2),
	.w4(32'h3bfa8cd1),
	.w5(32'h3c24a297),
	.w6(32'h3c3eb5ed),
	.w7(32'hbafcbf4a),
	.w8(32'hbbbe9a58),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8ad4d),
	.w1(32'h39a049de),
	.w2(32'h3b6855ca),
	.w3(32'hbc9d1e65),
	.w4(32'h3ca0f99e),
	.w5(32'h3c437828),
	.w6(32'hbd04de6e),
	.w7(32'h3bd7acc0),
	.w8(32'h3c981758),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a0dc3),
	.w1(32'hbb442dff),
	.w2(32'hb96c8df3),
	.w3(32'hbabb32ff),
	.w4(32'h3bf3f25a),
	.w5(32'h3bb3e286),
	.w6(32'hbb23ff48),
	.w7(32'h3af6db2f),
	.w8(32'h3b942507),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae64cd1),
	.w1(32'h3a7c3ab5),
	.w2(32'h3ae1f000),
	.w3(32'h3a2022ce),
	.w4(32'hb9b5d045),
	.w5(32'h3b1a88a3),
	.w6(32'h3a7a8c55),
	.w7(32'hba0e2265),
	.w8(32'h3b1ec64d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc936db5),
	.w1(32'hbbb05351),
	.w2(32'h3c11deea),
	.w3(32'hbb6716e1),
	.w4(32'h3c8c4938),
	.w5(32'h3beefa86),
	.w6(32'hb89c2fa6),
	.w7(32'h3c5d28ed),
	.w8(32'h39298239),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9442cf),
	.w1(32'h3a1bc1e5),
	.w2(32'h3a78f564),
	.w3(32'h3b3ca051),
	.w4(32'h3ae6a386),
	.w5(32'h3b3a97d4),
	.w6(32'h3b333086),
	.w7(32'h3b3503b2),
	.w8(32'h39751bed),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1a3dcf),
	.w1(32'hbc68eee7),
	.w2(32'hbaa00e5e),
	.w3(32'hbcf177eb),
	.w4(32'h3cbb5df5),
	.w5(32'h3c9d40e9),
	.w6(32'hbc98a4d6),
	.w7(32'h3c9a4b60),
	.w8(32'h3cd56fe3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52678e),
	.w1(32'hbb601dd5),
	.w2(32'h3af26673),
	.w3(32'hbb2d9d51),
	.w4(32'h3b831a70),
	.w5(32'hba817566),
	.w6(32'hbb78162a),
	.w7(32'h3b8d31d1),
	.w8(32'h3b907de4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b56b0),
	.w1(32'h3ad57a55),
	.w2(32'h3a42b131),
	.w3(32'h3ac56485),
	.w4(32'h3a5b2ff4),
	.w5(32'h3ac59306),
	.w6(32'h3b0bf5c0),
	.w7(32'h3b05f1a1),
	.w8(32'h3aacc583),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa86b7c),
	.w1(32'hba91109e),
	.w2(32'hbae73c2e),
	.w3(32'hbabeddf4),
	.w4(32'hbb3a2d57),
	.w5(32'h3a00f978),
	.w6(32'hba63815e),
	.w7(32'hbbcbbf81),
	.w8(32'hbb10e001),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9f768),
	.w1(32'h3b9a3fa8),
	.w2(32'h3b9351c8),
	.w3(32'h3b31bd76),
	.w4(32'h3b3d5644),
	.w5(32'h396316c3),
	.w6(32'h3b36431a),
	.w7(32'h39a11e3b),
	.w8(32'hbbadb1c6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac98bac),
	.w1(32'h3b8afeb5),
	.w2(32'hbab82eb7),
	.w3(32'h3b13b2c5),
	.w4(32'h3b1269a9),
	.w5(32'hba3d8bd8),
	.w6(32'h3b4125e4),
	.w7(32'hba0ba2b2),
	.w8(32'hba8ab8cd),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3eaddd),
	.w1(32'h3aa6d8ef),
	.w2(32'hbb1caa12),
	.w3(32'h398ac423),
	.w4(32'h3a27dbe9),
	.w5(32'h3b4f7fbb),
	.w6(32'h3ba1ce84),
	.w7(32'hbb2bf9e5),
	.w8(32'hbac6ed6b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3b351),
	.w1(32'hb9c37ab1),
	.w2(32'h398efe7a),
	.w3(32'hbbddfdd7),
	.w4(32'hba0e7672),
	.w5(32'h3aac997f),
	.w6(32'hbb0e28b3),
	.w7(32'h3a02f506),
	.w8(32'hba0606b0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffa109),
	.w1(32'h3b53105e),
	.w2(32'h3b946817),
	.w3(32'hbc52cafc),
	.w4(32'hb8b3bb74),
	.w5(32'h3be27625),
	.w6(32'hbc641268),
	.w7(32'h3b22015a),
	.w8(32'h3bdfb995),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7b655),
	.w1(32'hbba31e30),
	.w2(32'hbbf460df),
	.w3(32'hbb2403ea),
	.w4(32'hbbbf3509),
	.w5(32'hba5deff6),
	.w6(32'h3b1aa168),
	.w7(32'hbc197283),
	.w8(32'hbb995a81),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13def8),
	.w1(32'h3aadbc25),
	.w2(32'h3b526d8d),
	.w3(32'hbac19fa6),
	.w4(32'h3b075fcf),
	.w5(32'h3b86fe46),
	.w6(32'hba364a4e),
	.w7(32'h3a8fc969),
	.w8(32'h3b95b7f1),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a9ed4),
	.w1(32'hbabf455b),
	.w2(32'h39b23731),
	.w3(32'h3b0c8f97),
	.w4(32'hbb11f728),
	.w5(32'hbadfe352),
	.w6(32'h3acc16e3),
	.w7(32'hbabcaeaa),
	.w8(32'hba91f23d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0f6c0),
	.w1(32'hba98f86c),
	.w2(32'hb9041fda),
	.w3(32'hbb40d7ad),
	.w4(32'h38cc6d79),
	.w5(32'h3b4d757d),
	.w6(32'hba73c9ea),
	.w7(32'hba358189),
	.w8(32'h3a351a18),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26edb7),
	.w1(32'hba3de5c7),
	.w2(32'h3a333ad5),
	.w3(32'h3ae845d3),
	.w4(32'h3a8f17cb),
	.w5(32'h3abb95ec),
	.w6(32'h3adbca58),
	.w7(32'h3adb51d9),
	.w8(32'h39e8c96d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec277f),
	.w1(32'h3a034456),
	.w2(32'h3a96263f),
	.w3(32'h3b3a6028),
	.w4(32'h39ef2c99),
	.w5(32'hb98095f0),
	.w6(32'h3b00ab62),
	.w7(32'h3ad3e2b0),
	.w8(32'h3a97e980),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39460ac4),
	.w1(32'h3b66cdf4),
	.w2(32'h3baf26b3),
	.w3(32'hba46eda5),
	.w4(32'h3b7f5a0c),
	.w5(32'h3c054a70),
	.w6(32'h3a7adbba),
	.w7(32'h3b254d9b),
	.w8(32'h3bba9de3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b069101),
	.w1(32'h39ffd74a),
	.w2(32'hb9fd5b1e),
	.w3(32'h3b6a72f6),
	.w4(32'h3a8c5908),
	.w5(32'hb9e3985d),
	.w6(32'h3b707fb2),
	.w7(32'h3a7ad533),
	.w8(32'h386bae66),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb448bd2),
	.w1(32'hbb2e1a1d),
	.w2(32'hb980594c),
	.w3(32'hbb25ac2f),
	.w4(32'hba58a762),
	.w5(32'hbabc4ddc),
	.w6(32'hbb008b0a),
	.w7(32'h3ae3856a),
	.w8(32'hbb59f6e0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28fd38),
	.w1(32'h3a4f9e2a),
	.w2(32'h37c6528f),
	.w3(32'hbbc8e87a),
	.w4(32'hbb62283a),
	.w5(32'hba14d57a),
	.w6(32'hba6e0cce),
	.w7(32'hba9fddca),
	.w8(32'h3aa28b97),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3242f8),
	.w1(32'hb9c087bf),
	.w2(32'hbaa26f1f),
	.w3(32'hb9c4cb14),
	.w4(32'hb9fe4351),
	.w5(32'h388c1f2d),
	.w6(32'hba2a93e7),
	.w7(32'hb9b7bf6c),
	.w8(32'hba36e0c5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84fac1),
	.w1(32'hba429616),
	.w2(32'hba508bb8),
	.w3(32'hb80c5f7e),
	.w4(32'h3a5b202c),
	.w5(32'hba5b4787),
	.w6(32'h3a250b0b),
	.w7(32'hbaeae910),
	.w8(32'hbad91738),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49a32e),
	.w1(32'hbb1eb4ba),
	.w2(32'hba996d16),
	.w3(32'h39a12e17),
	.w4(32'hbabb0f7c),
	.w5(32'hb925fffc),
	.w6(32'hb97e1238),
	.w7(32'hbb2bd901),
	.w8(32'hb9c8c607),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba901dc4),
	.w1(32'h39bdec57),
	.w2(32'hba1242eb),
	.w3(32'h39a58d94),
	.w4(32'hba2797fe),
	.w5(32'hbbc811c7),
	.w6(32'h39fe2709),
	.w7(32'hb9cd6eb1),
	.w8(32'hbb4318b5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967d20),
	.w1(32'h3b3cb31e),
	.w2(32'hbb53decc),
	.w3(32'h3afaba9a),
	.w4(32'hba651c7f),
	.w5(32'hbc5e211c),
	.w6(32'hbc445e2c),
	.w7(32'h3a6f3729),
	.w8(32'hbae318eb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78fc3d),
	.w1(32'h3a533d63),
	.w2(32'h3ab9a183),
	.w3(32'h38a7419c),
	.w4(32'hbb28fd0f),
	.w5(32'hbb2049b9),
	.w6(32'h3b75c8ad),
	.w7(32'hba52214e),
	.w8(32'hbbc0b50c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20ec8a),
	.w1(32'hbab4fe33),
	.w2(32'hbb145927),
	.w3(32'hba302fee),
	.w4(32'hbaad5ef0),
	.w5(32'hbb0b9ed3),
	.w6(32'h3a47bad4),
	.w7(32'hb98377f5),
	.w8(32'hbb215177),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb99ee),
	.w1(32'hbc0399b4),
	.w2(32'hbbb35c3c),
	.w3(32'hb891af2d),
	.w4(32'hbb7367df),
	.w5(32'hbb594dbd),
	.w6(32'hbb37b0eb),
	.w7(32'hbb2c93a1),
	.w8(32'hbb0184c3),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02bf9f),
	.w1(32'hbb01ed94),
	.w2(32'hb82ce8c8),
	.w3(32'hbb465cc3),
	.w4(32'hbac80cf5),
	.w5(32'h3b8d8cd8),
	.w6(32'hbac48925),
	.w7(32'hbaeb0ed7),
	.w8(32'h3a66cb74),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbfaca),
	.w1(32'hb9cf99a7),
	.w2(32'hbaa81b53),
	.w3(32'h3afed56d),
	.w4(32'hbb2852e1),
	.w5(32'hbaea6415),
	.w6(32'h3b300395),
	.w7(32'hbae6ef65),
	.w8(32'hbb4bf483),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4bf52),
	.w1(32'hba05a5f6),
	.w2(32'hb92b947d),
	.w3(32'hbb046ea4),
	.w4(32'h39889d07),
	.w5(32'h3bd5648e),
	.w6(32'h3b2f06c4),
	.w7(32'hbb010869),
	.w8(32'h3b4a777b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac36fd),
	.w1(32'hba97f1c8),
	.w2(32'h3aec2804),
	.w3(32'h3a850cb0),
	.w4(32'hba63d365),
	.w5(32'hba6930ae),
	.w6(32'h3b3da643),
	.w7(32'h3aea71ce),
	.w8(32'hbbd659e5),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ac47d),
	.w1(32'hb9e01c95),
	.w2(32'h3aee6dcc),
	.w3(32'hbb70227c),
	.w4(32'hb990a368),
	.w5(32'h3ae0c1ea),
	.w6(32'hbb15cc69),
	.w7(32'h3a29e45d),
	.w8(32'h3b098f63),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba229d),
	.w1(32'hbacca081),
	.w2(32'h3902042d),
	.w3(32'h395cd4d4),
	.w4(32'h3b337773),
	.w5(32'h3babc69a),
	.w6(32'h3a8d8a1e),
	.w7(32'hbb10d3f5),
	.w8(32'h39036ed4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1ea3a),
	.w1(32'hbb4c3b94),
	.w2(32'hbb232c0b),
	.w3(32'hb8ff7267),
	.w4(32'h3b2cbd43),
	.w5(32'hba2c1fae),
	.w6(32'h3ae99a11),
	.w7(32'h3b84ff87),
	.w8(32'hbb3833b5),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb0c7a),
	.w1(32'h39befcbb),
	.w2(32'h3829df46),
	.w3(32'hbbd2cea9),
	.w4(32'h38eda926),
	.w5(32'h3b4885ff),
	.w6(32'hbc0d9032),
	.w7(32'hbb66f67c),
	.w8(32'h3b8c6d11),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba92ac9),
	.w1(32'h3a0edaf7),
	.w2(32'h3ba4dc57),
	.w3(32'hbb084b1d),
	.w4(32'h3b309fde),
	.w5(32'hba6daa88),
	.w6(32'h3b2b09ec),
	.w7(32'h3b062448),
	.w8(32'hbb91831f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5edec7),
	.w1(32'hb922cf84),
	.w2(32'h39be7e84),
	.w3(32'hbb159df9),
	.w4(32'hb9f2d299),
	.w5(32'h39d55161),
	.w6(32'hb9fab698),
	.w7(32'hba9d912f),
	.w8(32'h3a7fa454),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd6268),
	.w1(32'h3b1afc81),
	.w2(32'h3a61508c),
	.w3(32'h3a446595),
	.w4(32'hbb3b49fc),
	.w5(32'h3ab07555),
	.w6(32'h3bb9a903),
	.w7(32'hbb55a036),
	.w8(32'hbb026018),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a924c7c),
	.w1(32'h371c39ba),
	.w2(32'h3b1b299e),
	.w3(32'hba8b47ac),
	.w4(32'hb91b64ec),
	.w5(32'h3b045b3f),
	.w6(32'h3a568717),
	.w7(32'h3a267647),
	.w8(32'h3af50e6d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2f5a4),
	.w1(32'h3afde6e5),
	.w2(32'h3aeeed6e),
	.w3(32'h3a96144f),
	.w4(32'h3b00e485),
	.w5(32'hba0d6cfe),
	.w6(32'hb75ba06c),
	.w7(32'h3b11826a),
	.w8(32'h3ad4dcf0),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a532164),
	.w1(32'hb933bbd2),
	.w2(32'hb9c78207),
	.w3(32'hbaf00b79),
	.w4(32'hba5b80c5),
	.w5(32'hbb123ad1),
	.w6(32'hba9598ff),
	.w7(32'hbaf6ea2f),
	.w8(32'hbb223683),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacdef9),
	.w1(32'hbae54874),
	.w2(32'h3abe11b0),
	.w3(32'hbb56a185),
	.w4(32'h3a876141),
	.w5(32'h3aa84b4f),
	.w6(32'hbada7f39),
	.w7(32'h3a75ed44),
	.w8(32'h3b261f4a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4688c),
	.w1(32'hbaa9e8f1),
	.w2(32'h3abb106d),
	.w3(32'hbbc92789),
	.w4(32'h3a1f8d28),
	.w5(32'h3ba78848),
	.w6(32'hbb6ef3d3),
	.w7(32'h3b39bc26),
	.w8(32'h3be7ed12),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29387b),
	.w1(32'h3acdb2c1),
	.w2(32'h3a688f10),
	.w3(32'hba6697ea),
	.w4(32'hba04629b),
	.w5(32'hbb3c16b4),
	.w6(32'h39fce566),
	.w7(32'h38aa3f54),
	.w8(32'hbb46f0e8),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5511a9),
	.w1(32'h3a8c6afe),
	.w2(32'h3ab17136),
	.w3(32'hbaeecc0e),
	.w4(32'h3aefaf5f),
	.w5(32'h3aa10351),
	.w6(32'hba8acbde),
	.w7(32'h3b3dc522),
	.w8(32'h3b376463),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43f1d3),
	.w1(32'hba6925ee),
	.w2(32'h39359fbd),
	.w3(32'h3ac41eff),
	.w4(32'hb9265eae),
	.w5(32'hbb5e01cc),
	.w6(32'h3ba44815),
	.w7(32'hba0ed496),
	.w8(32'hbb9509fb),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1d78a),
	.w1(32'hb9a7947a),
	.w2(32'hbabb81f5),
	.w3(32'h3ae709a4),
	.w4(32'h3a3cf540),
	.w5(32'hbb65cb3e),
	.w6(32'hba00d767),
	.w7(32'hbaf0a501),
	.w8(32'hbb8f90e0),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42246f),
	.w1(32'hbbb71e71),
	.w2(32'hbb8e03c9),
	.w3(32'hbb5da786),
	.w4(32'h3b1202d4),
	.w5(32'hbb00e31a),
	.w6(32'h3935d0be),
	.w7(32'h3abdb8d7),
	.w8(32'hbbc0f947),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87940a),
	.w1(32'h3a86a628),
	.w2(32'h3aa6df4c),
	.w3(32'hbb8cf075),
	.w4(32'hbb5578cf),
	.w5(32'h3bf5f365),
	.w6(32'h3b065f83),
	.w7(32'hbbac266a),
	.w8(32'h3abcc2ac),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba94bd7),
	.w1(32'h3b96d3fd),
	.w2(32'h3b6fc09d),
	.w3(32'h3b4ac5a3),
	.w4(32'h3b891c42),
	.w5(32'h3b995deb),
	.w6(32'h3bacb420),
	.w7(32'h3b74f991),
	.w8(32'h3b2d85a0),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21b127),
	.w1(32'hbb547f6a),
	.w2(32'hbb96d3c2),
	.w3(32'h3b9b2cb3),
	.w4(32'hb9262b70),
	.w5(32'h3ae98ae6),
	.w6(32'h3bc74b37),
	.w7(32'h3a2e43f2),
	.w8(32'hb9cc6548),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbac307),
	.w1(32'hb8f2f05b),
	.w2(32'h3b41eea5),
	.w3(32'hbbb1397e),
	.w4(32'hba8fb3f3),
	.w5(32'h3bc14333),
	.w6(32'hbb9fe5e3),
	.w7(32'h3b069390),
	.w8(32'h3be992c5),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fdb9e),
	.w1(32'hba95fce5),
	.w2(32'h3a9e3f30),
	.w3(32'h3a26b575),
	.w4(32'hba2fd031),
	.w5(32'h3b6737ee),
	.w6(32'h3a9c3210),
	.w7(32'hbaffb499),
	.w8(32'h3b27cd3e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb41c6a),
	.w1(32'h3ab5e857),
	.w2(32'h3b434ce8),
	.w3(32'h3a70708f),
	.w4(32'h39519349),
	.w5(32'h3a3ea829),
	.w6(32'h3aca4c94),
	.w7(32'hb9f7b20a),
	.w8(32'h3aae995f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb116d23),
	.w1(32'h3a0c6b0e),
	.w2(32'h3a4dca0d),
	.w3(32'h39302378),
	.w4(32'h3b72dafa),
	.w5(32'h399aeb07),
	.w6(32'h3a93255c),
	.w7(32'h3b6fbe0b),
	.w8(32'hbac0dc39),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ef6ba),
	.w1(32'h3876d58e),
	.w2(32'h3998d0bd),
	.w3(32'hb99f006d),
	.w4(32'hb960f2c2),
	.w5(32'h3b10cede),
	.w6(32'h38ecb5a0),
	.w7(32'hb8222204),
	.w8(32'h3a8e9cc1),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97fcbb),
	.w1(32'hba2444ac),
	.w2(32'h383b7e87),
	.w3(32'h399a2f05),
	.w4(32'hbaea00e8),
	.w5(32'hbb0d34ff),
	.w6(32'h3ad81ba8),
	.w7(32'hba790f9c),
	.w8(32'hbb82202f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b800d),
	.w1(32'hb9f4988d),
	.w2(32'hbaffc57d),
	.w3(32'hba52288c),
	.w4(32'hba5cb7d0),
	.w5(32'hbab798eb),
	.w6(32'hbaf30314),
	.w7(32'hba9bc7ce),
	.w8(32'h3a0faa4c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7fd3f),
	.w1(32'h3ac2530e),
	.w2(32'h3ac3bae4),
	.w3(32'hba6e7def),
	.w4(32'hbb01c121),
	.w5(32'h3b085197),
	.w6(32'hb9fcf228),
	.w7(32'hbad9c782),
	.w8(32'h3b42aabc),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12ffb8),
	.w1(32'h3ab3d08b),
	.w2(32'h3a3b3e22),
	.w3(32'h3a40cb93),
	.w4(32'h3ac6ceb7),
	.w5(32'h3a7cf11f),
	.w6(32'h3af23513),
	.w7(32'h3b03c055),
	.w8(32'h3b2ffcd7),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09a463),
	.w1(32'h3a97d96c),
	.w2(32'hbb0c45e7),
	.w3(32'h3bf475f7),
	.w4(32'hbb97bf84),
	.w5(32'hbbd4b6e3),
	.w6(32'h3bb1134f),
	.w7(32'hbb4fff40),
	.w8(32'hbbd547b0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a987cf1),
	.w1(32'h3a80dddc),
	.w2(32'h3a712e62),
	.w3(32'hba5af5e9),
	.w4(32'h3a7c4b14),
	.w5(32'h3abaa806),
	.w6(32'hb9eaae72),
	.w7(32'h3aafa3b1),
	.w8(32'h3a293982),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1679e),
	.w1(32'hbb434244),
	.w2(32'hbb2e4da6),
	.w3(32'hba0bd43f),
	.w4(32'hbaf46633),
	.w5(32'hbb714d5f),
	.w6(32'h36a35014),
	.w7(32'hbab47f70),
	.w8(32'hbb33906f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93446a),
	.w1(32'hba82f98d),
	.w2(32'hba46030c),
	.w3(32'hbb65b8a5),
	.w4(32'h38d691ca),
	.w5(32'h3b1c59e1),
	.w6(32'hbab17765),
	.w7(32'h3a4c40c7),
	.w8(32'h3b35b62b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf416a6),
	.w1(32'h3bcb9e98),
	.w2(32'h3b92eb21),
	.w3(32'hbb789557),
	.w4(32'h3becacf5),
	.w5(32'hbacf8a89),
	.w6(32'hbc16200b),
	.w7(32'h3c17e004),
	.w8(32'h3aaa4281),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2ffd8),
	.w1(32'h3ac7ba90),
	.w2(32'hba0e6ff1),
	.w3(32'h3b7a650b),
	.w4(32'hb9bb2d7f),
	.w5(32'hbaa81141),
	.w6(32'h3bad936a),
	.w7(32'h3b191750),
	.w8(32'h3a96fed4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12a41b),
	.w1(32'h3b08e0bc),
	.w2(32'h3a426fb1),
	.w3(32'h38cfa0ab),
	.w4(32'h3a8d5ab3),
	.w5(32'h3b60e773),
	.w6(32'h3b47551e),
	.w7(32'h3a874d88),
	.w8(32'h3b0093e6),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae72eb),
	.w1(32'h3b0ec005),
	.w2(32'h3b269c9e),
	.w3(32'h39be602d),
	.w4(32'hbb350319),
	.w5(32'h3a86b860),
	.w6(32'h3aaf474f),
	.w7(32'hbb2d464a),
	.w8(32'h39c54428),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb86cf),
	.w1(32'hba7c7b1a),
	.w2(32'h3b183ea7),
	.w3(32'h3abec897),
	.w4(32'hb9a9b08b),
	.w5(32'hb88fe878),
	.w6(32'h3adb4b06),
	.w7(32'hbac023bb),
	.w8(32'hbb78f682),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a982f),
	.w1(32'h3b18f7e3),
	.w2(32'hbacbf383),
	.w3(32'hb940232a),
	.w4(32'h3b43068e),
	.w5(32'hbb3849b1),
	.w6(32'h3ac9bd94),
	.w7(32'h3b364b8b),
	.w8(32'h39c7d4f5),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba34095),
	.w1(32'h3af96a0f),
	.w2(32'h3986632f),
	.w3(32'h3a9c16ee),
	.w4(32'h3b472612),
	.w5(32'hbaa568b3),
	.w6(32'h3b1cb985),
	.w7(32'h3b885573),
	.w8(32'hbb66789b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49febd),
	.w1(32'h3b5bcac1),
	.w2(32'h3b6de935),
	.w3(32'h3aa51780),
	.w4(32'h3b8ab9c5),
	.w5(32'h3b45f5be),
	.w6(32'h391cc764),
	.w7(32'h3ba1ad85),
	.w8(32'h3b7dad12),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba465a51),
	.w1(32'h3b38d140),
	.w2(32'h3b64efdd),
	.w3(32'h3b49ab97),
	.w4(32'h3a97e636),
	.w5(32'h3b96b7c1),
	.w6(32'h3bd79809),
	.w7(32'h3b06de5f),
	.w8(32'h3ae3317b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2eb35),
	.w1(32'h3af4371a),
	.w2(32'h3ae90feb),
	.w3(32'h3b0bdf95),
	.w4(32'h3a81fe4d),
	.w5(32'h3aa44c34),
	.w6(32'h3b3638f1),
	.w7(32'h3ad6d14c),
	.w8(32'h3afda804),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3aba2),
	.w1(32'h399551e9),
	.w2(32'h3ad9f699),
	.w3(32'h3b0806bb),
	.w4(32'h39ffe332),
	.w5(32'hb921e6c0),
	.w6(32'h3b38f727),
	.w7(32'h3aba68b3),
	.w8(32'h3a1881c5),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae04a02),
	.w1(32'hbb3b382a),
	.w2(32'hbb44b65e),
	.w3(32'hba56d96a),
	.w4(32'hbb151463),
	.w5(32'hbb216150),
	.w6(32'h3a1f5a32),
	.w7(32'hbb0275bf),
	.w8(32'hbb37104a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b9f7f),
	.w1(32'h3a8d47a6),
	.w2(32'hbafd6bfa),
	.w3(32'h38afd920),
	.w4(32'hbb2d0196),
	.w5(32'h393c275f),
	.w6(32'h39fa26ed),
	.w7(32'hbb9f2819),
	.w8(32'hbb2f3c10),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29b6f8),
	.w1(32'h3b0f3e53),
	.w2(32'h3ae4a9ce),
	.w3(32'hb96453ad),
	.w4(32'h3a8b876f),
	.w5(32'h3b430f9e),
	.w6(32'h39903bd6),
	.w7(32'h3aee4180),
	.w8(32'h3b54126e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45911f),
	.w1(32'h38262e8a),
	.w2(32'h3ad64d74),
	.w3(32'h3af190b0),
	.w4(32'hb9f3a586),
	.w5(32'h3b1f89b0),
	.w6(32'h3b155015),
	.w7(32'hbab69209),
	.w8(32'h3a24ddfd),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a821511),
	.w1(32'hb9f44444),
	.w2(32'h3afbd727),
	.w3(32'hbab4938d),
	.w4(32'hbb1293cc),
	.w5(32'h3ba2eb40),
	.w6(32'hb99707f3),
	.w7(32'hbb7aee35),
	.w8(32'h3a2a9268),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e637e),
	.w1(32'h39b061c4),
	.w2(32'h39af4534),
	.w3(32'h3ad2302b),
	.w4(32'h3bc48923),
	.w5(32'h3a4dfa6f),
	.w6(32'h39e38368),
	.w7(32'h3b0c8453),
	.w8(32'hbb8b0cc0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d2195),
	.w1(32'hbc07ab8c),
	.w2(32'h3aec70bd),
	.w3(32'hbc70e0f7),
	.w4(32'h3b5da241),
	.w5(32'h3bd48fc2),
	.w6(32'hbbedf201),
	.w7(32'h3be7b328),
	.w8(32'h3b9e8edc),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb460f13),
	.w1(32'hbb3347ba),
	.w2(32'hbb32bb6d),
	.w3(32'hbb4b57d1),
	.w4(32'hbb8fa023),
	.w5(32'hbb77b244),
	.w6(32'hbad6c984),
	.w7(32'hbb6328bb),
	.w8(32'hbb58acc9),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30576c),
	.w1(32'hb93f9560),
	.w2(32'hbb71a0b7),
	.w3(32'h3adcd207),
	.w4(32'h3b924d98),
	.w5(32'hbbc8b0fb),
	.w6(32'h38b5dd5e),
	.w7(32'h3b12f3df),
	.w8(32'hbc15fcdb),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a809cc0),
	.w1(32'h3a9d96c5),
	.w2(32'h3bacc68e),
	.w3(32'hbb99fe85),
	.w4(32'h3a73d3ff),
	.w5(32'h3c9bc075),
	.w6(32'h3c02c8b5),
	.w7(32'hbb817550),
	.w8(32'h3b0f6245),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84bc86),
	.w1(32'hba8c231f),
	.w2(32'h3ada80ce),
	.w3(32'hb7b8e6ee),
	.w4(32'h39a76742),
	.w5(32'h3b7c0c69),
	.w6(32'hba31ccf3),
	.w7(32'hb93116bf),
	.w8(32'hbaa22092),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01fc9a),
	.w1(32'hb9fc2cff),
	.w2(32'hba17640e),
	.w3(32'h3a5496d0),
	.w4(32'hba675ff1),
	.w5(32'hb9b97bcb),
	.w6(32'h3a12ba1d),
	.w7(32'hba7d9d3e),
	.w8(32'hb9ddaeed),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b999a),
	.w1(32'hb753c81a),
	.w2(32'hba3d9029),
	.w3(32'hb986f26e),
	.w4(32'h3a48efe4),
	.w5(32'hbaa33453),
	.w6(32'h3a78b26d),
	.w7(32'h3a38f2f9),
	.w8(32'hba70c1f6),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8858f3),
	.w1(32'h3ad3dc4a),
	.w2(32'h3a135387),
	.w3(32'hbb10a2eb),
	.w4(32'h3a40c544),
	.w5(32'h3a4f4766),
	.w6(32'hba823824),
	.w7(32'h3b126a9f),
	.w8(32'h3aa9dca1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990e440),
	.w1(32'h3b1d4f54),
	.w2(32'h3bb0ac86),
	.w3(32'h3aaa3f0b),
	.w4(32'h3b7838b7),
	.w5(32'h3a70f56f),
	.w6(32'h3a446c6c),
	.w7(32'h3b988de3),
	.w8(32'hba1cab10),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5ee07),
	.w1(32'h39d33e1d),
	.w2(32'h3a3e6301),
	.w3(32'h3ad316f5),
	.w4(32'h3ad2a0f3),
	.w5(32'h3a41d4dd),
	.w6(32'h3abb8db9),
	.w7(32'h3b57c58e),
	.w8(32'h3b0e5c89),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cd6a1),
	.w1(32'hbb0506e8),
	.w2(32'hb9ab08cd),
	.w3(32'hbbacdc80),
	.w4(32'hbb84c9af),
	.w5(32'hb93e5d07),
	.w6(32'hbabe4492),
	.w7(32'hbb2adba6),
	.w8(32'hba962849),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a7c5a),
	.w1(32'h3b5b1b59),
	.w2(32'h3b39fcec),
	.w3(32'hba1f538a),
	.w4(32'h3b5ce840),
	.w5(32'h3b66ede2),
	.w6(32'hbada133e),
	.w7(32'h3b52da79),
	.w8(32'h3b3430a3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14db94),
	.w1(32'h3a9289cb),
	.w2(32'h3ac8267d),
	.w3(32'h3a447f79),
	.w4(32'h3aede66b),
	.w5(32'hbb20d5dd),
	.w6(32'h3b2a03de),
	.w7(32'h3b05d164),
	.w8(32'hbbb309d9),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbc8a4),
	.w1(32'hbba3417e),
	.w2(32'hba9cc2a6),
	.w3(32'hbbd6ec79),
	.w4(32'hbac3b529),
	.w5(32'hba2f0271),
	.w6(32'hbbc6dc67),
	.w7(32'hb87418f8),
	.w8(32'h3adacd53),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82e3bd),
	.w1(32'hbaae2fb5),
	.w2(32'hba388c44),
	.w3(32'hbabffe2f),
	.w4(32'hbab22272),
	.w5(32'h391f7fd6),
	.w6(32'hba1e49e7),
	.w7(32'hb9db38ae),
	.w8(32'hb9a1e717),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89ca5a),
	.w1(32'h3adf6dd7),
	.w2(32'hbb49b1b8),
	.w3(32'hbb0b7057),
	.w4(32'h3a8a14a5),
	.w5(32'hba95ae81),
	.w6(32'hba2e9815),
	.w7(32'h3a1cc38e),
	.w8(32'hbaed3059),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90692eb),
	.w1(32'hb9e7048f),
	.w2(32'hb9c365db),
	.w3(32'hba9806ef),
	.w4(32'hbaad5535),
	.w5(32'hba20b54d),
	.w6(32'hba04fe99),
	.w7(32'hba823dea),
	.w8(32'h392e8c01),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb158b11),
	.w1(32'h3a50fb74),
	.w2(32'hb9a303a6),
	.w3(32'hba2c4c85),
	.w4(32'hb7f63e84),
	.w5(32'hbafc0013),
	.w6(32'hbacc5c82),
	.w7(32'hb8f8188d),
	.w8(32'hb9eaf20c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2506d5),
	.w1(32'hb9715b2b),
	.w2(32'h3a6609c3),
	.w3(32'hbb5a9790),
	.w4(32'hbab6fde0),
	.w5(32'h3b732f8a),
	.w6(32'hb9731ada),
	.w7(32'hbb424962),
	.w8(32'h3aceadbb),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb948b633),
	.w1(32'h3a9b4b79),
	.w2(32'h3a72be87),
	.w3(32'hbb0bc632),
	.w4(32'hbaaa65ed),
	.w5(32'h3a9454f3),
	.w6(32'hba793445),
	.w7(32'hba6f252a),
	.w8(32'h39948b66),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba412539),
	.w1(32'h39e19555),
	.w2(32'h39444846),
	.w3(32'hbaad181f),
	.w4(32'hb97d7a23),
	.w5(32'hba7d960d),
	.w6(32'hba6f57f3),
	.w7(32'hbac00b26),
	.w8(32'hba1720fd),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cc920),
	.w1(32'h3a5d3384),
	.w2(32'h3bbab5ff),
	.w3(32'hbbbe26cf),
	.w4(32'hbb279747),
	.w5(32'h3c10b0f0),
	.w6(32'hba1109aa),
	.w7(32'hbaea2fbc),
	.w8(32'h3ba1dec7),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27b588),
	.w1(32'h393e38e2),
	.w2(32'hbab95862),
	.w3(32'hba35a95a),
	.w4(32'hbaba5c38),
	.w5(32'hbb1cbc48),
	.w6(32'h3b03f1f5),
	.w7(32'hb9789114),
	.w8(32'hbb1c6220),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d2e46),
	.w1(32'h3ad8dce9),
	.w2(32'h3ba6f65e),
	.w3(32'hbb91d929),
	.w4(32'h3b310f1d),
	.w5(32'h3b510894),
	.w6(32'hbb6870d5),
	.w7(32'h3b3d65f6),
	.w8(32'h3b38d6c6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b796306),
	.w1(32'hb9c68835),
	.w2(32'hb9e1e325),
	.w3(32'h3b3526eb),
	.w4(32'hba00fbc3),
	.w5(32'hb601acae),
	.w6(32'h3b2daa9f),
	.w7(32'hb817b950),
	.w8(32'hba60f71d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b738e2),
	.w1(32'hba1267ab),
	.w2(32'hb83299e5),
	.w3(32'hb8ae7a88),
	.w4(32'hba5380b1),
	.w5(32'hba257f0d),
	.w6(32'h3a0b3f78),
	.w7(32'hb9847693),
	.w8(32'hb9a8834f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd17cfd),
	.w1(32'hbb256156),
	.w2(32'hb9f27143),
	.w3(32'hba17c511),
	.w4(32'h3b7d6ea0),
	.w5(32'hb8eb2bf2),
	.w6(32'hbbe4532a),
	.w7(32'h3b718487),
	.w8(32'h3b298917),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98d658),
	.w1(32'h3a33cfd7),
	.w2(32'hba594de7),
	.w3(32'h3a2976e5),
	.w4(32'h3b3b74bd),
	.w5(32'hba326ec5),
	.w6(32'hbb930df7),
	.w7(32'h3ab8528f),
	.w8(32'hbb30cf3f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ef141),
	.w1(32'hbab245a8),
	.w2(32'hba41fcbe),
	.w3(32'hbb77b381),
	.w4(32'hbb2d81f9),
	.w5(32'h3b4c787c),
	.w6(32'hbb0af6e6),
	.w7(32'hbaef2c0f),
	.w8(32'h3a88575e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e86b2),
	.w1(32'hbc083e6c),
	.w2(32'h3b239738),
	.w3(32'hbbb3c3a2),
	.w4(32'h3ba742a1),
	.w5(32'h3c17c2e8),
	.w6(32'h3bc91d1e),
	.w7(32'hbab07a14),
	.w8(32'hbbf82dca),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac02451),
	.w1(32'hb8c8e51e),
	.w2(32'hba826614),
	.w3(32'hba2e8070),
	.w4(32'hba7f1457),
	.w5(32'hbb27c674),
	.w6(32'h38c0f255),
	.w7(32'hbb11bdaa),
	.w8(32'hb9b11dce),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10e625),
	.w1(32'h3a3eb0ca),
	.w2(32'hbad5f24a),
	.w3(32'hb972c69c),
	.w4(32'hb9af7ba3),
	.w5(32'hba4ac4f9),
	.w6(32'h39bbdcb0),
	.w7(32'hb9a3cacd),
	.w8(32'hbae3d6ff),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc833920),
	.w1(32'h3a9e2176),
	.w2(32'h3c73729f),
	.w3(32'hbc13a6ab),
	.w4(32'h3c88346b),
	.w5(32'h3be19e8a),
	.w6(32'hbca22c75),
	.w7(32'h3c6434fa),
	.w8(32'h3c2a8dc7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad4d37),
	.w1(32'hbac282ee),
	.w2(32'hbb020598),
	.w3(32'h3b4b5724),
	.w4(32'hba83be3c),
	.w5(32'hbb3c71b8),
	.w6(32'h3886f56d),
	.w7(32'h3961d477),
	.w8(32'hbbecbd4e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4888fe),
	.w1(32'hba09fc31),
	.w2(32'h3bced059),
	.w3(32'hbbd52af2),
	.w4(32'h3c1f1970),
	.w5(32'h3bb94fcb),
	.w6(32'hbc174559),
	.w7(32'h3c197efa),
	.w8(32'h3b618b5e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcdcf6),
	.w1(32'h3b0f84e1),
	.w2(32'h3aea299f),
	.w3(32'h3b338fe8),
	.w4(32'hb85b4cd3),
	.w5(32'h38f475a1),
	.w6(32'h3ad83417),
	.w7(32'h3a995bc6),
	.w8(32'h3a17e5c9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3384c),
	.w1(32'h3aa4f4fd),
	.w2(32'h39b40b92),
	.w3(32'hbaf8561f),
	.w4(32'hba81370b),
	.w5(32'h3b2f210e),
	.w6(32'h3a34698f),
	.w7(32'hbb675fc9),
	.w8(32'hba3f9332),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44fbc3),
	.w1(32'hb80d435f),
	.w2(32'hb994c323),
	.w3(32'hb9915bf1),
	.w4(32'h39164330),
	.w5(32'h3a1f4b23),
	.w6(32'hba86d260),
	.w7(32'h3ab00850),
	.w8(32'h3a9473b6),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b3dc5),
	.w1(32'hb995266a),
	.w2(32'hbab2d94e),
	.w3(32'h3a9fa426),
	.w4(32'hbaa5c9f6),
	.w5(32'hb99c6ea2),
	.w6(32'h3949dc2a),
	.w7(32'hb89e6a4d),
	.w8(32'hba95664d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba131db7),
	.w1(32'hb989c714),
	.w2(32'hbaba6ba8),
	.w3(32'hbb270c3a),
	.w4(32'hbb5fe715),
	.w5(32'hbb00c977),
	.w6(32'hbaf66f70),
	.w7(32'hbb080047),
	.w8(32'hba65f29d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990146f),
	.w1(32'hbace902f),
	.w2(32'hb95cffc2),
	.w3(32'hb78b3907),
	.w4(32'hbaf73aa5),
	.w5(32'hb8e86472),
	.w6(32'h3a1bb00e),
	.w7(32'hba23046f),
	.w8(32'h39db340e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac61ee1),
	.w1(32'h3aeef018),
	.w2(32'hb9c1acde),
	.w3(32'h3a8b155f),
	.w4(32'h3aac9e9a),
	.w5(32'hbac97548),
	.w6(32'hba0068bd),
	.w7(32'h3aee5cce),
	.w8(32'hba9356a0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369efe41),
	.w1(32'h3b3d8bc7),
	.w2(32'h3b448392),
	.w3(32'h3af7c4b4),
	.w4(32'h3b22ee0f),
	.w5(32'h393fa048),
	.w6(32'hbb3424c1),
	.w7(32'h3add33b6),
	.w8(32'h3ad4a4a6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8d8f4),
	.w1(32'h3941869c),
	.w2(32'h39d3207a),
	.w3(32'hba9c360b),
	.w4(32'hbaa83850),
	.w5(32'hba27d290),
	.w6(32'hbad2830b),
	.w7(32'hb74ddc41),
	.w8(32'h3a8b0dc7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a04c6b),
	.w1(32'hba8b0ce8),
	.w2(32'hbac9aabd),
	.w3(32'hbad47b18),
	.w4(32'hba32a985),
	.w5(32'h37f9a0d0),
	.w6(32'hba54c408),
	.w7(32'hb91c18ee),
	.w8(32'h3922127a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49b1cc),
	.w1(32'hbb85c43f),
	.w2(32'h3be52b26),
	.w3(32'hbc129ac4),
	.w4(32'h3c116c8b),
	.w5(32'hb989ac83),
	.w6(32'hbc84a4f8),
	.w7(32'h3c6a0464),
	.w8(32'hbb0f7f5b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c061c),
	.w1(32'hb69fdc1a),
	.w2(32'h3adc9155),
	.w3(32'hbad2018e),
	.w4(32'h3a5406f9),
	.w5(32'h399cfa4a),
	.w6(32'hba67b61c),
	.w7(32'h3b29ef6b),
	.w8(32'hba83a1ae),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8a412),
	.w1(32'h3a473b0e),
	.w2(32'h3ac3531c),
	.w3(32'hbac05e19),
	.w4(32'h39dc0059),
	.w5(32'h3a1deffc),
	.w6(32'h38abda4d),
	.w7(32'hb7e68598),
	.w8(32'h3a4a63fc),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedc661),
	.w1(32'hb91fa515),
	.w2(32'h3a10aef6),
	.w3(32'h3a850e9c),
	.w4(32'h37946016),
	.w5(32'h38e515f0),
	.w6(32'h3a7c4f01),
	.w7(32'h3a4c71f8),
	.w8(32'hbae58c75),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ba91f),
	.w1(32'h3944f4d0),
	.w2(32'hb89edc7d),
	.w3(32'h3a4d6930),
	.w4(32'h3a24e20b),
	.w5(32'h3761fd51),
	.w6(32'h3a52799b),
	.w7(32'h3a14f609),
	.w8(32'h38af26ca),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991a313),
	.w1(32'h38cf86b3),
	.w2(32'h3983292f),
	.w3(32'hb999e6b2),
	.w4(32'h3a86c106),
	.w5(32'hb9f3df53),
	.w6(32'h37be5319),
	.w7(32'h3aa3dd57),
	.w8(32'h393ab80d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915944f),
	.w1(32'hb9a7e830),
	.w2(32'hb9b27785),
	.w3(32'h3a693e4d),
	.w4(32'h38f65881),
	.w5(32'hba563dc9),
	.w6(32'hba2cc955),
	.w7(32'hb910e4de),
	.w8(32'h39dedd40),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e43b62),
	.w1(32'hba44d2d7),
	.w2(32'hba083d7d),
	.w3(32'h3a0ad561),
	.w4(32'hba46658c),
	.w5(32'hba98a2aa),
	.w6(32'h3aa24d93),
	.w7(32'hbab56709),
	.w8(32'hbab2ddec),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9921a2d),
	.w1(32'h3adfc318),
	.w2(32'h3b1957a9),
	.w3(32'hba8a596c),
	.w4(32'hb9a1edfc),
	.w5(32'h3b29b87c),
	.w6(32'hbac0063c),
	.w7(32'hba596037),
	.w8(32'h3a98b17c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc802a9),
	.w1(32'h3b1fb313),
	.w2(32'hba422b6e),
	.w3(32'h39cff7db),
	.w4(32'hbaa8118b),
	.w5(32'h3b73cc14),
	.w6(32'h3bd056db),
	.w7(32'hbbb0721f),
	.w8(32'hbbced112),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1777e0),
	.w1(32'hbb260701),
	.w2(32'hbb2fb0cc),
	.w3(32'h3a85abf4),
	.w4(32'hbb35db99),
	.w5(32'hbb135380),
	.w6(32'h3af554e4),
	.w7(32'h3affbfc2),
	.w8(32'hbb3af021),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d5589),
	.w1(32'hbb734967),
	.w2(32'hbaa07502),
	.w3(32'hbae6cb29),
	.w4(32'hbb25dc17),
	.w5(32'hbaa952b0),
	.w6(32'h3b6112e0),
	.w7(32'hbac65e62),
	.w8(32'hbb9f340c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a328158),
	.w1(32'h3a9e453a),
	.w2(32'h3b1e6f02),
	.w3(32'h3a37bd26),
	.w4(32'h3afaf0f2),
	.w5(32'h3b61c51c),
	.w6(32'h39891fd9),
	.w7(32'h3b172cac),
	.w8(32'h3b50727a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c4575),
	.w1(32'h3a470031),
	.w2(32'h36a4ec4b),
	.w3(32'h3abf1907),
	.w4(32'h37e63237),
	.w5(32'h387d4990),
	.w6(32'h3abe3ff3),
	.w7(32'h3a7373ec),
	.w8(32'hb9bea85c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a117227),
	.w1(32'hba9f34e6),
	.w2(32'hb9d6e1ba),
	.w3(32'h38a85969),
	.w4(32'hb9b92018),
	.w5(32'h3afe9c15),
	.w6(32'h3a0ccc20),
	.w7(32'hba8ab540),
	.w8(32'h3a1b021c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87f7358),
	.w1(32'h3a372849),
	.w2(32'h3a2ad07b),
	.w3(32'h3887e099),
	.w4(32'hb9c3059d),
	.w5(32'hba6ed7e7),
	.w6(32'h37611dc2),
	.w7(32'hba78894a),
	.w8(32'hbb321f0b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89361a),
	.w1(32'h38777406),
	.w2(32'hbab53499),
	.w3(32'h3b367ab9),
	.w4(32'hbb977436),
	.w5(32'hbb48b9dc),
	.w6(32'h3b897866),
	.w7(32'hbad5f06a),
	.w8(32'hbb800bf1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a85f5),
	.w1(32'hbacfad71),
	.w2(32'hbb3821cc),
	.w3(32'hba7d709b),
	.w4(32'hbb054e53),
	.w5(32'hbafdce52),
	.w6(32'hb9a72585),
	.w7(32'hbad32a3c),
	.w8(32'hbad0c7e6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92870e),
	.w1(32'h3aa362cd),
	.w2(32'h388fc13d),
	.w3(32'h3aaf475f),
	.w4(32'h3a9b2fbd),
	.w5(32'h3a18d248),
	.w6(32'h3a925c12),
	.w7(32'h3a9fd3f5),
	.w8(32'h389cb0af),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d0dca),
	.w1(32'hbaa47aea),
	.w2(32'hbaf07075),
	.w3(32'hbb95d700),
	.w4(32'hba9e9416),
	.w5(32'hbb0923b5),
	.w6(32'hbadb2401),
	.w7(32'hbac5fef8),
	.w8(32'h3ad9e509),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c63370),
	.w1(32'hbaaa4fd5),
	.w2(32'hbafad728),
	.w3(32'hb902316c),
	.w4(32'hbaa9470e),
	.w5(32'hb98a0484),
	.w6(32'h39fbc0ca),
	.w7(32'hba648152),
	.w8(32'hba254973),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ad6ce),
	.w1(32'hb995ea8c),
	.w2(32'h3a3da0b1),
	.w3(32'hba1c2ecc),
	.w4(32'h3a4e30ae),
	.w5(32'h3b083e20),
	.w6(32'h3a43f8f3),
	.w7(32'h3aab8155),
	.w8(32'h3aa2c869),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeddd99),
	.w1(32'hbad032e6),
	.w2(32'hbab6e0be),
	.w3(32'h3b262324),
	.w4(32'hbab84f15),
	.w5(32'hbb291a96),
	.w6(32'h3b1269f2),
	.w7(32'hbac599cd),
	.w8(32'hbb334325),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4788dc),
	.w1(32'hbb93c3f8),
	.w2(32'hbbbad008),
	.w3(32'hbb6510e2),
	.w4(32'hbc2d157f),
	.w5(32'h3b4f88b7),
	.w6(32'h3b15ea67),
	.w7(32'hbc7be13f),
	.w8(32'hbc144997),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aa4908),
	.w1(32'hbaca7448),
	.w2(32'hbb4679eb),
	.w3(32'hb8e2dd71),
	.w4(32'hbb72018e),
	.w5(32'hbb884a14),
	.w6(32'hb908ca3a),
	.w7(32'hbb2dac07),
	.w8(32'hbb7f5546),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0659c3),
	.w1(32'hbae24896),
	.w2(32'hbadcaa4c),
	.w3(32'hbc0e9571),
	.w4(32'hb97086b5),
	.w5(32'h3a970865),
	.w6(32'hbbda3837),
	.w7(32'h3a95785b),
	.w8(32'h3b8e7b67),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule