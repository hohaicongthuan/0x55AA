module layer_10_featuremap_198(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373f81ac),
	.w1(32'h35a9ab5a),
	.w2(32'hb62311f0),
	.w3(32'h37d220cb),
	.w4(32'h37ab61a2),
	.w5(32'h372da79e),
	.w6(32'h38761a58),
	.w7(32'h37ff58c3),
	.w8(32'h37dacf9a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a723972),
	.w1(32'h3b1d3c93),
	.w2(32'h3b4868b8),
	.w3(32'h3af784a5),
	.w4(32'h3b0831ce),
	.w5(32'h398a693f),
	.w6(32'h3b191693),
	.w7(32'h399a831e),
	.w8(32'hba067e71),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371bf5d6),
	.w1(32'h3696c15a),
	.w2(32'h373fa29c),
	.w3(32'h3714d8ae),
	.w4(32'h36b0d408),
	.w5(32'h370ae23e),
	.w6(32'h37866707),
	.w7(32'h3787583d),
	.w8(32'h3790e86c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364e13aa),
	.w1(32'h3a32d2ff),
	.w2(32'hb99f5b16),
	.w3(32'h379357e6),
	.w4(32'h399719f8),
	.w5(32'h38f40a5a),
	.w6(32'h39219201),
	.w7(32'h3a074a79),
	.w8(32'h39975ecb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0299d3),
	.w1(32'h3a00ffdc),
	.w2(32'hb6528f16),
	.w3(32'h3a2ac56a),
	.w4(32'h3a18d4d9),
	.w5(32'h391c153a),
	.w6(32'h3a2c2bdd),
	.w7(32'h3a29aef2),
	.w8(32'h39aeaa76),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8165642),
	.w1(32'hb85efce0),
	.w2(32'hb73c0314),
	.w3(32'h36e005b5),
	.w4(32'hb79031f2),
	.w5(32'hb6c9094a),
	.w6(32'h378a65c5),
	.w7(32'h3738c6d5),
	.w8(32'h37fa02ec),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54e70b),
	.w1(32'h3b00565d),
	.w2(32'h39ebf99a),
	.w3(32'h3b169881),
	.w4(32'h3ad7fd5b),
	.w5(32'hb9c3cfc3),
	.w6(32'h3aab7f1e),
	.w7(32'hb9f0ee30),
	.w8(32'hbb682e0e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab790b),
	.w1(32'hbb8bd22b),
	.w2(32'hbbe0e353),
	.w3(32'hbc3255b6),
	.w4(32'hbc061c07),
	.w5(32'hbb67e25a),
	.w6(32'hbbfad9e2),
	.w7(32'hbbd15331),
	.w8(32'hbb34b56a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba052cb8),
	.w1(32'hba817d31),
	.w2(32'hbab0bbef),
	.w3(32'hba261849),
	.w4(32'hba491c93),
	.w5(32'hba738c6b),
	.w6(32'hb98bcd1d),
	.w7(32'hba2cfe9f),
	.w8(32'hbaabe12d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0634fa),
	.w1(32'hba01cb44),
	.w2(32'hb9aad935),
	.w3(32'hbb2b6b57),
	.w4(32'hba5c6c8f),
	.w5(32'hbac43cac),
	.w6(32'hbad92e8b),
	.w7(32'hbb17da82),
	.w8(32'hbb81d769),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ffd8f6),
	.w1(32'hb6873c72),
	.w2(32'hba42479b),
	.w3(32'hb9230dfd),
	.w4(32'hb8044f80),
	.w5(32'hba896080),
	.w6(32'h39dffbb8),
	.w7(32'h39ef3e94),
	.w8(32'hba162755),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f7af6),
	.w1(32'h3b53a8de),
	.w2(32'hba56daa1),
	.w3(32'h3b3493d7),
	.w4(32'h3b938bb1),
	.w5(32'h3b1fef30),
	.w6(32'h3ae243a5),
	.w7(32'h3b83ae6f),
	.w8(32'h3a1a7089),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec6194),
	.w1(32'h398b3fb4),
	.w2(32'hb82f7d6f),
	.w3(32'hbb2f91e6),
	.w4(32'hbaf9c20d),
	.w5(32'hba957413),
	.w6(32'hb9d11ab1),
	.w7(32'hbac89e81),
	.w8(32'hbb0f31c7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03d934),
	.w1(32'h3aaf1cda),
	.w2(32'h392c5d2c),
	.w3(32'h39d7f179),
	.w4(32'hb86505f9),
	.w5(32'hb91b2232),
	.w6(32'h39c7b143),
	.w7(32'hb9ad4d06),
	.w8(32'hba116d0d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2198dd),
	.w1(32'h3a165394),
	.w2(32'h39d4ea83),
	.w3(32'h3a44f8b7),
	.w4(32'h3aab284d),
	.w5(32'h3a95ed0a),
	.w6(32'h3af6ff17),
	.w7(32'h3b098dc7),
	.w8(32'h3a9885ec),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886e9e4),
	.w1(32'h3a16f7f3),
	.w2(32'h390a966a),
	.w3(32'hbae282fb),
	.w4(32'hba62c906),
	.w5(32'hb9f10f98),
	.w6(32'hbb877806),
	.w7(32'hbbc377e2),
	.w8(32'hbb108ed5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b71b80),
	.w1(32'h39092dd9),
	.w2(32'h394763d7),
	.w3(32'hb921c62f),
	.w4(32'h3792115d),
	.w5(32'h38fedd78),
	.w6(32'hb8e68883),
	.w7(32'h391b1947),
	.w8(32'h39b292f2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76db49),
	.w1(32'hbc255e85),
	.w2(32'hbc51bb06),
	.w3(32'hbc2d1013),
	.w4(32'hbc194690),
	.w5(32'hbbf9bfd2),
	.w6(32'hbc140c18),
	.w7(32'hbc2767c9),
	.w8(32'hbbd3bdd0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba08e1),
	.w1(32'hbb479ced),
	.w2(32'hbb857e0c),
	.w3(32'hbb9826c7),
	.w4(32'hbb8b4711),
	.w5(32'hbb2986c9),
	.w6(32'hbb856cf8),
	.w7(32'hbb905028),
	.w8(32'hbb346fff),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb739b6d1),
	.w1(32'h3711c892),
	.w2(32'h37db3355),
	.w3(32'h37be66b7),
	.w4(32'h37b88cf1),
	.w5(32'h37ba39f7),
	.w6(32'h37e7f97d),
	.w7(32'h378cda30),
	.w8(32'hb780e3bd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5ae5e89),
	.w1(32'hb8b5e385),
	.w2(32'h36afc9b7),
	.w3(32'hb7444d20),
	.w4(32'hb90ed589),
	.w5(32'hb83503a7),
	.w6(32'hb6b6214f),
	.w7(32'hb839d2e1),
	.w8(32'h38c6f77f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a806120),
	.w1(32'h3aa22f25),
	.w2(32'h3a14067f),
	.w3(32'h3ad5fd71),
	.w4(32'h3aee0628),
	.w5(32'h3a150459),
	.w6(32'h3ae1b473),
	.w7(32'h3ada0dad),
	.w8(32'h3a51e1d5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987f218),
	.w1(32'hbc0b0b64),
	.w2(32'hbc99719d),
	.w3(32'hbc17b4f7),
	.w4(32'hbba26e78),
	.w5(32'hbc321801),
	.w6(32'hbc6bbf56),
	.w7(32'hbbb7d1e6),
	.w8(32'hbc451cf7),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28fdc4),
	.w1(32'h3a72db5d),
	.w2(32'h3b2db666),
	.w3(32'h3a578e62),
	.w4(32'h3ab199b2),
	.w5(32'h3a83ca3e),
	.w6(32'h3aa3c613),
	.w7(32'h3a04d175),
	.w8(32'hba3608c7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb144787),
	.w1(32'h3ade2ee9),
	.w2(32'h3b5e6dcd),
	.w3(32'h3a6418ae),
	.w4(32'h3b7dc3c3),
	.w5(32'h3b29de21),
	.w6(32'h3b025b4e),
	.w7(32'h3a7165e0),
	.w8(32'h39c94e7c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a5c2e),
	.w1(32'h3a2dabff),
	.w2(32'h39eae555),
	.w3(32'hb77bf7cd),
	.w4(32'h3975baea),
	.w5(32'h3988806c),
	.w6(32'hb9490d8b),
	.w7(32'h399f0c1b),
	.w8(32'h396e31fd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3803b757),
	.w1(32'hb3b0d753),
	.w2(32'h39039d9e),
	.w3(32'h3893bcbe),
	.w4(32'h3863d5f3),
	.w5(32'h3923d054),
	.w6(32'h392603a8),
	.w7(32'h38eddd4c),
	.w8(32'h398aad82),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95ad00),
	.w1(32'h3b330be6),
	.w2(32'h3b100f72),
	.w3(32'h3afc1231),
	.w4(32'h3b97d980),
	.w5(32'h3af85844),
	.w6(32'h3b79c45f),
	.w7(32'h3af493d1),
	.w8(32'h39e6a5af),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a533d93),
	.w1(32'h3a48fce0),
	.w2(32'h3a7a0cca),
	.w3(32'h3abe32ba),
	.w4(32'h3ad99bf8),
	.w5(32'h3ad65c70),
	.w6(32'h3b1e3e94),
	.w7(32'h3b28cda9),
	.w8(32'h3b2a888f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed1f17),
	.w1(32'h3b60386c),
	.w2(32'h3b6a39b0),
	.w3(32'h3aeb3987),
	.w4(32'h3b2c3a8e),
	.w5(32'h3abb0b94),
	.w6(32'h3b864fc8),
	.w7(32'h3ae96795),
	.w8(32'hb9ee5493),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3829ec26),
	.w1(32'h3841d710),
	.w2(32'h38d26c58),
	.w3(32'h388ad1da),
	.w4(32'h38a2bb5d),
	.w5(32'h38f8ae90),
	.w6(32'h38c7a3cf),
	.w7(32'h390a19ef),
	.w8(32'h392d71f5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82aa788),
	.w1(32'h39611969),
	.w2(32'h39941fea),
	.w3(32'h37cf66a3),
	.w4(32'h39cb6be4),
	.w5(32'h39c8548a),
	.w6(32'h39626caf),
	.w7(32'h3a0dda35),
	.w8(32'h39e11cc4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa04c2d),
	.w1(32'h3a5f94b3),
	.w2(32'h3a0167e3),
	.w3(32'h3a08ce9c),
	.w4(32'h3a406f6b),
	.w5(32'h3a444c17),
	.w6(32'h39f2c7bc),
	.w7(32'h3a083843),
	.w8(32'hb9847fd9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa47028),
	.w1(32'h39141433),
	.w2(32'h3a7cd848),
	.w3(32'hba6352d9),
	.w4(32'hba0ba4d2),
	.w5(32'h38f00572),
	.w6(32'hba48f9b0),
	.w7(32'hba98adef),
	.w8(32'hba7b8961),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c1448c),
	.w1(32'hb905d38d),
	.w2(32'h38c33f0c),
	.w3(32'hb91f21f5),
	.w4(32'h37216d25),
	.w5(32'h39680906),
	.w6(32'h3935d95e),
	.w7(32'hb9deedaa),
	.w8(32'hb9966316),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ab45a),
	.w1(32'h3aacbc8c),
	.w2(32'h3a0fa711),
	.w3(32'hba8bcefd),
	.w4(32'h388ae131),
	.w5(32'h38dba73b),
	.w6(32'h38fa5430),
	.w7(32'h3a8f56f5),
	.w8(32'hb9af0df3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a08a0f),
	.w1(32'h3b8f27ab),
	.w2(32'hbb9413f6),
	.w3(32'hb9535764),
	.w4(32'h3abe85b4),
	.w5(32'h3a93daa5),
	.w6(32'hbb3a21da),
	.w7(32'h3b141edd),
	.w8(32'hba7b6133),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb554373),
	.w1(32'h3bb751f3),
	.w2(32'h3bcc6c66),
	.w3(32'h3b943b65),
	.w4(32'h3c3abf7b),
	.w5(32'h3ba4bdb7),
	.w6(32'h3bdf787a),
	.w7(32'h3c07aa06),
	.w8(32'h3b8b3565),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab216c3),
	.w1(32'h3bdb16fb),
	.w2(32'h3b7acb4b),
	.w3(32'h3bfa0010),
	.w4(32'h3c16d083),
	.w5(32'h3a80f4a3),
	.w6(32'h3c1fd4fb),
	.w7(32'h3b9762c8),
	.w8(32'hb95b3122),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d97e89),
	.w1(32'h3ab64743),
	.w2(32'h3a450a2c),
	.w3(32'h3a8cda7a),
	.w4(32'h3aab175e),
	.w5(32'h39f5c9fa),
	.w6(32'h3aa55dc3),
	.w7(32'h3a72d1d6),
	.w8(32'h39c84062),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de0c00),
	.w1(32'hb99518a8),
	.w2(32'hba0117cd),
	.w3(32'hb9b4bc01),
	.w4(32'hb9a836c7),
	.w5(32'hba0d6f71),
	.w6(32'hb99d667e),
	.w7(32'hb9058840),
	.w8(32'hb9e7317c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3916a490),
	.w1(32'h386cd545),
	.w2(32'h3945db8b),
	.w3(32'h3942bee9),
	.w4(32'h38f330a1),
	.w5(32'h3930179b),
	.w6(32'h3952a6f6),
	.w7(32'hb78b9468),
	.w8(32'h395f53a6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b8c51),
	.w1(32'h3a799528),
	.w2(32'h3ad2bcbd),
	.w3(32'h39d823e9),
	.w4(32'h3aca5a11),
	.w5(32'h3a8527c0),
	.w6(32'hb9a26f31),
	.w7(32'h3a267b7e),
	.w8(32'h374aa00f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956ef1d),
	.w1(32'hba04bcc0),
	.w2(32'hbae0c93f),
	.w3(32'hbbb85f65),
	.w4(32'hbb4fa287),
	.w5(32'hbb2e55ee),
	.w6(32'hbb9a28e2),
	.w7(32'hbba06b75),
	.w8(32'hbb2d3fa3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0524da),
	.w1(32'h3a0e1ee5),
	.w2(32'h3a83e75f),
	.w3(32'hb9ac0b33),
	.w4(32'h3abf2ef1),
	.w5(32'h35350d18),
	.w6(32'h3aa51cb9),
	.w7(32'h3a93e80e),
	.w8(32'hba04b12a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb125da8),
	.w1(32'h39160327),
	.w2(32'h3b00726c),
	.w3(32'hba8e6b74),
	.w4(32'hba16077b),
	.w5(32'hba8e7c1b),
	.w6(32'hba10fc65),
	.w7(32'hba5367a2),
	.w8(32'hbad927f5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb355b5e),
	.w1(32'hbac45adc),
	.w2(32'hbb058c44),
	.w3(32'hbb25f95d),
	.w4(32'hbb0e1625),
	.w5(32'hbaf985cb),
	.w6(32'hbba0840a),
	.w7(32'hbb7c4d0c),
	.w8(32'hbb48299e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c04c6),
	.w1(32'hbbf5539e),
	.w2(32'hbc74e899),
	.w3(32'hbc3fb1b5),
	.w4(32'hbc3c7faf),
	.w5(32'hbc0f32cd),
	.w6(32'hbc4e77f1),
	.w7(32'hbc35071e),
	.w8(32'hbbf4f39e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ed318),
	.w1(32'hb8bf0620),
	.w2(32'hba523c22),
	.w3(32'h394fa2d2),
	.w4(32'hb8bbe928),
	.w5(32'hb9e1e81c),
	.w6(32'hb7929409),
	.w7(32'hb98ba547),
	.w8(32'hb9b615ab),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e76eb8),
	.w1(32'hbaa42123),
	.w2(32'hbb042831),
	.w3(32'hbad0bf98),
	.w4(32'hbb0ca70e),
	.w5(32'hbb0f9f54),
	.w6(32'hbb1192e2),
	.w7(32'hbb408b8f),
	.w8(32'hbb42e9db),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa43368),
	.w1(32'h39c0bdf9),
	.w2(32'hb9ccfadc),
	.w3(32'h3a83654d),
	.w4(32'h399704a0),
	.w5(32'hb926b0cd),
	.w6(32'h3a5d92d5),
	.w7(32'h396ca71a),
	.w8(32'hb9165b5f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3134c),
	.w1(32'hb9e36494),
	.w2(32'hbac91519),
	.w3(32'hbaf790e9),
	.w4(32'hb8835f8f),
	.w5(32'hba9f9b78),
	.w6(32'hba5df1b8),
	.w7(32'hb9eb6ea0),
	.w8(32'hbb223479),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22e251),
	.w1(32'hba95ca84),
	.w2(32'hbabd7be2),
	.w3(32'hba5635d4),
	.w4(32'hba972df6),
	.w5(32'hba8b9788),
	.w6(32'hbab61720),
	.w7(32'hba9779e3),
	.w8(32'hba88777f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2589cc),
	.w1(32'hbbdf7ade),
	.w2(32'hbc1180d9),
	.w3(32'hbc05288b),
	.w4(32'hbbdf5ea8),
	.w5(32'hbb1ab28c),
	.w6(32'hbbaeae19),
	.w7(32'hbbcda8ea),
	.w8(32'hbb49237c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51f868),
	.w1(32'hba3cfb6a),
	.w2(32'hbaaa9099),
	.w3(32'hba2aba51),
	.w4(32'hb959e032),
	.w5(32'hba43ad43),
	.w6(32'hb9771ad6),
	.w7(32'hb98194ca),
	.w8(32'hb96307d4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921b343),
	.w1(32'h38a91bf1),
	.w2(32'hb4c92c51),
	.w3(32'h391f5853),
	.w4(32'h3879b2b8),
	.w5(32'hb7ec36a6),
	.w6(32'h379dac3e),
	.w7(32'hb6203ce1),
	.w8(32'hb8531865),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6518eda),
	.w1(32'hb739f83d),
	.w2(32'h37196a22),
	.w3(32'h37c1d168),
	.w4(32'h369b2870),
	.w5(32'h3765203c),
	.w6(32'h38279867),
	.w7(32'h37e525fb),
	.w8(32'h38077e0e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385253d6),
	.w1(32'hb930ca52),
	.w2(32'hb81a1b41),
	.w3(32'h3956014a),
	.w4(32'h385dc7aa),
	.w5(32'hb8579216),
	.w6(32'h39a18c16),
	.w7(32'h38911338),
	.w8(32'h38422f69),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2309c0),
	.w1(32'h3a761ce6),
	.w2(32'h3a147d6d),
	.w3(32'h3a699cf7),
	.w4(32'h3a84342a),
	.w5(32'h39970041),
	.w6(32'h39f84466),
	.w7(32'h3a4e77b3),
	.w8(32'h3836ead9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954a2e7),
	.w1(32'h38b0e317),
	.w2(32'h393d3f1b),
	.w3(32'h39959ef2),
	.w4(32'h38165ea2),
	.w5(32'hb6ae2530),
	.w6(32'h3a5e0de6),
	.w7(32'h39856134),
	.w8(32'hb905c20e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86d910),
	.w1(32'hbb068972),
	.w2(32'hbb535843),
	.w3(32'hbb6cadf4),
	.w4(32'hbb123a9f),
	.w5(32'hbaeb7c9f),
	.w6(32'hbb2cfd70),
	.w7(32'hbafd29b8),
	.w8(32'hbabffca5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e0c8b),
	.w1(32'hbb320171),
	.w2(32'hbb402329),
	.w3(32'hbbcb7165),
	.w4(32'hbaf227b9),
	.w5(32'hbb490708),
	.w6(32'hbb907628),
	.w7(32'hbb3fe4c8),
	.w8(32'hbb552454),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8275d58),
	.w1(32'hb7736fc4),
	.w2(32'h3627f4cf),
	.w3(32'hb7ee7f12),
	.w4(32'h381b5548),
	.w5(32'h3898a3d6),
	.w6(32'hb7e1f288),
	.w7(32'h374e7129),
	.w8(32'h38b6fd60),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36074a16),
	.w1(32'hb736676c),
	.w2(32'h37b5225e),
	.w3(32'hb72664d4),
	.w4(32'hb7909f75),
	.w5(32'h37986f4e),
	.w6(32'h34cbdf45),
	.w7(32'hb6833816),
	.w8(32'h37fe3e1d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce031e),
	.w1(32'h39296866),
	.w2(32'h3980a5d8),
	.w3(32'h394e4510),
	.w4(32'h39480234),
	.w5(32'h3929d1ea),
	.w6(32'h39928d83),
	.w7(32'h3953c73f),
	.w8(32'h399c4a5c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e1b82e),
	.w1(32'hb7931165),
	.w2(32'h387fbc42),
	.w3(32'h383145c2),
	.w4(32'h37ee87d9),
	.w5(32'h389f67b5),
	.w6(32'h38a7e188),
	.w7(32'h3893b717),
	.w8(32'h390f172c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b061694),
	.w1(32'hba2bd02a),
	.w2(32'hbad01b79),
	.w3(32'h39c17d3d),
	.w4(32'h3a80c1de),
	.w5(32'h3b1e9629),
	.w6(32'hbaabc33a),
	.w7(32'hbb75fe3e),
	.w8(32'hbad9fc19),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb184164),
	.w1(32'h38b4334a),
	.w2(32'h3a849373),
	.w3(32'h3a8f318c),
	.w4(32'hba25469a),
	.w5(32'hbb260beb),
	.w6(32'hba628e52),
	.w7(32'hba909755),
	.w8(32'hbb867e65),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb543684),
	.w1(32'hbba17078),
	.w2(32'hbbcef759),
	.w3(32'hbb68ea8c),
	.w4(32'hbaaa5d33),
	.w5(32'hbb885177),
	.w6(32'hbb76ccf9),
	.w7(32'hbb5f86c9),
	.w8(32'hbb8b050c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb426b48),
	.w1(32'h3b3ded7d),
	.w2(32'h3bb145d8),
	.w3(32'h3b5c0984),
	.w4(32'h3bcb2984),
	.w5(32'h3b2d7713),
	.w6(32'h3bb0bf3f),
	.w7(32'h3b5398bd),
	.w8(32'h3a1e2471),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dc555f),
	.w1(32'hb704db02),
	.w2(32'h37d307dd),
	.w3(32'h37093e43),
	.w4(32'hb7d069db),
	.w5(32'h3786b3ee),
	.w6(32'h37680756),
	.w7(32'hb6d988df),
	.w8(32'h38248c10),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c427d3),
	.w1(32'h36ab0886),
	.w2(32'h38e7256a),
	.w3(32'h372a6617),
	.w4(32'hb6035e34),
	.w5(32'h38c54b30),
	.w6(32'h384109a9),
	.w7(32'h37f1374d),
	.w8(32'h39040320),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3605e2bf),
	.w1(32'hb8735d3e),
	.w2(32'h38a0a04d),
	.w3(32'hb798be7f),
	.w4(32'hb8356ae6),
	.w5(32'h381354ce),
	.w6(32'h381d7f7b),
	.w7(32'hb83ca715),
	.w8(32'h37ed389d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08c243),
	.w1(32'hba85cfb7),
	.w2(32'hbafb9f46),
	.w3(32'hba822436),
	.w4(32'hba8a5501),
	.w5(32'hba4dcf7a),
	.w6(32'hbad7dfec),
	.w7(32'hbb180c7f),
	.w8(32'hbad09533),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3888a28d),
	.w1(32'hb5f63901),
	.w2(32'h379b02f2),
	.w3(32'h38a00c62),
	.w4(32'hb801d0e9),
	.w5(32'hb65db1e9),
	.w6(32'h38cb5bd0),
	.w7(32'hb81972c8),
	.w8(32'h389a3bcc),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1cbee),
	.w1(32'hbb9ee938),
	.w2(32'hbbe0db90),
	.w3(32'hbb5b8e8d),
	.w4(32'hbb960f2e),
	.w5(32'hbaef65a7),
	.w6(32'hbb9d0290),
	.w7(32'hbb812403),
	.w8(32'hba5ec785),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2f211),
	.w1(32'hbb83c0bb),
	.w2(32'hbbf02117),
	.w3(32'hbbb93a7f),
	.w4(32'hbc0fe656),
	.w5(32'hbb897617),
	.w6(32'hbc108b65),
	.w7(32'hbbf5c63f),
	.w8(32'hbb483b06),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb410f87),
	.w1(32'h3aba4f76),
	.w2(32'h3af5b9d5),
	.w3(32'hbaa864e7),
	.w4(32'h39d9a384),
	.w5(32'hba9fa573),
	.w6(32'h3a48523f),
	.w7(32'h38e72794),
	.w8(32'hba83911d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c8b98),
	.w1(32'hbaa64c4e),
	.w2(32'hbb0089a5),
	.w3(32'hbac4b62e),
	.w4(32'hba7564be),
	.w5(32'hba8b87ca),
	.w6(32'hbaa3f704),
	.w7(32'hbb1406de),
	.w8(32'hbafa71ee),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f788d2),
	.w1(32'hba8b87fb),
	.w2(32'hba1373da),
	.w3(32'h3a1409cf),
	.w4(32'h3a07ec1e),
	.w5(32'h3a887ba5),
	.w6(32'h380467fd),
	.w7(32'hbacf6940),
	.w8(32'hbad45440),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80d762),
	.w1(32'hba17f7de),
	.w2(32'hb9c13754),
	.w3(32'hb8f111fc),
	.w4(32'h3a63887f),
	.w5(32'h38f5e149),
	.w6(32'hb88c5b65),
	.w7(32'hb9f6ddd4),
	.w8(32'hba00b84a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f438d),
	.w1(32'hbb25456a),
	.w2(32'hbba58f3f),
	.w3(32'hbb45070a),
	.w4(32'hbb419692),
	.w5(32'hbb2848dd),
	.w6(32'hbb845961),
	.w7(32'hbb81f43d),
	.w8(32'hbb3bf87b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80c0b4b),
	.w1(32'hb7252b26),
	.w2(32'h37fcd394),
	.w3(32'hb801a2c0),
	.w4(32'h37168a1a),
	.w5(32'h383df695),
	.w6(32'hb4e0f637),
	.w7(32'h3810244a),
	.w8(32'h3874b9c9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3803c690),
	.w1(32'h38254072),
	.w2(32'h38875056),
	.w3(32'h37ee2f17),
	.w4(32'h38048239),
	.w5(32'h383a02f2),
	.w6(32'h37093c37),
	.w7(32'hb6f0cf38),
	.w8(32'h38185053),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b3d860),
	.w1(32'h38c77bac),
	.w2(32'h39c2b7e4),
	.w3(32'h392d642a),
	.w4(32'h396ca1d5),
	.w5(32'h396dd1ab),
	.w6(32'h39b1876c),
	.w7(32'h394d4323),
	.w8(32'h3940c90d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f56dfc),
	.w1(32'hb8d2d0b3),
	.w2(32'hb807931b),
	.w3(32'h390c2b99),
	.w4(32'hb80bf17a),
	.w5(32'h3840d1c6),
	.w6(32'h394a05da),
	.w7(32'h382c1ce2),
	.w8(32'h38e7c1a8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6cda8),
	.w1(32'h3ac5304c),
	.w2(32'h3b2c2039),
	.w3(32'h3b04e49f),
	.w4(32'h3b85b348),
	.w5(32'h3b2081d2),
	.w6(32'h3aefcd18),
	.w7(32'h3a79962b),
	.w8(32'h3a3341d9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08176c),
	.w1(32'hb90aa1b4),
	.w2(32'h381d3b1c),
	.w3(32'hb98f4659),
	.w4(32'hb6c12df4),
	.w5(32'h37118f82),
	.w6(32'hb826a178),
	.w7(32'h398dff32),
	.w8(32'h39b416b2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01b5bb),
	.w1(32'hbac14bca),
	.w2(32'hba554a05),
	.w3(32'hb90f8655),
	.w4(32'hb99a63ff),
	.w5(32'hba483a74),
	.w6(32'h3a2305ba),
	.w7(32'hb821e5bc),
	.w8(32'hb915e6af),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eaf16),
	.w1(32'hbc05c536),
	.w2(32'hbc25da5a),
	.w3(32'hbc3a5cea),
	.w4(32'hbc288a22),
	.w5(32'hbba4a808),
	.w6(32'hbc6dc353),
	.w7(32'hbc35f3c8),
	.w8(32'hbb9aed2f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fe20e),
	.w1(32'h3b03f60c),
	.w2(32'h39bbc5ba),
	.w3(32'h3b3893b6),
	.w4(32'h3b6d0bb3),
	.w5(32'h3adaa40d),
	.w6(32'h3ab31ace),
	.w7(32'h3b1055a3),
	.w8(32'h3a9834bb),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4dfc43),
	.w1(32'h3a9d2c6f),
	.w2(32'hbb2c70bf),
	.w3(32'hb98e77dc),
	.w4(32'h3addedf8),
	.w5(32'h3a513d6a),
	.w6(32'h38eb640c),
	.w7(32'h3b35e1f6),
	.w8(32'hba8469ee),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a4638),
	.w1(32'h3b1f3eb6),
	.w2(32'h3afc2b72),
	.w3(32'h3b4f6e76),
	.w4(32'h3b702ac4),
	.w5(32'h3a96173d),
	.w6(32'h3b2f7966),
	.w7(32'h3b3270f6),
	.w8(32'h3a874e4f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbb100),
	.w1(32'hbb3b91e5),
	.w2(32'hbb2dc3ef),
	.w3(32'hbaecf5d5),
	.w4(32'hba94f189),
	.w5(32'h398ab364),
	.w6(32'hbaf5a0b8),
	.w7(32'hbb82e606),
	.w8(32'hbb2c31a7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ddb72),
	.w1(32'h38a05fdf),
	.w2(32'h3aabf937),
	.w3(32'h3b31b727),
	.w4(32'h3b429d07),
	.w5(32'h3b0a4976),
	.w6(32'h3b0340f4),
	.w7(32'hb8a203a3),
	.w8(32'hba74c99a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e7cd7),
	.w1(32'h3ae482f1),
	.w2(32'h3a065b55),
	.w3(32'h3b2950df),
	.w4(32'h3b5c5f6a),
	.w5(32'h3ad8f2b8),
	.w6(32'h3b3dfa5f),
	.w7(32'h3b0d7743),
	.w8(32'h3af73fdd),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa18606),
	.w1(32'hb9208e8e),
	.w2(32'h398ddbd6),
	.w3(32'h3a63b409),
	.w4(32'hb9c34b42),
	.w5(32'hb7c40833),
	.w6(32'hb98f595f),
	.w7(32'hb9baf4a4),
	.w8(32'h3a5be4d9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa776fd),
	.w1(32'hbad9e7f7),
	.w2(32'hbb792115),
	.w3(32'hbb599599),
	.w4(32'hbb73ac06),
	.w5(32'hbb275122),
	.w6(32'hbb586f38),
	.w7(32'hbb88900a),
	.w8(32'hbba67fec),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba601b24),
	.w1(32'h3a595725),
	.w2(32'hbaabaa40),
	.w3(32'h3b095167),
	.w4(32'h3b8d619e),
	.w5(32'h3b19c126),
	.w6(32'h3a5895e5),
	.w7(32'hbaca54cd),
	.w8(32'hbb607193),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c6e71),
	.w1(32'hbb5d37b1),
	.w2(32'hbc456870),
	.w3(32'hbc0d7321),
	.w4(32'hbc07eadb),
	.w5(32'hbb89ad9f),
	.w6(32'hbc3903ac),
	.w7(32'hbb9df158),
	.w8(32'hbaa5635f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c9254),
	.w1(32'h3c11ee9a),
	.w2(32'h39ed65ea),
	.w3(32'h3c145c62),
	.w4(32'h3c695157),
	.w5(32'h3b365170),
	.w6(32'h3b9eba26),
	.w7(32'h3be20b9e),
	.w8(32'hbb13bc00),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b85f2),
	.w1(32'h3b085580),
	.w2(32'h3b8876a6),
	.w3(32'hba87fd66),
	.w4(32'hb9d5d436),
	.w5(32'h3a1a9995),
	.w6(32'h3a1e702a),
	.w7(32'hb9fca69c),
	.w8(32'hba8a5a2d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b17044),
	.w1(32'h39fe2a46),
	.w2(32'hbbd9f016),
	.w3(32'h3aee81f6),
	.w4(32'h3b0addea),
	.w5(32'h385c29b9),
	.w6(32'hba57d98f),
	.w7(32'h3a893759),
	.w8(32'hbb442221),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ca394),
	.w1(32'h3a925cd4),
	.w2(32'hb9757d32),
	.w3(32'h3afeb7c3),
	.w4(32'h3a95fb75),
	.w5(32'h3a0a689c),
	.w6(32'h3b11a2e0),
	.w7(32'h3a8c95a9),
	.w8(32'h3a8befc6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf425cd),
	.w1(32'hbc2c22a4),
	.w2(32'hbcafd2bd),
	.w3(32'hbc2cf787),
	.w4(32'hbc470612),
	.w5(32'hbc0e4ce4),
	.w6(32'hbc5653ed),
	.w7(32'hbc33ee54),
	.w8(32'hbb98bd9d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf93ab),
	.w1(32'h3a73d42c),
	.w2(32'h399efb27),
	.w3(32'h3a119a0c),
	.w4(32'h3a670706),
	.w5(32'hbaad49fc),
	.w6(32'h3a9d30c8),
	.w7(32'h3b38be54),
	.w8(32'hba2a93b7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39928160),
	.w1(32'h3979d8b7),
	.w2(32'hb86254d5),
	.w3(32'h39c6faf5),
	.w4(32'h39a2e7af),
	.w5(32'hb836499b),
	.w6(32'h39b06cba),
	.w7(32'h395c3880),
	.w8(32'h3858c422),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76397c),
	.w1(32'hb9d5f9bc),
	.w2(32'hb9f6ae5c),
	.w3(32'hb99df3c6),
	.w4(32'h39c14b88),
	.w5(32'h3804cef8),
	.w6(32'hbaf65dee),
	.w7(32'hbaab3ee0),
	.w8(32'hb9832ff4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b307b8f),
	.w1(32'h3b4b4463),
	.w2(32'h3ab35e68),
	.w3(32'hba9ce553),
	.w4(32'hbabb6bdd),
	.w5(32'hba964624),
	.w6(32'hbb1ac0c2),
	.w7(32'hbb1a18cb),
	.w8(32'hbb2421a3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25a9d2),
	.w1(32'hb9d6129b),
	.w2(32'h39266aa9),
	.w3(32'hba1a8a67),
	.w4(32'hba45ceff),
	.w5(32'hbacc4da8),
	.w6(32'h3ac33020),
	.w7(32'hba22bab8),
	.w8(32'hbae8fb3d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaa8e4),
	.w1(32'hba1f477c),
	.w2(32'hbb639e3e),
	.w3(32'h3a66064d),
	.w4(32'hb9a06e3d),
	.w5(32'hbb65cebd),
	.w6(32'h3afddc74),
	.w7(32'hb9c9a72c),
	.w8(32'hbacb6a5e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d065b),
	.w1(32'h3a76cf56),
	.w2(32'hb901568c),
	.w3(32'h38c15a55),
	.w4(32'h3a37b613),
	.w5(32'hbac835c0),
	.w6(32'h370ba8c1),
	.w7(32'hba918177),
	.w8(32'hbb314619),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03c9d8),
	.w1(32'h3ad8ba71),
	.w2(32'h3b034933),
	.w3(32'hbb573d03),
	.w4(32'h3a5338fc),
	.w5(32'h3a2ef60f),
	.w6(32'h37eb3d78),
	.w7(32'h3b9c929d),
	.w8(32'h3b2f4374),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6446ec),
	.w1(32'hbaec134e),
	.w2(32'hbb41dc1f),
	.w3(32'hbadf0ba0),
	.w4(32'hbb160ee2),
	.w5(32'hbb202746),
	.w6(32'hbb96b2a4),
	.w7(32'hbb6439de),
	.w8(32'hbb4084ca),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9245f3),
	.w1(32'h394163b9),
	.w2(32'h3a427565),
	.w3(32'hba08dbea),
	.w4(32'hb880039f),
	.w5(32'hb9d673cb),
	.w6(32'h3a533c4a),
	.w7(32'h398eaec7),
	.w8(32'hba38bb8a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99cc9ec),
	.w1(32'hb8ddbf8a),
	.w2(32'hb8c412c2),
	.w3(32'hb968b9cc),
	.w4(32'hb908616e),
	.w5(32'hb916d2c2),
	.w6(32'hb8e402db),
	.w7(32'hb90bf6dd),
	.w8(32'hb8df1be5),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67edd8e),
	.w1(32'hb83545c1),
	.w2(32'hb968b651),
	.w3(32'h3849f0eb),
	.w4(32'h37383a72),
	.w5(32'hb7d99f3d),
	.w6(32'hb70a5094),
	.w7(32'hb93d19ef),
	.w8(32'hb818e9d0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e90f6),
	.w1(32'hb7d1feab),
	.w2(32'hb862e384),
	.w3(32'h38340693),
	.w4(32'h37283567),
	.w5(32'hb7965f08),
	.w6(32'h38a1e74b),
	.w7(32'h3886a41e),
	.w8(32'h38509415),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39261096),
	.w1(32'h3a1c37a1),
	.w2(32'h3a8530bc),
	.w3(32'h38fea961),
	.w4(32'h3a04b174),
	.w5(32'h3a3d5de1),
	.w6(32'h39159528),
	.w7(32'h391f1713),
	.w8(32'h38e65d72),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85d4323),
	.w1(32'h3ad42592),
	.w2(32'h3b593e78),
	.w3(32'h3a943b03),
	.w4(32'h3af978a7),
	.w5(32'h3b2549ef),
	.w6(32'h3b03f01c),
	.w7(32'h3ae9f8fa),
	.w8(32'h3aeab826),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb822635f),
	.w1(32'h398059a6),
	.w2(32'hba121364),
	.w3(32'h3a28049c),
	.w4(32'h3a789e34),
	.w5(32'hb8a4c62a),
	.w6(32'h3a8a8dda),
	.w7(32'h3a80ae87),
	.w8(32'h38ffe728),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2bf3e),
	.w1(32'hba97d289),
	.w2(32'hbacee9c3),
	.w3(32'hbb0e5f20),
	.w4(32'hbabda262),
	.w5(32'hb9961264),
	.w6(32'hbb140298),
	.w7(32'hba3c51cf),
	.w8(32'hba649b0f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4957f0),
	.w1(32'h3b4f45d6),
	.w2(32'h3b1ba17b),
	.w3(32'h3a6a5a8b),
	.w4(32'h3b2edcbd),
	.w5(32'hbab35242),
	.w6(32'h3b1b6595),
	.w7(32'hb9f58c41),
	.w8(32'hbb680170),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397aeed7),
	.w1(32'h3974c221),
	.w2(32'h38e5bf59),
	.w3(32'h3942b378),
	.w4(32'h3895089e),
	.w5(32'hb8811ea5),
	.w6(32'h390bebf4),
	.w7(32'hb84bd872),
	.w8(32'hb820642f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39290bdf),
	.w1(32'h393aff9b),
	.w2(32'hb8ea5c9e),
	.w3(32'h3950074b),
	.w4(32'h38f69472),
	.w5(32'hb96fff44),
	.w6(32'h392b4794),
	.w7(32'h38be845c),
	.w8(32'hb9820616),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e240fa),
	.w1(32'h381c1696),
	.w2(32'h38af319a),
	.w3(32'h379f3125),
	.w4(32'h3862d713),
	.w5(32'h38ad856c),
	.w6(32'h3710d927),
	.w7(32'h386403db),
	.w8(32'h38d8ef12),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c6982),
	.w1(32'h3a6ff983),
	.w2(32'h3a561a81),
	.w3(32'h3a280df3),
	.w4(32'h39b34cb6),
	.w5(32'hb91196c3),
	.w6(32'h3a433a9a),
	.w7(32'h3964885e),
	.w8(32'hb9ef0e2f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3906602f),
	.w1(32'h3a6ac1ef),
	.w2(32'hba8032e8),
	.w3(32'hbab4110e),
	.w4(32'hbafc6291),
	.w5(32'hbb2c13f1),
	.w6(32'hbb0a3a63),
	.w7(32'h39a38844),
	.w8(32'hbb3d1563),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a233775),
	.w1(32'hba802db4),
	.w2(32'hbac73187),
	.w3(32'hbb20362f),
	.w4(32'hbb05e1ef),
	.w5(32'hb82a6101),
	.w6(32'hba972bd2),
	.w7(32'hbb2d03bc),
	.w8(32'hba320440),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64c5a5e),
	.w1(32'hba753e5f),
	.w2(32'hbae61add),
	.w3(32'hb99c2fa5),
	.w4(32'hba315fba),
	.w5(32'hba49fc30),
	.w6(32'hba7ae2c2),
	.w7(32'hba69706f),
	.w8(32'hba4920e0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb129e7f),
	.w1(32'hbaba7a5b),
	.w2(32'hba25e468),
	.w3(32'hbb1e8371),
	.w4(32'hbacce62b),
	.w5(32'hba65458d),
	.w6(32'hba874002),
	.w7(32'hb9bd6e8b),
	.w8(32'hb8d914dd),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03f46d),
	.w1(32'h39b8b615),
	.w2(32'h39611a0c),
	.w3(32'h394bb7d4),
	.w4(32'h39eb8eab),
	.w5(32'hb7146050),
	.w6(32'h39bcdbe1),
	.w7(32'h39533c8e),
	.w8(32'h385909e2),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80e39c2),
	.w1(32'hb992ffc6),
	.w2(32'hb9ce0d81),
	.w3(32'hbaccd9e5),
	.w4(32'hba5a6d81),
	.w5(32'hb7a594c7),
	.w6(32'hba8ff3eb),
	.w7(32'hbab8e297),
	.w8(32'hb9da766b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0c6b9),
	.w1(32'h3aa4275b),
	.w2(32'h3b593cd9),
	.w3(32'hb5e53022),
	.w4(32'h3b1bb26b),
	.w5(32'h3b004572),
	.w6(32'hb93f22b2),
	.w7(32'hb655a35a),
	.w8(32'h3a203bea),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa65a84),
	.w1(32'hbbc289c5),
	.w2(32'hbc054a00),
	.w3(32'hbbb3d560),
	.w4(32'hbb88f23d),
	.w5(32'hbb174980),
	.w6(32'hbbd3d53c),
	.w7(32'hbbbfc6cd),
	.w8(32'hbb9a4139),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba439bb0),
	.w1(32'h3a5c0fee),
	.w2(32'h3a98f3d3),
	.w3(32'h3aed1132),
	.w4(32'h3a89ba86),
	.w5(32'hba36aebc),
	.w6(32'h3af0681c),
	.w7(32'h3a5ea84d),
	.w8(32'hb83bcc9a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17afee),
	.w1(32'hba8d95e6),
	.w2(32'hbb691552),
	.w3(32'hba12588f),
	.w4(32'h3a545338),
	.w5(32'hbad09db4),
	.w6(32'hbab1fe3a),
	.w7(32'hbadbda6e),
	.w8(32'hbb64e884),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72e549),
	.w1(32'hbb623494),
	.w2(32'hbbaac29c),
	.w3(32'hbb39bf4d),
	.w4(32'hbaf926a4),
	.w5(32'hba8bbe08),
	.w6(32'hbb37d55d),
	.w7(32'hb9d6333b),
	.w8(32'hba547bd9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5e96a),
	.w1(32'h3a882010),
	.w2(32'h3ad57905),
	.w3(32'hba043aa1),
	.w4(32'h371b659f),
	.w5(32'h3982d63b),
	.w6(32'hb94ed636),
	.w7(32'h39d45362),
	.w8(32'h3ab0a05a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73a1a3),
	.w1(32'h37c2e331),
	.w2(32'hba294689),
	.w3(32'h389f30a0),
	.w4(32'hba7b7643),
	.w5(32'hb9f49970),
	.w6(32'h3893d71e),
	.w7(32'hba16b954),
	.w8(32'hbaca1599),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67980c0),
	.w1(32'h39b1a792),
	.w2(32'h38105965),
	.w3(32'hb98e554d),
	.w4(32'h38ac7312),
	.w5(32'hb8b87008),
	.w6(32'hb91b3035),
	.w7(32'hb8bb32cc),
	.w8(32'hb9bb7c45),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cd962),
	.w1(32'h3b1d028b),
	.w2(32'h3ad1b916),
	.w3(32'h3b855cad),
	.w4(32'h3b7b4b12),
	.w5(32'hba406148),
	.w6(32'h3ba50eb0),
	.w7(32'h3b42c222),
	.w8(32'hbb161c0c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba195fc6),
	.w1(32'hb929f574),
	.w2(32'hba8388cb),
	.w3(32'hba8c3fb8),
	.w4(32'hb86a6379),
	.w5(32'hba0beff4),
	.w6(32'hba915552),
	.w7(32'hb8c5634f),
	.w8(32'hb975e3af),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f9112c),
	.w1(32'hb813250b),
	.w2(32'hb7ee4826),
	.w3(32'h37bc549b),
	.w4(32'hb82f7a34),
	.w5(32'hb7a20510),
	.w6(32'h37238963),
	.w7(32'h37dc0ca2),
	.w8(32'hb6bb511a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81e714c),
	.w1(32'hb8929325),
	.w2(32'hb70fb5c7),
	.w3(32'h3861e4da),
	.w4(32'h37916d60),
	.w5(32'hb70a9146),
	.w6(32'h3752a218),
	.w7(32'hb707abed),
	.w8(32'h385de840),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa470cc),
	.w1(32'h39cae25b),
	.w2(32'h3a262acf),
	.w3(32'hba345a9f),
	.w4(32'hb9618ffb),
	.w5(32'hb94d1d04),
	.w6(32'h39eb41f5),
	.w7(32'h3a065483),
	.w8(32'h399b83c6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a183088),
	.w1(32'h3aca1159),
	.w2(32'hbaaa856a),
	.w3(32'h3b348cb5),
	.w4(32'h3ab5a07b),
	.w5(32'hb9952353),
	.w6(32'h3a7ecf2c),
	.w7(32'h39af1f76),
	.w8(32'h37c43f88),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56fea1),
	.w1(32'h3a10c331),
	.w2(32'h3b0f165e),
	.w3(32'hbb7dea59),
	.w4(32'hbb05209f),
	.w5(32'hb8f99924),
	.w6(32'hba83152a),
	.w7(32'hbaf22e1b),
	.w8(32'hba23434b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8169522),
	.w1(32'hb81c7261),
	.w2(32'hb7844fd1),
	.w3(32'hb8406b53),
	.w4(32'hb80ebc75),
	.w5(32'hb6add875),
	.w6(32'hb79fd49a),
	.w7(32'hb781d9e9),
	.w8(32'h374ac5ec),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fcee1),
	.w1(32'h38c17da7),
	.w2(32'h3a186732),
	.w3(32'hbaaaaa15),
	.w4(32'hba80733f),
	.w5(32'h39c92beb),
	.w6(32'hba7abd4d),
	.w7(32'hbb1c8485),
	.w8(32'hbb140984),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fb34c),
	.w1(32'hb939af43),
	.w2(32'h3aa056b8),
	.w3(32'hba1fc4dd),
	.w4(32'hbaf76a4e),
	.w5(32'hbabb0a4d),
	.w6(32'h389b6cbb),
	.w7(32'hbb2e5f04),
	.w8(32'hbb1886fa),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad753d6),
	.w1(32'hbafe50f1),
	.w2(32'hbbc69a1f),
	.w3(32'hbada81db),
	.w4(32'hba82f1fd),
	.w5(32'hbb1b86ae),
	.w6(32'hbb76c8d4),
	.w7(32'hbb200622),
	.w8(32'hbb673845),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb2e42),
	.w1(32'h3a23a883),
	.w2(32'hba14bf48),
	.w3(32'h3aa65b0d),
	.w4(32'h3b4998c7),
	.w5(32'h3985ddbe),
	.w6(32'h3b7b3c62),
	.w7(32'h3a87c353),
	.w8(32'h3880b6e2),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86c51f),
	.w1(32'h3ab95eaa),
	.w2(32'h3a9509ef),
	.w3(32'h3adad6c3),
	.w4(32'h3acdab47),
	.w5(32'hb9119142),
	.w6(32'h3af08bf9),
	.w7(32'h39f07cb7),
	.w8(32'hba3b0637),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b065095),
	.w1(32'h3aee21e3),
	.w2(32'h3a9224d5),
	.w3(32'h3b6b926f),
	.w4(32'h3b329494),
	.w5(32'h3ab71003),
	.w6(32'h3b156db5),
	.w7(32'h3b12be17),
	.w8(32'h3af8ff68),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6a3bb),
	.w1(32'hba389e7b),
	.w2(32'hbb010ba6),
	.w3(32'hba333516),
	.w4(32'hb9dfe695),
	.w5(32'hbb1fdca7),
	.w6(32'h39e44f02),
	.w7(32'h3a583a8d),
	.w8(32'hbaf76281),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3853bf94),
	.w1(32'h3b4e8ea8),
	.w2(32'h3b13e6c3),
	.w3(32'h3b4983d0),
	.w4(32'h3b9ecb05),
	.w5(32'h3b29ebcd),
	.w6(32'h3b5b02c4),
	.w7(32'h3ad79c10),
	.w8(32'h3a4e50c1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa7056),
	.w1(32'h3af5d326),
	.w2(32'h3ad6e9e2),
	.w3(32'h3abaeba6),
	.w4(32'h3b0d7a3a),
	.w5(32'h3abf204f),
	.w6(32'h3a99ff69),
	.w7(32'h3aabb549),
	.w8(32'h3a9a9f9e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37fe6f),
	.w1(32'hbabb5ea5),
	.w2(32'hbaff5c69),
	.w3(32'hba72e9d7),
	.w4(32'hba5db9ba),
	.w5(32'hb98869a4),
	.w6(32'hbadfb1b2),
	.w7(32'hba6a0114),
	.w8(32'hb9b17fdc),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fb4721),
	.w1(32'h39078333),
	.w2(32'h393e0b61),
	.w3(32'h39b90d4f),
	.w4(32'h39c920e6),
	.w5(32'h39563cbd),
	.w6(32'h3957dd22),
	.w7(32'h39660804),
	.w8(32'h383e026f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b68ff),
	.w1(32'hbabf359a),
	.w2(32'hbada1491),
	.w3(32'hbad86977),
	.w4(32'hbaaba412),
	.w5(32'hb9671b10),
	.w6(32'hbb1207c3),
	.w7(32'hbaac68fc),
	.w8(32'hba829066),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949be6b),
	.w1(32'h386f34ef),
	.w2(32'h37ae86c7),
	.w3(32'h3a4f59af),
	.w4(32'h3a3eb7f5),
	.w5(32'h3998e0c5),
	.w6(32'h390892ea),
	.w7(32'h3a2b9a13),
	.w8(32'h38a0b69a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2b86a),
	.w1(32'h381d1a63),
	.w2(32'h3a34fc29),
	.w3(32'hba110dd9),
	.w4(32'h3a313d09),
	.w5(32'h39052805),
	.w6(32'h3a6b0c3c),
	.w7(32'h3ae00295),
	.w8(32'h3a22097b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397daffd),
	.w1(32'h39b05bdf),
	.w2(32'hb98695a6),
	.w3(32'h392435c3),
	.w4(32'h39d1ec25),
	.w5(32'hb9009fe8),
	.w6(32'h39a233ea),
	.w7(32'h3a15cb9a),
	.w8(32'h380ce93a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e52fb),
	.w1(32'h39dd500d),
	.w2(32'h384adb2c),
	.w3(32'h3b6179e7),
	.w4(32'h38d6ab7c),
	.w5(32'hba22369f),
	.w6(32'h3b4a569c),
	.w7(32'hba5ff400),
	.w8(32'hbb3aef89),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a16ea3),
	.w1(32'h39b287e2),
	.w2(32'h399a0b48),
	.w3(32'h398d229c),
	.w4(32'h39a6a3a1),
	.w5(32'h39c89b78),
	.w6(32'h399884da),
	.w7(32'h39a4ddfa),
	.w8(32'h39ede27d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39becb94),
	.w1(32'hb8da4a89),
	.w2(32'hb9d69179),
	.w3(32'h39a59dcd),
	.w4(32'h3978f7ba),
	.w5(32'hb8949cc3),
	.w6(32'h39899945),
	.w7(32'h38d34967),
	.w8(32'hb95e0b5f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7ba3d),
	.w1(32'h3abaeea2),
	.w2(32'hb935e923),
	.w3(32'h3b41743a),
	.w4(32'h3b4906a2),
	.w5(32'h395af903),
	.w6(32'h3b3a749e),
	.w7(32'h3b4e70f0),
	.w8(32'h3a64795c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a397e54),
	.w1(32'h39006bbc),
	.w2(32'hbb48c6d8),
	.w3(32'hbb190dc7),
	.w4(32'hbb242be2),
	.w5(32'hbb272590),
	.w6(32'hbbe5bd93),
	.w7(32'hbb880f18),
	.w8(32'hbb9b4533),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f64f79),
	.w1(32'h3a1f1d66),
	.w2(32'h3a117099),
	.w3(32'h3a74f16d),
	.w4(32'h3a9350e2),
	.w5(32'h39a91942),
	.w6(32'h3a96ce2d),
	.w7(32'h3ab4e7e1),
	.w8(32'h3a0d76a7),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954ea1b),
	.w1(32'h3b0cbebc),
	.w2(32'h385f1367),
	.w3(32'h3ae1fe84),
	.w4(32'h3afd4050),
	.w5(32'hba959d31),
	.w6(32'h3b1ceed1),
	.w7(32'h3a4dddde),
	.w8(32'hba83d2f9),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a423698),
	.w1(32'h3a720ddd),
	.w2(32'h39d023b7),
	.w3(32'h3a7f913d),
	.w4(32'h3a8de997),
	.w5(32'h3972eb06),
	.w6(32'h39d515ee),
	.w7(32'h39097740),
	.w8(32'h385e72bb),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e6c94),
	.w1(32'h3a2e026b),
	.w2(32'hb99be596),
	.w3(32'hbb0014f8),
	.w4(32'h3a22faf6),
	.w5(32'h37ec885d),
	.w6(32'hb93f9ed4),
	.w7(32'hb9b28d28),
	.w8(32'h3a36e7cb),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae971b2),
	.w1(32'hbad011d1),
	.w2(32'hbb35180e),
	.w3(32'hba80edf5),
	.w4(32'hb982fc78),
	.w5(32'hba94fd44),
	.w6(32'hbb04df93),
	.w7(32'hbaad5538),
	.w8(32'hbad926b6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d66caf),
	.w1(32'hbb1851b0),
	.w2(32'hbb6de62b),
	.w3(32'hbb82dff6),
	.w4(32'hbb604a50),
	.w5(32'hbb18337a),
	.w6(32'hbba70a57),
	.w7(32'hbbc50d84),
	.w8(32'hbba6f2de),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20d6fa),
	.w1(32'h3a36a24d),
	.w2(32'h3a0dcb23),
	.w3(32'h3a3ffbba),
	.w4(32'h3a88f767),
	.w5(32'h3a41f601),
	.w6(32'h3a451a8c),
	.w7(32'h3ab82c10),
	.w8(32'h3a9bf358),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397ce488),
	.w1(32'hba725a2c),
	.w2(32'hbad46ae8),
	.w3(32'h3a020cb6),
	.w4(32'h3a01328a),
	.w5(32'hb9480699),
	.w6(32'h3a82b2fe),
	.w7(32'h39c46fbb),
	.w8(32'hba5e8bf2),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c682b6),
	.w1(32'h36eca8f7),
	.w2(32'h3865af21),
	.w3(32'h37b14736),
	.w4(32'hb5a83298),
	.w5(32'h381d9f2b),
	.w6(32'h38524343),
	.w7(32'h374d7bba),
	.w8(32'h3874861d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3777204f),
	.w1(32'h39a118e7),
	.w2(32'h39a7acb0),
	.w3(32'hb98c5e1c),
	.w4(32'h39a3a7ad),
	.w5(32'h399dae5e),
	.w6(32'hb9153f44),
	.w7(32'h392996e2),
	.w8(32'h37d03b03),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3891d990),
	.w1(32'hb8235625),
	.w2(32'h3845149c),
	.w3(32'h39e0c54c),
	.w4(32'h399d87fc),
	.w5(32'hb56e5bfc),
	.w6(32'h39983e39),
	.w7(32'hb8c3f708),
	.w8(32'hb8bd3450),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0528b3),
	.w1(32'hba2360d9),
	.w2(32'hba8a0434),
	.w3(32'hbb078bde),
	.w4(32'hba7b0817),
	.w5(32'hbac895b0),
	.w6(32'hbb21aaee),
	.w7(32'hbb71a44f),
	.w8(32'hbb0a5046),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f0ae50),
	.w1(32'hb65c7c1c),
	.w2(32'h372d2a9c),
	.w3(32'hb72cb593),
	.w4(32'hb72701c6),
	.w5(32'h36e185ec),
	.w6(32'hb6e4e0ee),
	.w7(32'hb71dc5b5),
	.w8(32'h379f515e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a1919),
	.w1(32'hb8e31af6),
	.w2(32'hb98c09b9),
	.w3(32'hb8c51d38),
	.w4(32'hb8dfc313),
	.w5(32'hb9937103),
	.w6(32'hb8be0dd6),
	.w7(32'hb92aa6a3),
	.w8(32'hb9aa3bd1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ce0b7),
	.w1(32'h395a30c6),
	.w2(32'h3a67e311),
	.w3(32'h38fdccc6),
	.w4(32'h3a4a80a3),
	.w5(32'h3a3d8e6b),
	.w6(32'h38f131e5),
	.w7(32'hb8008236),
	.w8(32'h3a48570c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a6828),
	.w1(32'hbaac8440),
	.w2(32'hba84aa03),
	.w3(32'h3b0c7380),
	.w4(32'h3aac703b),
	.w5(32'hb88647cf),
	.w6(32'h3ad2c311),
	.w7(32'hb88b926f),
	.w8(32'hbab12ba6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c9333),
	.w1(32'h3abd41d7),
	.w2(32'hb9a91d5e),
	.w3(32'hba8137cf),
	.w4(32'h3aa7823a),
	.w5(32'h3adfd098),
	.w6(32'hbb1b375b),
	.w7(32'h3ad8bb44),
	.w8(32'h3a33465d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0f906),
	.w1(32'hbb05b264),
	.w2(32'hbb080842),
	.w3(32'hba92e401),
	.w4(32'hba62eee1),
	.w5(32'hbafbf4d6),
	.w6(32'hba7f795c),
	.w7(32'hba124463),
	.w8(32'hba40fda7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed1712),
	.w1(32'hbbd16658),
	.w2(32'hbb60a36d),
	.w3(32'hbbee3cd1),
	.w4(32'hbbe05dee),
	.w5(32'hbb4f449e),
	.w6(32'hbb30d4f2),
	.w7(32'hbb2b898f),
	.w8(32'hbae86f4f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadad2cf),
	.w1(32'h3b106373),
	.w2(32'h3b22982e),
	.w3(32'h3b9fd23f),
	.w4(32'h3bf3644c),
	.w5(32'h3aa5771a),
	.w6(32'h3bc48990),
	.w7(32'h3ad445a2),
	.w8(32'hbaf1daf4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab91d7a),
	.w1(32'h3a8cabff),
	.w2(32'hb9933b09),
	.w3(32'h3a4be60e),
	.w4(32'h3a11fc46),
	.w5(32'h3503fa64),
	.w6(32'h39f41367),
	.w7(32'h398c02f6),
	.w8(32'hba34a54f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83f49b5),
	.w1(32'hb85922d4),
	.w2(32'hb811bb6b),
	.w3(32'hb8c3a033),
	.w4(32'hb8e143ff),
	.w5(32'hb8a906ee),
	.w6(32'hb87f62e9),
	.w7(32'hb8bddf8c),
	.w8(32'hb89a2e5a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b094e),
	.w1(32'hba009ccc),
	.w2(32'hba35f874),
	.w3(32'hb9accfe0),
	.w4(32'hb9c99e6a),
	.w5(32'hba20e3d0),
	.w6(32'hb9df7c4f),
	.w7(32'hb9bc69a6),
	.w8(32'hba1682fa),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38312bb2),
	.w1(32'h35b77615),
	.w2(32'h38543dae),
	.w3(32'h380f152a),
	.w4(32'h3743b77e),
	.w5(32'h38348627),
	.w6(32'h368cfc7f),
	.w7(32'h37a53bf0),
	.w8(32'h3885db43),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b009473),
	.w1(32'h3b1f0892),
	.w2(32'h379237dc),
	.w3(32'h3a88c4f6),
	.w4(32'h3a75cfae),
	.w5(32'hba130733),
	.w6(32'h39de2ced),
	.w7(32'h3a51b709),
	.w8(32'hbabaf82d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918de6e),
	.w1(32'hba919994),
	.w2(32'hbaedfbd1),
	.w3(32'h3a83bfd9),
	.w4(32'h3970fd08),
	.w5(32'hb92e8b32),
	.w6(32'h3a22e0db),
	.w7(32'hbae80769),
	.w8(32'hbb0a69ab),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae29ffa),
	.w1(32'h3ada0919),
	.w2(32'h3b3d57d8),
	.w3(32'hba30eedf),
	.w4(32'h3a6ef0a1),
	.w5(32'h3af9a69b),
	.w6(32'h3a1f15e3),
	.w7(32'h3a5b2511),
	.w8(32'h3b2d8d65),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8648d7),
	.w1(32'hba56c18d),
	.w2(32'hb8e1e21e),
	.w3(32'hb9fb3c75),
	.w4(32'hb902624a),
	.w5(32'h39a474b7),
	.w6(32'hb9c9cdfe),
	.w7(32'h34cf0400),
	.w8(32'h390804c3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e8f66),
	.w1(32'h3a2f13ca),
	.w2(32'hbaf73ff0),
	.w3(32'hbb043e83),
	.w4(32'hba9f77b4),
	.w5(32'hbb2fa2be),
	.w6(32'hb9ff514a),
	.w7(32'hba41dc48),
	.w8(32'hbb606f44),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1162c),
	.w1(32'hba12216a),
	.w2(32'h39beab3f),
	.w3(32'hba948266),
	.w4(32'hb924fefe),
	.w5(32'h384e58d1),
	.w6(32'hba17fd7d),
	.w7(32'h3a5b9505),
	.w8(32'h3a8b6087),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f38446),
	.w1(32'h37dc6c23),
	.w2(32'h388ea5bd),
	.w3(32'h36e181a2),
	.w4(32'h37e40419),
	.w5(32'h388d2808),
	.w6(32'h37eab877),
	.w7(32'h3823bbb5),
	.w8(32'h38aa8a0c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a52c82),
	.w1(32'hbaa2a7be),
	.w2(32'hbad41acf),
	.w3(32'hbb11da35),
	.w4(32'hbb19bf81),
	.w5(32'hba61f0ef),
	.w6(32'hbb05a581),
	.w7(32'hb9618a57),
	.w8(32'h39caa364),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377b6d63),
	.w1(32'hb7f544df),
	.w2(32'h38f0c8b1),
	.w3(32'h38035128),
	.w4(32'hb726f6ae),
	.w5(32'h38dd499d),
	.w6(32'h38cb9d86),
	.w7(32'h37d890df),
	.w8(32'h391960b3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e88f1),
	.w1(32'h3a9079ee),
	.w2(32'hba7b50fb),
	.w3(32'hbb31daa2),
	.w4(32'hb838fbdc),
	.w5(32'hbaa3d5ff),
	.w6(32'hbaa9dfb3),
	.w7(32'h3a3c3486),
	.w8(32'hba81f996),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba567480),
	.w1(32'h3ad0ff04),
	.w2(32'h3b0c3d6f),
	.w3(32'h3b0487a6),
	.w4(32'h3b8b76f4),
	.w5(32'h3b4854fb),
	.w6(32'h3b3b5725),
	.w7(32'h3adef85e),
	.w8(32'h3acd3e9d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f6ccb9),
	.w1(32'h3a853ec0),
	.w2(32'h3a1f4661),
	.w3(32'h3abca51a),
	.w4(32'h3ac49636),
	.w5(32'hb9c57bca),
	.w6(32'h3b1a8c02),
	.w7(32'h3ab82d61),
	.w8(32'hb9bd056c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394810d5),
	.w1(32'h39cfa984),
	.w2(32'hb7b3fe40),
	.w3(32'h3a0a683c),
	.w4(32'h3a40f987),
	.w5(32'hb905e8c2),
	.w6(32'h392fc535),
	.w7(32'h397bb211),
	.w8(32'hb94b395b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a038343),
	.w1(32'h3b121b79),
	.w2(32'h3acc9262),
	.w3(32'h3b24136e),
	.w4(32'h3b24b7c3),
	.w5(32'hb9bca816),
	.w6(32'h3b77829d),
	.w7(32'h3b0e2f9c),
	.w8(32'h39af8b6b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d81a5),
	.w1(32'hba4131ab),
	.w2(32'hba1e773e),
	.w3(32'hbb3eaf98),
	.w4(32'hbb131e51),
	.w5(32'hba7a0a85),
	.w6(32'hbb332a68),
	.w7(32'hbb351a8b),
	.w8(32'hbabfc25e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96b300),
	.w1(32'h39c60453),
	.w2(32'h3ade0302),
	.w3(32'hbb9276d8),
	.w4(32'hbb03a847),
	.w5(32'h39ae7e86),
	.w6(32'hbad623d5),
	.w7(32'hbb2c0b86),
	.w8(32'hba506b40),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e1b3fc),
	.w1(32'hb7eb28cb),
	.w2(32'hb7a12941),
	.w3(32'h38a30601),
	.w4(32'h38ae75d4),
	.w5(32'h3873e80e),
	.w6(32'h38db5a20),
	.w7(32'h38ffbdef),
	.w8(32'h3850528e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38874831),
	.w1(32'h36831841),
	.w2(32'h35fd5894),
	.w3(32'hb910ee51),
	.w4(32'hb93a7317),
	.w5(32'hb77900d8),
	.w6(32'h38cd5cc8),
	.w7(32'h37a6eff7),
	.w8(32'h386cd7b6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e8a52),
	.w1(32'h3ae145c2),
	.w2(32'h3afda6c2),
	.w3(32'h3a4a0a90),
	.w4(32'h39a21a6a),
	.w5(32'hbacca1ef),
	.w6(32'h39dac67f),
	.w7(32'h39a5d640),
	.w8(32'hba55c7f6),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd9eb9),
	.w1(32'hbb440b89),
	.w2(32'hbb61a6ea),
	.w3(32'hbb3107b5),
	.w4(32'hbb69f6f2),
	.w5(32'hbb0cf5c9),
	.w6(32'hbbca48a5),
	.w7(32'hbb82985b),
	.w8(32'hbba00bd1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb256126),
	.w1(32'hb98e0c05),
	.w2(32'h3ae0d52a),
	.w3(32'hbaa21f13),
	.w4(32'hb8873522),
	.w5(32'h390bb15b),
	.w6(32'hb707e626),
	.w7(32'h3a2a8fa8),
	.w8(32'hb9e8996f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b2b88),
	.w1(32'h38f05ce8),
	.w2(32'hb97c70fc),
	.w3(32'h3aa4c44d),
	.w4(32'h3b59ab2d),
	.w5(32'h3b67e68d),
	.w6(32'h3aa26216),
	.w7(32'h39639d64),
	.w8(32'hba2419fc),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37df291c),
	.w1(32'hb9077e7e),
	.w2(32'h3880308e),
	.w3(32'hb8ce3c08),
	.w4(32'hb9a04df0),
	.w5(32'hb93d3ef1),
	.w6(32'hb9470ff6),
	.w7(32'hb9deac56),
	.w8(32'hb9c56970),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b54b2b),
	.w1(32'hb9e78880),
	.w2(32'hb9b38f00),
	.w3(32'hba73aff2),
	.w4(32'hba327cd8),
	.w5(32'hb984cad0),
	.w6(32'hba50aafe),
	.w7(32'hba2bf8b3),
	.w8(32'hb9a01b4e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39969bd2),
	.w1(32'h3ba45ec8),
	.w2(32'hba9d94ab),
	.w3(32'hbaa0741c),
	.w4(32'h39b80a39),
	.w5(32'hbaad0cf9),
	.w6(32'hbb0148e0),
	.w7(32'h3b22b895),
	.w8(32'hbae8775e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb23b10),
	.w1(32'hbbcd8b86),
	.w2(32'hbba1cd4b),
	.w3(32'hbc0a4635),
	.w4(32'hbbb1a22d),
	.w5(32'hbab44412),
	.w6(32'hbb9e9993),
	.w7(32'hbb677343),
	.w8(32'hbaab7429),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395134cd),
	.w1(32'h39c4ec53),
	.w2(32'hbb50268a),
	.w3(32'hbb14e8e4),
	.w4(32'hbb60443f),
	.w5(32'hbb037bc6),
	.w6(32'hbbac7a0a),
	.w7(32'hbb80d92c),
	.w8(32'hbb62a938),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28598d),
	.w1(32'h3ab9085b),
	.w2(32'h3a934f8d),
	.w3(32'h39bb518e),
	.w4(32'h3b12b20d),
	.w5(32'h3a8d165f),
	.w6(32'h3ab0b1df),
	.w7(32'h3ad7a70b),
	.w8(32'h3a3ee0f1),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fbd0d),
	.w1(32'hba5c5ba3),
	.w2(32'h3a1b9dd8),
	.w3(32'hba754ed4),
	.w4(32'h3ac875d1),
	.w5(32'h3a02058d),
	.w6(32'hb82a5bfe),
	.w7(32'hba3b6ec0),
	.w8(32'hb9c03191),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bd1fff),
	.w1(32'h37f9d6d1),
	.w2(32'h3877495a),
	.w3(32'h380864a4),
	.w4(32'h382ce532),
	.w5(32'h3873d7c0),
	.w6(32'h38621c3b),
	.w7(32'h38641cf4),
	.w8(32'h389e7e74),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36edeb5f),
	.w1(32'h36c9f589),
	.w2(32'h37e551cc),
	.w3(32'h36a58c35),
	.w4(32'h36583193),
	.w5(32'h37e31271),
	.w6(32'h376fc4dd),
	.w7(32'h3716273f),
	.w8(32'h380c098c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be1631),
	.w1(32'h399504bb),
	.w2(32'h38f1c0af),
	.w3(32'hb66e64f6),
	.w4(32'h3a1907f3),
	.w5(32'h36dd24fc),
	.w6(32'h3790441a),
	.w7(32'h355da1c8),
	.w8(32'hba1bcc86),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb623d1b9),
	.w1(32'hb761fdb4),
	.w2(32'h37ee3bfa),
	.w3(32'hb7158da0),
	.w4(32'hb72a5e80),
	.w5(32'h37e89758),
	.w6(32'h37addbaa),
	.w7(32'hb4c46f40),
	.w8(32'h37945aa9),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ea486),
	.w1(32'h3a9596bc),
	.w2(32'hb83f8ebc),
	.w3(32'h3a63b95e),
	.w4(32'h3a188113),
	.w5(32'hb9cbc0bf),
	.w6(32'h38b24edf),
	.w7(32'hb641223d),
	.w8(32'hba74a4a9),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d0bc2),
	.w1(32'hbad51c4c),
	.w2(32'hbb6cff85),
	.w3(32'hbabadca5),
	.w4(32'hbad1eb0d),
	.w5(32'hbb244c36),
	.w6(32'hbaf7701e),
	.w7(32'hba57f6e7),
	.w8(32'hbb9d0212),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba683670),
	.w1(32'h38a4a48c),
	.w2(32'hb9faa42e),
	.w3(32'h36c1ba3d),
	.w4(32'h39992e19),
	.w5(32'hba026ed7),
	.w6(32'h3a443223),
	.w7(32'h38b9bf09),
	.w8(32'hbaae7ba4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385b79b1),
	.w1(32'h38cde713),
	.w2(32'h385c96f2),
	.w3(32'h38562515),
	.w4(32'h38c6f0e0),
	.w5(32'h3887fdcf),
	.w6(32'h38924e80),
	.w7(32'h386c1575),
	.w8(32'h3867a7a8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba360ea0),
	.w1(32'hba914aa4),
	.w2(32'hbbddc8f8),
	.w3(32'hbbdd261f),
	.w4(32'hbb9d54b9),
	.w5(32'hbb3763c2),
	.w6(32'hbbe145f9),
	.w7(32'hbb6c2d89),
	.w8(32'hbb710823),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a0889),
	.w1(32'hba3bc1b2),
	.w2(32'hba5e60dd),
	.w3(32'hbab2be17),
	.w4(32'hba9a9f7a),
	.w5(32'hb9bb9f96),
	.w6(32'hba86fd51),
	.w7(32'hbacd1560),
	.w8(32'hbac28d89),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb782a4b2),
	.w1(32'h38583384),
	.w2(32'hb76b2e79),
	.w3(32'hb83533cb),
	.w4(32'hb713b839),
	.w5(32'hb8b9f17e),
	.w6(32'hb89000a9),
	.w7(32'hb81f16aa),
	.w8(32'hb8b0c2c6),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7cd92),
	.w1(32'hbb00e27e),
	.w2(32'hbb275359),
	.w3(32'hbb21d6d2),
	.w4(32'hbb0b5187),
	.w5(32'hbabae3ed),
	.w6(32'hbb290e9e),
	.w7(32'hbaf8745c),
	.w8(32'hbb0dfaf8),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1d3e0),
	.w1(32'h39aa111f),
	.w2(32'h39a86a3c),
	.w3(32'h39b47788),
	.w4(32'h3965efa2),
	.w5(32'h3979d660),
	.w6(32'h395d9488),
	.w7(32'h3943cb37),
	.w8(32'h39363251),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c26ca9),
	.w1(32'h39668dc4),
	.w2(32'hb8e8dbc7),
	.w3(32'h393b3b5f),
	.w4(32'hb38e133e),
	.w5(32'hb8b2aa5a),
	.w6(32'hb96f2fb8),
	.w7(32'hb9ae4c5d),
	.w8(32'hb894d793),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bda40c),
	.w1(32'h3802f4b2),
	.w2(32'h37251884),
	.w3(32'h379dc60c),
	.w4(32'h37865c81),
	.w5(32'h37dacf9f),
	.w6(32'h37f36c1b),
	.w7(32'h382319f5),
	.w8(32'h383f918e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383b6066),
	.w1(32'h3841230b),
	.w2(32'h388c8b3f),
	.w3(32'h388f754d),
	.w4(32'h38360c12),
	.w5(32'h3840dae6),
	.w6(32'h38a73ab4),
	.w7(32'h38b8a71d),
	.w8(32'h38c852e8),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6d72c),
	.w1(32'h3a6a1022),
	.w2(32'h3a79d245),
	.w3(32'hba2d1eed),
	.w4(32'h3a8a13fa),
	.w5(32'h3a95eb77),
	.w6(32'h39967c9f),
	.w7(32'h3a8b4b23),
	.w8(32'h3a40c222),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb863455c),
	.w1(32'hba845c2f),
	.w2(32'hbb017c72),
	.w3(32'hb9d9b647),
	.w4(32'h3a32c55b),
	.w5(32'h392f9ec9),
	.w6(32'hbafba35b),
	.w7(32'hbb4ce2a1),
	.w8(32'hbb1e242f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb9806),
	.w1(32'hbb1cbb57),
	.w2(32'hbb1ad94c),
	.w3(32'hbaf2ad8e),
	.w4(32'hbaaca0aa),
	.w5(32'hb95d89b7),
	.w6(32'hb9a46dfe),
	.w7(32'hba13362d),
	.w8(32'hba81ee3c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba836b45),
	.w1(32'hbad2881a),
	.w2(32'hbaa47d2b),
	.w3(32'hbb47b8b4),
	.w4(32'hba8c1332),
	.w5(32'h3a03b842),
	.w6(32'hbaed3a11),
	.w7(32'hbaee172d),
	.w8(32'hbab1e52d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7731b),
	.w1(32'h3a0e845c),
	.w2(32'h39967552),
	.w3(32'h39ff3c78),
	.w4(32'h3a180588),
	.w5(32'h398a2ba9),
	.w6(32'h39c455c4),
	.w7(32'h3a092f92),
	.w8(32'h399b6595),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939602e),
	.w1(32'h3886a41b),
	.w2(32'h38213305),
	.w3(32'h38af660d),
	.w4(32'hb8fbb6a4),
	.w5(32'hb9243f8d),
	.w6(32'h3730c61b),
	.w7(32'hb8db37eb),
	.w8(32'hb96c7198),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81f597e),
	.w1(32'hb7d3be58),
	.w2(32'hb76fa6cc),
	.w3(32'hb892cf8d),
	.w4(32'hb8aafc19),
	.w5(32'hb800c0c2),
	.w6(32'hb855dc74),
	.w7(32'hb712f11c),
	.w8(32'h37dd9f90),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb695dab6),
	.w1(32'hb843b977),
	.w2(32'hb843fb05),
	.w3(32'h3806d2e3),
	.w4(32'h37a4181e),
	.w5(32'h3620ddfc),
	.w6(32'h3839d4bf),
	.w7(32'h378f3c7c),
	.w8(32'h36058a89),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904b703),
	.w1(32'hbad87e50),
	.w2(32'hbb3e6048),
	.w3(32'hbada5406),
	.w4(32'hbb2c8d62),
	.w5(32'hbb2594cb),
	.w6(32'hbacd2872),
	.w7(32'hbb19ed53),
	.w8(32'hbaf2248b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f0005),
	.w1(32'hba4b7cbc),
	.w2(32'hba4ee558),
	.w3(32'hba4617b8),
	.w4(32'hba83408f),
	.w5(32'hba84155b),
	.w6(32'hba6a64aa),
	.w7(32'hba9ff3c4),
	.w8(32'hbaa325ea),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b3a0d),
	.w1(32'h3a79f533),
	.w2(32'h3a4baf67),
	.w3(32'h3aaaa95f),
	.w4(32'h3aebbbf4),
	.w5(32'h3a880a73),
	.w6(32'h3a9e1119),
	.w7(32'h3a9d8cc4),
	.w8(32'h3a2462fb),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb970bb9e),
	.w1(32'h39a191d8),
	.w2(32'hb6dedb91),
	.w3(32'hb8a4983a),
	.w4(32'h3927e083),
	.w5(32'h371f21a9),
	.w6(32'hb9879f1b),
	.w7(32'h395cce67),
	.w8(32'h3a3d527a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8150ae7),
	.w1(32'hb92511af),
	.w2(32'hb9022890),
	.w3(32'h37e58b69),
	.w4(32'hb8e78fc5),
	.w5(32'hb90ed868),
	.w6(32'h36954965),
	.w7(32'hb918a690),
	.w8(32'hb90fdbc9),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987f78d),
	.w1(32'hb8972af5),
	.w2(32'hba9033d0),
	.w3(32'hb907317f),
	.w4(32'hb9b8faab),
	.w5(32'hba7c78d3),
	.w6(32'h38ce8fbb),
	.w7(32'hb9b6ce2f),
	.w8(32'hba9ac254),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901b36b),
	.w1(32'h38241435),
	.w2(32'hb8d004a9),
	.w3(32'hb8b5732d),
	.w4(32'hb94c23e1),
	.w5(32'hb9004a9b),
	.w6(32'h39056d64),
	.w7(32'hb951d854),
	.w8(32'hb8e7e18d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba8137),
	.w1(32'hbb1bc7ee),
	.w2(32'hbbab5265),
	.w3(32'hbadf73b9),
	.w4(32'hb948a577),
	.w5(32'hbace14f6),
	.w6(32'hbbc69659),
	.w7(32'hbbbaacc5),
	.w8(32'hbb0cddd8),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921c4cf),
	.w1(32'hbacacc13),
	.w2(32'hba743d82),
	.w3(32'h38792247),
	.w4(32'hbaf0a755),
	.w5(32'hbaac08d7),
	.w6(32'hbad6fe1a),
	.w7(32'hba9f0d5d),
	.w8(32'hbaa712b6),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813697),
	.w1(32'hba957635),
	.w2(32'h3a1f0604),
	.w3(32'hbb8269c1),
	.w4(32'hb8739333),
	.w5(32'h3a380480),
	.w6(32'hba75bb5b),
	.w7(32'h3ad582e6),
	.w8(32'h3b06459f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule