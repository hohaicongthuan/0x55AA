module layer_8_featuremap_79(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe731a8),
	.w1(32'hbbb0ce49),
	.w2(32'h3a9a4232),
	.w3(32'h3a394159),
	.w4(32'hbb5701c4),
	.w5(32'hba1cd4a9),
	.w6(32'h39b1789f),
	.w7(32'h3b43a05f),
	.w8(32'h3ae1abcc),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11a59c),
	.w1(32'h3a82e6f6),
	.w2(32'h39f1a5be),
	.w3(32'h3b372662),
	.w4(32'h3b10f485),
	.w5(32'h3a7487a0),
	.w6(32'hba3b084f),
	.w7(32'hb9a41204),
	.w8(32'h3a220ba8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c6d21),
	.w1(32'h3b19f3ec),
	.w2(32'h3ac6d5e8),
	.w3(32'h3b5b131c),
	.w4(32'h3b4a1cf8),
	.w5(32'h3a99ba18),
	.w6(32'hba38624e),
	.w7(32'hb88c9f77),
	.w8(32'h3928e588),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9c0a7),
	.w1(32'hba3dc02b),
	.w2(32'h391a2404),
	.w3(32'hbc025893),
	.w4(32'hbb7ddde6),
	.w5(32'hb8bcba04),
	.w6(32'h3b39fb2f),
	.w7(32'h3abf07c9),
	.w8(32'h3b382645),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b696dac),
	.w1(32'h3b2ae71e),
	.w2(32'h3b004a9d),
	.w3(32'h3b53f6cc),
	.w4(32'h3b506390),
	.w5(32'h3b0ae778),
	.w6(32'h3af7da45),
	.w7(32'h3af82f3e),
	.w8(32'h3b47361b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc95120),
	.w1(32'h3bdcdd32),
	.w2(32'h39986483),
	.w3(32'h3816690a),
	.w4(32'h3b34f606),
	.w5(32'hbb532e51),
	.w6(32'h3b2714d6),
	.w7(32'hba188aeb),
	.w8(32'hbc0539f7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35341d),
	.w1(32'hb9929c43),
	.w2(32'hb9e8d2a5),
	.w3(32'h3a1a49f5),
	.w4(32'h38d448b8),
	.w5(32'hb8cfbe5d),
	.w6(32'hba44dbe3),
	.w7(32'hb9b1296f),
	.w8(32'h3a0d1426),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b3cba),
	.w1(32'h3ab1995d),
	.w2(32'h3b8f5bf6),
	.w3(32'hbb069b45),
	.w4(32'hbb267e7e),
	.w5(32'h3aac4839),
	.w6(32'hbaaabc24),
	.w7(32'h3935278a),
	.w8(32'h3aa57029),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6af29a),
	.w1(32'h3b37eeaa),
	.w2(32'h3b40969a),
	.w3(32'h3b7cab9b),
	.w4(32'h3b59403a),
	.w5(32'h3b4c2615),
	.w6(32'h3aa57d05),
	.w7(32'h3afeabb9),
	.w8(32'h3b63bebe),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d7dfe),
	.w1(32'hbbff0836),
	.w2(32'hbb2a7f72),
	.w3(32'hbbf4fc48),
	.w4(32'hbb8cca57),
	.w5(32'hb984e0cf),
	.w6(32'hbb919d8c),
	.w7(32'hbbc06d48),
	.w8(32'hba80aaad),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada00a6),
	.w1(32'h3afc0bef),
	.w2(32'h3ba65025),
	.w3(32'h3ae50f2e),
	.w4(32'hba6cd21a),
	.w5(32'h3b3ea79a),
	.w6(32'h3baf9ec7),
	.w7(32'h3bb208d7),
	.w8(32'h3b9c4024),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2cb9f),
	.w1(32'hbbeaded1),
	.w2(32'hbb2e7d3a),
	.w3(32'h3a30303f),
	.w4(32'h39ecddf4),
	.w5(32'hb93ca3a8),
	.w6(32'h3b1c561e),
	.w7(32'h3b830bae),
	.w8(32'h3ad888a0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87bb7c),
	.w1(32'h3b90ab45),
	.w2(32'h3b2a5f86),
	.w3(32'h3af5f467),
	.w4(32'h3b415d8a),
	.w5(32'h3b0d3995),
	.w6(32'h3a092a7c),
	.w7(32'h3ae3e27a),
	.w8(32'h3b5b56a9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984704a),
	.w1(32'h3a144058),
	.w2(32'h3b057dd1),
	.w3(32'h39579dc1),
	.w4(32'h3acbb9a0),
	.w5(32'h3a462217),
	.w6(32'h3b1a739d),
	.w7(32'h3b801733),
	.w8(32'h3ac0172d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a018cab),
	.w1(32'h39848bbb),
	.w2(32'h3a4e3b28),
	.w3(32'h39e14382),
	.w4(32'h3a1a9d36),
	.w5(32'h3912fcb8),
	.w6(32'h3a3c5e53),
	.w7(32'h3ad7c58a),
	.w8(32'hba7a8ab1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd6de1),
	.w1(32'hb95fd25d),
	.w2(32'hb8ce92b9),
	.w3(32'hb848d75d),
	.w4(32'h38ae45cd),
	.w5(32'hb8b781ff),
	.w6(32'hba2e70ea),
	.w7(32'hba4b558a),
	.w8(32'hba6c2715),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac769e0),
	.w1(32'hbb2d1d63),
	.w2(32'hba501f82),
	.w3(32'hbb508b66),
	.w4(32'hb7f0a644),
	.w5(32'h3a3284a4),
	.w6(32'hbaf85644),
	.w7(32'hbb307e00),
	.w8(32'hbad22ddc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba917b4c),
	.w1(32'hbb460169),
	.w2(32'h3a300874),
	.w3(32'h3b045dde),
	.w4(32'h3a7ccae5),
	.w5(32'hba769e92),
	.w6(32'h398fa0ea),
	.w7(32'h3b4ff120),
	.w8(32'h3a9c2a36),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccbc7f6),
	.w1(32'hbc5e7f7e),
	.w2(32'h3ba40376),
	.w3(32'h3bd59dd5),
	.w4(32'hbc3813a3),
	.w5(32'h3b3f8057),
	.w6(32'h3c72e197),
	.w7(32'h3c625f0e),
	.w8(32'h3bedee0a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab5eac),
	.w1(32'h39c8bdf4),
	.w2(32'hba7cfca3),
	.w3(32'h3bb374af),
	.w4(32'h399a0725),
	.w5(32'hbb100d49),
	.w6(32'h3b1211b1),
	.w7(32'h3a2d8912),
	.w8(32'hba9ce15d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dd172),
	.w1(32'h3ab6afae),
	.w2(32'h3b19694c),
	.w3(32'h3beaf83d),
	.w4(32'h3b995b2b),
	.w5(32'h3af08d9e),
	.w6(32'h3b474e11),
	.w7(32'h3b76733c),
	.w8(32'h3b3495e9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0e6ff),
	.w1(32'h3b9d7c5e),
	.w2(32'h3b66c843),
	.w3(32'h3b56efd2),
	.w4(32'h3b89fe0c),
	.w5(32'h3b60037a),
	.w6(32'hbadebe89),
	.w7(32'h3931555d),
	.w8(32'hb9e266a1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc39b42),
	.w1(32'hbb9f5bd2),
	.w2(32'h3c5f0ece),
	.w3(32'h3b2c1497),
	.w4(32'hbbb2746f),
	.w5(32'h3bef40bb),
	.w6(32'h3b674640),
	.w7(32'h3bd82a66),
	.w8(32'h3c271dce),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36ea94),
	.w1(32'h3a56e810),
	.w2(32'hb890e785),
	.w3(32'h3b41f490),
	.w4(32'h3acdf81e),
	.w5(32'h39e6396f),
	.w6(32'hba1bf44a),
	.w7(32'hbb08fbe3),
	.w8(32'hbc30618d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbde94a),
	.w1(32'hbbb4c87b),
	.w2(32'hbbb2b8f8),
	.w3(32'hbb23d785),
	.w4(32'hb9be9011),
	.w5(32'hb925b58e),
	.w6(32'hbbede154),
	.w7(32'hbbe0d556),
	.w8(32'hb8f593df),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb640370),
	.w1(32'hbbc4b82e),
	.w2(32'hba80f8a1),
	.w3(32'h3b898429),
	.w4(32'h39323f65),
	.w5(32'h3b039e4e),
	.w6(32'h3c1270cd),
	.w7(32'h3bc97d2b),
	.w8(32'h3b4b61b1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99c485),
	.w1(32'hba0494b9),
	.w2(32'h399b6848),
	.w3(32'hba12d110),
	.w4(32'hba26ddf4),
	.w5(32'h3ac7ab01),
	.w6(32'h3ab69a58),
	.w7(32'h3addec8d),
	.w8(32'hba59eb6a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb40f67),
	.w1(32'hbcd74f91),
	.w2(32'hbc77a6fd),
	.w3(32'h3cbe66ab),
	.w4(32'h3b677eb3),
	.w5(32'hbc8fd5f4),
	.w6(32'h3d2d8e24),
	.w7(32'h3cf4c42a),
	.w8(32'h3c867573),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd81e9d),
	.w1(32'hbb1bf494),
	.w2(32'h3a0ce3c9),
	.w3(32'hb88c2123),
	.w4(32'hbad91f65),
	.w5(32'hbb8e6a35),
	.w6(32'h3c13d5e2),
	.w7(32'h3bd68261),
	.w8(32'h3b091d18),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afad3a1),
	.w1(32'h3ab5f6c2),
	.w2(32'h3a8a785f),
	.w3(32'h3a919e51),
	.w4(32'h3aa5d6cc),
	.w5(32'h3a7fd410),
	.w6(32'h38fe5b71),
	.w7(32'h39c102a9),
	.w8(32'h3a9aa810),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61bebe),
	.w1(32'h3c15b83d),
	.w2(32'h3b802afd),
	.w3(32'hbad9d6aa),
	.w4(32'h3a83ac36),
	.w5(32'hbaba9d02),
	.w6(32'hba51b2e8),
	.w7(32'hba013dfb),
	.w8(32'hbb88c4b2),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3969e70e),
	.w1(32'hba1739d8),
	.w2(32'h39e6d1aa),
	.w3(32'h3b68bec5),
	.w4(32'h3b2aa7db),
	.w5(32'h3b751b02),
	.w6(32'hbb51cc64),
	.w7(32'hbaa61a5c),
	.w8(32'h38932436),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cf514),
	.w1(32'h3b84af75),
	.w2(32'h3b2ea098),
	.w3(32'h3a490051),
	.w4(32'h3b881318),
	.w5(32'h3b5af2a4),
	.w6(32'h3a9db974),
	.w7(32'h3a8dbe9c),
	.w8(32'h3b7e0b9e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e072e),
	.w1(32'h3b0f816c),
	.w2(32'hba10a46c),
	.w3(32'h3b1e8f86),
	.w4(32'h3b4da380),
	.w5(32'h3bc03cae),
	.w6(32'h3ba527f7),
	.w7(32'h3b85cff9),
	.w8(32'h3b20189c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73c0f6),
	.w1(32'h3b696993),
	.w2(32'h3b26fc87),
	.w3(32'h3b1d218a),
	.w4(32'h3b9303f5),
	.w5(32'h3b61466d),
	.w6(32'hbb7944c6),
	.w7(32'hba87d017),
	.w8(32'hbb0308f0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48e9da),
	.w1(32'hbbd12fda),
	.w2(32'hbabaaef8),
	.w3(32'h3b860199),
	.w4(32'hbb11d632),
	.w5(32'hbb0effcd),
	.w6(32'h3b4af751),
	.w7(32'h3b410f93),
	.w8(32'hbac21418),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c0810),
	.w1(32'hbad429d0),
	.w2(32'hbb0eaf5e),
	.w3(32'h3956b556),
	.w4(32'h3a5b5654),
	.w5(32'hb97ac588),
	.w6(32'hbb16962a),
	.w7(32'hbb30d25d),
	.w8(32'h3a08612f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ad75b),
	.w1(32'h3b48aadc),
	.w2(32'h3b39dca3),
	.w3(32'h3b8458ee),
	.w4(32'h3b8798cb),
	.w5(32'h3b401436),
	.w6(32'h3b0b1174),
	.w7(32'h3b42dccf),
	.w8(32'h3ba712cd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92a1af),
	.w1(32'h39c679c9),
	.w2(32'h3aa043be),
	.w3(32'h3aa18685),
	.w4(32'h3a6e1923),
	.w5(32'h39b6de63),
	.w6(32'h3a831102),
	.w7(32'h3b3b79fa),
	.w8(32'hbb2ac57a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82afc7),
	.w1(32'hba3c8e3b),
	.w2(32'hba56c157),
	.w3(32'h390983e8),
	.w4(32'h39f59e45),
	.w5(32'h3a5bcdf4),
	.w6(32'hbb2105b1),
	.w7(32'hbaf9dacd),
	.w8(32'hb933bffa),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20c895),
	.w1(32'hbbe407f6),
	.w2(32'hb96c5097),
	.w3(32'hb9de3ef9),
	.w4(32'h3aff27a9),
	.w5(32'h3b30cbd5),
	.w6(32'h3c86e1a0),
	.w7(32'h3caeb9de),
	.w8(32'h3bb11b87),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dca6b),
	.w1(32'hbb884ded),
	.w2(32'h39866dd3),
	.w3(32'hbc0d1679),
	.w4(32'hbc2900d3),
	.w5(32'hbb1d8640),
	.w6(32'h3ab2ccae),
	.w7(32'hba38601a),
	.w8(32'hbc72f6ac),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc160dce),
	.w1(32'hbc1f7f78),
	.w2(32'h3b039aa5),
	.w3(32'hbbb08710),
	.w4(32'hbbd2bc44),
	.w5(32'hbc8f6026),
	.w6(32'hbc92762b),
	.w7(32'h3c0b2075),
	.w8(32'hbb5eeabe),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1269f9),
	.w1(32'hbb7e053c),
	.w2(32'h3bd3770d),
	.w3(32'hbc47d744),
	.w4(32'hbc7a7c1c),
	.w5(32'hbb64f936),
	.w6(32'h3c15ffd1),
	.w7(32'h3bedd4e9),
	.w8(32'h3a3e9636),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c23b7),
	.w1(32'hbbab6c04),
	.w2(32'h3bf1fe45),
	.w3(32'hbc91c683),
	.w4(32'hbca5d8bd),
	.w5(32'hbb376986),
	.w6(32'h3c3147cd),
	.w7(32'h3c17e535),
	.w8(32'h3a7f0302),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a2a77),
	.w1(32'hbc3e4490),
	.w2(32'hbb8188b8),
	.w3(32'hbc61733c),
	.w4(32'hbc85b4a3),
	.w5(32'hbb786400),
	.w6(32'hbbe9e752),
	.w7(32'hbb8a0192),
	.w8(32'h3bd957a3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1be973),
	.w1(32'hb9fc8a54),
	.w2(32'h3c686cf1),
	.w3(32'hbc07a29e),
	.w4(32'hbb7e462e),
	.w5(32'h3bd10b17),
	.w6(32'hba744386),
	.w7(32'hba73cf20),
	.w8(32'hbb4f725d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8babc6),
	.w1(32'hbc0e063d),
	.w2(32'hbbd1ba83),
	.w3(32'hbc54059b),
	.w4(32'hbcc8399b),
	.w5(32'hbc0c02c3),
	.w6(32'hbb8ec832),
	.w7(32'hbbdfa66f),
	.w8(32'h3b815e9c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e01b5),
	.w1(32'hb9feae5a),
	.w2(32'hbcc4e35b),
	.w3(32'h3d0b9112),
	.w4(32'h3cfef9e1),
	.w5(32'h3b93ad61),
	.w6(32'hbceee9f0),
	.w7(32'hbd057447),
	.w8(32'hbaaf872f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc855a3b),
	.w1(32'hbb867b53),
	.w2(32'h3b80254a),
	.w3(32'hbca38b90),
	.w4(32'hbc8e08d0),
	.w5(32'hbabd2b16),
	.w6(32'h3c3ddafd),
	.w7(32'h3c3d22b1),
	.w8(32'h3aa11d69),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41b45a),
	.w1(32'h3ba9089c),
	.w2(32'h3bc5f296),
	.w3(32'hbb4d5ec0),
	.w4(32'hba86a94c),
	.w5(32'h3a16535d),
	.w6(32'h3bf6f685),
	.w7(32'h3bdbcef2),
	.w8(32'hbbd0dc76),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95ec1f),
	.w1(32'hbc0a074a),
	.w2(32'h3c580e11),
	.w3(32'hbcabf767),
	.w4(32'hbcce8685),
	.w5(32'hbbc0ec39),
	.w6(32'h3ce21c7f),
	.w7(32'h3c91d11a),
	.w8(32'h3cb7d433),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ca6fe),
	.w1(32'hbb2e26ce),
	.w2(32'h3b76ffd0),
	.w3(32'hbcb7940c),
	.w4(32'hbbff987c),
	.w5(32'h3be4ae79),
	.w6(32'hbb4df660),
	.w7(32'hbc0b738b),
	.w8(32'hbb47fab1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8565ef),
	.w1(32'hbbd90f27),
	.w2(32'hbc4c9de2),
	.w3(32'h3b46d997),
	.w4(32'h3bdc64aa),
	.w5(32'h39d40f38),
	.w6(32'hbca40963),
	.w7(32'hbca264f5),
	.w8(32'hbc01ddaa),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2dcf9),
	.w1(32'hbbf331c3),
	.w2(32'h3c4ba169),
	.w3(32'h3c10ab0d),
	.w4(32'hbc52a3c7),
	.w5(32'h3aa33ba3),
	.w6(32'hbc316391),
	.w7(32'h3c8b288c),
	.w8(32'hbc0494e7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67d40f),
	.w1(32'hbc82bc21),
	.w2(32'h3ae77c55),
	.w3(32'hbb97e081),
	.w4(32'hbc1db84f),
	.w5(32'hbb8b9a3f),
	.w6(32'hbc913453),
	.w7(32'hbc7cc4c7),
	.w8(32'h3b8010e5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bae48),
	.w1(32'hbb66d12c),
	.w2(32'h3bc8666d),
	.w3(32'hbbb5f89b),
	.w4(32'hbc138c27),
	.w5(32'h3c424cb4),
	.w6(32'h3af9c732),
	.w7(32'h3b3e6c4e),
	.w8(32'hbc514efe),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6b5b1),
	.w1(32'hbc98f8b3),
	.w2(32'hba94bac1),
	.w3(32'hbc32c60f),
	.w4(32'hbca8b1dd),
	.w5(32'hbbd3d5e1),
	.w6(32'hbc1e0391),
	.w7(32'h3be8c966),
	.w8(32'h3c1f4473),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2905e),
	.w1(32'hbb9f8d59),
	.w2(32'hbbd3696d),
	.w3(32'hbb7d6e79),
	.w4(32'hbbe319ba),
	.w5(32'hbbc1f8cd),
	.w6(32'h3c06829b),
	.w7(32'h3a094c86),
	.w8(32'h3c07c774),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc117b94),
	.w1(32'hbbebe242),
	.w2(32'h3b81087f),
	.w3(32'hbc6cfff8),
	.w4(32'hbbaafa37),
	.w5(32'hbb2c0cac),
	.w6(32'hbbc610a0),
	.w7(32'h3c466ada),
	.w8(32'h3bf10fa1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8500b9),
	.w1(32'hbb2c4fc6),
	.w2(32'hbbca6171),
	.w3(32'h3bb1d49f),
	.w4(32'hbc14a837),
	.w5(32'h3b888cdf),
	.w6(32'h3a29adfc),
	.w7(32'hb9bcd6fa),
	.w8(32'hbbbcbe8e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f8ea0),
	.w1(32'hbbb734fb),
	.w2(32'hbb37679f),
	.w3(32'hbc7ee983),
	.w4(32'hbc25af22),
	.w5(32'hb99b2c0d),
	.w6(32'hbabb57dc),
	.w7(32'h3b5155f5),
	.w8(32'h3a577ec7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd2454d),
	.w1(32'hbbe158c9),
	.w2(32'h3bfd98a4),
	.w3(32'hbcb8665b),
	.w4(32'hbc6f4376),
	.w5(32'hbae62c04),
	.w6(32'h3c84aea0),
	.w7(32'h3c976490),
	.w8(32'hbba764d5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43ac5b),
	.w1(32'hbc752cea),
	.w2(32'hbc8503be),
	.w3(32'hbc7cfe07),
	.w4(32'hbd008fa7),
	.w5(32'hbcc38a8f),
	.w6(32'hbcb48116),
	.w7(32'hbc3f9746),
	.w8(32'h3a7c94ca),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39ca08),
	.w1(32'hb992bfab),
	.w2(32'h3b475ca1),
	.w3(32'hbbe077bf),
	.w4(32'hbc34fc8f),
	.w5(32'hbb130189),
	.w6(32'h3bb75e1b),
	.w7(32'h3b6064d1),
	.w8(32'hb99eca70),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fce54),
	.w1(32'hba737488),
	.w2(32'h3bb84e00),
	.w3(32'hbb94c9de),
	.w4(32'hbbc77a1a),
	.w5(32'h3a3fd3f8),
	.w6(32'h3be536ef),
	.w7(32'h3bc944b0),
	.w8(32'h3ac77cd2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8695d),
	.w1(32'h3ae7f078),
	.w2(32'h3b7acb3e),
	.w3(32'hbbdfcdea),
	.w4(32'hbb86fe0c),
	.w5(32'hba9fca52),
	.w6(32'h3bce10c7),
	.w7(32'h3bacac67),
	.w8(32'h39ba0d56),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77f8f4),
	.w1(32'hbc207a39),
	.w2(32'hbc0d7d38),
	.w3(32'hbb886e63),
	.w4(32'hbb871288),
	.w5(32'h3b2f7892),
	.w6(32'h3b9f4c36),
	.w7(32'hbb35f335),
	.w8(32'hbb8f7230),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0825f1),
	.w1(32'hbaaae718),
	.w2(32'h3b8bbf87),
	.w3(32'hbc61c741),
	.w4(32'hbc4ade9d),
	.w5(32'hbb4964b3),
	.w6(32'h3bd4f515),
	.w7(32'h3bbf5767),
	.w8(32'h3c35129b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdfbc18),
	.w1(32'hbb7c170a),
	.w2(32'h3cd6a02b),
	.w3(32'hbd1a8db7),
	.w4(32'hbd38a797),
	.w5(32'hbc51879b),
	.w6(32'h3d6ae45f),
	.w7(32'h3d49b993),
	.w8(32'h3c0d0871),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd47b03),
	.w1(32'hbaa4fcdf),
	.w2(32'h3b1e0235),
	.w3(32'hbc146590),
	.w4(32'hbbfd4250),
	.w5(32'hbaec570f),
	.w6(32'h3b264599),
	.w7(32'h3ae8ce6a),
	.w8(32'hbb25402f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13a7b2),
	.w1(32'hbabc53fb),
	.w2(32'h3b878a7f),
	.w3(32'hbc4bf937),
	.w4(32'hbc3c7d66),
	.w5(32'hbb4d3bdc),
	.w6(32'h3c047993),
	.w7(32'h3c01d1f9),
	.w8(32'h3908b2a7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d547e),
	.w1(32'hbab538d5),
	.w2(32'h3b74948a),
	.w3(32'hbc5013e6),
	.w4(32'hbc2b942d),
	.w5(32'hbb5e5606),
	.w6(32'h3ba3df87),
	.w7(32'h3b8cd356),
	.w8(32'h3c556b7d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc895f32),
	.w1(32'hbc8b4560),
	.w2(32'hbbdda08b),
	.w3(32'hbc7b9f40),
	.w4(32'hbc87253a),
	.w5(32'hbbf5f52d),
	.w6(32'hba9c289c),
	.w7(32'hbc2ac28f),
	.w8(32'hbb9f23a9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26b2b8),
	.w1(32'hbb843db4),
	.w2(32'hb94a9647),
	.w3(32'hbc7a70b7),
	.w4(32'hbc64bbd9),
	.w5(32'hbbb865f9),
	.w6(32'h3b8e8ab4),
	.w7(32'h3b5b2553),
	.w8(32'hbb6b1c2e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb5af6),
	.w1(32'hbaa05607),
	.w2(32'h3b89f82c),
	.w3(32'hbc17992c),
	.w4(32'hbc1bf50b),
	.w5(32'hbb20b40f),
	.w6(32'h3bb7a457),
	.w7(32'h3b47801e),
	.w8(32'hbb95dc10),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15144d),
	.w1(32'hbb667a67),
	.w2(32'h3a065a8b),
	.w3(32'hbc4f4a34),
	.w4(32'hbc2d37d1),
	.w5(32'hbb5884dd),
	.w6(32'h3ae501c2),
	.w7(32'h3ae93774),
	.w8(32'h3c5dbb97),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd120498),
	.w1(32'hbb7ba8c0),
	.w2(32'h3cacff97),
	.w3(32'hbd15ae6d),
	.w4(32'hbd1aa41d),
	.w5(32'hbc19d8fa),
	.w6(32'h3d88b160),
	.w7(32'h3d6cab8b),
	.w8(32'h3c0bbc21),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce0eed7),
	.w1(32'hbc0c587c),
	.w2(32'h3c6ed6d8),
	.w3(32'hbce64e15),
	.w4(32'hbce9d5d8),
	.w5(32'hbb9ce806),
	.w6(32'h3cbe5049),
	.w7(32'h3c9b4031),
	.w8(32'h3a30b63a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb151dfa),
	.w1(32'hbb95153b),
	.w2(32'h3b3667bd),
	.w3(32'hbb73656b),
	.w4(32'hbc064ac4),
	.w5(32'h3b0a8c39),
	.w6(32'h3b4ba4fa),
	.w7(32'h3b272059),
	.w8(32'h3cbc3dea),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01eaec),
	.w1(32'h3b9e2d91),
	.w2(32'hbbd3de01),
	.w3(32'hbc9a9b34),
	.w4(32'hbc69f9ed),
	.w5(32'hbc0b8132),
	.w6(32'h3c2e6767),
	.w7(32'h3aa58627),
	.w8(32'hbb086d11),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79392c),
	.w1(32'h3a89c99b),
	.w2(32'h3b9eea73),
	.w3(32'hbc5cfd39),
	.w4(32'hbc4ed97f),
	.w5(32'hbb94e280),
	.w6(32'h3b191fe4),
	.w7(32'h3a8da72c),
	.w8(32'h3adbc57d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc588e08),
	.w1(32'hbba91622),
	.w2(32'h3ba5d03c),
	.w3(32'hbc9fe04d),
	.w4(32'hbca4f254),
	.w5(32'hbb6b64be),
	.w6(32'h3c40e2a2),
	.w7(32'h3c33a57e),
	.w8(32'h3cf36792),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd7745),
	.w1(32'hbc75d65a),
	.w2(32'hbbd6bd24),
	.w3(32'hbba96fff),
	.w4(32'h3c6185df),
	.w5(32'h3bed269a),
	.w6(32'h3c7a8770),
	.w7(32'h3b1f266b),
	.w8(32'hbc084d4e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb57a50),
	.w1(32'hbc56ff4d),
	.w2(32'hbbb83f59),
	.w3(32'hbab95af0),
	.w4(32'hbc0796a4),
	.w5(32'hbbddb76a),
	.w6(32'hb95e4622),
	.w7(32'hba98f2da),
	.w8(32'h3bdc6292),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8965bd),
	.w1(32'hbbb3212d),
	.w2(32'h3bc8dbe2),
	.w3(32'hbcb568ad),
	.w4(32'hbc949f09),
	.w5(32'hbbadd582),
	.w6(32'h3c3f4525),
	.w7(32'h3c10138c),
	.w8(32'h3bd8b43e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc68f2),
	.w1(32'hbb3a43ac),
	.w2(32'hbd0f0e83),
	.w3(32'h3d34fd18),
	.w4(32'h3d1fb704),
	.w5(32'h3b83fea7),
	.w6(32'hbd1eea96),
	.w7(32'hbd394ae7),
	.w8(32'h3aa9b7b0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb957489),
	.w1(32'hba2665de),
	.w2(32'hba866935),
	.w3(32'hbc0420dc),
	.w4(32'hbc6b691f),
	.w5(32'hbb76606d),
	.w6(32'h3bc1ce78),
	.w7(32'hbaa80706),
	.w8(32'h3ad55582),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c3201),
	.w1(32'hbc17543e),
	.w2(32'hbbdf4128),
	.w3(32'hbca45c83),
	.w4(32'hbc255e4d),
	.w5(32'hbc0212e0),
	.w6(32'hbb478ced),
	.w7(32'h3ac89cd6),
	.w8(32'h3a90c5c8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe097d),
	.w1(32'hbb6ccd5d),
	.w2(32'hbd0799d2),
	.w3(32'h3d2518a4),
	.w4(32'h3d0eceec),
	.w5(32'h3b3c951a),
	.w6(32'hbd12d839),
	.w7(32'hbd2cf1e9),
	.w8(32'h3a91e9c7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9144c7),
	.w1(32'hbb87d5f8),
	.w2(32'hbcf06ba5),
	.w3(32'h3d096135),
	.w4(32'h3ce917e5),
	.w5(32'h39e10626),
	.w6(32'hbd064c1e),
	.w7(32'hbd1988f6),
	.w8(32'hbbe9da56),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d97eb7),
	.w1(32'hbb7977a3),
	.w2(32'hbc24ad97),
	.w3(32'hbab3c7fe),
	.w4(32'h3b18339f),
	.w5(32'hbb8e572b),
	.w6(32'hbc40ab0c),
	.w7(32'hbc3dd1c4),
	.w8(32'h3c78c29e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be84c6d),
	.w1(32'hbb669dc9),
	.w2(32'h3bb5c8c4),
	.w3(32'hbc6ade1b),
	.w4(32'hbcc75f5a),
	.w5(32'h3c3b983e),
	.w6(32'hbb8a2056),
	.w7(32'hbc75ddfa),
	.w8(32'h399bca3c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0996c),
	.w1(32'hba31e579),
	.w2(32'h3b86eed3),
	.w3(32'hbb9dfb9f),
	.w4(32'hbb92d80f),
	.w5(32'hba5ad1ea),
	.w6(32'h3bdba8df),
	.w7(32'h3bca780f),
	.w8(32'hbb755d44),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b976868),
	.w1(32'hbb92a0bd),
	.w2(32'hbc076dc5),
	.w3(32'hbb147b20),
	.w4(32'hbb91525c),
	.w5(32'hbc1e3f85),
	.w6(32'h39401060),
	.w7(32'hbb5f649b),
	.w8(32'hbc6cde9a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56bb27),
	.w1(32'hbc9bc4d0),
	.w2(32'hbca7efcf),
	.w3(32'hbcaae546),
	.w4(32'hbcb23b47),
	.w5(32'hbce57a25),
	.w6(32'hbcb3e734),
	.w7(32'hbc81f2b4),
	.w8(32'hbc6492c4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3509db),
	.w1(32'hbb78dc8f),
	.w2(32'hbbb341ba),
	.w3(32'hbacdb630),
	.w4(32'hbba4ea22),
	.w5(32'hbbbc3078),
	.w6(32'hbb841e8f),
	.w7(32'hbbb53fc6),
	.w8(32'hbb127478),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f1301),
	.w1(32'hbb240397),
	.w2(32'hb96a15e1),
	.w3(32'h3bacdf57),
	.w4(32'h3c347674),
	.w5(32'hbbb45f99),
	.w6(32'hbc30dd30),
	.w7(32'hbb961fe3),
	.w8(32'h3c40a39e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccbed5b),
	.w1(32'h3a99943d),
	.w2(32'h3c954672),
	.w3(32'hbd07449d),
	.w4(32'hbcfceb6a),
	.w5(32'hbbe5409a),
	.w6(32'h3d4e6ef5),
	.w7(32'h3d2ca66c),
	.w8(32'h39b30aae),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed02bf),
	.w1(32'hbb12352d),
	.w2(32'h3b97e984),
	.w3(32'hbc47e08c),
	.w4(32'hbc760f8e),
	.w5(32'hbb38a4ea),
	.w6(32'h3ba30f21),
	.w7(32'h3b66e300),
	.w8(32'h3ba53e77),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe72854),
	.w1(32'hbc30bd7b),
	.w2(32'hbbc9456c),
	.w3(32'hbc75213d),
	.w4(32'hbc162bda),
	.w5(32'hbba1d92b),
	.w6(32'hbc1f136b),
	.w7(32'h3b630452),
	.w8(32'hba102f55),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87dabd),
	.w1(32'h3afb333a),
	.w2(32'h3bb580a6),
	.w3(32'hbc02c964),
	.w4(32'hbbd25da6),
	.w5(32'hbae80c86),
	.w6(32'h3bd75a4b),
	.w7(32'h3bba2caf),
	.w8(32'hbb2ba44e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0a7ee3),
	.w1(32'hbba2f113),
	.w2(32'h3ca8f8f1),
	.w3(32'hbd47dd59),
	.w4(32'hbd43d052),
	.w5(32'hbc5435ab),
	.w6(32'h3d4c26e9),
	.w7(32'h3d35596b),
	.w8(32'hbba9f882),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9ea8a),
	.w1(32'hbbc2e546),
	.w2(32'hbc2c4fa2),
	.w3(32'hbbb519b2),
	.w4(32'hbaab61e6),
	.w5(32'hbbf9ac32),
	.w6(32'hbc6abeb1),
	.w7(32'hbc4d4714),
	.w8(32'h3a6d126b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d2400),
	.w1(32'hba2a7a25),
	.w2(32'hbc55e5fc),
	.w3(32'h3c803fa4),
	.w4(32'h3c6d0eaa),
	.w5(32'h3a90e37a),
	.w6(32'hbc9c5cc3),
	.w7(32'hbca77a82),
	.w8(32'hbadf1722),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1a1d2),
	.w1(32'hbb3100dc),
	.w2(32'h3b572895),
	.w3(32'h3ad2e64c),
	.w4(32'hbb8214b5),
	.w5(32'hbae838da),
	.w6(32'h3bcde9c7),
	.w7(32'h3b8bee84),
	.w8(32'h3b0b07eb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1feddb),
	.w1(32'hba38bc3a),
	.w2(32'hba9d5f63),
	.w3(32'hbae2c216),
	.w4(32'hb9645474),
	.w5(32'hb9f31feb),
	.w6(32'h3b26717b),
	.w7(32'hb9a632b0),
	.w8(32'h3af5bed1),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37148b),
	.w1(32'h3ac8986d),
	.w2(32'h3a266326),
	.w3(32'h38375572),
	.w4(32'hba6de4b1),
	.w5(32'hba98078c),
	.w6(32'hbae3b7ee),
	.w7(32'hbab0e703),
	.w8(32'hbacf7b18),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b3496),
	.w1(32'hba8289a4),
	.w2(32'hbaa4690b),
	.w3(32'hbb09490c),
	.w4(32'hbaec84ce),
	.w5(32'hbafaf2cb),
	.w6(32'hbb7d0256),
	.w7(32'hbb57b2d6),
	.w8(32'hbaeb8b41),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ac2fe),
	.w1(32'h3ab1fe6b),
	.w2(32'h3acd81d2),
	.w3(32'h3a950b4b),
	.w4(32'h3b08b142),
	.w5(32'h3b13caff),
	.w6(32'h3ae92f5b),
	.w7(32'h3abe105a),
	.w8(32'h39a1decb),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d5f43),
	.w1(32'hbabc711d),
	.w2(32'hbadc6d5d),
	.w3(32'h3b1aceae),
	.w4(32'h3a411e6d),
	.w5(32'h3b0151f0),
	.w6(32'hbac1e50c),
	.w7(32'hbaab7894),
	.w8(32'hbb8604b3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3d7c3),
	.w1(32'hbb14f993),
	.w2(32'hbb091d48),
	.w3(32'hbacb28ca),
	.w4(32'hba5bcb8e),
	.w5(32'hba9a71a0),
	.w6(32'hbaa72dd7),
	.w7(32'hba0187b7),
	.w8(32'hba25754e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8438c4),
	.w1(32'h3b8c64ae),
	.w2(32'h3b708818),
	.w3(32'hba2fa06f),
	.w4(32'h3b3cda3a),
	.w5(32'h3b53f74e),
	.w6(32'hbb9d027a),
	.w7(32'hbb0dbe26),
	.w8(32'hbad2f184),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39164ecf),
	.w1(32'h39deed3f),
	.w2(32'h3a947d2a),
	.w3(32'h3a6a51a1),
	.w4(32'h3a90c90d),
	.w5(32'h3aa7f61d),
	.w6(32'h3a766d7e),
	.w7(32'h3ab4d4dd),
	.w8(32'h39ab9e97),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba235f9e),
	.w1(32'hba8b1bd6),
	.w2(32'hba9b9844),
	.w3(32'hb9c2b52a),
	.w4(32'hba9f8538),
	.w5(32'hba8fef06),
	.w6(32'hb9d2e3b2),
	.w7(32'hba3d1485),
	.w8(32'hb902772b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397131db),
	.w1(32'h39940b84),
	.w2(32'hb97a8599),
	.w3(32'h3a4d090f),
	.w4(32'h399056dd),
	.w5(32'h39758f7b),
	.w6(32'h3a95f8fb),
	.w7(32'h3aa14ac7),
	.w8(32'hbaf081da),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba554cc2),
	.w1(32'h3a4a6b33),
	.w2(32'hbb94faca),
	.w3(32'hba8ac62f),
	.w4(32'h3aaf5f35),
	.w5(32'hbb34e616),
	.w6(32'hba86f5d8),
	.w7(32'hbbacbe4d),
	.w8(32'h3b5cb8a6),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbb1e1),
	.w1(32'hbb3a2433),
	.w2(32'h3a293c58),
	.w3(32'hba0f5970),
	.w4(32'hbb0e3122),
	.w5(32'h39573168),
	.w6(32'h3b7d2b70),
	.w7(32'h3b7cd298),
	.w8(32'hba9858fc),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04be0d),
	.w1(32'h38315823),
	.w2(32'hb9d33ccf),
	.w3(32'h3a056b56),
	.w4(32'h38dec1bb),
	.w5(32'h3a1ee1fa),
	.w6(32'hba373380),
	.w7(32'hbaae2fe8),
	.w8(32'h3ad9dcb8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6f090),
	.w1(32'h3a2ff1f3),
	.w2(32'hb8938aea),
	.w3(32'hb8dd83e9),
	.w4(32'hba8d3417),
	.w5(32'h396c5cfa),
	.w6(32'h3a5a76bf),
	.w7(32'h38b7d1c5),
	.w8(32'h3a115ced),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a956648),
	.w1(32'h3a6c7e25),
	.w2(32'h3b8509af),
	.w3(32'hbbb25334),
	.w4(32'hbb894353),
	.w5(32'hba663b90),
	.w6(32'hbc2d33ad),
	.w7(32'hbbfbd2ca),
	.w8(32'hbb3b5434),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57d17c),
	.w1(32'h399334ca),
	.w2(32'h39df864d),
	.w3(32'h3bafc1de),
	.w4(32'h3b8504ad),
	.w5(32'h3b763ba8),
	.w6(32'h3bd8527e),
	.w7(32'h3bae94e4),
	.w8(32'h3a4da785),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85dc9e),
	.w1(32'hb9953666),
	.w2(32'hb6fff9f3),
	.w3(32'hba0bfc02),
	.w4(32'h3a115344),
	.w5(32'h39d73e43),
	.w6(32'hba79cc5f),
	.w7(32'hba7e3fb4),
	.w8(32'h3a9de8f1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0de69a),
	.w1(32'h3bc5a12a),
	.w2(32'h3a91762e),
	.w3(32'hb897e264),
	.w4(32'h3b3bc546),
	.w5(32'hb9096d32),
	.w6(32'h3a5d1bb9),
	.w7(32'hbb4124b5),
	.w8(32'hbb9910dc),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0f24a),
	.w1(32'h3b646dc1),
	.w2(32'h3b35996d),
	.w3(32'h3b06d4b8),
	.w4(32'h3b7060a2),
	.w5(32'h3b704e6c),
	.w6(32'hbaafd87d),
	.w7(32'h3970480c),
	.w8(32'h3ad648c0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23f54f),
	.w1(32'hbae045a3),
	.w2(32'hbb1ea303),
	.w3(32'hbb05e7cf),
	.w4(32'hbadaa3cc),
	.w5(32'hbb7a14a2),
	.w6(32'hbb306104),
	.w7(32'hbb0b4e2b),
	.w8(32'hbb8f16dd),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03870b),
	.w1(32'hbb14e271),
	.w2(32'hba36a0f2),
	.w3(32'hb9d898d6),
	.w4(32'hba668e93),
	.w5(32'hba69c7c0),
	.w6(32'hba9c47db),
	.w7(32'hbaa9a327),
	.w8(32'hba3d0bd4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb077708),
	.w1(32'hbb255dd9),
	.w2(32'hbaa5e299),
	.w3(32'hbb43335e),
	.w4(32'hbb97f480),
	.w5(32'hbb756f0b),
	.w6(32'hba3e8726),
	.w7(32'hbb85370a),
	.w8(32'h3a8a2f4c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule